library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(10239 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);
    signal layer1_outputs : std_logic_vector(10239 downto 0);
    signal layer2_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= inputs(106);
    layer0_outputs(1) <= (inputs(108)) xor (inputs(107));
    layer0_outputs(2) <= not(inputs(104));
    layer0_outputs(3) <= inputs(116);
    layer0_outputs(4) <= not((inputs(154)) and (inputs(119)));
    layer0_outputs(5) <= inputs(128);
    layer0_outputs(6) <= not(inputs(189)) or (inputs(61));
    layer0_outputs(7) <= (inputs(32)) and not (inputs(113));
    layer0_outputs(8) <= not(inputs(80)) or (inputs(254));
    layer0_outputs(9) <= not(inputs(82));
    layer0_outputs(10) <= not((inputs(111)) xor (inputs(154)));
    layer0_outputs(11) <= (inputs(72)) xor (inputs(118));
    layer0_outputs(12) <= (inputs(45)) and not (inputs(152));
    layer0_outputs(13) <= inputs(183);
    layer0_outputs(14) <= inputs(22);
    layer0_outputs(15) <= inputs(126);
    layer0_outputs(16) <= not((inputs(204)) xor (inputs(114)));
    layer0_outputs(17) <= not((inputs(59)) or (inputs(79)));
    layer0_outputs(18) <= not(inputs(69));
    layer0_outputs(19) <= not(inputs(101));
    layer0_outputs(20) <= not((inputs(223)) or (inputs(172)));
    layer0_outputs(21) <= not(inputs(24));
    layer0_outputs(22) <= (inputs(156)) or (inputs(128));
    layer0_outputs(23) <= inputs(3);
    layer0_outputs(24) <= (inputs(62)) or (inputs(126));
    layer0_outputs(25) <= not((inputs(198)) or (inputs(48)));
    layer0_outputs(26) <= '0';
    layer0_outputs(27) <= (inputs(160)) or (inputs(185));
    layer0_outputs(28) <= '1';
    layer0_outputs(29) <= not(inputs(120)) or (inputs(243));
    layer0_outputs(30) <= not(inputs(56));
    layer0_outputs(31) <= (inputs(86)) and (inputs(119));
    layer0_outputs(32) <= (inputs(167)) and not (inputs(101));
    layer0_outputs(33) <= not(inputs(123));
    layer0_outputs(34) <= not(inputs(113));
    layer0_outputs(35) <= (inputs(232)) and (inputs(152));
    layer0_outputs(36) <= inputs(7);
    layer0_outputs(37) <= not(inputs(27));
    layer0_outputs(38) <= not((inputs(127)) or (inputs(82)));
    layer0_outputs(39) <= not((inputs(117)) and (inputs(11)));
    layer0_outputs(40) <= not(inputs(189)) or (inputs(61));
    layer0_outputs(41) <= not(inputs(23)) or (inputs(82));
    layer0_outputs(42) <= not(inputs(133)) or (inputs(18));
    layer0_outputs(43) <= not((inputs(66)) or (inputs(36)));
    layer0_outputs(44) <= not((inputs(219)) or (inputs(206)));
    layer0_outputs(45) <= not(inputs(66)) or (inputs(178));
    layer0_outputs(46) <= not(inputs(187)) or (inputs(250));
    layer0_outputs(47) <= (inputs(233)) and not (inputs(18));
    layer0_outputs(48) <= not((inputs(157)) or (inputs(135)));
    layer0_outputs(49) <= (inputs(74)) and not (inputs(23));
    layer0_outputs(50) <= (inputs(140)) and (inputs(125));
    layer0_outputs(51) <= not(inputs(18));
    layer0_outputs(52) <= inputs(246);
    layer0_outputs(53) <= not(inputs(115)) or (inputs(49));
    layer0_outputs(54) <= (inputs(8)) and not (inputs(226));
    layer0_outputs(55) <= not((inputs(216)) or (inputs(158)));
    layer0_outputs(56) <= not((inputs(98)) or (inputs(167)));
    layer0_outputs(57) <= not((inputs(23)) or (inputs(109)));
    layer0_outputs(58) <= inputs(158);
    layer0_outputs(59) <= not(inputs(244)) or (inputs(13));
    layer0_outputs(60) <= not(inputs(219));
    layer0_outputs(61) <= inputs(14);
    layer0_outputs(62) <= (inputs(191)) and (inputs(252));
    layer0_outputs(63) <= (inputs(21)) and not (inputs(98));
    layer0_outputs(64) <= not(inputs(75)) or (inputs(204));
    layer0_outputs(65) <= inputs(75);
    layer0_outputs(66) <= inputs(166);
    layer0_outputs(67) <= '1';
    layer0_outputs(68) <= inputs(248);
    layer0_outputs(69) <= (inputs(23)) and (inputs(137));
    layer0_outputs(70) <= not(inputs(22));
    layer0_outputs(71) <= (inputs(207)) or (inputs(35));
    layer0_outputs(72) <= not((inputs(198)) or (inputs(185)));
    layer0_outputs(73) <= (inputs(6)) or (inputs(251));
    layer0_outputs(74) <= (inputs(33)) or (inputs(234));
    layer0_outputs(75) <= (inputs(246)) or (inputs(65));
    layer0_outputs(76) <= inputs(60);
    layer0_outputs(77) <= inputs(30);
    layer0_outputs(78) <= not(inputs(200)) or (inputs(77));
    layer0_outputs(79) <= inputs(243);
    layer0_outputs(80) <= not((inputs(131)) xor (inputs(128)));
    layer0_outputs(81) <= not(inputs(24));
    layer0_outputs(82) <= (inputs(217)) and not (inputs(194));
    layer0_outputs(83) <= (inputs(88)) and not (inputs(189));
    layer0_outputs(84) <= inputs(74);
    layer0_outputs(85) <= not(inputs(193));
    layer0_outputs(86) <= not(inputs(125));
    layer0_outputs(87) <= inputs(77);
    layer0_outputs(88) <= not((inputs(100)) xor (inputs(89)));
    layer0_outputs(89) <= not((inputs(253)) or (inputs(107)));
    layer0_outputs(90) <= not(inputs(150));
    layer0_outputs(91) <= not(inputs(169));
    layer0_outputs(92) <= (inputs(13)) or (inputs(244));
    layer0_outputs(93) <= not((inputs(232)) or (inputs(145)));
    layer0_outputs(94) <= not(inputs(226));
    layer0_outputs(95) <= not(inputs(195));
    layer0_outputs(96) <= '0';
    layer0_outputs(97) <= inputs(73);
    layer0_outputs(98) <= not(inputs(149)) or (inputs(33));
    layer0_outputs(99) <= not((inputs(225)) or (inputs(166)));
    layer0_outputs(100) <= (inputs(127)) and not (inputs(87));
    layer0_outputs(101) <= (inputs(103)) or (inputs(162));
    layer0_outputs(102) <= not(inputs(179)) or (inputs(78));
    layer0_outputs(103) <= not(inputs(127));
    layer0_outputs(104) <= not(inputs(18));
    layer0_outputs(105) <= not(inputs(69));
    layer0_outputs(106) <= not(inputs(69));
    layer0_outputs(107) <= not(inputs(6));
    layer0_outputs(108) <= (inputs(104)) and not (inputs(137));
    layer0_outputs(109) <= not((inputs(0)) or (inputs(4)));
    layer0_outputs(110) <= '1';
    layer0_outputs(111) <= not(inputs(131));
    layer0_outputs(112) <= not((inputs(149)) or (inputs(210)));
    layer0_outputs(113) <= not(inputs(93));
    layer0_outputs(114) <= not(inputs(16));
    layer0_outputs(115) <= not((inputs(178)) or (inputs(221)));
    layer0_outputs(116) <= inputs(97);
    layer0_outputs(117) <= not(inputs(137));
    layer0_outputs(118) <= not((inputs(57)) or (inputs(49)));
    layer0_outputs(119) <= (inputs(11)) and (inputs(14));
    layer0_outputs(120) <= inputs(177);
    layer0_outputs(121) <= inputs(193);
    layer0_outputs(122) <= inputs(91);
    layer0_outputs(123) <= not(inputs(173));
    layer0_outputs(124) <= not((inputs(135)) xor (inputs(31)));
    layer0_outputs(125) <= (inputs(57)) or (inputs(177));
    layer0_outputs(126) <= not((inputs(242)) or (inputs(36)));
    layer0_outputs(127) <= (inputs(164)) or (inputs(64));
    layer0_outputs(128) <= '0';
    layer0_outputs(129) <= not((inputs(205)) xor (inputs(122)));
    layer0_outputs(130) <= not(inputs(195));
    layer0_outputs(131) <= not((inputs(96)) or (inputs(125)));
    layer0_outputs(132) <= inputs(115);
    layer0_outputs(133) <= inputs(211);
    layer0_outputs(134) <= (inputs(211)) and not (inputs(99));
    layer0_outputs(135) <= not(inputs(150));
    layer0_outputs(136) <= not((inputs(70)) and (inputs(189)));
    layer0_outputs(137) <= inputs(99);
    layer0_outputs(138) <= (inputs(74)) xor (inputs(125));
    layer0_outputs(139) <= not(inputs(150));
    layer0_outputs(140) <= inputs(151);
    layer0_outputs(141) <= not((inputs(60)) or (inputs(121)));
    layer0_outputs(142) <= (inputs(187)) xor (inputs(172));
    layer0_outputs(143) <= not((inputs(138)) and (inputs(172)));
    layer0_outputs(144) <= inputs(5);
    layer0_outputs(145) <= not(inputs(120));
    layer0_outputs(146) <= not(inputs(111)) or (inputs(80));
    layer0_outputs(147) <= not(inputs(136)) or (inputs(28));
    layer0_outputs(148) <= inputs(116);
    layer0_outputs(149) <= (inputs(185)) or (inputs(178));
    layer0_outputs(150) <= inputs(201);
    layer0_outputs(151) <= not(inputs(195));
    layer0_outputs(152) <= not(inputs(100));
    layer0_outputs(153) <= (inputs(43)) and not (inputs(254));
    layer0_outputs(154) <= (inputs(117)) xor (inputs(183));
    layer0_outputs(155) <= (inputs(8)) and (inputs(200));
    layer0_outputs(156) <= (inputs(116)) or (inputs(132));
    layer0_outputs(157) <= inputs(157);
    layer0_outputs(158) <= not(inputs(111));
    layer0_outputs(159) <= (inputs(119)) and not (inputs(62));
    layer0_outputs(160) <= not(inputs(44));
    layer0_outputs(161) <= not((inputs(246)) or (inputs(159)));
    layer0_outputs(162) <= '1';
    layer0_outputs(163) <= not(inputs(200)) or (inputs(112));
    layer0_outputs(164) <= not((inputs(119)) or (inputs(214)));
    layer0_outputs(165) <= not((inputs(158)) or (inputs(222)));
    layer0_outputs(166) <= inputs(81);
    layer0_outputs(167) <= not((inputs(83)) or (inputs(76)));
    layer0_outputs(168) <= inputs(109);
    layer0_outputs(169) <= not((inputs(30)) or (inputs(5)));
    layer0_outputs(170) <= not((inputs(207)) and (inputs(31)));
    layer0_outputs(171) <= inputs(57);
    layer0_outputs(172) <= '1';
    layer0_outputs(173) <= inputs(229);
    layer0_outputs(174) <= (inputs(252)) or (inputs(140));
    layer0_outputs(175) <= (inputs(32)) or (inputs(183));
    layer0_outputs(176) <= not(inputs(28)) or (inputs(229));
    layer0_outputs(177) <= not((inputs(84)) and (inputs(203)));
    layer0_outputs(178) <= inputs(161);
    layer0_outputs(179) <= (inputs(219)) xor (inputs(16));
    layer0_outputs(180) <= not(inputs(107)) or (inputs(227));
    layer0_outputs(181) <= (inputs(40)) xor (inputs(95));
    layer0_outputs(182) <= not((inputs(210)) or (inputs(228)));
    layer0_outputs(183) <= (inputs(134)) and (inputs(194));
    layer0_outputs(184) <= (inputs(151)) and not (inputs(95));
    layer0_outputs(185) <= not((inputs(79)) xor (inputs(159)));
    layer0_outputs(186) <= (inputs(9)) and not (inputs(218));
    layer0_outputs(187) <= (inputs(170)) and not (inputs(11));
    layer0_outputs(188) <= inputs(230);
    layer0_outputs(189) <= inputs(227);
    layer0_outputs(190) <= (inputs(216)) or (inputs(184));
    layer0_outputs(191) <= not((inputs(83)) or (inputs(69)));
    layer0_outputs(192) <= inputs(177);
    layer0_outputs(193) <= not(inputs(231));
    layer0_outputs(194) <= (inputs(204)) or (inputs(39));
    layer0_outputs(195) <= (inputs(101)) and not (inputs(196));
    layer0_outputs(196) <= not(inputs(42));
    layer0_outputs(197) <= '0';
    layer0_outputs(198) <= not((inputs(66)) or (inputs(100)));
    layer0_outputs(199) <= (inputs(66)) or (inputs(255));
    layer0_outputs(200) <= (inputs(115)) and not (inputs(186));
    layer0_outputs(201) <= (inputs(176)) and not (inputs(247));
    layer0_outputs(202) <= (inputs(234)) or (inputs(175));
    layer0_outputs(203) <= inputs(55);
    layer0_outputs(204) <= not(inputs(235));
    layer0_outputs(205) <= (inputs(128)) or (inputs(171));
    layer0_outputs(206) <= not(inputs(3)) or (inputs(153));
    layer0_outputs(207) <= '0';
    layer0_outputs(208) <= not(inputs(70)) or (inputs(94));
    layer0_outputs(209) <= not(inputs(136));
    layer0_outputs(210) <= (inputs(230)) or (inputs(47));
    layer0_outputs(211) <= not((inputs(91)) or (inputs(60)));
    layer0_outputs(212) <= (inputs(54)) or (inputs(110));
    layer0_outputs(213) <= not((inputs(222)) and (inputs(225)));
    layer0_outputs(214) <= (inputs(35)) and not (inputs(224));
    layer0_outputs(215) <= not(inputs(103)) or (inputs(114));
    layer0_outputs(216) <= (inputs(49)) or (inputs(254));
    layer0_outputs(217) <= '1';
    layer0_outputs(218) <= not((inputs(20)) xor (inputs(10)));
    layer0_outputs(219) <= (inputs(9)) xor (inputs(220));
    layer0_outputs(220) <= (inputs(64)) or (inputs(157));
    layer0_outputs(221) <= not(inputs(52)) or (inputs(63));
    layer0_outputs(222) <= '0';
    layer0_outputs(223) <= not((inputs(79)) or (inputs(116)));
    layer0_outputs(224) <= not(inputs(71));
    layer0_outputs(225) <= inputs(166);
    layer0_outputs(226) <= inputs(174);
    layer0_outputs(227) <= (inputs(10)) and not (inputs(156));
    layer0_outputs(228) <= (inputs(0)) and not (inputs(30));
    layer0_outputs(229) <= (inputs(231)) and not (inputs(134));
    layer0_outputs(230) <= '0';
    layer0_outputs(231) <= (inputs(219)) xor (inputs(191));
    layer0_outputs(232) <= not((inputs(111)) or (inputs(108)));
    layer0_outputs(233) <= not((inputs(39)) or (inputs(176)));
    layer0_outputs(234) <= not(inputs(110));
    layer0_outputs(235) <= not((inputs(26)) xor (inputs(49)));
    layer0_outputs(236) <= inputs(216);
    layer0_outputs(237) <= inputs(102);
    layer0_outputs(238) <= (inputs(248)) or (inputs(65));
    layer0_outputs(239) <= '1';
    layer0_outputs(240) <= not(inputs(193)) or (inputs(142));
    layer0_outputs(241) <= not(inputs(11));
    layer0_outputs(242) <= not(inputs(105));
    layer0_outputs(243) <= (inputs(232)) and not (inputs(8));
    layer0_outputs(244) <= '0';
    layer0_outputs(245) <= inputs(250);
    layer0_outputs(246) <= not(inputs(163)) or (inputs(203));
    layer0_outputs(247) <= not(inputs(92));
    layer0_outputs(248) <= (inputs(26)) and not (inputs(18));
    layer0_outputs(249) <= not(inputs(11));
    layer0_outputs(250) <= (inputs(9)) or (inputs(6));
    layer0_outputs(251) <= (inputs(248)) and not (inputs(17));
    layer0_outputs(252) <= (inputs(4)) and not (inputs(151));
    layer0_outputs(253) <= (inputs(204)) or (inputs(232));
    layer0_outputs(254) <= (inputs(26)) xor (inputs(48));
    layer0_outputs(255) <= inputs(86);
    layer0_outputs(256) <= (inputs(161)) and (inputs(192));
    layer0_outputs(257) <= (inputs(24)) and not (inputs(130));
    layer0_outputs(258) <= not(inputs(62));
    layer0_outputs(259) <= (inputs(107)) or (inputs(7));
    layer0_outputs(260) <= (inputs(8)) or (inputs(99));
    layer0_outputs(261) <= not((inputs(170)) or (inputs(88)));
    layer0_outputs(262) <= not(inputs(197));
    layer0_outputs(263) <= not((inputs(133)) xor (inputs(173)));
    layer0_outputs(264) <= not(inputs(218));
    layer0_outputs(265) <= (inputs(178)) and not (inputs(236));
    layer0_outputs(266) <= not(inputs(125)) or (inputs(249));
    layer0_outputs(267) <= (inputs(7)) and not (inputs(65));
    layer0_outputs(268) <= inputs(40);
    layer0_outputs(269) <= (inputs(60)) and (inputs(211));
    layer0_outputs(270) <= '0';
    layer0_outputs(271) <= inputs(189);
    layer0_outputs(272) <= inputs(234);
    layer0_outputs(273) <= (inputs(197)) and not (inputs(70));
    layer0_outputs(274) <= not((inputs(153)) or (inputs(181)));
    layer0_outputs(275) <= not(inputs(184));
    layer0_outputs(276) <= not(inputs(22));
    layer0_outputs(277) <= (inputs(81)) and not (inputs(218));
    layer0_outputs(278) <= (inputs(42)) and not (inputs(168));
    layer0_outputs(279) <= inputs(157);
    layer0_outputs(280) <= not(inputs(165));
    layer0_outputs(281) <= not((inputs(172)) or (inputs(186)));
    layer0_outputs(282) <= (inputs(160)) xor (inputs(162));
    layer0_outputs(283) <= inputs(252);
    layer0_outputs(284) <= (inputs(64)) or (inputs(254));
    layer0_outputs(285) <= not(inputs(75));
    layer0_outputs(286) <= inputs(165);
    layer0_outputs(287) <= not(inputs(7));
    layer0_outputs(288) <= not((inputs(132)) xor (inputs(50)));
    layer0_outputs(289) <= (inputs(107)) and not (inputs(152));
    layer0_outputs(290) <= not(inputs(41));
    layer0_outputs(291) <= (inputs(40)) and not (inputs(155));
    layer0_outputs(292) <= (inputs(200)) xor (inputs(232));
    layer0_outputs(293) <= not((inputs(95)) or (inputs(59)));
    layer0_outputs(294) <= (inputs(75)) and not (inputs(239));
    layer0_outputs(295) <= (inputs(57)) or (inputs(3));
    layer0_outputs(296) <= inputs(63);
    layer0_outputs(297) <= (inputs(91)) or (inputs(14));
    layer0_outputs(298) <= (inputs(9)) or (inputs(233));
    layer0_outputs(299) <= not(inputs(199));
    layer0_outputs(300) <= not((inputs(220)) xor (inputs(127)));
    layer0_outputs(301) <= not(inputs(147));
    layer0_outputs(302) <= inputs(161);
    layer0_outputs(303) <= '1';
    layer0_outputs(304) <= (inputs(157)) and not (inputs(169));
    layer0_outputs(305) <= not((inputs(128)) or (inputs(83)));
    layer0_outputs(306) <= (inputs(255)) xor (inputs(83));
    layer0_outputs(307) <= (inputs(122)) and not (inputs(219));
    layer0_outputs(308) <= not(inputs(156)) or (inputs(108));
    layer0_outputs(309) <= (inputs(90)) and not (inputs(190));
    layer0_outputs(310) <= inputs(102);
    layer0_outputs(311) <= not(inputs(245));
    layer0_outputs(312) <= not(inputs(227)) or (inputs(73));
    layer0_outputs(313) <= (inputs(156)) and not (inputs(242));
    layer0_outputs(314) <= not((inputs(172)) or (inputs(255)));
    layer0_outputs(315) <= not((inputs(30)) and (inputs(204)));
    layer0_outputs(316) <= not((inputs(125)) or (inputs(127)));
    layer0_outputs(317) <= not(inputs(37)) or (inputs(141));
    layer0_outputs(318) <= inputs(6);
    layer0_outputs(319) <= not(inputs(250)) or (inputs(38));
    layer0_outputs(320) <= not((inputs(154)) or (inputs(175)));
    layer0_outputs(321) <= not(inputs(147)) or (inputs(109));
    layer0_outputs(322) <= not((inputs(23)) xor (inputs(80)));
    layer0_outputs(323) <= (inputs(243)) and not (inputs(43));
    layer0_outputs(324) <= '0';
    layer0_outputs(325) <= not(inputs(181));
    layer0_outputs(326) <= inputs(79);
    layer0_outputs(327) <= '0';
    layer0_outputs(328) <= not(inputs(80));
    layer0_outputs(329) <= (inputs(164)) and not (inputs(32));
    layer0_outputs(330) <= not(inputs(84));
    layer0_outputs(331) <= (inputs(245)) or (inputs(49));
    layer0_outputs(332) <= not(inputs(59));
    layer0_outputs(333) <= not(inputs(103));
    layer0_outputs(334) <= not((inputs(136)) xor (inputs(184)));
    layer0_outputs(335) <= '0';
    layer0_outputs(336) <= inputs(136);
    layer0_outputs(337) <= not(inputs(230));
    layer0_outputs(338) <= '1';
    layer0_outputs(339) <= inputs(129);
    layer0_outputs(340) <= not(inputs(90)) or (inputs(14));
    layer0_outputs(341) <= (inputs(43)) or (inputs(170));
    layer0_outputs(342) <= not((inputs(28)) or (inputs(108)));
    layer0_outputs(343) <= (inputs(126)) and not (inputs(242));
    layer0_outputs(344) <= (inputs(113)) or (inputs(208));
    layer0_outputs(345) <= not((inputs(168)) or (inputs(253)));
    layer0_outputs(346) <= inputs(60);
    layer0_outputs(347) <= inputs(180);
    layer0_outputs(348) <= (inputs(254)) or (inputs(137));
    layer0_outputs(349) <= not(inputs(17)) or (inputs(216));
    layer0_outputs(350) <= not((inputs(25)) xor (inputs(103)));
    layer0_outputs(351) <= not((inputs(12)) xor (inputs(46)));
    layer0_outputs(352) <= (inputs(98)) or (inputs(8));
    layer0_outputs(353) <= (inputs(97)) or (inputs(247));
    layer0_outputs(354) <= not((inputs(254)) or (inputs(14)));
    layer0_outputs(355) <= (inputs(2)) or (inputs(44));
    layer0_outputs(356) <= not(inputs(140));
    layer0_outputs(357) <= '0';
    layer0_outputs(358) <= not((inputs(137)) and (inputs(64)));
    layer0_outputs(359) <= (inputs(82)) and (inputs(158));
    layer0_outputs(360) <= (inputs(233)) and not (inputs(1));
    layer0_outputs(361) <= not(inputs(115)) or (inputs(56));
    layer0_outputs(362) <= (inputs(192)) or (inputs(157));
    layer0_outputs(363) <= not(inputs(72)) or (inputs(107));
    layer0_outputs(364) <= (inputs(56)) xor (inputs(80));
    layer0_outputs(365) <= not(inputs(174));
    layer0_outputs(366) <= inputs(228);
    layer0_outputs(367) <= '1';
    layer0_outputs(368) <= not((inputs(172)) and (inputs(157)));
    layer0_outputs(369) <= not((inputs(5)) xor (inputs(162)));
    layer0_outputs(370) <= inputs(47);
    layer0_outputs(371) <= not(inputs(246));
    layer0_outputs(372) <= not(inputs(147));
    layer0_outputs(373) <= not(inputs(142));
    layer0_outputs(374) <= inputs(6);
    layer0_outputs(375) <= '1';
    layer0_outputs(376) <= '1';
    layer0_outputs(377) <= not(inputs(51));
    layer0_outputs(378) <= not((inputs(65)) or (inputs(119)));
    layer0_outputs(379) <= not(inputs(194)) or (inputs(63));
    layer0_outputs(380) <= not((inputs(159)) and (inputs(102)));
    layer0_outputs(381) <= not(inputs(25));
    layer0_outputs(382) <= not(inputs(167)) or (inputs(187));
    layer0_outputs(383) <= not(inputs(145));
    layer0_outputs(384) <= not(inputs(230)) or (inputs(95));
    layer0_outputs(385) <= not(inputs(119));
    layer0_outputs(386) <= not(inputs(83)) or (inputs(94));
    layer0_outputs(387) <= not(inputs(153)) or (inputs(112));
    layer0_outputs(388) <= (inputs(71)) and not (inputs(138));
    layer0_outputs(389) <= not(inputs(67));
    layer0_outputs(390) <= not(inputs(107));
    layer0_outputs(391) <= (inputs(139)) and not (inputs(235));
    layer0_outputs(392) <= inputs(88);
    layer0_outputs(393) <= not((inputs(42)) or (inputs(218)));
    layer0_outputs(394) <= inputs(8);
    layer0_outputs(395) <= (inputs(213)) and not (inputs(157));
    layer0_outputs(396) <= (inputs(247)) and (inputs(71));
    layer0_outputs(397) <= '1';
    layer0_outputs(398) <= (inputs(156)) xor (inputs(143));
    layer0_outputs(399) <= not((inputs(55)) or (inputs(237)));
    layer0_outputs(400) <= (inputs(235)) or (inputs(224));
    layer0_outputs(401) <= (inputs(213)) or (inputs(16));
    layer0_outputs(402) <= not((inputs(158)) or (inputs(231)));
    layer0_outputs(403) <= not(inputs(226)) or (inputs(141));
    layer0_outputs(404) <= not(inputs(85));
    layer0_outputs(405) <= not((inputs(102)) or (inputs(158)));
    layer0_outputs(406) <= inputs(249);
    layer0_outputs(407) <= not(inputs(99)) or (inputs(227));
    layer0_outputs(408) <= not((inputs(161)) or (inputs(175)));
    layer0_outputs(409) <= (inputs(128)) and not (inputs(46));
    layer0_outputs(410) <= (inputs(73)) xor (inputs(6));
    layer0_outputs(411) <= '0';
    layer0_outputs(412) <= (inputs(131)) and not (inputs(239));
    layer0_outputs(413) <= (inputs(244)) and not (inputs(145));
    layer0_outputs(414) <= not((inputs(40)) or (inputs(56)));
    layer0_outputs(415) <= (inputs(41)) or (inputs(10));
    layer0_outputs(416) <= not(inputs(234));
    layer0_outputs(417) <= not(inputs(98));
    layer0_outputs(418) <= (inputs(171)) and not (inputs(136));
    layer0_outputs(419) <= not(inputs(227));
    layer0_outputs(420) <= inputs(228);
    layer0_outputs(421) <= not((inputs(98)) or (inputs(132)));
    layer0_outputs(422) <= (inputs(51)) and not (inputs(75));
    layer0_outputs(423) <= inputs(75);
    layer0_outputs(424) <= (inputs(102)) or (inputs(245));
    layer0_outputs(425) <= inputs(31);
    layer0_outputs(426) <= not(inputs(83));
    layer0_outputs(427) <= not(inputs(60)) or (inputs(191));
    layer0_outputs(428) <= (inputs(64)) or (inputs(186));
    layer0_outputs(429) <= not((inputs(36)) or (inputs(243)));
    layer0_outputs(430) <= not((inputs(80)) or (inputs(195)));
    layer0_outputs(431) <= (inputs(176)) or (inputs(199));
    layer0_outputs(432) <= inputs(40);
    layer0_outputs(433) <= not(inputs(195)) or (inputs(77));
    layer0_outputs(434) <= inputs(112);
    layer0_outputs(435) <= not(inputs(177));
    layer0_outputs(436) <= not(inputs(134)) or (inputs(129));
    layer0_outputs(437) <= (inputs(21)) xor (inputs(225));
    layer0_outputs(438) <= (inputs(146)) and (inputs(102));
    layer0_outputs(439) <= not(inputs(176)) or (inputs(85));
    layer0_outputs(440) <= (inputs(171)) and not (inputs(66));
    layer0_outputs(441) <= inputs(166);
    layer0_outputs(442) <= not(inputs(243));
    layer0_outputs(443) <= not(inputs(209));
    layer0_outputs(444) <= not(inputs(120));
    layer0_outputs(445) <= (inputs(73)) and not (inputs(192));
    layer0_outputs(446) <= not(inputs(151));
    layer0_outputs(447) <= not(inputs(195));
    layer0_outputs(448) <= '1';
    layer0_outputs(449) <= inputs(81);
    layer0_outputs(450) <= not(inputs(39)) or (inputs(222));
    layer0_outputs(451) <= inputs(240);
    layer0_outputs(452) <= not((inputs(197)) xor (inputs(75)));
    layer0_outputs(453) <= (inputs(4)) and not (inputs(78));
    layer0_outputs(454) <= not((inputs(178)) or (inputs(65)));
    layer0_outputs(455) <= (inputs(89)) and not (inputs(13));
    layer0_outputs(456) <= inputs(92);
    layer0_outputs(457) <= inputs(229);
    layer0_outputs(458) <= (inputs(85)) or (inputs(160));
    layer0_outputs(459) <= (inputs(254)) and not (inputs(45));
    layer0_outputs(460) <= inputs(89);
    layer0_outputs(461) <= not(inputs(26)) or (inputs(74));
    layer0_outputs(462) <= not((inputs(85)) xor (inputs(129)));
    layer0_outputs(463) <= not(inputs(36)) or (inputs(234));
    layer0_outputs(464) <= '1';
    layer0_outputs(465) <= not(inputs(111));
    layer0_outputs(466) <= inputs(162);
    layer0_outputs(467) <= not(inputs(74)) or (inputs(32));
    layer0_outputs(468) <= not(inputs(170));
    layer0_outputs(469) <= not((inputs(229)) xor (inputs(205)));
    layer0_outputs(470) <= not(inputs(219)) or (inputs(165));
    layer0_outputs(471) <= inputs(105);
    layer0_outputs(472) <= inputs(253);
    layer0_outputs(473) <= (inputs(31)) and not (inputs(117));
    layer0_outputs(474) <= not(inputs(61)) or (inputs(241));
    layer0_outputs(475) <= (inputs(23)) or (inputs(65));
    layer0_outputs(476) <= (inputs(182)) and not (inputs(185));
    layer0_outputs(477) <= (inputs(159)) or (inputs(98));
    layer0_outputs(478) <= not((inputs(64)) or (inputs(71)));
    layer0_outputs(479) <= (inputs(42)) and not (inputs(96));
    layer0_outputs(480) <= not((inputs(232)) or (inputs(133)));
    layer0_outputs(481) <= inputs(232);
    layer0_outputs(482) <= (inputs(3)) or (inputs(200));
    layer0_outputs(483) <= not(inputs(20));
    layer0_outputs(484) <= not(inputs(185)) or (inputs(249));
    layer0_outputs(485) <= (inputs(168)) xor (inputs(216));
    layer0_outputs(486) <= (inputs(2)) and (inputs(29));
    layer0_outputs(487) <= (inputs(13)) or (inputs(43));
    layer0_outputs(488) <= not((inputs(95)) or (inputs(44)));
    layer0_outputs(489) <= not((inputs(167)) and (inputs(26)));
    layer0_outputs(490) <= (inputs(152)) and not (inputs(222));
    layer0_outputs(491) <= (inputs(38)) and not (inputs(187));
    layer0_outputs(492) <= not((inputs(216)) or (inputs(230)));
    layer0_outputs(493) <= (inputs(170)) or (inputs(197));
    layer0_outputs(494) <= not(inputs(14));
    layer0_outputs(495) <= not(inputs(152));
    layer0_outputs(496) <= inputs(4);
    layer0_outputs(497) <= not(inputs(65)) or (inputs(202));
    layer0_outputs(498) <= not((inputs(114)) or (inputs(106)));
    layer0_outputs(499) <= (inputs(27)) or (inputs(143));
    layer0_outputs(500) <= inputs(199);
    layer0_outputs(501) <= (inputs(60)) or (inputs(79));
    layer0_outputs(502) <= (inputs(107)) xor (inputs(154));
    layer0_outputs(503) <= '0';
    layer0_outputs(504) <= (inputs(47)) and not (inputs(69));
    layer0_outputs(505) <= not((inputs(177)) or (inputs(21)));
    layer0_outputs(506) <= not((inputs(70)) and (inputs(235)));
    layer0_outputs(507) <= not((inputs(206)) xor (inputs(190)));
    layer0_outputs(508) <= not((inputs(212)) or (inputs(188)));
    layer0_outputs(509) <= inputs(30);
    layer0_outputs(510) <= (inputs(254)) or (inputs(224));
    layer0_outputs(511) <= not((inputs(235)) and (inputs(174)));
    layer0_outputs(512) <= not((inputs(223)) or (inputs(23)));
    layer0_outputs(513) <= (inputs(123)) and not (inputs(132));
    layer0_outputs(514) <= not(inputs(68)) or (inputs(194));
    layer0_outputs(515) <= inputs(116);
    layer0_outputs(516) <= not(inputs(69)) or (inputs(40));
    layer0_outputs(517) <= not(inputs(121)) or (inputs(21));
    layer0_outputs(518) <= (inputs(87)) or (inputs(118));
    layer0_outputs(519) <= not(inputs(18)) or (inputs(36));
    layer0_outputs(520) <= not((inputs(45)) or (inputs(83)));
    layer0_outputs(521) <= (inputs(241)) and not (inputs(75));
    layer0_outputs(522) <= (inputs(219)) xor (inputs(122));
    layer0_outputs(523) <= (inputs(118)) xor (inputs(86));
    layer0_outputs(524) <= (inputs(234)) and not (inputs(90));
    layer0_outputs(525) <= (inputs(180)) and not (inputs(128));
    layer0_outputs(526) <= not(inputs(240)) or (inputs(185));
    layer0_outputs(527) <= '1';
    layer0_outputs(528) <= not((inputs(95)) xor (inputs(245)));
    layer0_outputs(529) <= not(inputs(179));
    layer0_outputs(530) <= (inputs(149)) and (inputs(19));
    layer0_outputs(531) <= inputs(119);
    layer0_outputs(532) <= (inputs(10)) and not (inputs(149));
    layer0_outputs(533) <= (inputs(202)) or (inputs(102));
    layer0_outputs(534) <= not(inputs(121)) or (inputs(196));
    layer0_outputs(535) <= not((inputs(33)) and (inputs(238)));
    layer0_outputs(536) <= '1';
    layer0_outputs(537) <= not(inputs(16)) or (inputs(209));
    layer0_outputs(538) <= (inputs(29)) and not (inputs(87));
    layer0_outputs(539) <= (inputs(193)) or (inputs(133));
    layer0_outputs(540) <= not((inputs(161)) or (inputs(213)));
    layer0_outputs(541) <= '1';
    layer0_outputs(542) <= not((inputs(149)) or (inputs(182)));
    layer0_outputs(543) <= '1';
    layer0_outputs(544) <= '1';
    layer0_outputs(545) <= '0';
    layer0_outputs(546) <= '0';
    layer0_outputs(547) <= not(inputs(119)) or (inputs(144));
    layer0_outputs(548) <= not(inputs(166)) or (inputs(93));
    layer0_outputs(549) <= not((inputs(234)) xor (inputs(200)));
    layer0_outputs(550) <= inputs(100);
    layer0_outputs(551) <= (inputs(166)) or (inputs(28));
    layer0_outputs(552) <= (inputs(24)) and (inputs(174));
    layer0_outputs(553) <= inputs(196);
    layer0_outputs(554) <= not((inputs(21)) or (inputs(204)));
    layer0_outputs(555) <= inputs(212);
    layer0_outputs(556) <= not(inputs(16)) or (inputs(32));
    layer0_outputs(557) <= not((inputs(173)) or (inputs(41)));
    layer0_outputs(558) <= not(inputs(255)) or (inputs(137));
    layer0_outputs(559) <= inputs(191);
    layer0_outputs(560) <= (inputs(104)) and not (inputs(147));
    layer0_outputs(561) <= (inputs(239)) and (inputs(128));
    layer0_outputs(562) <= '0';
    layer0_outputs(563) <= not((inputs(160)) and (inputs(3)));
    layer0_outputs(564) <= (inputs(193)) xor (inputs(180));
    layer0_outputs(565) <= inputs(98);
    layer0_outputs(566) <= not((inputs(189)) xor (inputs(101)));
    layer0_outputs(567) <= not((inputs(60)) or (inputs(108)));
    layer0_outputs(568) <= not(inputs(174)) or (inputs(32));
    layer0_outputs(569) <= inputs(194);
    layer0_outputs(570) <= inputs(78);
    layer0_outputs(571) <= (inputs(117)) or (inputs(168));
    layer0_outputs(572) <= (inputs(253)) xor (inputs(177));
    layer0_outputs(573) <= not((inputs(190)) or (inputs(43)));
    layer0_outputs(574) <= (inputs(193)) or (inputs(32));
    layer0_outputs(575) <= inputs(102);
    layer0_outputs(576) <= (inputs(226)) and not (inputs(36));
    layer0_outputs(577) <= inputs(203);
    layer0_outputs(578) <= not(inputs(64));
    layer0_outputs(579) <= not(inputs(44)) or (inputs(83));
    layer0_outputs(580) <= not((inputs(64)) or (inputs(111)));
    layer0_outputs(581) <= not((inputs(91)) or (inputs(113)));
    layer0_outputs(582) <= inputs(115);
    layer0_outputs(583) <= inputs(114);
    layer0_outputs(584) <= (inputs(51)) and not (inputs(114));
    layer0_outputs(585) <= inputs(5);
    layer0_outputs(586) <= not((inputs(170)) or (inputs(17)));
    layer0_outputs(587) <= (inputs(210)) and not (inputs(125));
    layer0_outputs(588) <= (inputs(104)) xor (inputs(166));
    layer0_outputs(589) <= not(inputs(98)) or (inputs(64));
    layer0_outputs(590) <= (inputs(19)) xor (inputs(11));
    layer0_outputs(591) <= not(inputs(26));
    layer0_outputs(592) <= not(inputs(129)) or (inputs(101));
    layer0_outputs(593) <= (inputs(22)) or (inputs(172));
    layer0_outputs(594) <= (inputs(73)) or (inputs(104));
    layer0_outputs(595) <= inputs(196);
    layer0_outputs(596) <= inputs(253);
    layer0_outputs(597) <= not((inputs(206)) and (inputs(37)));
    layer0_outputs(598) <= (inputs(177)) and not (inputs(46));
    layer0_outputs(599) <= not(inputs(177)) or (inputs(33));
    layer0_outputs(600) <= inputs(105);
    layer0_outputs(601) <= not((inputs(1)) or (inputs(77)));
    layer0_outputs(602) <= (inputs(126)) or (inputs(169));
    layer0_outputs(603) <= not(inputs(69)) or (inputs(0));
    layer0_outputs(604) <= (inputs(200)) and not (inputs(38));
    layer0_outputs(605) <= not(inputs(231));
    layer0_outputs(606) <= not(inputs(149));
    layer0_outputs(607) <= not((inputs(127)) or (inputs(130)));
    layer0_outputs(608) <= (inputs(95)) or (inputs(176));
    layer0_outputs(609) <= inputs(188);
    layer0_outputs(610) <= (inputs(21)) xor (inputs(141));
    layer0_outputs(611) <= inputs(176);
    layer0_outputs(612) <= '0';
    layer0_outputs(613) <= inputs(99);
    layer0_outputs(614) <= (inputs(103)) and not (inputs(110));
    layer0_outputs(615) <= not(inputs(156)) or (inputs(32));
    layer0_outputs(616) <= not((inputs(24)) xor (inputs(246)));
    layer0_outputs(617) <= not((inputs(127)) or (inputs(71)));
    layer0_outputs(618) <= not(inputs(70));
    layer0_outputs(619) <= (inputs(242)) or (inputs(111));
    layer0_outputs(620) <= not(inputs(189));
    layer0_outputs(621) <= not((inputs(80)) xor (inputs(163)));
    layer0_outputs(622) <= not((inputs(8)) or (inputs(4)));
    layer0_outputs(623) <= (inputs(180)) and not (inputs(253));
    layer0_outputs(624) <= (inputs(187)) and (inputs(57));
    layer0_outputs(625) <= inputs(88);
    layer0_outputs(626) <= (inputs(167)) and not (inputs(180));
    layer0_outputs(627) <= not(inputs(174));
    layer0_outputs(628) <= not(inputs(38)) or (inputs(23));
    layer0_outputs(629) <= (inputs(237)) and (inputs(245));
    layer0_outputs(630) <= (inputs(80)) and (inputs(76));
    layer0_outputs(631) <= inputs(36);
    layer0_outputs(632) <= (inputs(125)) xor (inputs(171));
    layer0_outputs(633) <= not((inputs(174)) or (inputs(56)));
    layer0_outputs(634) <= (inputs(66)) xor (inputs(105));
    layer0_outputs(635) <= not(inputs(58));
    layer0_outputs(636) <= not((inputs(21)) and (inputs(88)));
    layer0_outputs(637) <= (inputs(147)) and not (inputs(243));
    layer0_outputs(638) <= (inputs(90)) or (inputs(45));
    layer0_outputs(639) <= not(inputs(203)) or (inputs(7));
    layer0_outputs(640) <= (inputs(2)) and not (inputs(56));
    layer0_outputs(641) <= (inputs(111)) or (inputs(252));
    layer0_outputs(642) <= inputs(142);
    layer0_outputs(643) <= not(inputs(162)) or (inputs(185));
    layer0_outputs(644) <= (inputs(43)) and not (inputs(17));
    layer0_outputs(645) <= not((inputs(65)) or (inputs(25)));
    layer0_outputs(646) <= not(inputs(58)) or (inputs(70));
    layer0_outputs(647) <= (inputs(149)) or (inputs(196));
    layer0_outputs(648) <= inputs(20);
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= (inputs(219)) and (inputs(161));
    layer0_outputs(651) <= inputs(248);
    layer0_outputs(652) <= inputs(69);
    layer0_outputs(653) <= (inputs(129)) or (inputs(131));
    layer0_outputs(654) <= not(inputs(121)) or (inputs(242));
    layer0_outputs(655) <= inputs(130);
    layer0_outputs(656) <= not(inputs(141));
    layer0_outputs(657) <= (inputs(143)) or (inputs(248));
    layer0_outputs(658) <= not(inputs(233)) or (inputs(120));
    layer0_outputs(659) <= not((inputs(165)) or (inputs(191)));
    layer0_outputs(660) <= not((inputs(66)) xor (inputs(88)));
    layer0_outputs(661) <= (inputs(159)) xor (inputs(69));
    layer0_outputs(662) <= not((inputs(189)) and (inputs(231)));
    layer0_outputs(663) <= (inputs(246)) or (inputs(236));
    layer0_outputs(664) <= not(inputs(16)) or (inputs(3));
    layer0_outputs(665) <= not((inputs(163)) xor (inputs(79)));
    layer0_outputs(666) <= not((inputs(164)) or (inputs(190)));
    layer0_outputs(667) <= not(inputs(249)) or (inputs(79));
    layer0_outputs(668) <= not((inputs(53)) or (inputs(158)));
    layer0_outputs(669) <= not(inputs(90)) or (inputs(163));
    layer0_outputs(670) <= (inputs(199)) and not (inputs(88));
    layer0_outputs(671) <= inputs(91);
    layer0_outputs(672) <= not(inputs(227)) or (inputs(72));
    layer0_outputs(673) <= not((inputs(17)) xor (inputs(238)));
    layer0_outputs(674) <= not(inputs(16)) or (inputs(223));
    layer0_outputs(675) <= not(inputs(191)) or (inputs(172));
    layer0_outputs(676) <= not((inputs(168)) and (inputs(219)));
    layer0_outputs(677) <= inputs(211);
    layer0_outputs(678) <= inputs(11);
    layer0_outputs(679) <= not((inputs(105)) and (inputs(146)));
    layer0_outputs(680) <= not(inputs(127));
    layer0_outputs(681) <= not((inputs(48)) xor (inputs(156)));
    layer0_outputs(682) <= (inputs(58)) and not (inputs(13));
    layer0_outputs(683) <= (inputs(173)) or (inputs(172));
    layer0_outputs(684) <= not((inputs(161)) or (inputs(123)));
    layer0_outputs(685) <= not(inputs(119));
    layer0_outputs(686) <= inputs(254);
    layer0_outputs(687) <= not(inputs(234)) or (inputs(25));
    layer0_outputs(688) <= (inputs(207)) xor (inputs(36));
    layer0_outputs(689) <= inputs(97);
    layer0_outputs(690) <= inputs(136);
    layer0_outputs(691) <= not(inputs(38)) or (inputs(141));
    layer0_outputs(692) <= (inputs(160)) or (inputs(245));
    layer0_outputs(693) <= not((inputs(255)) xor (inputs(153)));
    layer0_outputs(694) <= '1';
    layer0_outputs(695) <= not((inputs(146)) or (inputs(143)));
    layer0_outputs(696) <= not(inputs(88));
    layer0_outputs(697) <= inputs(235);
    layer0_outputs(698) <= not((inputs(143)) or (inputs(50)));
    layer0_outputs(699) <= (inputs(175)) and (inputs(170));
    layer0_outputs(700) <= '1';
    layer0_outputs(701) <= not((inputs(217)) or (inputs(201)));
    layer0_outputs(702) <= inputs(3);
    layer0_outputs(703) <= (inputs(151)) and not (inputs(52));
    layer0_outputs(704) <= (inputs(215)) and not (inputs(65));
    layer0_outputs(705) <= not(inputs(4));
    layer0_outputs(706) <= not((inputs(231)) or (inputs(98)));
    layer0_outputs(707) <= (inputs(163)) and not (inputs(239));
    layer0_outputs(708) <= not(inputs(39));
    layer0_outputs(709) <= not(inputs(20));
    layer0_outputs(710) <= not((inputs(159)) or (inputs(20)));
    layer0_outputs(711) <= inputs(179);
    layer0_outputs(712) <= (inputs(38)) and not (inputs(70));
    layer0_outputs(713) <= (inputs(5)) and not (inputs(243));
    layer0_outputs(714) <= (inputs(159)) or (inputs(50));
    layer0_outputs(715) <= (inputs(169)) and (inputs(205));
    layer0_outputs(716) <= inputs(84);
    layer0_outputs(717) <= (inputs(220)) and (inputs(215));
    layer0_outputs(718) <= inputs(105);
    layer0_outputs(719) <= not(inputs(183));
    layer0_outputs(720) <= inputs(171);
    layer0_outputs(721) <= inputs(116);
    layer0_outputs(722) <= not(inputs(78));
    layer0_outputs(723) <= not(inputs(171));
    layer0_outputs(724) <= inputs(78);
    layer0_outputs(725) <= (inputs(232)) or (inputs(32));
    layer0_outputs(726) <= not(inputs(153));
    layer0_outputs(727) <= '0';
    layer0_outputs(728) <= '1';
    layer0_outputs(729) <= not((inputs(244)) and (inputs(211)));
    layer0_outputs(730) <= inputs(127);
    layer0_outputs(731) <= not(inputs(41)) or (inputs(119));
    layer0_outputs(732) <= inputs(168);
    layer0_outputs(733) <= not((inputs(247)) or (inputs(18)));
    layer0_outputs(734) <= inputs(66);
    layer0_outputs(735) <= not(inputs(123));
    layer0_outputs(736) <= not(inputs(227)) or (inputs(239));
    layer0_outputs(737) <= inputs(232);
    layer0_outputs(738) <= not((inputs(30)) or (inputs(188)));
    layer0_outputs(739) <= inputs(97);
    layer0_outputs(740) <= (inputs(124)) and (inputs(246));
    layer0_outputs(741) <= not((inputs(172)) or (inputs(79)));
    layer0_outputs(742) <= '0';
    layer0_outputs(743) <= (inputs(133)) and (inputs(17));
    layer0_outputs(744) <= (inputs(171)) and not (inputs(135));
    layer0_outputs(745) <= not(inputs(111));
    layer0_outputs(746) <= not(inputs(236));
    layer0_outputs(747) <= not((inputs(112)) or (inputs(211)));
    layer0_outputs(748) <= '1';
    layer0_outputs(749) <= '0';
    layer0_outputs(750) <= not((inputs(20)) or (inputs(47)));
    layer0_outputs(751) <= (inputs(150)) and not (inputs(92));
    layer0_outputs(752) <= not((inputs(73)) and (inputs(52)));
    layer0_outputs(753) <= not((inputs(137)) xor (inputs(251)));
    layer0_outputs(754) <= not(inputs(249)) or (inputs(49));
    layer0_outputs(755) <= inputs(24);
    layer0_outputs(756) <= not(inputs(68)) or (inputs(175));
    layer0_outputs(757) <= (inputs(38)) or (inputs(27));
    layer0_outputs(758) <= (inputs(53)) and not (inputs(182));
    layer0_outputs(759) <= not((inputs(126)) xor (inputs(155)));
    layer0_outputs(760) <= (inputs(173)) or (inputs(46));
    layer0_outputs(761) <= (inputs(210)) and not (inputs(189));
    layer0_outputs(762) <= not(inputs(162)) or (inputs(56));
    layer0_outputs(763) <= (inputs(33)) or (inputs(109));
    layer0_outputs(764) <= (inputs(220)) xor (inputs(141));
    layer0_outputs(765) <= not((inputs(76)) xor (inputs(253)));
    layer0_outputs(766) <= not((inputs(235)) or (inputs(158)));
    layer0_outputs(767) <= (inputs(221)) or (inputs(192));
    layer0_outputs(768) <= (inputs(204)) and (inputs(195));
    layer0_outputs(769) <= (inputs(156)) and not (inputs(40));
    layer0_outputs(770) <= not(inputs(92));
    layer0_outputs(771) <= not(inputs(212)) or (inputs(48));
    layer0_outputs(772) <= not(inputs(244)) or (inputs(181));
    layer0_outputs(773) <= not(inputs(96));
    layer0_outputs(774) <= not(inputs(53)) or (inputs(87));
    layer0_outputs(775) <= (inputs(218)) and not (inputs(36));
    layer0_outputs(776) <= not((inputs(229)) xor (inputs(159)));
    layer0_outputs(777) <= (inputs(138)) or (inputs(110));
    layer0_outputs(778) <= '0';
    layer0_outputs(779) <= inputs(125);
    layer0_outputs(780) <= not((inputs(113)) xor (inputs(117)));
    layer0_outputs(781) <= not(inputs(91));
    layer0_outputs(782) <= not(inputs(166));
    layer0_outputs(783) <= inputs(131);
    layer0_outputs(784) <= not(inputs(87));
    layer0_outputs(785) <= (inputs(246)) or (inputs(226));
    layer0_outputs(786) <= not(inputs(157)) or (inputs(35));
    layer0_outputs(787) <= not((inputs(168)) xor (inputs(69)));
    layer0_outputs(788) <= (inputs(95)) or (inputs(123));
    layer0_outputs(789) <= (inputs(230)) and not (inputs(120));
    layer0_outputs(790) <= not((inputs(220)) or (inputs(136)));
    layer0_outputs(791) <= not((inputs(151)) or (inputs(148)));
    layer0_outputs(792) <= not(inputs(49)) or (inputs(5));
    layer0_outputs(793) <= not((inputs(235)) or (inputs(86)));
    layer0_outputs(794) <= (inputs(37)) and not (inputs(8));
    layer0_outputs(795) <= '1';
    layer0_outputs(796) <= (inputs(178)) or (inputs(173));
    layer0_outputs(797) <= (inputs(40)) and not (inputs(144));
    layer0_outputs(798) <= '0';
    layer0_outputs(799) <= inputs(70);
    layer0_outputs(800) <= not((inputs(20)) xor (inputs(100)));
    layer0_outputs(801) <= not(inputs(135)) or (inputs(18));
    layer0_outputs(802) <= '1';
    layer0_outputs(803) <= (inputs(12)) or (inputs(208));
    layer0_outputs(804) <= '0';
    layer0_outputs(805) <= not((inputs(135)) or (inputs(192)));
    layer0_outputs(806) <= '0';
    layer0_outputs(807) <= inputs(251);
    layer0_outputs(808) <= not(inputs(180));
    layer0_outputs(809) <= not(inputs(223)) or (inputs(175));
    layer0_outputs(810) <= (inputs(115)) and not (inputs(119));
    layer0_outputs(811) <= inputs(121);
    layer0_outputs(812) <= not((inputs(73)) or (inputs(196)));
    layer0_outputs(813) <= not((inputs(123)) or (inputs(189)));
    layer0_outputs(814) <= inputs(158);
    layer0_outputs(815) <= not(inputs(128));
    layer0_outputs(816) <= not((inputs(233)) or (inputs(211)));
    layer0_outputs(817) <= inputs(49);
    layer0_outputs(818) <= not(inputs(52)) or (inputs(185));
    layer0_outputs(819) <= not(inputs(17));
    layer0_outputs(820) <= not(inputs(118)) or (inputs(18));
    layer0_outputs(821) <= not(inputs(120)) or (inputs(55));
    layer0_outputs(822) <= not((inputs(87)) or (inputs(99)));
    layer0_outputs(823) <= (inputs(144)) or (inputs(158));
    layer0_outputs(824) <= (inputs(182)) and not (inputs(63));
    layer0_outputs(825) <= '1';
    layer0_outputs(826) <= not(inputs(44));
    layer0_outputs(827) <= inputs(120);
    layer0_outputs(828) <= '1';
    layer0_outputs(829) <= not(inputs(109));
    layer0_outputs(830) <= not((inputs(86)) or (inputs(251)));
    layer0_outputs(831) <= not(inputs(248));
    layer0_outputs(832) <= (inputs(85)) or (inputs(178));
    layer0_outputs(833) <= (inputs(213)) and not (inputs(37));
    layer0_outputs(834) <= (inputs(209)) xor (inputs(219));
    layer0_outputs(835) <= (inputs(204)) and not (inputs(233));
    layer0_outputs(836) <= not(inputs(162));
    layer0_outputs(837) <= (inputs(2)) or (inputs(158));
    layer0_outputs(838) <= not(inputs(172));
    layer0_outputs(839) <= (inputs(251)) or (inputs(23));
    layer0_outputs(840) <= inputs(147);
    layer0_outputs(841) <= not(inputs(120));
    layer0_outputs(842) <= not((inputs(174)) xor (inputs(53)));
    layer0_outputs(843) <= not(inputs(169)) or (inputs(117));
    layer0_outputs(844) <= not(inputs(231));
    layer0_outputs(845) <= (inputs(233)) xor (inputs(229));
    layer0_outputs(846) <= not((inputs(58)) or (inputs(206)));
    layer0_outputs(847) <= not(inputs(172)) or (inputs(246));
    layer0_outputs(848) <= not(inputs(58)) or (inputs(251));
    layer0_outputs(849) <= (inputs(209)) or (inputs(224));
    layer0_outputs(850) <= not(inputs(2));
    layer0_outputs(851) <= not(inputs(21));
    layer0_outputs(852) <= not(inputs(39)) or (inputs(211));
    layer0_outputs(853) <= '1';
    layer0_outputs(854) <= (inputs(34)) or (inputs(136));
    layer0_outputs(855) <= not((inputs(122)) xor (inputs(220)));
    layer0_outputs(856) <= '0';
    layer0_outputs(857) <= (inputs(107)) or (inputs(175));
    layer0_outputs(858) <= not(inputs(120));
    layer0_outputs(859) <= (inputs(248)) and not (inputs(93));
    layer0_outputs(860) <= not((inputs(178)) or (inputs(32)));
    layer0_outputs(861) <= not((inputs(196)) or (inputs(211)));
    layer0_outputs(862) <= not((inputs(139)) and (inputs(245)));
    layer0_outputs(863) <= not(inputs(70));
    layer0_outputs(864) <= not(inputs(183));
    layer0_outputs(865) <= inputs(135);
    layer0_outputs(866) <= inputs(42);
    layer0_outputs(867) <= not(inputs(218));
    layer0_outputs(868) <= (inputs(8)) and not (inputs(222));
    layer0_outputs(869) <= (inputs(9)) and not (inputs(16));
    layer0_outputs(870) <= not((inputs(188)) or (inputs(180)));
    layer0_outputs(871) <= not(inputs(11)) or (inputs(72));
    layer0_outputs(872) <= not((inputs(15)) and (inputs(110)));
    layer0_outputs(873) <= not(inputs(248)) or (inputs(214));
    layer0_outputs(874) <= (inputs(212)) and not (inputs(98));
    layer0_outputs(875) <= inputs(160);
    layer0_outputs(876) <= not((inputs(219)) or (inputs(245)));
    layer0_outputs(877) <= not((inputs(238)) xor (inputs(230)));
    layer0_outputs(878) <= not(inputs(211));
    layer0_outputs(879) <= '0';
    layer0_outputs(880) <= (inputs(47)) and (inputs(207));
    layer0_outputs(881) <= (inputs(114)) and (inputs(182));
    layer0_outputs(882) <= (inputs(44)) and not (inputs(71));
    layer0_outputs(883) <= (inputs(48)) xor (inputs(10));
    layer0_outputs(884) <= (inputs(93)) and not (inputs(192));
    layer0_outputs(885) <= not(inputs(26)) or (inputs(164));
    layer0_outputs(886) <= inputs(232);
    layer0_outputs(887) <= (inputs(155)) or (inputs(246));
    layer0_outputs(888) <= not(inputs(86)) or (inputs(157));
    layer0_outputs(889) <= (inputs(200)) and (inputs(159));
    layer0_outputs(890) <= not((inputs(177)) or (inputs(199)));
    layer0_outputs(891) <= not((inputs(223)) or (inputs(168)));
    layer0_outputs(892) <= '0';
    layer0_outputs(893) <= (inputs(170)) xor (inputs(181));
    layer0_outputs(894) <= not((inputs(84)) or (inputs(239)));
    layer0_outputs(895) <= not(inputs(28)) or (inputs(163));
    layer0_outputs(896) <= not(inputs(206));
    layer0_outputs(897) <= not(inputs(93)) or (inputs(12));
    layer0_outputs(898) <= '1';
    layer0_outputs(899) <= (inputs(252)) or (inputs(137));
    layer0_outputs(900) <= (inputs(8)) or (inputs(190));
    layer0_outputs(901) <= not(inputs(133));
    layer0_outputs(902) <= not(inputs(104));
    layer0_outputs(903) <= (inputs(102)) and not (inputs(155));
    layer0_outputs(904) <= (inputs(155)) xor (inputs(2));
    layer0_outputs(905) <= inputs(144);
    layer0_outputs(906) <= (inputs(207)) xor (inputs(23));
    layer0_outputs(907) <= not((inputs(233)) and (inputs(190)));
    layer0_outputs(908) <= not(inputs(88));
    layer0_outputs(909) <= (inputs(172)) or (inputs(47));
    layer0_outputs(910) <= not(inputs(250));
    layer0_outputs(911) <= (inputs(165)) or (inputs(108));
    layer0_outputs(912) <= '1';
    layer0_outputs(913) <= inputs(113);
    layer0_outputs(914) <= not(inputs(35));
    layer0_outputs(915) <= (inputs(195)) and not (inputs(113));
    layer0_outputs(916) <= not((inputs(81)) xor (inputs(14)));
    layer0_outputs(917) <= not(inputs(156));
    layer0_outputs(918) <= not((inputs(162)) or (inputs(175)));
    layer0_outputs(919) <= (inputs(128)) or (inputs(214));
    layer0_outputs(920) <= not(inputs(55));
    layer0_outputs(921) <= not(inputs(211)) or (inputs(0));
    layer0_outputs(922) <= inputs(212);
    layer0_outputs(923) <= not(inputs(73));
    layer0_outputs(924) <= not((inputs(67)) or (inputs(170)));
    layer0_outputs(925) <= not((inputs(34)) xor (inputs(115)));
    layer0_outputs(926) <= not(inputs(211)) or (inputs(109));
    layer0_outputs(927) <= '0';
    layer0_outputs(928) <= inputs(229);
    layer0_outputs(929) <= inputs(88);
    layer0_outputs(930) <= not(inputs(240)) or (inputs(55));
    layer0_outputs(931) <= not((inputs(53)) and (inputs(96)));
    layer0_outputs(932) <= not(inputs(125));
    layer0_outputs(933) <= not((inputs(116)) xor (inputs(57)));
    layer0_outputs(934) <= (inputs(178)) and not (inputs(214));
    layer0_outputs(935) <= not(inputs(71));
    layer0_outputs(936) <= not((inputs(212)) or (inputs(137)));
    layer0_outputs(937) <= not((inputs(13)) xor (inputs(199)));
    layer0_outputs(938) <= (inputs(136)) or (inputs(178));
    layer0_outputs(939) <= inputs(162);
    layer0_outputs(940) <= not(inputs(8)) or (inputs(212));
    layer0_outputs(941) <= not((inputs(53)) or (inputs(76)));
    layer0_outputs(942) <= not(inputs(170));
    layer0_outputs(943) <= (inputs(169)) and not (inputs(95));
    layer0_outputs(944) <= (inputs(121)) and not (inputs(19));
    layer0_outputs(945) <= inputs(33);
    layer0_outputs(946) <= not((inputs(192)) xor (inputs(152)));
    layer0_outputs(947) <= inputs(60);
    layer0_outputs(948) <= (inputs(52)) and not (inputs(0));
    layer0_outputs(949) <= (inputs(229)) xor (inputs(238));
    layer0_outputs(950) <= '0';
    layer0_outputs(951) <= inputs(215);
    layer0_outputs(952) <= (inputs(180)) and (inputs(124));
    layer0_outputs(953) <= not((inputs(221)) or (inputs(54)));
    layer0_outputs(954) <= not((inputs(248)) xor (inputs(176)));
    layer0_outputs(955) <= not((inputs(174)) or (inputs(218)));
    layer0_outputs(956) <= (inputs(216)) or (inputs(201));
    layer0_outputs(957) <= inputs(84);
    layer0_outputs(958) <= (inputs(57)) and (inputs(155));
    layer0_outputs(959) <= not(inputs(88));
    layer0_outputs(960) <= not((inputs(68)) or (inputs(134)));
    layer0_outputs(961) <= not((inputs(80)) xor (inputs(1)));
    layer0_outputs(962) <= (inputs(56)) or (inputs(20));
    layer0_outputs(963) <= '0';
    layer0_outputs(964) <= inputs(229);
    layer0_outputs(965) <= '0';
    layer0_outputs(966) <= not(inputs(194));
    layer0_outputs(967) <= not((inputs(61)) or (inputs(164)));
    layer0_outputs(968) <= not(inputs(96)) or (inputs(141));
    layer0_outputs(969) <= not((inputs(250)) or (inputs(118)));
    layer0_outputs(970) <= not((inputs(87)) or (inputs(84)));
    layer0_outputs(971) <= inputs(41);
    layer0_outputs(972) <= (inputs(238)) or (inputs(184));
    layer0_outputs(973) <= not(inputs(140));
    layer0_outputs(974) <= (inputs(228)) and not (inputs(64));
    layer0_outputs(975) <= inputs(144);
    layer0_outputs(976) <= inputs(152);
    layer0_outputs(977) <= not(inputs(107));
    layer0_outputs(978) <= (inputs(110)) and not (inputs(241));
    layer0_outputs(979) <= (inputs(16)) xor (inputs(55));
    layer0_outputs(980) <= inputs(7);
    layer0_outputs(981) <= (inputs(89)) and not (inputs(94));
    layer0_outputs(982) <= not(inputs(218)) or (inputs(103));
    layer0_outputs(983) <= (inputs(68)) xor (inputs(148));
    layer0_outputs(984) <= not(inputs(77));
    layer0_outputs(985) <= not(inputs(129));
    layer0_outputs(986) <= (inputs(67)) and not (inputs(127));
    layer0_outputs(987) <= not(inputs(249));
    layer0_outputs(988) <= inputs(122);
    layer0_outputs(989) <= not(inputs(5));
    layer0_outputs(990) <= not(inputs(188)) or (inputs(16));
    layer0_outputs(991) <= (inputs(163)) and not (inputs(47));
    layer0_outputs(992) <= (inputs(7)) and not (inputs(66));
    layer0_outputs(993) <= inputs(77);
    layer0_outputs(994) <= (inputs(15)) or (inputs(166));
    layer0_outputs(995) <= (inputs(205)) xor (inputs(165));
    layer0_outputs(996) <= not((inputs(196)) and (inputs(230)));
    layer0_outputs(997) <= not((inputs(169)) or (inputs(25)));
    layer0_outputs(998) <= (inputs(166)) and not (inputs(33));
    layer0_outputs(999) <= inputs(227);
    layer0_outputs(1000) <= (inputs(52)) or (inputs(122));
    layer0_outputs(1001) <= inputs(173);
    layer0_outputs(1002) <= not((inputs(194)) xor (inputs(203)));
    layer0_outputs(1003) <= not(inputs(233));
    layer0_outputs(1004) <= not(inputs(103));
    layer0_outputs(1005) <= inputs(209);
    layer0_outputs(1006) <= inputs(170);
    layer0_outputs(1007) <= (inputs(121)) or (inputs(251));
    layer0_outputs(1008) <= '1';
    layer0_outputs(1009) <= (inputs(54)) or (inputs(116));
    layer0_outputs(1010) <= inputs(131);
    layer0_outputs(1011) <= not(inputs(220));
    layer0_outputs(1012) <= (inputs(172)) xor (inputs(192));
    layer0_outputs(1013) <= (inputs(40)) or (inputs(63));
    layer0_outputs(1014) <= not((inputs(166)) and (inputs(197)));
    layer0_outputs(1015) <= not((inputs(151)) or (inputs(35)));
    layer0_outputs(1016) <= (inputs(242)) or (inputs(217));
    layer0_outputs(1017) <= not(inputs(177)) or (inputs(239));
    layer0_outputs(1018) <= '1';
    layer0_outputs(1019) <= (inputs(196)) or (inputs(204));
    layer0_outputs(1020) <= not(inputs(26));
    layer0_outputs(1021) <= inputs(184);
    layer0_outputs(1022) <= inputs(160);
    layer0_outputs(1023) <= (inputs(169)) or (inputs(29));
    layer0_outputs(1024) <= '0';
    layer0_outputs(1025) <= not(inputs(101));
    layer0_outputs(1026) <= not((inputs(176)) and (inputs(6)));
    layer0_outputs(1027) <= inputs(230);
    layer0_outputs(1028) <= not(inputs(153));
    layer0_outputs(1029) <= inputs(34);
    layer0_outputs(1030) <= not((inputs(69)) or (inputs(186)));
    layer0_outputs(1031) <= (inputs(60)) xor (inputs(208));
    layer0_outputs(1032) <= inputs(208);
    layer0_outputs(1033) <= (inputs(84)) and not (inputs(95));
    layer0_outputs(1034) <= not((inputs(121)) and (inputs(144)));
    layer0_outputs(1035) <= not(inputs(102)) or (inputs(99));
    layer0_outputs(1036) <= inputs(174);
    layer0_outputs(1037) <= (inputs(134)) or (inputs(19));
    layer0_outputs(1038) <= (inputs(130)) or (inputs(71));
    layer0_outputs(1039) <= (inputs(116)) xor (inputs(161));
    layer0_outputs(1040) <= (inputs(9)) and not (inputs(253));
    layer0_outputs(1041) <= (inputs(207)) xor (inputs(253));
    layer0_outputs(1042) <= '1';
    layer0_outputs(1043) <= (inputs(167)) or (inputs(187));
    layer0_outputs(1044) <= not(inputs(56));
    layer0_outputs(1045) <= not(inputs(84));
    layer0_outputs(1046) <= not(inputs(192)) or (inputs(15));
    layer0_outputs(1047) <= inputs(143);
    layer0_outputs(1048) <= inputs(89);
    layer0_outputs(1049) <= not((inputs(137)) or (inputs(105)));
    layer0_outputs(1050) <= not((inputs(79)) or (inputs(92)));
    layer0_outputs(1051) <= not((inputs(172)) or (inputs(250)));
    layer0_outputs(1052) <= not((inputs(196)) or (inputs(174)));
    layer0_outputs(1053) <= (inputs(93)) and not (inputs(3));
    layer0_outputs(1054) <= not(inputs(107)) or (inputs(215));
    layer0_outputs(1055) <= inputs(226);
    layer0_outputs(1056) <= not(inputs(199));
    layer0_outputs(1057) <= (inputs(134)) or (inputs(65));
    layer0_outputs(1058) <= (inputs(74)) or (inputs(65));
    layer0_outputs(1059) <= not(inputs(198));
    layer0_outputs(1060) <= (inputs(53)) or (inputs(124));
    layer0_outputs(1061) <= inputs(82);
    layer0_outputs(1062) <= (inputs(123)) and not (inputs(149));
    layer0_outputs(1063) <= (inputs(235)) and (inputs(165));
    layer0_outputs(1064) <= inputs(169);
    layer0_outputs(1065) <= (inputs(78)) xor (inputs(44));
    layer0_outputs(1066) <= '0';
    layer0_outputs(1067) <= inputs(132);
    layer0_outputs(1068) <= not(inputs(121));
    layer0_outputs(1069) <= (inputs(153)) or (inputs(161));
    layer0_outputs(1070) <= '0';
    layer0_outputs(1071) <= (inputs(237)) and not (inputs(206));
    layer0_outputs(1072) <= inputs(134);
    layer0_outputs(1073) <= inputs(59);
    layer0_outputs(1074) <= not(inputs(244)) or (inputs(58));
    layer0_outputs(1075) <= '0';
    layer0_outputs(1076) <= (inputs(104)) xor (inputs(134));
    layer0_outputs(1077) <= not(inputs(187));
    layer0_outputs(1078) <= (inputs(24)) or (inputs(7));
    layer0_outputs(1079) <= not((inputs(62)) or (inputs(16)));
    layer0_outputs(1080) <= not(inputs(236));
    layer0_outputs(1081) <= '0';
    layer0_outputs(1082) <= not((inputs(127)) or (inputs(251)));
    layer0_outputs(1083) <= (inputs(102)) or (inputs(94));
    layer0_outputs(1084) <= not((inputs(25)) or (inputs(34)));
    layer0_outputs(1085) <= (inputs(17)) and not (inputs(186));
    layer0_outputs(1086) <= not(inputs(101));
    layer0_outputs(1087) <= not((inputs(114)) or (inputs(132)));
    layer0_outputs(1088) <= '1';
    layer0_outputs(1089) <= (inputs(50)) or (inputs(101));
    layer0_outputs(1090) <= not(inputs(161));
    layer0_outputs(1091) <= (inputs(43)) xor (inputs(58));
    layer0_outputs(1092) <= (inputs(189)) and not (inputs(21));
    layer0_outputs(1093) <= not((inputs(48)) and (inputs(87)));
    layer0_outputs(1094) <= inputs(130);
    layer0_outputs(1095) <= not((inputs(80)) xor (inputs(228)));
    layer0_outputs(1096) <= (inputs(40)) and (inputs(40));
    layer0_outputs(1097) <= (inputs(205)) and not (inputs(111));
    layer0_outputs(1098) <= (inputs(5)) and not (inputs(86));
    layer0_outputs(1099) <= (inputs(85)) and not (inputs(41));
    layer0_outputs(1100) <= (inputs(38)) xor (inputs(61));
    layer0_outputs(1101) <= (inputs(230)) and not (inputs(175));
    layer0_outputs(1102) <= not(inputs(122));
    layer0_outputs(1103) <= not(inputs(185));
    layer0_outputs(1104) <= inputs(58);
    layer0_outputs(1105) <= not((inputs(92)) xor (inputs(74)));
    layer0_outputs(1106) <= not(inputs(168)) or (inputs(102));
    layer0_outputs(1107) <= not((inputs(171)) or (inputs(197)));
    layer0_outputs(1108) <= (inputs(140)) and not (inputs(81));
    layer0_outputs(1109) <= (inputs(72)) and not (inputs(191));
    layer0_outputs(1110) <= not(inputs(66));
    layer0_outputs(1111) <= not((inputs(152)) and (inputs(9)));
    layer0_outputs(1112) <= not(inputs(120)) or (inputs(178));
    layer0_outputs(1113) <= (inputs(101)) or (inputs(84));
    layer0_outputs(1114) <= not((inputs(133)) xor (inputs(151)));
    layer0_outputs(1115) <= not((inputs(64)) or (inputs(50)));
    layer0_outputs(1116) <= (inputs(111)) or (inputs(61));
    layer0_outputs(1117) <= inputs(53);
    layer0_outputs(1118) <= not(inputs(153)) or (inputs(194));
    layer0_outputs(1119) <= not(inputs(83)) or (inputs(51));
    layer0_outputs(1120) <= not(inputs(232));
    layer0_outputs(1121) <= (inputs(204)) and not (inputs(216));
    layer0_outputs(1122) <= (inputs(27)) and (inputs(229));
    layer0_outputs(1123) <= (inputs(84)) and not (inputs(3));
    layer0_outputs(1124) <= not(inputs(23));
    layer0_outputs(1125) <= (inputs(31)) or (inputs(250));
    layer0_outputs(1126) <= not(inputs(149)) or (inputs(82));
    layer0_outputs(1127) <= (inputs(240)) or (inputs(182));
    layer0_outputs(1128) <= (inputs(124)) or (inputs(111));
    layer0_outputs(1129) <= (inputs(81)) xor (inputs(131));
    layer0_outputs(1130) <= not(inputs(94));
    layer0_outputs(1131) <= not((inputs(81)) or (inputs(15)));
    layer0_outputs(1132) <= inputs(183);
    layer0_outputs(1133) <= not(inputs(122));
    layer0_outputs(1134) <= not(inputs(145));
    layer0_outputs(1135) <= not(inputs(67)) or (inputs(55));
    layer0_outputs(1136) <= not(inputs(157));
    layer0_outputs(1137) <= not((inputs(193)) or (inputs(171)));
    layer0_outputs(1138) <= not(inputs(117));
    layer0_outputs(1139) <= (inputs(20)) or (inputs(32));
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= inputs(136);
    layer0_outputs(1142) <= not((inputs(187)) or (inputs(164)));
    layer0_outputs(1143) <= inputs(247);
    layer0_outputs(1144) <= not(inputs(207));
    layer0_outputs(1145) <= (inputs(139)) and not (inputs(240));
    layer0_outputs(1146) <= not((inputs(23)) and (inputs(224)));
    layer0_outputs(1147) <= (inputs(252)) or (inputs(29));
    layer0_outputs(1148) <= (inputs(204)) and (inputs(152));
    layer0_outputs(1149) <= not(inputs(252)) or (inputs(63));
    layer0_outputs(1150) <= inputs(239);
    layer0_outputs(1151) <= (inputs(254)) and not (inputs(169));
    layer0_outputs(1152) <= not(inputs(168));
    layer0_outputs(1153) <= not((inputs(15)) or (inputs(19)));
    layer0_outputs(1154) <= (inputs(113)) and not (inputs(54));
    layer0_outputs(1155) <= '0';
    layer0_outputs(1156) <= (inputs(229)) and (inputs(225));
    layer0_outputs(1157) <= (inputs(122)) or (inputs(251));
    layer0_outputs(1158) <= not((inputs(23)) or (inputs(62)));
    layer0_outputs(1159) <= inputs(182);
    layer0_outputs(1160) <= (inputs(9)) or (inputs(191));
    layer0_outputs(1161) <= inputs(218);
    layer0_outputs(1162) <= not(inputs(50));
    layer0_outputs(1163) <= not((inputs(168)) or (inputs(110)));
    layer0_outputs(1164) <= not(inputs(120));
    layer0_outputs(1165) <= not(inputs(78));
    layer0_outputs(1166) <= (inputs(100)) or (inputs(43));
    layer0_outputs(1167) <= not((inputs(99)) or (inputs(147)));
    layer0_outputs(1168) <= not(inputs(198));
    layer0_outputs(1169) <= inputs(30);
    layer0_outputs(1170) <= not(inputs(231)) or (inputs(238));
    layer0_outputs(1171) <= not(inputs(89));
    layer0_outputs(1172) <= (inputs(144)) xor (inputs(254));
    layer0_outputs(1173) <= not(inputs(229)) or (inputs(166));
    layer0_outputs(1174) <= (inputs(179)) or (inputs(50));
    layer0_outputs(1175) <= (inputs(216)) and (inputs(72));
    layer0_outputs(1176) <= not((inputs(141)) and (inputs(54)));
    layer0_outputs(1177) <= not((inputs(65)) or (inputs(206)));
    layer0_outputs(1178) <= not(inputs(102));
    layer0_outputs(1179) <= inputs(203);
    layer0_outputs(1180) <= inputs(46);
    layer0_outputs(1181) <= not(inputs(129)) or (inputs(166));
    layer0_outputs(1182) <= not((inputs(199)) or (inputs(156)));
    layer0_outputs(1183) <= not(inputs(168));
    layer0_outputs(1184) <= not((inputs(112)) xor (inputs(86)));
    layer0_outputs(1185) <= not(inputs(143)) or (inputs(96));
    layer0_outputs(1186) <= inputs(51);
    layer0_outputs(1187) <= inputs(76);
    layer0_outputs(1188) <= (inputs(203)) or (inputs(126));
    layer0_outputs(1189) <= not((inputs(40)) or (inputs(88)));
    layer0_outputs(1190) <= inputs(145);
    layer0_outputs(1191) <= not((inputs(252)) or (inputs(208)));
    layer0_outputs(1192) <= '0';
    layer0_outputs(1193) <= (inputs(71)) xor (inputs(134));
    layer0_outputs(1194) <= not((inputs(144)) xor (inputs(112)));
    layer0_outputs(1195) <= not(inputs(48));
    layer0_outputs(1196) <= not(inputs(206));
    layer0_outputs(1197) <= (inputs(15)) and not (inputs(92));
    layer0_outputs(1198) <= inputs(89);
    layer0_outputs(1199) <= (inputs(85)) and not (inputs(215));
    layer0_outputs(1200) <= (inputs(216)) or (inputs(149));
    layer0_outputs(1201) <= (inputs(153)) and not (inputs(60));
    layer0_outputs(1202) <= not(inputs(78));
    layer0_outputs(1203) <= (inputs(217)) and not (inputs(219));
    layer0_outputs(1204) <= not(inputs(99)) or (inputs(242));
    layer0_outputs(1205) <= not((inputs(214)) or (inputs(251)));
    layer0_outputs(1206) <= not(inputs(179)) or (inputs(162));
    layer0_outputs(1207) <= (inputs(46)) or (inputs(31));
    layer0_outputs(1208) <= not(inputs(91)) or (inputs(12));
    layer0_outputs(1209) <= (inputs(157)) and not (inputs(32));
    layer0_outputs(1210) <= not(inputs(232));
    layer0_outputs(1211) <= inputs(92);
    layer0_outputs(1212) <= (inputs(84)) and not (inputs(165));
    layer0_outputs(1213) <= (inputs(127)) xor (inputs(110));
    layer0_outputs(1214) <= not((inputs(158)) and (inputs(68)));
    layer0_outputs(1215) <= not(inputs(243));
    layer0_outputs(1216) <= (inputs(128)) and not (inputs(253));
    layer0_outputs(1217) <= (inputs(110)) and not (inputs(54));
    layer0_outputs(1218) <= not(inputs(231));
    layer0_outputs(1219) <= inputs(200);
    layer0_outputs(1220) <= not(inputs(238));
    layer0_outputs(1221) <= (inputs(163)) and not (inputs(90));
    layer0_outputs(1222) <= not(inputs(73));
    layer0_outputs(1223) <= not((inputs(29)) xor (inputs(128)));
    layer0_outputs(1224) <= (inputs(156)) and not (inputs(230));
    layer0_outputs(1225) <= inputs(183);
    layer0_outputs(1226) <= not((inputs(247)) and (inputs(102)));
    layer0_outputs(1227) <= not(inputs(26));
    layer0_outputs(1228) <= not(inputs(15)) or (inputs(33));
    layer0_outputs(1229) <= not((inputs(78)) xor (inputs(16)));
    layer0_outputs(1230) <= not(inputs(153)) or (inputs(187));
    layer0_outputs(1231) <= inputs(69);
    layer0_outputs(1232) <= (inputs(165)) and not (inputs(152));
    layer0_outputs(1233) <= not((inputs(62)) and (inputs(119)));
    layer0_outputs(1234) <= (inputs(36)) and not (inputs(16));
    layer0_outputs(1235) <= (inputs(90)) xor (inputs(180));
    layer0_outputs(1236) <= not(inputs(143));
    layer0_outputs(1237) <= not((inputs(3)) or (inputs(186)));
    layer0_outputs(1238) <= (inputs(32)) or (inputs(135));
    layer0_outputs(1239) <= (inputs(197)) xor (inputs(1));
    layer0_outputs(1240) <= not(inputs(245));
    layer0_outputs(1241) <= inputs(42);
    layer0_outputs(1242) <= not((inputs(219)) or (inputs(149)));
    layer0_outputs(1243) <= not(inputs(106));
    layer0_outputs(1244) <= '1';
    layer0_outputs(1245) <= not((inputs(143)) xor (inputs(133)));
    layer0_outputs(1246) <= inputs(129);
    layer0_outputs(1247) <= (inputs(35)) and not (inputs(53));
    layer0_outputs(1248) <= (inputs(70)) xor (inputs(68));
    layer0_outputs(1249) <= not(inputs(220));
    layer0_outputs(1250) <= inputs(253);
    layer0_outputs(1251) <= not((inputs(238)) xor (inputs(253)));
    layer0_outputs(1252) <= inputs(32);
    layer0_outputs(1253) <= not(inputs(246)) or (inputs(207));
    layer0_outputs(1254) <= inputs(250);
    layer0_outputs(1255) <= not(inputs(62)) or (inputs(248));
    layer0_outputs(1256) <= inputs(100);
    layer0_outputs(1257) <= (inputs(151)) or (inputs(101));
    layer0_outputs(1258) <= not((inputs(185)) and (inputs(143)));
    layer0_outputs(1259) <= not((inputs(74)) xor (inputs(63)));
    layer0_outputs(1260) <= (inputs(26)) and (inputs(216));
    layer0_outputs(1261) <= (inputs(33)) and (inputs(33));
    layer0_outputs(1262) <= (inputs(92)) or (inputs(224));
    layer0_outputs(1263) <= not(inputs(91)) or (inputs(121));
    layer0_outputs(1264) <= not(inputs(231)) or (inputs(15));
    layer0_outputs(1265) <= inputs(209);
    layer0_outputs(1266) <= not((inputs(162)) or (inputs(197)));
    layer0_outputs(1267) <= '0';
    layer0_outputs(1268) <= not(inputs(205));
    layer0_outputs(1269) <= not(inputs(100));
    layer0_outputs(1270) <= not((inputs(61)) or (inputs(55)));
    layer0_outputs(1271) <= (inputs(61)) or (inputs(187));
    layer0_outputs(1272) <= not((inputs(59)) or (inputs(17)));
    layer0_outputs(1273) <= not(inputs(90)) or (inputs(117));
    layer0_outputs(1274) <= not((inputs(141)) or (inputs(83)));
    layer0_outputs(1275) <= '1';
    layer0_outputs(1276) <= not(inputs(128));
    layer0_outputs(1277) <= (inputs(248)) xor (inputs(128));
    layer0_outputs(1278) <= (inputs(189)) and not (inputs(48));
    layer0_outputs(1279) <= (inputs(135)) and not (inputs(126));
    layer0_outputs(1280) <= not((inputs(63)) or (inputs(56)));
    layer0_outputs(1281) <= inputs(145);
    layer0_outputs(1282) <= not((inputs(152)) and (inputs(29)));
    layer0_outputs(1283) <= not((inputs(224)) or (inputs(187)));
    layer0_outputs(1284) <= (inputs(200)) and (inputs(240));
    layer0_outputs(1285) <= inputs(106);
    layer0_outputs(1286) <= '1';
    layer0_outputs(1287) <= '0';
    layer0_outputs(1288) <= (inputs(115)) and not (inputs(104));
    layer0_outputs(1289) <= (inputs(105)) and not (inputs(112));
    layer0_outputs(1290) <= inputs(41);
    layer0_outputs(1291) <= not((inputs(185)) and (inputs(215)));
    layer0_outputs(1292) <= not(inputs(66));
    layer0_outputs(1293) <= inputs(201);
    layer0_outputs(1294) <= inputs(180);
    layer0_outputs(1295) <= (inputs(111)) or (inputs(48));
    layer0_outputs(1296) <= not(inputs(150));
    layer0_outputs(1297) <= (inputs(58)) xor (inputs(45));
    layer0_outputs(1298) <= (inputs(65)) or (inputs(197));
    layer0_outputs(1299) <= not((inputs(93)) or (inputs(238)));
    layer0_outputs(1300) <= inputs(140);
    layer0_outputs(1301) <= not(inputs(211));
    layer0_outputs(1302) <= not(inputs(92)) or (inputs(3));
    layer0_outputs(1303) <= not(inputs(176)) or (inputs(73));
    layer0_outputs(1304) <= (inputs(101)) and not (inputs(17));
    layer0_outputs(1305) <= (inputs(77)) and not (inputs(25));
    layer0_outputs(1306) <= '0';
    layer0_outputs(1307) <= not(inputs(233));
    layer0_outputs(1308) <= '1';
    layer0_outputs(1309) <= not(inputs(104)) or (inputs(246));
    layer0_outputs(1310) <= not((inputs(139)) and (inputs(116)));
    layer0_outputs(1311) <= not((inputs(159)) or (inputs(3)));
    layer0_outputs(1312) <= not((inputs(77)) or (inputs(95)));
    layer0_outputs(1313) <= not(inputs(130)) or (inputs(16));
    layer0_outputs(1314) <= '0';
    layer0_outputs(1315) <= not((inputs(73)) xor (inputs(173)));
    layer0_outputs(1316) <= inputs(77);
    layer0_outputs(1317) <= (inputs(19)) xor (inputs(190));
    layer0_outputs(1318) <= not(inputs(78));
    layer0_outputs(1319) <= not(inputs(56));
    layer0_outputs(1320) <= (inputs(102)) xor (inputs(82));
    layer0_outputs(1321) <= (inputs(205)) or (inputs(153));
    layer0_outputs(1322) <= not((inputs(203)) or (inputs(28)));
    layer0_outputs(1323) <= not((inputs(50)) or (inputs(205)));
    layer0_outputs(1324) <= '1';
    layer0_outputs(1325) <= (inputs(246)) or (inputs(204));
    layer0_outputs(1326) <= inputs(228);
    layer0_outputs(1327) <= inputs(213);
    layer0_outputs(1328) <= not((inputs(88)) or (inputs(59)));
    layer0_outputs(1329) <= not(inputs(134)) or (inputs(221));
    layer0_outputs(1330) <= not(inputs(181));
    layer0_outputs(1331) <= '1';
    layer0_outputs(1332) <= not(inputs(230)) or (inputs(6));
    layer0_outputs(1333) <= not((inputs(152)) xor (inputs(94)));
    layer0_outputs(1334) <= (inputs(84)) and not (inputs(228));
    layer0_outputs(1335) <= not(inputs(242)) or (inputs(132));
    layer0_outputs(1336) <= not((inputs(95)) or (inputs(170)));
    layer0_outputs(1337) <= not((inputs(75)) and (inputs(68)));
    layer0_outputs(1338) <= (inputs(7)) and not (inputs(171));
    layer0_outputs(1339) <= (inputs(120)) and not (inputs(35));
    layer0_outputs(1340) <= not((inputs(215)) and (inputs(117)));
    layer0_outputs(1341) <= not((inputs(83)) and (inputs(165)));
    layer0_outputs(1342) <= '1';
    layer0_outputs(1343) <= not((inputs(32)) and (inputs(145)));
    layer0_outputs(1344) <= not(inputs(247));
    layer0_outputs(1345) <= not((inputs(69)) or (inputs(45)));
    layer0_outputs(1346) <= not(inputs(96));
    layer0_outputs(1347) <= inputs(168);
    layer0_outputs(1348) <= not(inputs(95)) or (inputs(139));
    layer0_outputs(1349) <= inputs(98);
    layer0_outputs(1350) <= not((inputs(144)) xor (inputs(46)));
    layer0_outputs(1351) <= inputs(60);
    layer0_outputs(1352) <= (inputs(189)) or (inputs(226));
    layer0_outputs(1353) <= not(inputs(76));
    layer0_outputs(1354) <= inputs(250);
    layer0_outputs(1355) <= not(inputs(142));
    layer0_outputs(1356) <= inputs(223);
    layer0_outputs(1357) <= not((inputs(241)) or (inputs(154)));
    layer0_outputs(1358) <= '1';
    layer0_outputs(1359) <= (inputs(125)) or (inputs(73));
    layer0_outputs(1360) <= inputs(83);
    layer0_outputs(1361) <= (inputs(238)) and (inputs(156));
    layer0_outputs(1362) <= (inputs(141)) and (inputs(114));
    layer0_outputs(1363) <= (inputs(134)) or (inputs(105));
    layer0_outputs(1364) <= '1';
    layer0_outputs(1365) <= not(inputs(232));
    layer0_outputs(1366) <= (inputs(96)) or (inputs(71));
    layer0_outputs(1367) <= (inputs(217)) and (inputs(121));
    layer0_outputs(1368) <= (inputs(61)) and not (inputs(226));
    layer0_outputs(1369) <= not(inputs(68));
    layer0_outputs(1370) <= not(inputs(0)) or (inputs(221));
    layer0_outputs(1371) <= (inputs(96)) or (inputs(0));
    layer0_outputs(1372) <= not(inputs(159)) or (inputs(141));
    layer0_outputs(1373) <= (inputs(207)) and (inputs(125));
    layer0_outputs(1374) <= not(inputs(181)) or (inputs(71));
    layer0_outputs(1375) <= (inputs(96)) or (inputs(80));
    layer0_outputs(1376) <= not(inputs(167));
    layer0_outputs(1377) <= inputs(144);
    layer0_outputs(1378) <= not((inputs(80)) or (inputs(192)));
    layer0_outputs(1379) <= not(inputs(251)) or (inputs(248));
    layer0_outputs(1380) <= not(inputs(133));
    layer0_outputs(1381) <= not(inputs(197));
    layer0_outputs(1382) <= inputs(13);
    layer0_outputs(1383) <= (inputs(73)) or (inputs(12));
    layer0_outputs(1384) <= not((inputs(117)) or (inputs(24)));
    layer0_outputs(1385) <= (inputs(53)) or (inputs(114));
    layer0_outputs(1386) <= inputs(126);
    layer0_outputs(1387) <= not(inputs(211)) or (inputs(62));
    layer0_outputs(1388) <= not(inputs(19)) or (inputs(11));
    layer0_outputs(1389) <= not((inputs(133)) xor (inputs(161)));
    layer0_outputs(1390) <= not(inputs(163));
    layer0_outputs(1391) <= (inputs(7)) and not (inputs(136));
    layer0_outputs(1392) <= (inputs(194)) and not (inputs(228));
    layer0_outputs(1393) <= not(inputs(63)) or (inputs(200));
    layer0_outputs(1394) <= (inputs(208)) and not (inputs(110));
    layer0_outputs(1395) <= (inputs(84)) and not (inputs(72));
    layer0_outputs(1396) <= (inputs(194)) and (inputs(1));
    layer0_outputs(1397) <= inputs(102);
    layer0_outputs(1398) <= (inputs(45)) and not (inputs(10));
    layer0_outputs(1399) <= not((inputs(32)) xor (inputs(118)));
    layer0_outputs(1400) <= not((inputs(165)) or (inputs(104)));
    layer0_outputs(1401) <= (inputs(199)) and not (inputs(173));
    layer0_outputs(1402) <= inputs(244);
    layer0_outputs(1403) <= not((inputs(56)) or (inputs(160)));
    layer0_outputs(1404) <= inputs(243);
    layer0_outputs(1405) <= not(inputs(10)) or (inputs(237));
    layer0_outputs(1406) <= not((inputs(133)) xor (inputs(37)));
    layer0_outputs(1407) <= not(inputs(183));
    layer0_outputs(1408) <= '0';
    layer0_outputs(1409) <= inputs(131);
    layer0_outputs(1410) <= inputs(233);
    layer0_outputs(1411) <= (inputs(65)) or (inputs(204));
    layer0_outputs(1412) <= inputs(70);
    layer0_outputs(1413) <= (inputs(108)) or (inputs(42));
    layer0_outputs(1414) <= '1';
    layer0_outputs(1415) <= not(inputs(115)) or (inputs(41));
    layer0_outputs(1416) <= not((inputs(30)) and (inputs(156)));
    layer0_outputs(1417) <= (inputs(110)) or (inputs(153));
    layer0_outputs(1418) <= (inputs(27)) xor (inputs(58));
    layer0_outputs(1419) <= not((inputs(128)) xor (inputs(82)));
    layer0_outputs(1420) <= not(inputs(120));
    layer0_outputs(1421) <= '0';
    layer0_outputs(1422) <= not(inputs(134)) or (inputs(241));
    layer0_outputs(1423) <= '1';
    layer0_outputs(1424) <= '1';
    layer0_outputs(1425) <= not(inputs(60));
    layer0_outputs(1426) <= (inputs(46)) and not (inputs(124));
    layer0_outputs(1427) <= inputs(14);
    layer0_outputs(1428) <= not((inputs(126)) xor (inputs(18)));
    layer0_outputs(1429) <= not((inputs(166)) or (inputs(93)));
    layer0_outputs(1430) <= not(inputs(157)) or (inputs(34));
    layer0_outputs(1431) <= (inputs(111)) xor (inputs(157));
    layer0_outputs(1432) <= not((inputs(178)) or (inputs(226)));
    layer0_outputs(1433) <= (inputs(6)) or (inputs(57));
    layer0_outputs(1434) <= (inputs(100)) and (inputs(83));
    layer0_outputs(1435) <= inputs(28);
    layer0_outputs(1436) <= (inputs(231)) xor (inputs(199));
    layer0_outputs(1437) <= not(inputs(250));
    layer0_outputs(1438) <= (inputs(58)) xor (inputs(40));
    layer0_outputs(1439) <= inputs(162);
    layer0_outputs(1440) <= not(inputs(231));
    layer0_outputs(1441) <= not((inputs(186)) or (inputs(202)));
    layer0_outputs(1442) <= not(inputs(188)) or (inputs(22));
    layer0_outputs(1443) <= not(inputs(232));
    layer0_outputs(1444) <= (inputs(194)) and not (inputs(31));
    layer0_outputs(1445) <= not((inputs(107)) or (inputs(141)));
    layer0_outputs(1446) <= not((inputs(102)) xor (inputs(82)));
    layer0_outputs(1447) <= not(inputs(253));
    layer0_outputs(1448) <= (inputs(193)) or (inputs(236));
    layer0_outputs(1449) <= '1';
    layer0_outputs(1450) <= not(inputs(170));
    layer0_outputs(1451) <= inputs(223);
    layer0_outputs(1452) <= inputs(90);
    layer0_outputs(1453) <= inputs(100);
    layer0_outputs(1454) <= not((inputs(188)) xor (inputs(195)));
    layer0_outputs(1455) <= not(inputs(100));
    layer0_outputs(1456) <= not(inputs(218)) or (inputs(152));
    layer0_outputs(1457) <= not(inputs(152)) or (inputs(143));
    layer0_outputs(1458) <= '0';
    layer0_outputs(1459) <= (inputs(107)) xor (inputs(63));
    layer0_outputs(1460) <= inputs(147);
    layer0_outputs(1461) <= not((inputs(55)) or (inputs(20)));
    layer0_outputs(1462) <= (inputs(199)) and not (inputs(19));
    layer0_outputs(1463) <= (inputs(75)) xor (inputs(27));
    layer0_outputs(1464) <= (inputs(178)) and not (inputs(202));
    layer0_outputs(1465) <= not(inputs(223));
    layer0_outputs(1466) <= '0';
    layer0_outputs(1467) <= not(inputs(167));
    layer0_outputs(1468) <= not(inputs(155));
    layer0_outputs(1469) <= (inputs(89)) or (inputs(1));
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= inputs(4);
    layer0_outputs(1472) <= not((inputs(46)) or (inputs(196)));
    layer0_outputs(1473) <= (inputs(197)) and not (inputs(69));
    layer0_outputs(1474) <= inputs(233);
    layer0_outputs(1475) <= inputs(15);
    layer0_outputs(1476) <= (inputs(200)) and not (inputs(10));
    layer0_outputs(1477) <= (inputs(218)) or (inputs(172));
    layer0_outputs(1478) <= '0';
    layer0_outputs(1479) <= '0';
    layer0_outputs(1480) <= (inputs(183)) and not (inputs(12));
    layer0_outputs(1481) <= (inputs(254)) and not (inputs(131));
    layer0_outputs(1482) <= inputs(127);
    layer0_outputs(1483) <= not(inputs(102));
    layer0_outputs(1484) <= (inputs(135)) or (inputs(147));
    layer0_outputs(1485) <= not((inputs(73)) xor (inputs(36)));
    layer0_outputs(1486) <= not((inputs(79)) xor (inputs(201)));
    layer0_outputs(1487) <= not(inputs(221));
    layer0_outputs(1488) <= '1';
    layer0_outputs(1489) <= not(inputs(211));
    layer0_outputs(1490) <= not((inputs(222)) xor (inputs(126)));
    layer0_outputs(1491) <= (inputs(230)) and not (inputs(30));
    layer0_outputs(1492) <= '0';
    layer0_outputs(1493) <= inputs(141);
    layer0_outputs(1494) <= not(inputs(184)) or (inputs(60));
    layer0_outputs(1495) <= (inputs(212)) or (inputs(9));
    layer0_outputs(1496) <= (inputs(64)) or (inputs(156));
    layer0_outputs(1497) <= inputs(100);
    layer0_outputs(1498) <= (inputs(133)) or (inputs(67));
    layer0_outputs(1499) <= '1';
    layer0_outputs(1500) <= not((inputs(21)) or (inputs(105)));
    layer0_outputs(1501) <= (inputs(171)) and not (inputs(57));
    layer0_outputs(1502) <= (inputs(245)) or (inputs(97));
    layer0_outputs(1503) <= inputs(228);
    layer0_outputs(1504) <= inputs(115);
    layer0_outputs(1505) <= (inputs(176)) xor (inputs(117));
    layer0_outputs(1506) <= not(inputs(126)) or (inputs(25));
    layer0_outputs(1507) <= inputs(108);
    layer0_outputs(1508) <= not(inputs(211));
    layer0_outputs(1509) <= not(inputs(214)) or (inputs(35));
    layer0_outputs(1510) <= (inputs(181)) and not (inputs(1));
    layer0_outputs(1511) <= not((inputs(211)) or (inputs(211)));
    layer0_outputs(1512) <= not(inputs(247)) or (inputs(2));
    layer0_outputs(1513) <= inputs(85);
    layer0_outputs(1514) <= (inputs(201)) and not (inputs(44));
    layer0_outputs(1515) <= not((inputs(79)) xor (inputs(205)));
    layer0_outputs(1516) <= (inputs(183)) xor (inputs(169));
    layer0_outputs(1517) <= not(inputs(183)) or (inputs(225));
    layer0_outputs(1518) <= (inputs(237)) xor (inputs(48));
    layer0_outputs(1519) <= not((inputs(167)) or (inputs(148)));
    layer0_outputs(1520) <= not(inputs(62));
    layer0_outputs(1521) <= (inputs(100)) and (inputs(120));
    layer0_outputs(1522) <= (inputs(140)) xor (inputs(104));
    layer0_outputs(1523) <= (inputs(197)) or (inputs(182));
    layer0_outputs(1524) <= not(inputs(169));
    layer0_outputs(1525) <= (inputs(180)) and (inputs(111));
    layer0_outputs(1526) <= not(inputs(100)) or (inputs(48));
    layer0_outputs(1527) <= inputs(113);
    layer0_outputs(1528) <= inputs(27);
    layer0_outputs(1529) <= (inputs(110)) and not (inputs(248));
    layer0_outputs(1530) <= (inputs(206)) or (inputs(173));
    layer0_outputs(1531) <= (inputs(33)) and not (inputs(69));
    layer0_outputs(1532) <= not(inputs(92)) or (inputs(178));
    layer0_outputs(1533) <= (inputs(134)) and not (inputs(144));
    layer0_outputs(1534) <= not((inputs(31)) xor (inputs(217)));
    layer0_outputs(1535) <= (inputs(16)) or (inputs(73));
    layer0_outputs(1536) <= inputs(30);
    layer0_outputs(1537) <= not((inputs(242)) or (inputs(218)));
    layer0_outputs(1538) <= inputs(231);
    layer0_outputs(1539) <= not(inputs(142)) or (inputs(85));
    layer0_outputs(1540) <= '1';
    layer0_outputs(1541) <= not(inputs(70));
    layer0_outputs(1542) <= (inputs(76)) and not (inputs(116));
    layer0_outputs(1543) <= not(inputs(250));
    layer0_outputs(1544) <= '0';
    layer0_outputs(1545) <= not(inputs(255));
    layer0_outputs(1546) <= inputs(233);
    layer0_outputs(1547) <= (inputs(187)) or (inputs(24));
    layer0_outputs(1548) <= inputs(129);
    layer0_outputs(1549) <= not(inputs(145));
    layer0_outputs(1550) <= (inputs(105)) or (inputs(102));
    layer0_outputs(1551) <= inputs(202);
    layer0_outputs(1552) <= (inputs(193)) or (inputs(181));
    layer0_outputs(1553) <= not((inputs(156)) or (inputs(161)));
    layer0_outputs(1554) <= inputs(221);
    layer0_outputs(1555) <= not((inputs(253)) xor (inputs(219)));
    layer0_outputs(1556) <= (inputs(27)) or (inputs(18));
    layer0_outputs(1557) <= (inputs(215)) and not (inputs(87));
    layer0_outputs(1558) <= '0';
    layer0_outputs(1559) <= not((inputs(32)) or (inputs(219)));
    layer0_outputs(1560) <= inputs(131);
    layer0_outputs(1561) <= (inputs(229)) and not (inputs(151));
    layer0_outputs(1562) <= (inputs(2)) and not (inputs(212));
    layer0_outputs(1563) <= not((inputs(12)) and (inputs(217)));
    layer0_outputs(1564) <= not(inputs(212)) or (inputs(130));
    layer0_outputs(1565) <= '0';
    layer0_outputs(1566) <= inputs(150);
    layer0_outputs(1567) <= not(inputs(180));
    layer0_outputs(1568) <= not(inputs(64)) or (inputs(7));
    layer0_outputs(1569) <= not(inputs(165));
    layer0_outputs(1570) <= (inputs(144)) and (inputs(240));
    layer0_outputs(1571) <= not(inputs(32)) or (inputs(48));
    layer0_outputs(1572) <= not(inputs(231));
    layer0_outputs(1573) <= '1';
    layer0_outputs(1574) <= not(inputs(93));
    layer0_outputs(1575) <= inputs(190);
    layer0_outputs(1576) <= not(inputs(124)) or (inputs(222));
    layer0_outputs(1577) <= not((inputs(210)) or (inputs(253)));
    layer0_outputs(1578) <= not(inputs(113));
    layer0_outputs(1579) <= (inputs(12)) and not (inputs(159));
    layer0_outputs(1580) <= not(inputs(184));
    layer0_outputs(1581) <= not(inputs(10));
    layer0_outputs(1582) <= (inputs(191)) or (inputs(39));
    layer0_outputs(1583) <= not(inputs(125));
    layer0_outputs(1584) <= not(inputs(147));
    layer0_outputs(1585) <= inputs(131);
    layer0_outputs(1586) <= not(inputs(67));
    layer0_outputs(1587) <= not((inputs(194)) or (inputs(215)));
    layer0_outputs(1588) <= (inputs(220)) or (inputs(127));
    layer0_outputs(1589) <= '1';
    layer0_outputs(1590) <= not(inputs(91)) or (inputs(130));
    layer0_outputs(1591) <= inputs(15);
    layer0_outputs(1592) <= not(inputs(100)) or (inputs(165));
    layer0_outputs(1593) <= not(inputs(178));
    layer0_outputs(1594) <= not((inputs(77)) or (inputs(110)));
    layer0_outputs(1595) <= (inputs(120)) xor (inputs(192));
    layer0_outputs(1596) <= not((inputs(121)) or (inputs(102)));
    layer0_outputs(1597) <= inputs(127);
    layer0_outputs(1598) <= (inputs(90)) or (inputs(132));
    layer0_outputs(1599) <= not(inputs(215));
    layer0_outputs(1600) <= inputs(182);
    layer0_outputs(1601) <= (inputs(63)) or (inputs(188));
    layer0_outputs(1602) <= not(inputs(169));
    layer0_outputs(1603) <= not(inputs(25));
    layer0_outputs(1604) <= not((inputs(111)) or (inputs(49)));
    layer0_outputs(1605) <= not((inputs(221)) or (inputs(146)));
    layer0_outputs(1606) <= '0';
    layer0_outputs(1607) <= not(inputs(237)) or (inputs(58));
    layer0_outputs(1608) <= not((inputs(34)) and (inputs(48)));
    layer0_outputs(1609) <= (inputs(132)) xor (inputs(101));
    layer0_outputs(1610) <= not(inputs(203)) or (inputs(229));
    layer0_outputs(1611) <= not((inputs(231)) or (inputs(116)));
    layer0_outputs(1612) <= (inputs(161)) and not (inputs(168));
    layer0_outputs(1613) <= not(inputs(245));
    layer0_outputs(1614) <= (inputs(253)) and not (inputs(34));
    layer0_outputs(1615) <= inputs(0);
    layer0_outputs(1616) <= not((inputs(203)) or (inputs(53)));
    layer0_outputs(1617) <= not(inputs(110));
    layer0_outputs(1618) <= not((inputs(212)) or (inputs(236)));
    layer0_outputs(1619) <= not(inputs(70)) or (inputs(146));
    layer0_outputs(1620) <= '0';
    layer0_outputs(1621) <= not(inputs(212));
    layer0_outputs(1622) <= not(inputs(163));
    layer0_outputs(1623) <= (inputs(47)) or (inputs(203));
    layer0_outputs(1624) <= not((inputs(221)) xor (inputs(160)));
    layer0_outputs(1625) <= inputs(56);
    layer0_outputs(1626) <= not(inputs(217));
    layer0_outputs(1627) <= not(inputs(219));
    layer0_outputs(1628) <= (inputs(57)) or (inputs(142));
    layer0_outputs(1629) <= inputs(98);
    layer0_outputs(1630) <= (inputs(207)) xor (inputs(158));
    layer0_outputs(1631) <= (inputs(251)) or (inputs(210));
    layer0_outputs(1632) <= (inputs(140)) and not (inputs(178));
    layer0_outputs(1633) <= inputs(25);
    layer0_outputs(1634) <= (inputs(108)) xor (inputs(157));
    layer0_outputs(1635) <= (inputs(89)) xor (inputs(42));
    layer0_outputs(1636) <= not((inputs(23)) or (inputs(242)));
    layer0_outputs(1637) <= not((inputs(78)) or (inputs(162)));
    layer0_outputs(1638) <= (inputs(133)) and not (inputs(0));
    layer0_outputs(1639) <= inputs(113);
    layer0_outputs(1640) <= (inputs(23)) or (inputs(171));
    layer0_outputs(1641) <= (inputs(190)) and (inputs(129));
    layer0_outputs(1642) <= (inputs(28)) xor (inputs(206));
    layer0_outputs(1643) <= inputs(34);
    layer0_outputs(1644) <= (inputs(208)) xor (inputs(211));
    layer0_outputs(1645) <= not(inputs(198)) or (inputs(62));
    layer0_outputs(1646) <= not(inputs(91));
    layer0_outputs(1647) <= not((inputs(222)) or (inputs(100)));
    layer0_outputs(1648) <= inputs(235);
    layer0_outputs(1649) <= (inputs(173)) or (inputs(91));
    layer0_outputs(1650) <= not(inputs(90));
    layer0_outputs(1651) <= (inputs(44)) or (inputs(232));
    layer0_outputs(1652) <= not((inputs(150)) xor (inputs(72)));
    layer0_outputs(1653) <= not(inputs(146));
    layer0_outputs(1654) <= inputs(61);
    layer0_outputs(1655) <= not(inputs(213));
    layer0_outputs(1656) <= (inputs(134)) or (inputs(112));
    layer0_outputs(1657) <= (inputs(240)) or (inputs(45));
    layer0_outputs(1658) <= (inputs(169)) and not (inputs(6));
    layer0_outputs(1659) <= not(inputs(80));
    layer0_outputs(1660) <= inputs(200);
    layer0_outputs(1661) <= not((inputs(4)) or (inputs(77)));
    layer0_outputs(1662) <= (inputs(42)) and not (inputs(56));
    layer0_outputs(1663) <= '0';
    layer0_outputs(1664) <= not(inputs(163)) or (inputs(95));
    layer0_outputs(1665) <= not((inputs(95)) or (inputs(246)));
    layer0_outputs(1666) <= (inputs(135)) xor (inputs(242));
    layer0_outputs(1667) <= (inputs(156)) xor (inputs(143));
    layer0_outputs(1668) <= (inputs(49)) xor (inputs(236));
    layer0_outputs(1669) <= (inputs(16)) and not (inputs(60));
    layer0_outputs(1670) <= not(inputs(92)) or (inputs(241));
    layer0_outputs(1671) <= inputs(26);
    layer0_outputs(1672) <= '1';
    layer0_outputs(1673) <= (inputs(180)) xor (inputs(43));
    layer0_outputs(1674) <= (inputs(57)) or (inputs(29));
    layer0_outputs(1675) <= not((inputs(9)) or (inputs(27)));
    layer0_outputs(1676) <= not(inputs(82));
    layer0_outputs(1677) <= not(inputs(77)) or (inputs(240));
    layer0_outputs(1678) <= not(inputs(32));
    layer0_outputs(1679) <= not(inputs(85));
    layer0_outputs(1680) <= not(inputs(147));
    layer0_outputs(1681) <= (inputs(5)) xor (inputs(91));
    layer0_outputs(1682) <= '0';
    layer0_outputs(1683) <= not((inputs(207)) xor (inputs(221)));
    layer0_outputs(1684) <= not((inputs(11)) and (inputs(94)));
    layer0_outputs(1685) <= not((inputs(193)) or (inputs(214)));
    layer0_outputs(1686) <= not(inputs(123)) or (inputs(226));
    layer0_outputs(1687) <= inputs(111);
    layer0_outputs(1688) <= (inputs(246)) xor (inputs(198));
    layer0_outputs(1689) <= not((inputs(170)) and (inputs(139)));
    layer0_outputs(1690) <= inputs(30);
    layer0_outputs(1691) <= not((inputs(5)) and (inputs(137)));
    layer0_outputs(1692) <= inputs(181);
    layer0_outputs(1693) <= not((inputs(230)) or (inputs(244)));
    layer0_outputs(1694) <= not((inputs(206)) or (inputs(32)));
    layer0_outputs(1695) <= not((inputs(17)) and (inputs(196)));
    layer0_outputs(1696) <= not((inputs(42)) xor (inputs(220)));
    layer0_outputs(1697) <= not((inputs(91)) and (inputs(237)));
    layer0_outputs(1698) <= (inputs(195)) and not (inputs(124));
    layer0_outputs(1699) <= not(inputs(113));
    layer0_outputs(1700) <= (inputs(22)) and not (inputs(19));
    layer0_outputs(1701) <= inputs(0);
    layer0_outputs(1702) <= (inputs(105)) or (inputs(93));
    layer0_outputs(1703) <= not((inputs(184)) or (inputs(179)));
    layer0_outputs(1704) <= not(inputs(183)) or (inputs(106));
    layer0_outputs(1705) <= inputs(67);
    layer0_outputs(1706) <= (inputs(29)) xor (inputs(168));
    layer0_outputs(1707) <= (inputs(151)) and (inputs(9));
    layer0_outputs(1708) <= not(inputs(198)) or (inputs(62));
    layer0_outputs(1709) <= (inputs(241)) xor (inputs(195));
    layer0_outputs(1710) <= not((inputs(225)) or (inputs(68)));
    layer0_outputs(1711) <= not((inputs(157)) xor (inputs(221)));
    layer0_outputs(1712) <= (inputs(3)) and (inputs(48));
    layer0_outputs(1713) <= (inputs(167)) xor (inputs(5));
    layer0_outputs(1714) <= '1';
    layer0_outputs(1715) <= inputs(86);
    layer0_outputs(1716) <= inputs(201);
    layer0_outputs(1717) <= not(inputs(56));
    layer0_outputs(1718) <= inputs(200);
    layer0_outputs(1719) <= not((inputs(43)) xor (inputs(7)));
    layer0_outputs(1720) <= inputs(30);
    layer0_outputs(1721) <= (inputs(2)) and not (inputs(207));
    layer0_outputs(1722) <= (inputs(135)) and not (inputs(77));
    layer0_outputs(1723) <= (inputs(123)) and not (inputs(50));
    layer0_outputs(1724) <= not((inputs(234)) or (inputs(212)));
    layer0_outputs(1725) <= inputs(89);
    layer0_outputs(1726) <= (inputs(221)) and not (inputs(81));
    layer0_outputs(1727) <= not(inputs(191));
    layer0_outputs(1728) <= inputs(129);
    layer0_outputs(1729) <= not(inputs(139)) or (inputs(62));
    layer0_outputs(1730) <= inputs(174);
    layer0_outputs(1731) <= not(inputs(159));
    layer0_outputs(1732) <= (inputs(13)) xor (inputs(30));
    layer0_outputs(1733) <= not(inputs(137));
    layer0_outputs(1734) <= not(inputs(44));
    layer0_outputs(1735) <= inputs(192);
    layer0_outputs(1736) <= inputs(66);
    layer0_outputs(1737) <= inputs(122);
    layer0_outputs(1738) <= '1';
    layer0_outputs(1739) <= not(inputs(116));
    layer0_outputs(1740) <= not(inputs(131)) or (inputs(18));
    layer0_outputs(1741) <= inputs(46);
    layer0_outputs(1742) <= (inputs(183)) and not (inputs(183));
    layer0_outputs(1743) <= inputs(121);
    layer0_outputs(1744) <= inputs(149);
    layer0_outputs(1745) <= not(inputs(182));
    layer0_outputs(1746) <= inputs(59);
    layer0_outputs(1747) <= (inputs(133)) and (inputs(4));
    layer0_outputs(1748) <= not(inputs(12)) or (inputs(93));
    layer0_outputs(1749) <= not((inputs(61)) or (inputs(143)));
    layer0_outputs(1750) <= not(inputs(184)) or (inputs(128));
    layer0_outputs(1751) <= not((inputs(152)) or (inputs(1)));
    layer0_outputs(1752) <= not(inputs(13));
    layer0_outputs(1753) <= not(inputs(193));
    layer0_outputs(1754) <= not(inputs(78)) or (inputs(238));
    layer0_outputs(1755) <= (inputs(142)) or (inputs(173));
    layer0_outputs(1756) <= (inputs(213)) xor (inputs(248));
    layer0_outputs(1757) <= '0';
    layer0_outputs(1758) <= inputs(255);
    layer0_outputs(1759) <= inputs(116);
    layer0_outputs(1760) <= inputs(230);
    layer0_outputs(1761) <= (inputs(247)) and not (inputs(36));
    layer0_outputs(1762) <= not(inputs(49)) or (inputs(191));
    layer0_outputs(1763) <= not(inputs(235));
    layer0_outputs(1764) <= (inputs(103)) and (inputs(231));
    layer0_outputs(1765) <= (inputs(103)) or (inputs(224));
    layer0_outputs(1766) <= not(inputs(88));
    layer0_outputs(1767) <= inputs(134);
    layer0_outputs(1768) <= (inputs(96)) and not (inputs(34));
    layer0_outputs(1769) <= not(inputs(106)) or (inputs(196));
    layer0_outputs(1770) <= not(inputs(59));
    layer0_outputs(1771) <= not(inputs(37)) or (inputs(179));
    layer0_outputs(1772) <= not(inputs(84));
    layer0_outputs(1773) <= inputs(93);
    layer0_outputs(1774) <= (inputs(190)) and (inputs(119));
    layer0_outputs(1775) <= not(inputs(37)) or (inputs(251));
    layer0_outputs(1776) <= (inputs(70)) or (inputs(120));
    layer0_outputs(1777) <= not(inputs(169));
    layer0_outputs(1778) <= inputs(236);
    layer0_outputs(1779) <= (inputs(147)) and not (inputs(81));
    layer0_outputs(1780) <= not(inputs(67)) or (inputs(127));
    layer0_outputs(1781) <= inputs(161);
    layer0_outputs(1782) <= not(inputs(126)) or (inputs(152));
    layer0_outputs(1783) <= (inputs(156)) and not (inputs(82));
    layer0_outputs(1784) <= not((inputs(136)) and (inputs(169)));
    layer0_outputs(1785) <= (inputs(24)) xor (inputs(47));
    layer0_outputs(1786) <= (inputs(69)) or (inputs(79));
    layer0_outputs(1787) <= (inputs(50)) and not (inputs(0));
    layer0_outputs(1788) <= not((inputs(205)) xor (inputs(45)));
    layer0_outputs(1789) <= inputs(148);
    layer0_outputs(1790) <= inputs(176);
    layer0_outputs(1791) <= inputs(43);
    layer0_outputs(1792) <= not(inputs(84));
    layer0_outputs(1793) <= not(inputs(91));
    layer0_outputs(1794) <= not((inputs(93)) or (inputs(28)));
    layer0_outputs(1795) <= (inputs(88)) and not (inputs(181));
    layer0_outputs(1796) <= (inputs(168)) or (inputs(76));
    layer0_outputs(1797) <= not((inputs(189)) or (inputs(197)));
    layer0_outputs(1798) <= (inputs(76)) and not (inputs(136));
    layer0_outputs(1799) <= not(inputs(118));
    layer0_outputs(1800) <= not(inputs(66));
    layer0_outputs(1801) <= inputs(77);
    layer0_outputs(1802) <= not(inputs(74)) or (inputs(47));
    layer0_outputs(1803) <= not(inputs(74)) or (inputs(31));
    layer0_outputs(1804) <= not(inputs(189));
    layer0_outputs(1805) <= (inputs(248)) xor (inputs(200));
    layer0_outputs(1806) <= not(inputs(253)) or (inputs(127));
    layer0_outputs(1807) <= '1';
    layer0_outputs(1808) <= inputs(106);
    layer0_outputs(1809) <= not((inputs(59)) xor (inputs(88)));
    layer0_outputs(1810) <= (inputs(211)) or (inputs(42));
    layer0_outputs(1811) <= not((inputs(157)) xor (inputs(70)));
    layer0_outputs(1812) <= '0';
    layer0_outputs(1813) <= (inputs(148)) or (inputs(107));
    layer0_outputs(1814) <= not(inputs(52));
    layer0_outputs(1815) <= not(inputs(177));
    layer0_outputs(1816) <= inputs(89);
    layer0_outputs(1817) <= (inputs(150)) and not (inputs(45));
    layer0_outputs(1818) <= not((inputs(83)) and (inputs(98)));
    layer0_outputs(1819) <= (inputs(18)) or (inputs(202));
    layer0_outputs(1820) <= inputs(29);
    layer0_outputs(1821) <= inputs(179);
    layer0_outputs(1822) <= not((inputs(138)) xor (inputs(188)));
    layer0_outputs(1823) <= (inputs(193)) and (inputs(144));
    layer0_outputs(1824) <= (inputs(219)) and not (inputs(154));
    layer0_outputs(1825) <= inputs(112);
    layer0_outputs(1826) <= not(inputs(160));
    layer0_outputs(1827) <= not(inputs(49));
    layer0_outputs(1828) <= '1';
    layer0_outputs(1829) <= (inputs(88)) and not (inputs(49));
    layer0_outputs(1830) <= (inputs(27)) xor (inputs(78));
    layer0_outputs(1831) <= inputs(98);
    layer0_outputs(1832) <= (inputs(74)) xor (inputs(29));
    layer0_outputs(1833) <= inputs(211);
    layer0_outputs(1834) <= not(inputs(71));
    layer0_outputs(1835) <= not(inputs(208));
    layer0_outputs(1836) <= inputs(105);
    layer0_outputs(1837) <= not((inputs(115)) xor (inputs(31)));
    layer0_outputs(1838) <= not(inputs(247)) or (inputs(9));
    layer0_outputs(1839) <= not((inputs(188)) or (inputs(157)));
    layer0_outputs(1840) <= inputs(148);
    layer0_outputs(1841) <= not(inputs(27)) or (inputs(183));
    layer0_outputs(1842) <= (inputs(179)) or (inputs(204));
    layer0_outputs(1843) <= (inputs(151)) and not (inputs(226));
    layer0_outputs(1844) <= '0';
    layer0_outputs(1845) <= (inputs(231)) or (inputs(217));
    layer0_outputs(1846) <= (inputs(204)) or (inputs(201));
    layer0_outputs(1847) <= not(inputs(217)) or (inputs(84));
    layer0_outputs(1848) <= not((inputs(1)) and (inputs(23)));
    layer0_outputs(1849) <= not((inputs(173)) or (inputs(239)));
    layer0_outputs(1850) <= (inputs(50)) xor (inputs(112));
    layer0_outputs(1851) <= not(inputs(190)) or (inputs(32));
    layer0_outputs(1852) <= (inputs(235)) or (inputs(255));
    layer0_outputs(1853) <= inputs(25);
    layer0_outputs(1854) <= (inputs(114)) or (inputs(134));
    layer0_outputs(1855) <= inputs(80);
    layer0_outputs(1856) <= not(inputs(252)) or (inputs(113));
    layer0_outputs(1857) <= '1';
    layer0_outputs(1858) <= not((inputs(200)) and (inputs(122)));
    layer0_outputs(1859) <= inputs(162);
    layer0_outputs(1860) <= not((inputs(82)) xor (inputs(223)));
    layer0_outputs(1861) <= not(inputs(34)) or (inputs(235));
    layer0_outputs(1862) <= not(inputs(139));
    layer0_outputs(1863) <= (inputs(147)) and (inputs(154));
    layer0_outputs(1864) <= inputs(184);
    layer0_outputs(1865) <= inputs(34);
    layer0_outputs(1866) <= not(inputs(204));
    layer0_outputs(1867) <= not((inputs(74)) xor (inputs(64)));
    layer0_outputs(1868) <= '1';
    layer0_outputs(1869) <= inputs(253);
    layer0_outputs(1870) <= (inputs(229)) or (inputs(238));
    layer0_outputs(1871) <= inputs(173);
    layer0_outputs(1872) <= inputs(180);
    layer0_outputs(1873) <= (inputs(181)) xor (inputs(35));
    layer0_outputs(1874) <= not(inputs(52));
    layer0_outputs(1875) <= (inputs(126)) and not (inputs(35));
    layer0_outputs(1876) <= not((inputs(136)) or (inputs(61)));
    layer0_outputs(1877) <= not((inputs(237)) or (inputs(3)));
    layer0_outputs(1878) <= not(inputs(59));
    layer0_outputs(1879) <= not(inputs(167));
    layer0_outputs(1880) <= (inputs(33)) or (inputs(43));
    layer0_outputs(1881) <= not(inputs(246));
    layer0_outputs(1882) <= not((inputs(15)) xor (inputs(73)));
    layer0_outputs(1883) <= inputs(174);
    layer0_outputs(1884) <= inputs(196);
    layer0_outputs(1885) <= not(inputs(135)) or (inputs(96));
    layer0_outputs(1886) <= not((inputs(164)) or (inputs(197)));
    layer0_outputs(1887) <= not(inputs(96));
    layer0_outputs(1888) <= '0';
    layer0_outputs(1889) <= (inputs(181)) or (inputs(94));
    layer0_outputs(1890) <= not(inputs(61));
    layer0_outputs(1891) <= not(inputs(192));
    layer0_outputs(1892) <= not(inputs(185));
    layer0_outputs(1893) <= inputs(49);
    layer0_outputs(1894) <= (inputs(81)) xor (inputs(68));
    layer0_outputs(1895) <= inputs(213);
    layer0_outputs(1896) <= not((inputs(15)) xor (inputs(33)));
    layer0_outputs(1897) <= (inputs(149)) or (inputs(103));
    layer0_outputs(1898) <= (inputs(17)) xor (inputs(60));
    layer0_outputs(1899) <= inputs(189);
    layer0_outputs(1900) <= not(inputs(208));
    layer0_outputs(1901) <= not(inputs(252));
    layer0_outputs(1902) <= not((inputs(159)) or (inputs(113)));
    layer0_outputs(1903) <= inputs(122);
    layer0_outputs(1904) <= not((inputs(133)) or (inputs(55)));
    layer0_outputs(1905) <= not(inputs(111));
    layer0_outputs(1906) <= not(inputs(153));
    layer0_outputs(1907) <= not((inputs(80)) and (inputs(0)));
    layer0_outputs(1908) <= not((inputs(112)) or (inputs(125)));
    layer0_outputs(1909) <= (inputs(168)) and not (inputs(68));
    layer0_outputs(1910) <= (inputs(192)) or (inputs(49));
    layer0_outputs(1911) <= not((inputs(149)) or (inputs(174)));
    layer0_outputs(1912) <= (inputs(115)) xor (inputs(50));
    layer0_outputs(1913) <= not(inputs(224));
    layer0_outputs(1914) <= inputs(223);
    layer0_outputs(1915) <= not((inputs(48)) or (inputs(154)));
    layer0_outputs(1916) <= not((inputs(149)) or (inputs(237)));
    layer0_outputs(1917) <= inputs(182);
    layer0_outputs(1918) <= not(inputs(123)) or (inputs(146));
    layer0_outputs(1919) <= (inputs(205)) and not (inputs(64));
    layer0_outputs(1920) <= (inputs(12)) and not (inputs(26));
    layer0_outputs(1921) <= not(inputs(223));
    layer0_outputs(1922) <= not(inputs(141)) or (inputs(251));
    layer0_outputs(1923) <= (inputs(188)) xor (inputs(169));
    layer0_outputs(1924) <= not(inputs(36));
    layer0_outputs(1925) <= not(inputs(248));
    layer0_outputs(1926) <= '0';
    layer0_outputs(1927) <= not((inputs(86)) and (inputs(252)));
    layer0_outputs(1928) <= not(inputs(103)) or (inputs(58));
    layer0_outputs(1929) <= (inputs(76)) or (inputs(75));
    layer0_outputs(1930) <= not((inputs(62)) or (inputs(24)));
    layer0_outputs(1931) <= not((inputs(95)) xor (inputs(173)));
    layer0_outputs(1932) <= inputs(38);
    layer0_outputs(1933) <= (inputs(230)) or (inputs(173));
    layer0_outputs(1934) <= not(inputs(139)) or (inputs(177));
    layer0_outputs(1935) <= (inputs(149)) and not (inputs(123));
    layer0_outputs(1936) <= not(inputs(175));
    layer0_outputs(1937) <= '0';
    layer0_outputs(1938) <= not(inputs(140)) or (inputs(121));
    layer0_outputs(1939) <= (inputs(138)) and not (inputs(170));
    layer0_outputs(1940) <= not(inputs(184)) or (inputs(10));
    layer0_outputs(1941) <= not(inputs(176));
    layer0_outputs(1942) <= inputs(246);
    layer0_outputs(1943) <= (inputs(79)) or (inputs(97));
    layer0_outputs(1944) <= not(inputs(106)) or (inputs(98));
    layer0_outputs(1945) <= not((inputs(162)) or (inputs(232)));
    layer0_outputs(1946) <= not(inputs(169)) or (inputs(209));
    layer0_outputs(1947) <= not((inputs(144)) xor (inputs(32)));
    layer0_outputs(1948) <= not((inputs(49)) or (inputs(0)));
    layer0_outputs(1949) <= inputs(75);
    layer0_outputs(1950) <= (inputs(171)) and not (inputs(243));
    layer0_outputs(1951) <= '1';
    layer0_outputs(1952) <= not((inputs(231)) xor (inputs(151)));
    layer0_outputs(1953) <= not(inputs(99)) or (inputs(165));
    layer0_outputs(1954) <= (inputs(114)) or (inputs(116));
    layer0_outputs(1955) <= (inputs(125)) or (inputs(113));
    layer0_outputs(1956) <= not(inputs(60));
    layer0_outputs(1957) <= (inputs(203)) and not (inputs(4));
    layer0_outputs(1958) <= not(inputs(220)) or (inputs(232));
    layer0_outputs(1959) <= not(inputs(82)) or (inputs(221));
    layer0_outputs(1960) <= not((inputs(155)) or (inputs(222)));
    layer0_outputs(1961) <= not(inputs(213)) or (inputs(206));
    layer0_outputs(1962) <= (inputs(195)) or (inputs(213));
    layer0_outputs(1963) <= (inputs(68)) and not (inputs(136));
    layer0_outputs(1964) <= not((inputs(251)) or (inputs(154)));
    layer0_outputs(1965) <= (inputs(183)) and (inputs(139));
    layer0_outputs(1966) <= not(inputs(7));
    layer0_outputs(1967) <= not(inputs(245));
    layer0_outputs(1968) <= inputs(163);
    layer0_outputs(1969) <= (inputs(64)) or (inputs(16));
    layer0_outputs(1970) <= inputs(198);
    layer0_outputs(1971) <= (inputs(56)) and not (inputs(205));
    layer0_outputs(1972) <= (inputs(171)) xor (inputs(34));
    layer0_outputs(1973) <= inputs(104);
    layer0_outputs(1974) <= inputs(21);
    layer0_outputs(1975) <= (inputs(106)) xor (inputs(140));
    layer0_outputs(1976) <= not(inputs(101));
    layer0_outputs(1977) <= not(inputs(56)) or (inputs(136));
    layer0_outputs(1978) <= inputs(216);
    layer0_outputs(1979) <= (inputs(102)) or (inputs(247));
    layer0_outputs(1980) <= not(inputs(19));
    layer0_outputs(1981) <= not((inputs(212)) xor (inputs(190)));
    layer0_outputs(1982) <= inputs(95);
    layer0_outputs(1983) <= (inputs(226)) and not (inputs(126));
    layer0_outputs(1984) <= (inputs(110)) xor (inputs(36));
    layer0_outputs(1985) <= not(inputs(65));
    layer0_outputs(1986) <= (inputs(149)) and (inputs(194));
    layer0_outputs(1987) <= not(inputs(205)) or (inputs(112));
    layer0_outputs(1988) <= (inputs(83)) and not (inputs(123));
    layer0_outputs(1989) <= (inputs(130)) and not (inputs(210));
    layer0_outputs(1990) <= (inputs(85)) and (inputs(27));
    layer0_outputs(1991) <= inputs(94);
    layer0_outputs(1992) <= not((inputs(37)) or (inputs(13)));
    layer0_outputs(1993) <= not((inputs(1)) or (inputs(20)));
    layer0_outputs(1994) <= inputs(36);
    layer0_outputs(1995) <= inputs(23);
    layer0_outputs(1996) <= inputs(227);
    layer0_outputs(1997) <= inputs(68);
    layer0_outputs(1998) <= not(inputs(208));
    layer0_outputs(1999) <= not((inputs(54)) or (inputs(239)));
    layer0_outputs(2000) <= not(inputs(51));
    layer0_outputs(2001) <= inputs(70);
    layer0_outputs(2002) <= inputs(24);
    layer0_outputs(2003) <= (inputs(232)) and (inputs(25));
    layer0_outputs(2004) <= inputs(231);
    layer0_outputs(2005) <= not((inputs(104)) or (inputs(88)));
    layer0_outputs(2006) <= not((inputs(182)) and (inputs(191)));
    layer0_outputs(2007) <= '1';
    layer0_outputs(2008) <= not(inputs(105)) or (inputs(198));
    layer0_outputs(2009) <= inputs(177);
    layer0_outputs(2010) <= not((inputs(181)) or (inputs(214)));
    layer0_outputs(2011) <= not(inputs(178));
    layer0_outputs(2012) <= not(inputs(19)) or (inputs(128));
    layer0_outputs(2013) <= '1';
    layer0_outputs(2014) <= (inputs(92)) or (inputs(152));
    layer0_outputs(2015) <= not(inputs(216)) or (inputs(0));
    layer0_outputs(2016) <= not(inputs(107)) or (inputs(183));
    layer0_outputs(2017) <= not(inputs(203));
    layer0_outputs(2018) <= inputs(96);
    layer0_outputs(2019) <= not(inputs(102)) or (inputs(43));
    layer0_outputs(2020) <= not((inputs(228)) xor (inputs(198)));
    layer0_outputs(2021) <= (inputs(92)) and not (inputs(166));
    layer0_outputs(2022) <= not(inputs(143));
    layer0_outputs(2023) <= inputs(97);
    layer0_outputs(2024) <= inputs(9);
    layer0_outputs(2025) <= '1';
    layer0_outputs(2026) <= (inputs(206)) xor (inputs(123));
    layer0_outputs(2027) <= inputs(195);
    layer0_outputs(2028) <= not(inputs(91));
    layer0_outputs(2029) <= not(inputs(25));
    layer0_outputs(2030) <= not(inputs(187));
    layer0_outputs(2031) <= (inputs(228)) and (inputs(83));
    layer0_outputs(2032) <= (inputs(103)) xor (inputs(146));
    layer0_outputs(2033) <= (inputs(244)) and not (inputs(76));
    layer0_outputs(2034) <= not((inputs(192)) or (inputs(220)));
    layer0_outputs(2035) <= (inputs(137)) or (inputs(44));
    layer0_outputs(2036) <= not((inputs(81)) xor (inputs(71)));
    layer0_outputs(2037) <= not((inputs(31)) or (inputs(38)));
    layer0_outputs(2038) <= not((inputs(251)) and (inputs(142)));
    layer0_outputs(2039) <= (inputs(130)) or (inputs(201));
    layer0_outputs(2040) <= not((inputs(3)) and (inputs(226)));
    layer0_outputs(2041) <= not(inputs(74));
    layer0_outputs(2042) <= not(inputs(193)) or (inputs(108));
    layer0_outputs(2043) <= not((inputs(155)) or (inputs(57)));
    layer0_outputs(2044) <= (inputs(70)) or (inputs(37));
    layer0_outputs(2045) <= (inputs(90)) and (inputs(37));
    layer0_outputs(2046) <= not(inputs(147));
    layer0_outputs(2047) <= not(inputs(146));
    layer0_outputs(2048) <= not((inputs(34)) or (inputs(214)));
    layer0_outputs(2049) <= inputs(38);
    layer0_outputs(2050) <= not(inputs(197));
    layer0_outputs(2051) <= (inputs(194)) xor (inputs(8));
    layer0_outputs(2052) <= not(inputs(100));
    layer0_outputs(2053) <= inputs(53);
    layer0_outputs(2054) <= not(inputs(25)) or (inputs(115));
    layer0_outputs(2055) <= (inputs(7)) and not (inputs(129));
    layer0_outputs(2056) <= not((inputs(222)) or (inputs(43)));
    layer0_outputs(2057) <= not(inputs(107)) or (inputs(57));
    layer0_outputs(2058) <= inputs(166);
    layer0_outputs(2059) <= (inputs(15)) or (inputs(70));
    layer0_outputs(2060) <= not((inputs(185)) or (inputs(172)));
    layer0_outputs(2061) <= (inputs(136)) and not (inputs(203));
    layer0_outputs(2062) <= not(inputs(154));
    layer0_outputs(2063) <= not(inputs(215));
    layer0_outputs(2064) <= not((inputs(39)) or (inputs(38)));
    layer0_outputs(2065) <= (inputs(30)) or (inputs(36));
    layer0_outputs(2066) <= not(inputs(22));
    layer0_outputs(2067) <= not(inputs(211));
    layer0_outputs(2068) <= not((inputs(86)) or (inputs(67)));
    layer0_outputs(2069) <= inputs(210);
    layer0_outputs(2070) <= not((inputs(240)) or (inputs(65)));
    layer0_outputs(2071) <= (inputs(80)) and not (inputs(45));
    layer0_outputs(2072) <= not((inputs(229)) and (inputs(92)));
    layer0_outputs(2073) <= not(inputs(231));
    layer0_outputs(2074) <= not((inputs(222)) or (inputs(173)));
    layer0_outputs(2075) <= (inputs(47)) or (inputs(95));
    layer0_outputs(2076) <= not(inputs(129));
    layer0_outputs(2077) <= not(inputs(10));
    layer0_outputs(2078) <= not((inputs(35)) or (inputs(176)));
    layer0_outputs(2079) <= '1';
    layer0_outputs(2080) <= (inputs(236)) and not (inputs(75));
    layer0_outputs(2081) <= not((inputs(148)) and (inputs(110)));
    layer0_outputs(2082) <= (inputs(30)) xor (inputs(223));
    layer0_outputs(2083) <= not(inputs(230));
    layer0_outputs(2084) <= not((inputs(103)) or (inputs(176)));
    layer0_outputs(2085) <= (inputs(16)) xor (inputs(16));
    layer0_outputs(2086) <= not((inputs(50)) xor (inputs(22)));
    layer0_outputs(2087) <= not(inputs(202)) or (inputs(124));
    layer0_outputs(2088) <= not(inputs(233));
    layer0_outputs(2089) <= (inputs(59)) and (inputs(191));
    layer0_outputs(2090) <= (inputs(25)) and not (inputs(210));
    layer0_outputs(2091) <= not(inputs(91)) or (inputs(161));
    layer0_outputs(2092) <= not((inputs(61)) or (inputs(223)));
    layer0_outputs(2093) <= not(inputs(40));
    layer0_outputs(2094) <= (inputs(37)) xor (inputs(242));
    layer0_outputs(2095) <= (inputs(178)) or (inputs(91));
    layer0_outputs(2096) <= inputs(79);
    layer0_outputs(2097) <= (inputs(200)) and (inputs(123));
    layer0_outputs(2098) <= (inputs(248)) or (inputs(172));
    layer0_outputs(2099) <= inputs(178);
    layer0_outputs(2100) <= not(inputs(18));
    layer0_outputs(2101) <= (inputs(36)) or (inputs(187));
    layer0_outputs(2102) <= (inputs(66)) and not (inputs(254));
    layer0_outputs(2103) <= inputs(114);
    layer0_outputs(2104) <= (inputs(157)) and not (inputs(108));
    layer0_outputs(2105) <= not((inputs(237)) xor (inputs(25)));
    layer0_outputs(2106) <= inputs(236);
    layer0_outputs(2107) <= not(inputs(79));
    layer0_outputs(2108) <= '1';
    layer0_outputs(2109) <= inputs(203);
    layer0_outputs(2110) <= not((inputs(196)) xor (inputs(228)));
    layer0_outputs(2111) <= not(inputs(82));
    layer0_outputs(2112) <= (inputs(204)) or (inputs(195));
    layer0_outputs(2113) <= not((inputs(145)) or (inputs(150)));
    layer0_outputs(2114) <= not((inputs(137)) xor (inputs(205)));
    layer0_outputs(2115) <= (inputs(20)) or (inputs(27));
    layer0_outputs(2116) <= (inputs(71)) xor (inputs(40));
    layer0_outputs(2117) <= inputs(156);
    layer0_outputs(2118) <= inputs(234);
    layer0_outputs(2119) <= (inputs(10)) and not (inputs(64));
    layer0_outputs(2120) <= not((inputs(246)) or (inputs(225)));
    layer0_outputs(2121) <= inputs(55);
    layer0_outputs(2122) <= not((inputs(201)) xor (inputs(127)));
    layer0_outputs(2123) <= not(inputs(4)) or (inputs(28));
    layer0_outputs(2124) <= not((inputs(54)) or (inputs(222)));
    layer0_outputs(2125) <= not((inputs(64)) or (inputs(20)));
    layer0_outputs(2126) <= (inputs(72)) and (inputs(33));
    layer0_outputs(2127) <= (inputs(95)) and not (inputs(214));
    layer0_outputs(2128) <= not(inputs(230)) or (inputs(0));
    layer0_outputs(2129) <= (inputs(142)) or (inputs(174));
    layer0_outputs(2130) <= (inputs(252)) xor (inputs(171));
    layer0_outputs(2131) <= not((inputs(197)) or (inputs(116)));
    layer0_outputs(2132) <= inputs(213);
    layer0_outputs(2133) <= (inputs(143)) and not (inputs(50));
    layer0_outputs(2134) <= (inputs(187)) or (inputs(157));
    layer0_outputs(2135) <= (inputs(88)) and not (inputs(118));
    layer0_outputs(2136) <= not(inputs(243));
    layer0_outputs(2137) <= not(inputs(234));
    layer0_outputs(2138) <= not(inputs(37));
    layer0_outputs(2139) <= inputs(117);
    layer0_outputs(2140) <= not((inputs(17)) or (inputs(123)));
    layer0_outputs(2141) <= (inputs(98)) xor (inputs(170));
    layer0_outputs(2142) <= (inputs(58)) or (inputs(62));
    layer0_outputs(2143) <= not(inputs(55)) or (inputs(28));
    layer0_outputs(2144) <= not((inputs(111)) or (inputs(156)));
    layer0_outputs(2145) <= (inputs(44)) xor (inputs(88));
    layer0_outputs(2146) <= not(inputs(77));
    layer0_outputs(2147) <= (inputs(134)) or (inputs(207));
    layer0_outputs(2148) <= not(inputs(69));
    layer0_outputs(2149) <= '0';
    layer0_outputs(2150) <= not(inputs(252));
    layer0_outputs(2151) <= not(inputs(109)) or (inputs(42));
    layer0_outputs(2152) <= not(inputs(29));
    layer0_outputs(2153) <= inputs(114);
    layer0_outputs(2154) <= (inputs(69)) and not (inputs(226));
    layer0_outputs(2155) <= (inputs(177)) and not (inputs(142));
    layer0_outputs(2156) <= not(inputs(194)) or (inputs(45));
    layer0_outputs(2157) <= not(inputs(67));
    layer0_outputs(2158) <= not((inputs(64)) xor (inputs(121)));
    layer0_outputs(2159) <= not(inputs(22));
    layer0_outputs(2160) <= '0';
    layer0_outputs(2161) <= '0';
    layer0_outputs(2162) <= (inputs(105)) and not (inputs(42));
    layer0_outputs(2163) <= inputs(78);
    layer0_outputs(2164) <= (inputs(175)) and not (inputs(55));
    layer0_outputs(2165) <= (inputs(188)) or (inputs(144));
    layer0_outputs(2166) <= not((inputs(249)) and (inputs(57)));
    layer0_outputs(2167) <= not(inputs(74));
    layer0_outputs(2168) <= (inputs(13)) or (inputs(179));
    layer0_outputs(2169) <= '0';
    layer0_outputs(2170) <= (inputs(57)) xor (inputs(22));
    layer0_outputs(2171) <= (inputs(253)) or (inputs(189));
    layer0_outputs(2172) <= not(inputs(18)) or (inputs(74));
    layer0_outputs(2173) <= not((inputs(16)) or (inputs(60)));
    layer0_outputs(2174) <= not((inputs(253)) and (inputs(136)));
    layer0_outputs(2175) <= (inputs(116)) xor (inputs(249));
    layer0_outputs(2176) <= (inputs(171)) or (inputs(145));
    layer0_outputs(2177) <= not(inputs(7)) or (inputs(12));
    layer0_outputs(2178) <= (inputs(181)) xor (inputs(242));
    layer0_outputs(2179) <= inputs(59);
    layer0_outputs(2180) <= (inputs(59)) or (inputs(19));
    layer0_outputs(2181) <= (inputs(179)) xor (inputs(160));
    layer0_outputs(2182) <= not(inputs(98));
    layer0_outputs(2183) <= (inputs(227)) xor (inputs(211));
    layer0_outputs(2184) <= (inputs(133)) or (inputs(253));
    layer0_outputs(2185) <= not(inputs(23)) or (inputs(116));
    layer0_outputs(2186) <= '1';
    layer0_outputs(2187) <= not(inputs(214)) or (inputs(125));
    layer0_outputs(2188) <= not((inputs(37)) or (inputs(194)));
    layer0_outputs(2189) <= not((inputs(135)) or (inputs(35)));
    layer0_outputs(2190) <= not(inputs(102));
    layer0_outputs(2191) <= not(inputs(1)) or (inputs(154));
    layer0_outputs(2192) <= not((inputs(78)) or (inputs(151)));
    layer0_outputs(2193) <= not(inputs(210));
    layer0_outputs(2194) <= not(inputs(87)) or (inputs(185));
    layer0_outputs(2195) <= (inputs(62)) and not (inputs(224));
    layer0_outputs(2196) <= not((inputs(84)) or (inputs(180)));
    layer0_outputs(2197) <= not(inputs(130)) or (inputs(73));
    layer0_outputs(2198) <= (inputs(141)) or (inputs(131));
    layer0_outputs(2199) <= (inputs(250)) xor (inputs(53));
    layer0_outputs(2200) <= not((inputs(156)) xor (inputs(65)));
    layer0_outputs(2201) <= not((inputs(199)) and (inputs(102)));
    layer0_outputs(2202) <= not((inputs(165)) or (inputs(208)));
    layer0_outputs(2203) <= inputs(159);
    layer0_outputs(2204) <= (inputs(244)) and not (inputs(97));
    layer0_outputs(2205) <= not((inputs(126)) xor (inputs(6)));
    layer0_outputs(2206) <= not(inputs(40)) or (inputs(45));
    layer0_outputs(2207) <= not(inputs(125));
    layer0_outputs(2208) <= not(inputs(139)) or (inputs(199));
    layer0_outputs(2209) <= not(inputs(70)) or (inputs(253));
    layer0_outputs(2210) <= (inputs(56)) and not (inputs(209));
    layer0_outputs(2211) <= inputs(76);
    layer0_outputs(2212) <= not((inputs(13)) or (inputs(131)));
    layer0_outputs(2213) <= (inputs(116)) or (inputs(36));
    layer0_outputs(2214) <= not((inputs(87)) and (inputs(235)));
    layer0_outputs(2215) <= not((inputs(90)) xor (inputs(3)));
    layer0_outputs(2216) <= not(inputs(59));
    layer0_outputs(2217) <= not(inputs(209));
    layer0_outputs(2218) <= not(inputs(46));
    layer0_outputs(2219) <= (inputs(114)) or (inputs(112));
    layer0_outputs(2220) <= (inputs(237)) or (inputs(208));
    layer0_outputs(2221) <= not(inputs(102)) or (inputs(170));
    layer0_outputs(2222) <= not((inputs(82)) or (inputs(133)));
    layer0_outputs(2223) <= '0';
    layer0_outputs(2224) <= not((inputs(242)) and (inputs(15)));
    layer0_outputs(2225) <= not(inputs(133));
    layer0_outputs(2226) <= (inputs(85)) and not (inputs(189));
    layer0_outputs(2227) <= inputs(224);
    layer0_outputs(2228) <= not(inputs(86));
    layer0_outputs(2229) <= (inputs(226)) and not (inputs(237));
    layer0_outputs(2230) <= (inputs(9)) and (inputs(117));
    layer0_outputs(2231) <= (inputs(185)) or (inputs(79));
    layer0_outputs(2232) <= not(inputs(115)) or (inputs(123));
    layer0_outputs(2233) <= not(inputs(244));
    layer0_outputs(2234) <= inputs(91);
    layer0_outputs(2235) <= not(inputs(183)) or (inputs(67));
    layer0_outputs(2236) <= (inputs(141)) and (inputs(57));
    layer0_outputs(2237) <= inputs(40);
    layer0_outputs(2238) <= (inputs(12)) or (inputs(68));
    layer0_outputs(2239) <= inputs(107);
    layer0_outputs(2240) <= (inputs(117)) and not (inputs(125));
    layer0_outputs(2241) <= '0';
    layer0_outputs(2242) <= (inputs(129)) and (inputs(201));
    layer0_outputs(2243) <= inputs(83);
    layer0_outputs(2244) <= not(inputs(109));
    layer0_outputs(2245) <= inputs(93);
    layer0_outputs(2246) <= not(inputs(99));
    layer0_outputs(2247) <= (inputs(166)) xor (inputs(212));
    layer0_outputs(2248) <= (inputs(201)) xor (inputs(144));
    layer0_outputs(2249) <= not(inputs(178));
    layer0_outputs(2250) <= not(inputs(100));
    layer0_outputs(2251) <= inputs(173);
    layer0_outputs(2252) <= '1';
    layer0_outputs(2253) <= not(inputs(148));
    layer0_outputs(2254) <= (inputs(41)) and (inputs(219));
    layer0_outputs(2255) <= not(inputs(26)) or (inputs(178));
    layer0_outputs(2256) <= (inputs(204)) and not (inputs(245));
    layer0_outputs(2257) <= not((inputs(95)) xor (inputs(247)));
    layer0_outputs(2258) <= not(inputs(104));
    layer0_outputs(2259) <= not(inputs(212)) or (inputs(137));
    layer0_outputs(2260) <= not((inputs(101)) or (inputs(103)));
    layer0_outputs(2261) <= '0';
    layer0_outputs(2262) <= inputs(200);
    layer0_outputs(2263) <= not(inputs(94));
    layer0_outputs(2264) <= (inputs(102)) and not (inputs(175));
    layer0_outputs(2265) <= not(inputs(149)) or (inputs(240));
    layer0_outputs(2266) <= (inputs(92)) xor (inputs(28));
    layer0_outputs(2267) <= not((inputs(234)) xor (inputs(11)));
    layer0_outputs(2268) <= not((inputs(150)) or (inputs(106)));
    layer0_outputs(2269) <= inputs(162);
    layer0_outputs(2270) <= not(inputs(204)) or (inputs(14));
    layer0_outputs(2271) <= (inputs(98)) or (inputs(81));
    layer0_outputs(2272) <= (inputs(106)) or (inputs(48));
    layer0_outputs(2273) <= not(inputs(103));
    layer0_outputs(2274) <= (inputs(107)) and not (inputs(84));
    layer0_outputs(2275) <= (inputs(51)) xor (inputs(72));
    layer0_outputs(2276) <= not(inputs(82));
    layer0_outputs(2277) <= (inputs(75)) and (inputs(25));
    layer0_outputs(2278) <= not(inputs(209)) or (inputs(140));
    layer0_outputs(2279) <= (inputs(102)) and not (inputs(0));
    layer0_outputs(2280) <= inputs(169);
    layer0_outputs(2281) <= '0';
    layer0_outputs(2282) <= not(inputs(114));
    layer0_outputs(2283) <= not((inputs(237)) and (inputs(6)));
    layer0_outputs(2284) <= inputs(102);
    layer0_outputs(2285) <= (inputs(167)) and (inputs(251));
    layer0_outputs(2286) <= not(inputs(228));
    layer0_outputs(2287) <= (inputs(8)) and not (inputs(45));
    layer0_outputs(2288) <= (inputs(59)) or (inputs(211));
    layer0_outputs(2289) <= not(inputs(73)) or (inputs(13));
    layer0_outputs(2290) <= not((inputs(197)) xor (inputs(46)));
    layer0_outputs(2291) <= not((inputs(94)) or (inputs(26)));
    layer0_outputs(2292) <= not(inputs(35));
    layer0_outputs(2293) <= '1';
    layer0_outputs(2294) <= not((inputs(168)) or (inputs(164)));
    layer0_outputs(2295) <= not((inputs(144)) or (inputs(214)));
    layer0_outputs(2296) <= inputs(113);
    layer0_outputs(2297) <= not((inputs(113)) or (inputs(157)));
    layer0_outputs(2298) <= inputs(184);
    layer0_outputs(2299) <= (inputs(131)) and (inputs(142));
    layer0_outputs(2300) <= inputs(235);
    layer0_outputs(2301) <= not((inputs(10)) and (inputs(214)));
    layer0_outputs(2302) <= (inputs(77)) and not (inputs(106));
    layer0_outputs(2303) <= (inputs(21)) or (inputs(89));
    layer0_outputs(2304) <= (inputs(252)) xor (inputs(75));
    layer0_outputs(2305) <= inputs(46);
    layer0_outputs(2306) <= (inputs(195)) and not (inputs(47));
    layer0_outputs(2307) <= not(inputs(55));
    layer0_outputs(2308) <= not(inputs(166)) or (inputs(97));
    layer0_outputs(2309) <= not((inputs(247)) xor (inputs(46)));
    layer0_outputs(2310) <= not(inputs(99)) or (inputs(72));
    layer0_outputs(2311) <= (inputs(59)) and (inputs(99));
    layer0_outputs(2312) <= not((inputs(97)) xor (inputs(6)));
    layer0_outputs(2313) <= not((inputs(204)) and (inputs(182)));
    layer0_outputs(2314) <= inputs(153);
    layer0_outputs(2315) <= inputs(106);
    layer0_outputs(2316) <= '0';
    layer0_outputs(2317) <= not(inputs(181));
    layer0_outputs(2318) <= not((inputs(244)) or (inputs(254)));
    layer0_outputs(2319) <= (inputs(239)) and (inputs(240));
    layer0_outputs(2320) <= not((inputs(56)) or (inputs(241)));
    layer0_outputs(2321) <= not((inputs(127)) and (inputs(166)));
    layer0_outputs(2322) <= not(inputs(21)) or (inputs(254));
    layer0_outputs(2323) <= not((inputs(143)) and (inputs(160)));
    layer0_outputs(2324) <= (inputs(60)) or (inputs(111));
    layer0_outputs(2325) <= (inputs(170)) or (inputs(53));
    layer0_outputs(2326) <= (inputs(17)) or (inputs(65));
    layer0_outputs(2327) <= (inputs(90)) or (inputs(226));
    layer0_outputs(2328) <= inputs(245);
    layer0_outputs(2329) <= inputs(39);
    layer0_outputs(2330) <= not(inputs(80)) or (inputs(252));
    layer0_outputs(2331) <= inputs(46);
    layer0_outputs(2332) <= not(inputs(53)) or (inputs(229));
    layer0_outputs(2333) <= (inputs(32)) xor (inputs(206));
    layer0_outputs(2334) <= not(inputs(119)) or (inputs(111));
    layer0_outputs(2335) <= '1';
    layer0_outputs(2336) <= not((inputs(235)) or (inputs(66)));
    layer0_outputs(2337) <= (inputs(11)) and not (inputs(34));
    layer0_outputs(2338) <= not(inputs(232));
    layer0_outputs(2339) <= not((inputs(28)) or (inputs(134)));
    layer0_outputs(2340) <= (inputs(180)) or (inputs(195));
    layer0_outputs(2341) <= not(inputs(86)) or (inputs(154));
    layer0_outputs(2342) <= (inputs(121)) or (inputs(115));
    layer0_outputs(2343) <= not(inputs(108));
    layer0_outputs(2344) <= not(inputs(136)) or (inputs(146));
    layer0_outputs(2345) <= inputs(148);
    layer0_outputs(2346) <= (inputs(186)) xor (inputs(17));
    layer0_outputs(2347) <= (inputs(135)) or (inputs(223));
    layer0_outputs(2348) <= (inputs(91)) and not (inputs(141));
    layer0_outputs(2349) <= (inputs(205)) and not (inputs(159));
    layer0_outputs(2350) <= (inputs(122)) and not (inputs(160));
    layer0_outputs(2351) <= inputs(34);
    layer0_outputs(2352) <= not((inputs(190)) or (inputs(120)));
    layer0_outputs(2353) <= (inputs(221)) and not (inputs(128));
    layer0_outputs(2354) <= not((inputs(178)) and (inputs(146)));
    layer0_outputs(2355) <= '1';
    layer0_outputs(2356) <= not(inputs(172)) or (inputs(15));
    layer0_outputs(2357) <= inputs(147);
    layer0_outputs(2358) <= inputs(60);
    layer0_outputs(2359) <= not(inputs(173)) or (inputs(138));
    layer0_outputs(2360) <= '0';
    layer0_outputs(2361) <= not((inputs(78)) or (inputs(85)));
    layer0_outputs(2362) <= inputs(40);
    layer0_outputs(2363) <= '1';
    layer0_outputs(2364) <= not(inputs(22));
    layer0_outputs(2365) <= not((inputs(97)) xor (inputs(132)));
    layer0_outputs(2366) <= not(inputs(91));
    layer0_outputs(2367) <= not(inputs(194));
    layer0_outputs(2368) <= inputs(141);
    layer0_outputs(2369) <= not((inputs(48)) xor (inputs(223)));
    layer0_outputs(2370) <= (inputs(240)) and (inputs(36));
    layer0_outputs(2371) <= not((inputs(125)) xor (inputs(174)));
    layer0_outputs(2372) <= not((inputs(99)) and (inputs(66)));
    layer0_outputs(2373) <= (inputs(135)) xor (inputs(181));
    layer0_outputs(2374) <= not((inputs(178)) or (inputs(179)));
    layer0_outputs(2375) <= (inputs(187)) xor (inputs(157));
    layer0_outputs(2376) <= (inputs(4)) and (inputs(191));
    layer0_outputs(2377) <= (inputs(179)) xor (inputs(88));
    layer0_outputs(2378) <= not(inputs(205));
    layer0_outputs(2379) <= not((inputs(108)) or (inputs(190)));
    layer0_outputs(2380) <= not((inputs(34)) xor (inputs(179)));
    layer0_outputs(2381) <= (inputs(95)) or (inputs(233));
    layer0_outputs(2382) <= (inputs(98)) and not (inputs(43));
    layer0_outputs(2383) <= not((inputs(220)) and (inputs(199)));
    layer0_outputs(2384) <= not((inputs(86)) or (inputs(161)));
    layer0_outputs(2385) <= inputs(134);
    layer0_outputs(2386) <= '1';
    layer0_outputs(2387) <= not(inputs(179));
    layer0_outputs(2388) <= (inputs(185)) or (inputs(177));
    layer0_outputs(2389) <= not((inputs(242)) or (inputs(179)));
    layer0_outputs(2390) <= not((inputs(164)) xor (inputs(181)));
    layer0_outputs(2391) <= (inputs(141)) xor (inputs(205));
    layer0_outputs(2392) <= not(inputs(24)) or (inputs(222));
    layer0_outputs(2393) <= not((inputs(160)) or (inputs(141)));
    layer0_outputs(2394) <= not(inputs(84));
    layer0_outputs(2395) <= (inputs(200)) or (inputs(224));
    layer0_outputs(2396) <= not((inputs(92)) xor (inputs(74)));
    layer0_outputs(2397) <= '1';
    layer0_outputs(2398) <= (inputs(188)) or (inputs(246));
    layer0_outputs(2399) <= (inputs(192)) and not (inputs(152));
    layer0_outputs(2400) <= (inputs(120)) and not (inputs(233));
    layer0_outputs(2401) <= not((inputs(175)) xor (inputs(222)));
    layer0_outputs(2402) <= (inputs(159)) and not (inputs(149));
    layer0_outputs(2403) <= (inputs(225)) and not (inputs(253));
    layer0_outputs(2404) <= inputs(127);
    layer0_outputs(2405) <= (inputs(251)) or (inputs(80));
    layer0_outputs(2406) <= inputs(176);
    layer0_outputs(2407) <= (inputs(152)) and not (inputs(175));
    layer0_outputs(2408) <= not(inputs(161));
    layer0_outputs(2409) <= not(inputs(55)) or (inputs(0));
    layer0_outputs(2410) <= (inputs(36)) and not (inputs(47));
    layer0_outputs(2411) <= not(inputs(99)) or (inputs(1));
    layer0_outputs(2412) <= not(inputs(83));
    layer0_outputs(2413) <= (inputs(41)) and (inputs(6));
    layer0_outputs(2414) <= not((inputs(179)) xor (inputs(160)));
    layer0_outputs(2415) <= not(inputs(88));
    layer0_outputs(2416) <= not((inputs(199)) or (inputs(132)));
    layer0_outputs(2417) <= not(inputs(109));
    layer0_outputs(2418) <= inputs(163);
    layer0_outputs(2419) <= inputs(92);
    layer0_outputs(2420) <= (inputs(198)) xor (inputs(194));
    layer0_outputs(2421) <= (inputs(186)) and (inputs(130));
    layer0_outputs(2422) <= not(inputs(117));
    layer0_outputs(2423) <= (inputs(39)) or (inputs(193));
    layer0_outputs(2424) <= not((inputs(92)) xor (inputs(33)));
    layer0_outputs(2425) <= not((inputs(105)) or (inputs(47)));
    layer0_outputs(2426) <= not(inputs(13));
    layer0_outputs(2427) <= inputs(243);
    layer0_outputs(2428) <= '1';
    layer0_outputs(2429) <= not((inputs(158)) or (inputs(245)));
    layer0_outputs(2430) <= inputs(120);
    layer0_outputs(2431) <= inputs(14);
    layer0_outputs(2432) <= inputs(9);
    layer0_outputs(2433) <= inputs(171);
    layer0_outputs(2434) <= (inputs(224)) or (inputs(44));
    layer0_outputs(2435) <= (inputs(9)) and not (inputs(98));
    layer0_outputs(2436) <= inputs(137);
    layer0_outputs(2437) <= not(inputs(159)) or (inputs(148));
    layer0_outputs(2438) <= not((inputs(164)) or (inputs(115)));
    layer0_outputs(2439) <= not(inputs(214)) or (inputs(153));
    layer0_outputs(2440) <= not(inputs(23));
    layer0_outputs(2441) <= '1';
    layer0_outputs(2442) <= (inputs(20)) and not (inputs(223));
    layer0_outputs(2443) <= (inputs(57)) and (inputs(222));
    layer0_outputs(2444) <= not(inputs(135));
    layer0_outputs(2445) <= not(inputs(38)) or (inputs(33));
    layer0_outputs(2446) <= not(inputs(209)) or (inputs(136));
    layer0_outputs(2447) <= not((inputs(34)) or (inputs(11)));
    layer0_outputs(2448) <= not((inputs(121)) or (inputs(51)));
    layer0_outputs(2449) <= '0';
    layer0_outputs(2450) <= not(inputs(186)) or (inputs(122));
    layer0_outputs(2451) <= not(inputs(130));
    layer0_outputs(2452) <= not(inputs(92)) or (inputs(30));
    layer0_outputs(2453) <= not(inputs(48)) or (inputs(150));
    layer0_outputs(2454) <= not(inputs(179)) or (inputs(201));
    layer0_outputs(2455) <= (inputs(19)) and not (inputs(162));
    layer0_outputs(2456) <= not(inputs(143));
    layer0_outputs(2457) <= (inputs(236)) xor (inputs(113));
    layer0_outputs(2458) <= '0';
    layer0_outputs(2459) <= not(inputs(84));
    layer0_outputs(2460) <= (inputs(200)) and not (inputs(137));
    layer0_outputs(2461) <= not((inputs(109)) or (inputs(156)));
    layer0_outputs(2462) <= not((inputs(149)) or (inputs(115)));
    layer0_outputs(2463) <= not((inputs(36)) or (inputs(228)));
    layer0_outputs(2464) <= not(inputs(45));
    layer0_outputs(2465) <= not(inputs(251)) or (inputs(214));
    layer0_outputs(2466) <= not(inputs(77));
    layer0_outputs(2467) <= not(inputs(193));
    layer0_outputs(2468) <= (inputs(251)) or (inputs(135));
    layer0_outputs(2469) <= (inputs(218)) and not (inputs(12));
    layer0_outputs(2470) <= not(inputs(123));
    layer0_outputs(2471) <= (inputs(57)) xor (inputs(72));
    layer0_outputs(2472) <= not((inputs(77)) xor (inputs(79)));
    layer0_outputs(2473) <= '1';
    layer0_outputs(2474) <= (inputs(110)) or (inputs(57));
    layer0_outputs(2475) <= inputs(152);
    layer0_outputs(2476) <= not(inputs(227));
    layer0_outputs(2477) <= inputs(52);
    layer0_outputs(2478) <= (inputs(254)) and not (inputs(71));
    layer0_outputs(2479) <= not(inputs(21));
    layer0_outputs(2480) <= not((inputs(92)) or (inputs(18)));
    layer0_outputs(2481) <= not(inputs(230)) or (inputs(25));
    layer0_outputs(2482) <= inputs(25);
    layer0_outputs(2483) <= (inputs(241)) and not (inputs(114));
    layer0_outputs(2484) <= not((inputs(115)) or (inputs(69)));
    layer0_outputs(2485) <= (inputs(51)) and (inputs(101));
    layer0_outputs(2486) <= not(inputs(121));
    layer0_outputs(2487) <= (inputs(209)) or (inputs(9));
    layer0_outputs(2488) <= (inputs(155)) and not (inputs(71));
    layer0_outputs(2489) <= not((inputs(29)) xor (inputs(219)));
    layer0_outputs(2490) <= (inputs(192)) or (inputs(99));
    layer0_outputs(2491) <= not(inputs(110)) or (inputs(104));
    layer0_outputs(2492) <= (inputs(53)) and not (inputs(222));
    layer0_outputs(2493) <= not((inputs(211)) and (inputs(172)));
    layer0_outputs(2494) <= not((inputs(117)) xor (inputs(237)));
    layer0_outputs(2495) <= (inputs(51)) xor (inputs(109));
    layer0_outputs(2496) <= (inputs(75)) xor (inputs(78));
    layer0_outputs(2497) <= not((inputs(10)) xor (inputs(160)));
    layer0_outputs(2498) <= not(inputs(23)) or (inputs(249));
    layer0_outputs(2499) <= not((inputs(179)) or (inputs(46)));
    layer0_outputs(2500) <= (inputs(11)) or (inputs(59));
    layer0_outputs(2501) <= inputs(241);
    layer0_outputs(2502) <= '0';
    layer0_outputs(2503) <= (inputs(224)) xor (inputs(5));
    layer0_outputs(2504) <= (inputs(60)) or (inputs(176));
    layer0_outputs(2505) <= (inputs(51)) or (inputs(96));
    layer0_outputs(2506) <= (inputs(89)) or (inputs(126));
    layer0_outputs(2507) <= not((inputs(90)) and (inputs(19)));
    layer0_outputs(2508) <= inputs(7);
    layer0_outputs(2509) <= (inputs(115)) xor (inputs(5));
    layer0_outputs(2510) <= (inputs(28)) or (inputs(39));
    layer0_outputs(2511) <= (inputs(171)) or (inputs(14));
    layer0_outputs(2512) <= inputs(91);
    layer0_outputs(2513) <= (inputs(3)) xor (inputs(109));
    layer0_outputs(2514) <= (inputs(107)) and not (inputs(193));
    layer0_outputs(2515) <= (inputs(209)) and not (inputs(233));
    layer0_outputs(2516) <= (inputs(214)) and not (inputs(2));
    layer0_outputs(2517) <= (inputs(137)) and not (inputs(19));
    layer0_outputs(2518) <= not((inputs(217)) or (inputs(31)));
    layer0_outputs(2519) <= (inputs(54)) and not (inputs(255));
    layer0_outputs(2520) <= inputs(45);
    layer0_outputs(2521) <= (inputs(158)) and (inputs(103));
    layer0_outputs(2522) <= not(inputs(30));
    layer0_outputs(2523) <= not(inputs(148));
    layer0_outputs(2524) <= '1';
    layer0_outputs(2525) <= not(inputs(29));
    layer0_outputs(2526) <= (inputs(188)) and not (inputs(21));
    layer0_outputs(2527) <= not((inputs(220)) and (inputs(104)));
    layer0_outputs(2528) <= inputs(167);
    layer0_outputs(2529) <= not(inputs(18));
    layer0_outputs(2530) <= (inputs(151)) or (inputs(126));
    layer0_outputs(2531) <= (inputs(238)) and (inputs(200));
    layer0_outputs(2532) <= '0';
    layer0_outputs(2533) <= '1';
    layer0_outputs(2534) <= not(inputs(163));
    layer0_outputs(2535) <= not(inputs(135)) or (inputs(208));
    layer0_outputs(2536) <= not((inputs(167)) or (inputs(238)));
    layer0_outputs(2537) <= not((inputs(176)) xor (inputs(199)));
    layer0_outputs(2538) <= '0';
    layer0_outputs(2539) <= not((inputs(173)) xor (inputs(92)));
    layer0_outputs(2540) <= (inputs(90)) and not (inputs(218));
    layer0_outputs(2541) <= '0';
    layer0_outputs(2542) <= inputs(189);
    layer0_outputs(2543) <= (inputs(134)) xor (inputs(40));
    layer0_outputs(2544) <= inputs(205);
    layer0_outputs(2545) <= (inputs(123)) and not (inputs(83));
    layer0_outputs(2546) <= not((inputs(117)) or (inputs(162)));
    layer0_outputs(2547) <= not(inputs(38));
    layer0_outputs(2548) <= (inputs(250)) or (inputs(216));
    layer0_outputs(2549) <= not(inputs(144)) or (inputs(153));
    layer0_outputs(2550) <= (inputs(172)) xor (inputs(70));
    layer0_outputs(2551) <= inputs(25);
    layer0_outputs(2552) <= '1';
    layer0_outputs(2553) <= inputs(204);
    layer0_outputs(2554) <= not(inputs(146)) or (inputs(14));
    layer0_outputs(2555) <= not(inputs(161)) or (inputs(90));
    layer0_outputs(2556) <= not((inputs(182)) xor (inputs(0)));
    layer0_outputs(2557) <= inputs(214);
    layer0_outputs(2558) <= not((inputs(247)) or (inputs(21)));
    layer0_outputs(2559) <= not(inputs(27));
    layer0_outputs(2560) <= not(inputs(10));
    layer0_outputs(2561) <= inputs(253);
    layer0_outputs(2562) <= not((inputs(101)) and (inputs(101)));
    layer0_outputs(2563) <= not((inputs(253)) and (inputs(8)));
    layer0_outputs(2564) <= (inputs(150)) or (inputs(52));
    layer0_outputs(2565) <= not((inputs(173)) xor (inputs(79)));
    layer0_outputs(2566) <= (inputs(197)) and not (inputs(146));
    layer0_outputs(2567) <= not(inputs(135)) or (inputs(162));
    layer0_outputs(2568) <= not((inputs(102)) or (inputs(187)));
    layer0_outputs(2569) <= not((inputs(103)) or (inputs(130)));
    layer0_outputs(2570) <= not(inputs(154)) or (inputs(216));
    layer0_outputs(2571) <= not((inputs(67)) xor (inputs(51)));
    layer0_outputs(2572) <= not(inputs(20)) or (inputs(45));
    layer0_outputs(2573) <= (inputs(225)) or (inputs(41));
    layer0_outputs(2574) <= not(inputs(32)) or (inputs(149));
    layer0_outputs(2575) <= inputs(165);
    layer0_outputs(2576) <= not(inputs(136)) or (inputs(132));
    layer0_outputs(2577) <= (inputs(249)) or (inputs(177));
    layer0_outputs(2578) <= (inputs(211)) or (inputs(81));
    layer0_outputs(2579) <= not(inputs(24));
    layer0_outputs(2580) <= inputs(92);
    layer0_outputs(2581) <= not(inputs(45));
    layer0_outputs(2582) <= not((inputs(32)) or (inputs(202)));
    layer0_outputs(2583) <= inputs(162);
    layer0_outputs(2584) <= (inputs(137)) and not (inputs(28));
    layer0_outputs(2585) <= not(inputs(84));
    layer0_outputs(2586) <= '0';
    layer0_outputs(2587) <= (inputs(28)) and (inputs(51));
    layer0_outputs(2588) <= not(inputs(116));
    layer0_outputs(2589) <= not(inputs(217)) or (inputs(153));
    layer0_outputs(2590) <= not(inputs(158)) or (inputs(158));
    layer0_outputs(2591) <= (inputs(84)) and (inputs(158));
    layer0_outputs(2592) <= (inputs(106)) xor (inputs(77));
    layer0_outputs(2593) <= not((inputs(126)) and (inputs(196)));
    layer0_outputs(2594) <= inputs(22);
    layer0_outputs(2595) <= (inputs(160)) and not (inputs(5));
    layer0_outputs(2596) <= not((inputs(101)) or (inputs(162)));
    layer0_outputs(2597) <= not((inputs(205)) or (inputs(170)));
    layer0_outputs(2598) <= not(inputs(171)) or (inputs(34));
    layer0_outputs(2599) <= not(inputs(13));
    layer0_outputs(2600) <= inputs(212);
    layer0_outputs(2601) <= not((inputs(230)) xor (inputs(190)));
    layer0_outputs(2602) <= inputs(167);
    layer0_outputs(2603) <= not((inputs(190)) or (inputs(49)));
    layer0_outputs(2604) <= inputs(237);
    layer0_outputs(2605) <= not(inputs(94));
    layer0_outputs(2606) <= (inputs(195)) or (inputs(5));
    layer0_outputs(2607) <= inputs(12);
    layer0_outputs(2608) <= not(inputs(105));
    layer0_outputs(2609) <= not((inputs(10)) and (inputs(101)));
    layer0_outputs(2610) <= not((inputs(116)) and (inputs(152)));
    layer0_outputs(2611) <= (inputs(224)) and not (inputs(162));
    layer0_outputs(2612) <= (inputs(76)) and not (inputs(154));
    layer0_outputs(2613) <= (inputs(128)) and not (inputs(37));
    layer0_outputs(2614) <= not(inputs(151));
    layer0_outputs(2615) <= not(inputs(28)) or (inputs(10));
    layer0_outputs(2616) <= not(inputs(187)) or (inputs(238));
    layer0_outputs(2617) <= inputs(204);
    layer0_outputs(2618) <= not(inputs(57)) or (inputs(144));
    layer0_outputs(2619) <= not(inputs(59)) or (inputs(193));
    layer0_outputs(2620) <= not((inputs(160)) or (inputs(151)));
    layer0_outputs(2621) <= inputs(130);
    layer0_outputs(2622) <= not((inputs(214)) xor (inputs(247)));
    layer0_outputs(2623) <= inputs(141);
    layer0_outputs(2624) <= not(inputs(248)) or (inputs(64));
    layer0_outputs(2625) <= '0';
    layer0_outputs(2626) <= (inputs(72)) xor (inputs(13));
    layer0_outputs(2627) <= not(inputs(121));
    layer0_outputs(2628) <= not((inputs(106)) or (inputs(57)));
    layer0_outputs(2629) <= '1';
    layer0_outputs(2630) <= not((inputs(77)) xor (inputs(29)));
    layer0_outputs(2631) <= not(inputs(89));
    layer0_outputs(2632) <= (inputs(231)) and not (inputs(72));
    layer0_outputs(2633) <= inputs(188);
    layer0_outputs(2634) <= inputs(238);
    layer0_outputs(2635) <= not((inputs(50)) or (inputs(90)));
    layer0_outputs(2636) <= not(inputs(117)) or (inputs(93));
    layer0_outputs(2637) <= not(inputs(182));
    layer0_outputs(2638) <= inputs(70);
    layer0_outputs(2639) <= (inputs(200)) and not (inputs(97));
    layer0_outputs(2640) <= '1';
    layer0_outputs(2641) <= not((inputs(165)) or (inputs(81)));
    layer0_outputs(2642) <= not(inputs(64));
    layer0_outputs(2643) <= (inputs(188)) or (inputs(172));
    layer0_outputs(2644) <= (inputs(7)) and not (inputs(34));
    layer0_outputs(2645) <= not(inputs(35)) or (inputs(113));
    layer0_outputs(2646) <= (inputs(247)) and not (inputs(3));
    layer0_outputs(2647) <= not(inputs(133)) or (inputs(73));
    layer0_outputs(2648) <= inputs(208);
    layer0_outputs(2649) <= (inputs(229)) and not (inputs(145));
    layer0_outputs(2650) <= not((inputs(64)) and (inputs(21)));
    layer0_outputs(2651) <= inputs(216);
    layer0_outputs(2652) <= not(inputs(21));
    layer0_outputs(2653) <= '1';
    layer0_outputs(2654) <= inputs(30);
    layer0_outputs(2655) <= inputs(98);
    layer0_outputs(2656) <= not(inputs(84)) or (inputs(184));
    layer0_outputs(2657) <= (inputs(190)) and not (inputs(224));
    layer0_outputs(2658) <= not(inputs(105)) or (inputs(241));
    layer0_outputs(2659) <= not(inputs(246));
    layer0_outputs(2660) <= not(inputs(57));
    layer0_outputs(2661) <= '0';
    layer0_outputs(2662) <= (inputs(194)) or (inputs(176));
    layer0_outputs(2663) <= (inputs(32)) xor (inputs(90));
    layer0_outputs(2664) <= (inputs(71)) and (inputs(255));
    layer0_outputs(2665) <= not(inputs(180)) or (inputs(50));
    layer0_outputs(2666) <= (inputs(132)) xor (inputs(247));
    layer0_outputs(2667) <= not((inputs(191)) xor (inputs(110)));
    layer0_outputs(2668) <= not(inputs(157)) or (inputs(80));
    layer0_outputs(2669) <= not((inputs(131)) or (inputs(107)));
    layer0_outputs(2670) <= not(inputs(8));
    layer0_outputs(2671) <= not(inputs(67));
    layer0_outputs(2672) <= not((inputs(220)) xor (inputs(75)));
    layer0_outputs(2673) <= inputs(168);
    layer0_outputs(2674) <= not(inputs(246)) or (inputs(44));
    layer0_outputs(2675) <= (inputs(159)) and not (inputs(148));
    layer0_outputs(2676) <= (inputs(77)) and not (inputs(134));
    layer0_outputs(2677) <= inputs(87);
    layer0_outputs(2678) <= inputs(27);
    layer0_outputs(2679) <= (inputs(84)) and not (inputs(4));
    layer0_outputs(2680) <= (inputs(218)) xor (inputs(186));
    layer0_outputs(2681) <= not((inputs(191)) or (inputs(243)));
    layer0_outputs(2682) <= (inputs(215)) or (inputs(116));
    layer0_outputs(2683) <= '1';
    layer0_outputs(2684) <= not((inputs(240)) xor (inputs(245)));
    layer0_outputs(2685) <= not(inputs(193)) or (inputs(0));
    layer0_outputs(2686) <= not((inputs(24)) or (inputs(177)));
    layer0_outputs(2687) <= '0';
    layer0_outputs(2688) <= inputs(89);
    layer0_outputs(2689) <= not((inputs(34)) xor (inputs(125)));
    layer0_outputs(2690) <= (inputs(68)) and not (inputs(158));
    layer0_outputs(2691) <= (inputs(69)) or (inputs(111));
    layer0_outputs(2692) <= not(inputs(210)) or (inputs(17));
    layer0_outputs(2693) <= not(inputs(239)) or (inputs(105));
    layer0_outputs(2694) <= inputs(253);
    layer0_outputs(2695) <= inputs(171);
    layer0_outputs(2696) <= not(inputs(88));
    layer0_outputs(2697) <= not((inputs(171)) or (inputs(8)));
    layer0_outputs(2698) <= '1';
    layer0_outputs(2699) <= not((inputs(123)) and (inputs(233)));
    layer0_outputs(2700) <= not(inputs(173)) or (inputs(154));
    layer0_outputs(2701) <= not(inputs(112));
    layer0_outputs(2702) <= (inputs(40)) and not (inputs(180));
    layer0_outputs(2703) <= not((inputs(42)) or (inputs(19)));
    layer0_outputs(2704) <= not((inputs(202)) and (inputs(247)));
    layer0_outputs(2705) <= not(inputs(64)) or (inputs(78));
    layer0_outputs(2706) <= (inputs(39)) and (inputs(181));
    layer0_outputs(2707) <= '0';
    layer0_outputs(2708) <= (inputs(151)) and not (inputs(115));
    layer0_outputs(2709) <= not(inputs(161)) or (inputs(75));
    layer0_outputs(2710) <= not((inputs(55)) and (inputs(96)));
    layer0_outputs(2711) <= (inputs(77)) xor (inputs(19));
    layer0_outputs(2712) <= (inputs(119)) or (inputs(238));
    layer0_outputs(2713) <= not((inputs(14)) xor (inputs(64)));
    layer0_outputs(2714) <= (inputs(231)) and not (inputs(148));
    layer0_outputs(2715) <= (inputs(183)) or (inputs(128));
    layer0_outputs(2716) <= (inputs(123)) or (inputs(224));
    layer0_outputs(2717) <= inputs(161);
    layer0_outputs(2718) <= not((inputs(180)) xor (inputs(174)));
    layer0_outputs(2719) <= inputs(146);
    layer0_outputs(2720) <= not(inputs(227));
    layer0_outputs(2721) <= not(inputs(33)) or (inputs(237));
    layer0_outputs(2722) <= inputs(164);
    layer0_outputs(2723) <= not(inputs(27)) or (inputs(242));
    layer0_outputs(2724) <= not(inputs(37));
    layer0_outputs(2725) <= not((inputs(103)) and (inputs(99)));
    layer0_outputs(2726) <= not((inputs(211)) or (inputs(249)));
    layer0_outputs(2727) <= not((inputs(222)) and (inputs(10)));
    layer0_outputs(2728) <= '1';
    layer0_outputs(2729) <= (inputs(118)) and not (inputs(39));
    layer0_outputs(2730) <= '1';
    layer0_outputs(2731) <= not(inputs(53));
    layer0_outputs(2732) <= not(inputs(6)) or (inputs(171));
    layer0_outputs(2733) <= not((inputs(208)) or (inputs(191)));
    layer0_outputs(2734) <= not((inputs(161)) or (inputs(159)));
    layer0_outputs(2735) <= not(inputs(5));
    layer0_outputs(2736) <= (inputs(203)) and not (inputs(215));
    layer0_outputs(2737) <= (inputs(244)) or (inputs(113));
    layer0_outputs(2738) <= not((inputs(53)) xor (inputs(201)));
    layer0_outputs(2739) <= (inputs(60)) or (inputs(207));
    layer0_outputs(2740) <= not((inputs(9)) or (inputs(99)));
    layer0_outputs(2741) <= not((inputs(105)) and (inputs(25)));
    layer0_outputs(2742) <= not(inputs(146));
    layer0_outputs(2743) <= (inputs(164)) and not (inputs(176));
    layer0_outputs(2744) <= inputs(9);
    layer0_outputs(2745) <= not(inputs(83));
    layer0_outputs(2746) <= not(inputs(205)) or (inputs(83));
    layer0_outputs(2747) <= (inputs(194)) xor (inputs(174));
    layer0_outputs(2748) <= not((inputs(190)) xor (inputs(134)));
    layer0_outputs(2749) <= not(inputs(107));
    layer0_outputs(2750) <= not(inputs(168));
    layer0_outputs(2751) <= not(inputs(214)) or (inputs(49));
    layer0_outputs(2752) <= '0';
    layer0_outputs(2753) <= '1';
    layer0_outputs(2754) <= (inputs(69)) or (inputs(226));
    layer0_outputs(2755) <= (inputs(124)) and not (inputs(225));
    layer0_outputs(2756) <= '1';
    layer0_outputs(2757) <= inputs(131);
    layer0_outputs(2758) <= not(inputs(117));
    layer0_outputs(2759) <= not((inputs(252)) or (inputs(218)));
    layer0_outputs(2760) <= (inputs(243)) and not (inputs(44));
    layer0_outputs(2761) <= (inputs(148)) and (inputs(172));
    layer0_outputs(2762) <= (inputs(195)) or (inputs(147));
    layer0_outputs(2763) <= not(inputs(195));
    layer0_outputs(2764) <= (inputs(203)) or (inputs(173));
    layer0_outputs(2765) <= not(inputs(144));
    layer0_outputs(2766) <= inputs(196);
    layer0_outputs(2767) <= (inputs(104)) and not (inputs(84));
    layer0_outputs(2768) <= not((inputs(241)) or (inputs(13)));
    layer0_outputs(2769) <= not(inputs(211));
    layer0_outputs(2770) <= not(inputs(172)) or (inputs(191));
    layer0_outputs(2771) <= inputs(233);
    layer0_outputs(2772) <= (inputs(86)) or (inputs(71));
    layer0_outputs(2773) <= (inputs(42)) or (inputs(48));
    layer0_outputs(2774) <= not((inputs(26)) xor (inputs(45)));
    layer0_outputs(2775) <= not((inputs(181)) or (inputs(174)));
    layer0_outputs(2776) <= not((inputs(133)) and (inputs(216)));
    layer0_outputs(2777) <= (inputs(165)) xor (inputs(237));
    layer0_outputs(2778) <= not(inputs(162)) or (inputs(94));
    layer0_outputs(2779) <= '1';
    layer0_outputs(2780) <= (inputs(153)) xor (inputs(185));
    layer0_outputs(2781) <= inputs(239);
    layer0_outputs(2782) <= (inputs(67)) and not (inputs(245));
    layer0_outputs(2783) <= not(inputs(38)) or (inputs(130));
    layer0_outputs(2784) <= not(inputs(101)) or (inputs(62));
    layer0_outputs(2785) <= inputs(215);
    layer0_outputs(2786) <= inputs(19);
    layer0_outputs(2787) <= not(inputs(173));
    layer0_outputs(2788) <= not(inputs(130));
    layer0_outputs(2789) <= not((inputs(138)) and (inputs(225)));
    layer0_outputs(2790) <= not((inputs(108)) xor (inputs(42)));
    layer0_outputs(2791) <= (inputs(57)) and not (inputs(19));
    layer0_outputs(2792) <= (inputs(192)) and (inputs(28));
    layer0_outputs(2793) <= not(inputs(137)) or (inputs(101));
    layer0_outputs(2794) <= not((inputs(152)) and (inputs(87)));
    layer0_outputs(2795) <= not((inputs(6)) xor (inputs(55)));
    layer0_outputs(2796) <= not((inputs(193)) or (inputs(76)));
    layer0_outputs(2797) <= not(inputs(169)) or (inputs(104));
    layer0_outputs(2798) <= (inputs(170)) and not (inputs(78));
    layer0_outputs(2799) <= not(inputs(10));
    layer0_outputs(2800) <= not((inputs(79)) or (inputs(16)));
    layer0_outputs(2801) <= (inputs(82)) and (inputs(39));
    layer0_outputs(2802) <= (inputs(162)) xor (inputs(221));
    layer0_outputs(2803) <= (inputs(189)) and not (inputs(31));
    layer0_outputs(2804) <= not(inputs(239)) or (inputs(148));
    layer0_outputs(2805) <= inputs(180);
    layer0_outputs(2806) <= not((inputs(23)) and (inputs(42)));
    layer0_outputs(2807) <= (inputs(45)) and not (inputs(191));
    layer0_outputs(2808) <= not(inputs(209)) or (inputs(20));
    layer0_outputs(2809) <= not((inputs(98)) or (inputs(164)));
    layer0_outputs(2810) <= (inputs(103)) and (inputs(188));
    layer0_outputs(2811) <= not((inputs(188)) and (inputs(21)));
    layer0_outputs(2812) <= (inputs(159)) or (inputs(151));
    layer0_outputs(2813) <= '0';
    layer0_outputs(2814) <= not((inputs(173)) or (inputs(118)));
    layer0_outputs(2815) <= inputs(232);
    layer0_outputs(2816) <= '1';
    layer0_outputs(2817) <= not(inputs(12)) or (inputs(213));
    layer0_outputs(2818) <= not(inputs(134));
    layer0_outputs(2819) <= not(inputs(246));
    layer0_outputs(2820) <= not((inputs(128)) or (inputs(155)));
    layer0_outputs(2821) <= (inputs(208)) and not (inputs(159));
    layer0_outputs(2822) <= '0';
    layer0_outputs(2823) <= not(inputs(158)) or (inputs(162));
    layer0_outputs(2824) <= (inputs(114)) and (inputs(207));
    layer0_outputs(2825) <= not((inputs(117)) and (inputs(69)));
    layer0_outputs(2826) <= not((inputs(242)) xor (inputs(213)));
    layer0_outputs(2827) <= not(inputs(57));
    layer0_outputs(2828) <= not(inputs(39)) or (inputs(182));
    layer0_outputs(2829) <= (inputs(158)) or (inputs(127));
    layer0_outputs(2830) <= inputs(126);
    layer0_outputs(2831) <= not(inputs(159));
    layer0_outputs(2832) <= '0';
    layer0_outputs(2833) <= inputs(41);
    layer0_outputs(2834) <= (inputs(136)) and not (inputs(144));
    layer0_outputs(2835) <= inputs(44);
    layer0_outputs(2836) <= not((inputs(143)) xor (inputs(206)));
    layer0_outputs(2837) <= not(inputs(123));
    layer0_outputs(2838) <= not(inputs(25));
    layer0_outputs(2839) <= inputs(105);
    layer0_outputs(2840) <= not((inputs(209)) xor (inputs(246)));
    layer0_outputs(2841) <= not(inputs(168));
    layer0_outputs(2842) <= (inputs(124)) and not (inputs(173));
    layer0_outputs(2843) <= inputs(200);
    layer0_outputs(2844) <= (inputs(172)) or (inputs(242));
    layer0_outputs(2845) <= (inputs(127)) and not (inputs(253));
    layer0_outputs(2846) <= not(inputs(230)) or (inputs(191));
    layer0_outputs(2847) <= not(inputs(85));
    layer0_outputs(2848) <= '1';
    layer0_outputs(2849) <= (inputs(239)) xor (inputs(22));
    layer0_outputs(2850) <= not((inputs(152)) or (inputs(150)));
    layer0_outputs(2851) <= not(inputs(249));
    layer0_outputs(2852) <= not(inputs(193)) or (inputs(25));
    layer0_outputs(2853) <= not(inputs(91));
    layer0_outputs(2854) <= (inputs(134)) and not (inputs(55));
    layer0_outputs(2855) <= not((inputs(196)) or (inputs(22)));
    layer0_outputs(2856) <= not((inputs(178)) or (inputs(207)));
    layer0_outputs(2857) <= not(inputs(39));
    layer0_outputs(2858) <= (inputs(67)) and not (inputs(10));
    layer0_outputs(2859) <= not(inputs(23)) or (inputs(130));
    layer0_outputs(2860) <= not(inputs(25)) or (inputs(144));
    layer0_outputs(2861) <= not((inputs(11)) or (inputs(52)));
    layer0_outputs(2862) <= (inputs(65)) and not (inputs(10));
    layer0_outputs(2863) <= not((inputs(77)) and (inputs(211)));
    layer0_outputs(2864) <= (inputs(98)) or (inputs(44));
    layer0_outputs(2865) <= not(inputs(149)) or (inputs(40));
    layer0_outputs(2866) <= (inputs(218)) and not (inputs(215));
    layer0_outputs(2867) <= not(inputs(249)) or (inputs(46));
    layer0_outputs(2868) <= not(inputs(100)) or (inputs(18));
    layer0_outputs(2869) <= (inputs(240)) and not (inputs(33));
    layer0_outputs(2870) <= inputs(128);
    layer0_outputs(2871) <= not((inputs(243)) or (inputs(46)));
    layer0_outputs(2872) <= (inputs(117)) or (inputs(186));
    layer0_outputs(2873) <= inputs(107);
    layer0_outputs(2874) <= (inputs(60)) and not (inputs(71));
    layer0_outputs(2875) <= (inputs(182)) or (inputs(174));
    layer0_outputs(2876) <= not(inputs(101));
    layer0_outputs(2877) <= inputs(102);
    layer0_outputs(2878) <= (inputs(187)) and not (inputs(3));
    layer0_outputs(2879) <= not((inputs(31)) or (inputs(163)));
    layer0_outputs(2880) <= inputs(125);
    layer0_outputs(2881) <= not((inputs(81)) or (inputs(245)));
    layer0_outputs(2882) <= not((inputs(79)) and (inputs(15)));
    layer0_outputs(2883) <= not(inputs(163));
    layer0_outputs(2884) <= (inputs(104)) xor (inputs(222));
    layer0_outputs(2885) <= (inputs(49)) or (inputs(73));
    layer0_outputs(2886) <= not(inputs(64));
    layer0_outputs(2887) <= (inputs(255)) and not (inputs(185));
    layer0_outputs(2888) <= not(inputs(43));
    layer0_outputs(2889) <= not(inputs(61)) or (inputs(145));
    layer0_outputs(2890) <= '0';
    layer0_outputs(2891) <= inputs(204);
    layer0_outputs(2892) <= not(inputs(36));
    layer0_outputs(2893) <= (inputs(22)) or (inputs(190));
    layer0_outputs(2894) <= not((inputs(191)) or (inputs(142)));
    layer0_outputs(2895) <= not(inputs(103));
    layer0_outputs(2896) <= inputs(101);
    layer0_outputs(2897) <= (inputs(167)) or (inputs(149));
    layer0_outputs(2898) <= '0';
    layer0_outputs(2899) <= (inputs(169)) and not (inputs(103));
    layer0_outputs(2900) <= not((inputs(80)) xor (inputs(24)));
    layer0_outputs(2901) <= (inputs(150)) or (inputs(182));
    layer0_outputs(2902) <= not((inputs(203)) or (inputs(205)));
    layer0_outputs(2903) <= not((inputs(53)) or (inputs(7)));
    layer0_outputs(2904) <= not(inputs(59)) or (inputs(194));
    layer0_outputs(2905) <= inputs(229);
    layer0_outputs(2906) <= (inputs(50)) and not (inputs(182));
    layer0_outputs(2907) <= inputs(164);
    layer0_outputs(2908) <= not((inputs(40)) or (inputs(55)));
    layer0_outputs(2909) <= '1';
    layer0_outputs(2910) <= (inputs(230)) and (inputs(59));
    layer0_outputs(2911) <= not(inputs(131));
    layer0_outputs(2912) <= (inputs(80)) or (inputs(130));
    layer0_outputs(2913) <= not(inputs(24));
    layer0_outputs(2914) <= inputs(153);
    layer0_outputs(2915) <= not(inputs(26));
    layer0_outputs(2916) <= '0';
    layer0_outputs(2917) <= (inputs(207)) or (inputs(199));
    layer0_outputs(2918) <= not(inputs(149)) or (inputs(19));
    layer0_outputs(2919) <= not((inputs(20)) or (inputs(255)));
    layer0_outputs(2920) <= (inputs(205)) xor (inputs(61));
    layer0_outputs(2921) <= not(inputs(168));
    layer0_outputs(2922) <= inputs(99);
    layer0_outputs(2923) <= inputs(77);
    layer0_outputs(2924) <= not((inputs(3)) or (inputs(63)));
    layer0_outputs(2925) <= not((inputs(85)) and (inputs(183)));
    layer0_outputs(2926) <= (inputs(216)) or (inputs(21));
    layer0_outputs(2927) <= not(inputs(27)) or (inputs(26));
    layer0_outputs(2928) <= (inputs(15)) and not (inputs(66));
    layer0_outputs(2929) <= (inputs(47)) and not (inputs(238));
    layer0_outputs(2930) <= (inputs(254)) or (inputs(243));
    layer0_outputs(2931) <= not(inputs(219));
    layer0_outputs(2932) <= not(inputs(54)) or (inputs(15));
    layer0_outputs(2933) <= '0';
    layer0_outputs(2934) <= (inputs(174)) xor (inputs(18));
    layer0_outputs(2935) <= '0';
    layer0_outputs(2936) <= (inputs(197)) and not (inputs(83));
    layer0_outputs(2937) <= (inputs(96)) and not (inputs(72));
    layer0_outputs(2938) <= (inputs(165)) or (inputs(18));
    layer0_outputs(2939) <= inputs(229);
    layer0_outputs(2940) <= '0';
    layer0_outputs(2941) <= (inputs(37)) or (inputs(18));
    layer0_outputs(2942) <= (inputs(188)) and not (inputs(3));
    layer0_outputs(2943) <= (inputs(82)) and (inputs(162));
    layer0_outputs(2944) <= '1';
    layer0_outputs(2945) <= not(inputs(119)) or (inputs(139));
    layer0_outputs(2946) <= '0';
    layer0_outputs(2947) <= not(inputs(88)) or (inputs(224));
    layer0_outputs(2948) <= (inputs(231)) xor (inputs(3));
    layer0_outputs(2949) <= not(inputs(89)) or (inputs(102));
    layer0_outputs(2950) <= (inputs(12)) or (inputs(165));
    layer0_outputs(2951) <= inputs(193);
    layer0_outputs(2952) <= not((inputs(249)) or (inputs(173)));
    layer0_outputs(2953) <= not((inputs(202)) and (inputs(232)));
    layer0_outputs(2954) <= not(inputs(87)) or (inputs(148));
    layer0_outputs(2955) <= not(inputs(189));
    layer0_outputs(2956) <= inputs(148);
    layer0_outputs(2957) <= not(inputs(36));
    layer0_outputs(2958) <= inputs(106);
    layer0_outputs(2959) <= (inputs(115)) or (inputs(239));
    layer0_outputs(2960) <= inputs(23);
    layer0_outputs(2961) <= (inputs(133)) or (inputs(115));
    layer0_outputs(2962) <= not(inputs(151));
    layer0_outputs(2963) <= not((inputs(169)) xor (inputs(119)));
    layer0_outputs(2964) <= (inputs(15)) or (inputs(198));
    layer0_outputs(2965) <= (inputs(95)) or (inputs(127));
    layer0_outputs(2966) <= inputs(199);
    layer0_outputs(2967) <= (inputs(110)) xor (inputs(96));
    layer0_outputs(2968) <= (inputs(220)) and (inputs(233));
    layer0_outputs(2969) <= not(inputs(211)) or (inputs(64));
    layer0_outputs(2970) <= (inputs(194)) or (inputs(80));
    layer0_outputs(2971) <= (inputs(50)) and not (inputs(211));
    layer0_outputs(2972) <= (inputs(11)) xor (inputs(18));
    layer0_outputs(2973) <= not(inputs(51));
    layer0_outputs(2974) <= (inputs(154)) and (inputs(42));
    layer0_outputs(2975) <= inputs(109);
    layer0_outputs(2976) <= not((inputs(200)) or (inputs(67)));
    layer0_outputs(2977) <= inputs(253);
    layer0_outputs(2978) <= (inputs(43)) or (inputs(3));
    layer0_outputs(2979) <= not((inputs(62)) or (inputs(17)));
    layer0_outputs(2980) <= not((inputs(252)) and (inputs(244)));
    layer0_outputs(2981) <= not((inputs(220)) or (inputs(82)));
    layer0_outputs(2982) <= not((inputs(51)) xor (inputs(20)));
    layer0_outputs(2983) <= (inputs(147)) xor (inputs(193));
    layer0_outputs(2984) <= (inputs(98)) or (inputs(185));
    layer0_outputs(2985) <= not(inputs(66)) or (inputs(179));
    layer0_outputs(2986) <= inputs(147);
    layer0_outputs(2987) <= not(inputs(153));
    layer0_outputs(2988) <= (inputs(141)) or (inputs(84));
    layer0_outputs(2989) <= inputs(105);
    layer0_outputs(2990) <= not((inputs(141)) and (inputs(197)));
    layer0_outputs(2991) <= not(inputs(148));
    layer0_outputs(2992) <= not(inputs(103));
    layer0_outputs(2993) <= not((inputs(6)) or (inputs(156)));
    layer0_outputs(2994) <= not(inputs(247)) or (inputs(50));
    layer0_outputs(2995) <= not(inputs(164)) or (inputs(140));
    layer0_outputs(2996) <= not((inputs(195)) and (inputs(99)));
    layer0_outputs(2997) <= inputs(245);
    layer0_outputs(2998) <= (inputs(247)) xor (inputs(178));
    layer0_outputs(2999) <= not(inputs(232));
    layer0_outputs(3000) <= '1';
    layer0_outputs(3001) <= (inputs(85)) or (inputs(11));
    layer0_outputs(3002) <= (inputs(224)) and not (inputs(236));
    layer0_outputs(3003) <= inputs(133);
    layer0_outputs(3004) <= not(inputs(198));
    layer0_outputs(3005) <= (inputs(128)) and not (inputs(255));
    layer0_outputs(3006) <= (inputs(77)) and not (inputs(137));
    layer0_outputs(3007) <= (inputs(193)) and not (inputs(251));
    layer0_outputs(3008) <= not(inputs(221));
    layer0_outputs(3009) <= (inputs(22)) and not (inputs(246));
    layer0_outputs(3010) <= (inputs(125)) and not (inputs(239));
    layer0_outputs(3011) <= not(inputs(38)) or (inputs(131));
    layer0_outputs(3012) <= (inputs(255)) and not (inputs(226));
    layer0_outputs(3013) <= '0';
    layer0_outputs(3014) <= not((inputs(9)) or (inputs(224)));
    layer0_outputs(3015) <= (inputs(58)) and not (inputs(238));
    layer0_outputs(3016) <= (inputs(68)) and not (inputs(196));
    layer0_outputs(3017) <= not(inputs(231));
    layer0_outputs(3018) <= not(inputs(48));
    layer0_outputs(3019) <= (inputs(78)) and (inputs(209));
    layer0_outputs(3020) <= inputs(13);
    layer0_outputs(3021) <= not(inputs(124));
    layer0_outputs(3022) <= (inputs(244)) and not (inputs(238));
    layer0_outputs(3023) <= inputs(53);
    layer0_outputs(3024) <= not(inputs(97));
    layer0_outputs(3025) <= not((inputs(28)) and (inputs(143)));
    layer0_outputs(3026) <= not(inputs(50)) or (inputs(75));
    layer0_outputs(3027) <= inputs(110);
    layer0_outputs(3028) <= not(inputs(53)) or (inputs(94));
    layer0_outputs(3029) <= inputs(130);
    layer0_outputs(3030) <= (inputs(131)) and not (inputs(205));
    layer0_outputs(3031) <= not((inputs(81)) and (inputs(112)));
    layer0_outputs(3032) <= not(inputs(103)) or (inputs(145));
    layer0_outputs(3033) <= inputs(122);
    layer0_outputs(3034) <= inputs(227);
    layer0_outputs(3035) <= not((inputs(4)) and (inputs(39)));
    layer0_outputs(3036) <= not(inputs(17));
    layer0_outputs(3037) <= (inputs(119)) and not (inputs(19));
    layer0_outputs(3038) <= (inputs(31)) and (inputs(164));
    layer0_outputs(3039) <= (inputs(153)) or (inputs(101));
    layer0_outputs(3040) <= not((inputs(251)) or (inputs(156)));
    layer0_outputs(3041) <= inputs(48);
    layer0_outputs(3042) <= not(inputs(100));
    layer0_outputs(3043) <= not(inputs(41));
    layer0_outputs(3044) <= not((inputs(224)) or (inputs(198)));
    layer0_outputs(3045) <= not(inputs(28));
    layer0_outputs(3046) <= not(inputs(123));
    layer0_outputs(3047) <= not((inputs(7)) or (inputs(122)));
    layer0_outputs(3048) <= inputs(205);
    layer0_outputs(3049) <= (inputs(82)) xor (inputs(233));
    layer0_outputs(3050) <= not((inputs(95)) xor (inputs(166)));
    layer0_outputs(3051) <= (inputs(208)) xor (inputs(0));
    layer0_outputs(3052) <= not((inputs(76)) xor (inputs(14)));
    layer0_outputs(3053) <= inputs(10);
    layer0_outputs(3054) <= '1';
    layer0_outputs(3055) <= not(inputs(38)) or (inputs(210));
    layer0_outputs(3056) <= inputs(42);
    layer0_outputs(3057) <= not(inputs(103)) or (inputs(203));
    layer0_outputs(3058) <= not((inputs(104)) and (inputs(23)));
    layer0_outputs(3059) <= '0';
    layer0_outputs(3060) <= not(inputs(148));
    layer0_outputs(3061) <= '1';
    layer0_outputs(3062) <= not(inputs(154)) or (inputs(227));
    layer0_outputs(3063) <= not((inputs(157)) or (inputs(220)));
    layer0_outputs(3064) <= '1';
    layer0_outputs(3065) <= not(inputs(54)) or (inputs(159));
    layer0_outputs(3066) <= (inputs(222)) or (inputs(180));
    layer0_outputs(3067) <= not(inputs(170));
    layer0_outputs(3068) <= not(inputs(173));
    layer0_outputs(3069) <= (inputs(184)) and not (inputs(112));
    layer0_outputs(3070) <= inputs(137);
    layer0_outputs(3071) <= (inputs(97)) or (inputs(224));
    layer0_outputs(3072) <= not((inputs(46)) or (inputs(235)));
    layer0_outputs(3073) <= not(inputs(39)) or (inputs(238));
    layer0_outputs(3074) <= (inputs(104)) and not (inputs(196));
    layer0_outputs(3075) <= not(inputs(228));
    layer0_outputs(3076) <= (inputs(252)) and (inputs(240));
    layer0_outputs(3077) <= inputs(177);
    layer0_outputs(3078) <= (inputs(60)) and not (inputs(154));
    layer0_outputs(3079) <= (inputs(22)) and not (inputs(164));
    layer0_outputs(3080) <= not((inputs(23)) or (inputs(64)));
    layer0_outputs(3081) <= inputs(104);
    layer0_outputs(3082) <= not(inputs(101));
    layer0_outputs(3083) <= not(inputs(241)) or (inputs(232));
    layer0_outputs(3084) <= (inputs(227)) and not (inputs(65));
    layer0_outputs(3085) <= not(inputs(13));
    layer0_outputs(3086) <= inputs(147);
    layer0_outputs(3087) <= not((inputs(88)) or (inputs(28)));
    layer0_outputs(3088) <= (inputs(122)) and not (inputs(94));
    layer0_outputs(3089) <= not((inputs(100)) xor (inputs(129)));
    layer0_outputs(3090) <= inputs(245);
    layer0_outputs(3091) <= not((inputs(78)) or (inputs(110)));
    layer0_outputs(3092) <= (inputs(235)) or (inputs(80));
    layer0_outputs(3093) <= (inputs(61)) and (inputs(237));
    layer0_outputs(3094) <= not(inputs(15));
    layer0_outputs(3095) <= not((inputs(16)) or (inputs(42)));
    layer0_outputs(3096) <= '0';
    layer0_outputs(3097) <= inputs(162);
    layer0_outputs(3098) <= not((inputs(5)) or (inputs(180)));
    layer0_outputs(3099) <= (inputs(243)) or (inputs(219));
    layer0_outputs(3100) <= (inputs(188)) or (inputs(108));
    layer0_outputs(3101) <= (inputs(120)) and not (inputs(206));
    layer0_outputs(3102) <= (inputs(222)) and not (inputs(15));
    layer0_outputs(3103) <= inputs(183);
    layer0_outputs(3104) <= not(inputs(217));
    layer0_outputs(3105) <= '0';
    layer0_outputs(3106) <= not(inputs(181));
    layer0_outputs(3107) <= not((inputs(75)) and (inputs(10)));
    layer0_outputs(3108) <= not((inputs(77)) and (inputs(63)));
    layer0_outputs(3109) <= inputs(185);
    layer0_outputs(3110) <= inputs(184);
    layer0_outputs(3111) <= '1';
    layer0_outputs(3112) <= not(inputs(153)) or (inputs(67));
    layer0_outputs(3113) <= (inputs(245)) and not (inputs(20));
    layer0_outputs(3114) <= not((inputs(18)) or (inputs(14)));
    layer0_outputs(3115) <= (inputs(211)) and not (inputs(239));
    layer0_outputs(3116) <= (inputs(28)) xor (inputs(71));
    layer0_outputs(3117) <= not((inputs(252)) or (inputs(150)));
    layer0_outputs(3118) <= not((inputs(219)) or (inputs(224)));
    layer0_outputs(3119) <= (inputs(26)) or (inputs(21));
    layer0_outputs(3120) <= inputs(160);
    layer0_outputs(3121) <= not((inputs(190)) or (inputs(100)));
    layer0_outputs(3122) <= (inputs(78)) and not (inputs(219));
    layer0_outputs(3123) <= not(inputs(197));
    layer0_outputs(3124) <= not(inputs(162));
    layer0_outputs(3125) <= inputs(236);
    layer0_outputs(3126) <= inputs(119);
    layer0_outputs(3127) <= not(inputs(222)) or (inputs(143));
    layer0_outputs(3128) <= not(inputs(159));
    layer0_outputs(3129) <= (inputs(27)) and (inputs(20));
    layer0_outputs(3130) <= not((inputs(35)) xor (inputs(111)));
    layer0_outputs(3131) <= '1';
    layer0_outputs(3132) <= not(inputs(212)) or (inputs(239));
    layer0_outputs(3133) <= inputs(218);
    layer0_outputs(3134) <= not(inputs(142));
    layer0_outputs(3135) <= not(inputs(146)) or (inputs(61));
    layer0_outputs(3136) <= (inputs(30)) and not (inputs(2));
    layer0_outputs(3137) <= (inputs(240)) and (inputs(198));
    layer0_outputs(3138) <= (inputs(132)) and not (inputs(175));
    layer0_outputs(3139) <= not(inputs(91));
    layer0_outputs(3140) <= not((inputs(249)) or (inputs(233)));
    layer0_outputs(3141) <= inputs(3);
    layer0_outputs(3142) <= inputs(207);
    layer0_outputs(3143) <= not(inputs(89));
    layer0_outputs(3144) <= not((inputs(104)) or (inputs(206)));
    layer0_outputs(3145) <= not(inputs(2));
    layer0_outputs(3146) <= not(inputs(205));
    layer0_outputs(3147) <= (inputs(233)) and not (inputs(170));
    layer0_outputs(3148) <= not((inputs(176)) or (inputs(216)));
    layer0_outputs(3149) <= '0';
    layer0_outputs(3150) <= not((inputs(114)) or (inputs(162)));
    layer0_outputs(3151) <= inputs(221);
    layer0_outputs(3152) <= not(inputs(186));
    layer0_outputs(3153) <= inputs(106);
    layer0_outputs(3154) <= not(inputs(59));
    layer0_outputs(3155) <= (inputs(182)) and not (inputs(114));
    layer0_outputs(3156) <= not(inputs(66)) or (inputs(148));
    layer0_outputs(3157) <= not(inputs(168));
    layer0_outputs(3158) <= inputs(148);
    layer0_outputs(3159) <= inputs(181);
    layer0_outputs(3160) <= not(inputs(162));
    layer0_outputs(3161) <= inputs(178);
    layer0_outputs(3162) <= not(inputs(214));
    layer0_outputs(3163) <= not((inputs(89)) and (inputs(248)));
    layer0_outputs(3164) <= inputs(59);
    layer0_outputs(3165) <= not(inputs(119)) or (inputs(131));
    layer0_outputs(3166) <= not(inputs(145));
    layer0_outputs(3167) <= not(inputs(219)) or (inputs(228));
    layer0_outputs(3168) <= not(inputs(159));
    layer0_outputs(3169) <= inputs(70);
    layer0_outputs(3170) <= inputs(166);
    layer0_outputs(3171) <= (inputs(120)) and (inputs(87));
    layer0_outputs(3172) <= inputs(169);
    layer0_outputs(3173) <= inputs(90);
    layer0_outputs(3174) <= (inputs(144)) xor (inputs(223));
    layer0_outputs(3175) <= not((inputs(221)) or (inputs(238)));
    layer0_outputs(3176) <= '0';
    layer0_outputs(3177) <= (inputs(162)) or (inputs(221));
    layer0_outputs(3178) <= inputs(173);
    layer0_outputs(3179) <= not(inputs(169));
    layer0_outputs(3180) <= not(inputs(20));
    layer0_outputs(3181) <= (inputs(171)) and not (inputs(74));
    layer0_outputs(3182) <= not((inputs(152)) and (inputs(119)));
    layer0_outputs(3183) <= not(inputs(229)) or (inputs(61));
    layer0_outputs(3184) <= inputs(23);
    layer0_outputs(3185) <= not((inputs(17)) or (inputs(108)));
    layer0_outputs(3186) <= inputs(232);
    layer0_outputs(3187) <= (inputs(34)) xor (inputs(54));
    layer0_outputs(3188) <= '0';
    layer0_outputs(3189) <= '0';
    layer0_outputs(3190) <= (inputs(162)) and not (inputs(17));
    layer0_outputs(3191) <= not(inputs(147));
    layer0_outputs(3192) <= (inputs(122)) and not (inputs(86));
    layer0_outputs(3193) <= (inputs(6)) or (inputs(89));
    layer0_outputs(3194) <= not((inputs(249)) or (inputs(29)));
    layer0_outputs(3195) <= not((inputs(186)) or (inputs(237)));
    layer0_outputs(3196) <= not((inputs(60)) or (inputs(5)));
    layer0_outputs(3197) <= inputs(9);
    layer0_outputs(3198) <= (inputs(63)) xor (inputs(76));
    layer0_outputs(3199) <= not(inputs(223)) or (inputs(85));
    layer0_outputs(3200) <= (inputs(70)) xor (inputs(3));
    layer0_outputs(3201) <= (inputs(33)) or (inputs(38));
    layer0_outputs(3202) <= not((inputs(129)) or (inputs(142)));
    layer0_outputs(3203) <= (inputs(90)) and (inputs(151));
    layer0_outputs(3204) <= '1';
    layer0_outputs(3205) <= not(inputs(140)) or (inputs(206));
    layer0_outputs(3206) <= not(inputs(119)) or (inputs(118));
    layer0_outputs(3207) <= '1';
    layer0_outputs(3208) <= not(inputs(201));
    layer0_outputs(3209) <= '1';
    layer0_outputs(3210) <= not(inputs(48)) or (inputs(16));
    layer0_outputs(3211) <= not(inputs(88));
    layer0_outputs(3212) <= inputs(233);
    layer0_outputs(3213) <= inputs(45);
    layer0_outputs(3214) <= not(inputs(106));
    layer0_outputs(3215) <= inputs(38);
    layer0_outputs(3216) <= (inputs(73)) and (inputs(28));
    layer0_outputs(3217) <= inputs(25);
    layer0_outputs(3218) <= (inputs(103)) and not (inputs(40));
    layer0_outputs(3219) <= (inputs(126)) or (inputs(198));
    layer0_outputs(3220) <= (inputs(183)) and not (inputs(46));
    layer0_outputs(3221) <= inputs(126);
    layer0_outputs(3222) <= not(inputs(76));
    layer0_outputs(3223) <= inputs(54);
    layer0_outputs(3224) <= (inputs(18)) or (inputs(245));
    layer0_outputs(3225) <= '0';
    layer0_outputs(3226) <= (inputs(44)) and not (inputs(252));
    layer0_outputs(3227) <= not((inputs(144)) or (inputs(65)));
    layer0_outputs(3228) <= not(inputs(5)) or (inputs(149));
    layer0_outputs(3229) <= (inputs(138)) and not (inputs(199));
    layer0_outputs(3230) <= (inputs(77)) or (inputs(176));
    layer0_outputs(3231) <= inputs(44);
    layer0_outputs(3232) <= not((inputs(156)) and (inputs(252)));
    layer0_outputs(3233) <= (inputs(123)) or (inputs(172));
    layer0_outputs(3234) <= not((inputs(218)) or (inputs(226)));
    layer0_outputs(3235) <= (inputs(163)) or (inputs(98));
    layer0_outputs(3236) <= (inputs(217)) or (inputs(218));
    layer0_outputs(3237) <= inputs(186);
    layer0_outputs(3238) <= not((inputs(39)) and (inputs(254)));
    layer0_outputs(3239) <= '1';
    layer0_outputs(3240) <= (inputs(247)) or (inputs(67));
    layer0_outputs(3241) <= (inputs(91)) or (inputs(237));
    layer0_outputs(3242) <= (inputs(70)) xor (inputs(37));
    layer0_outputs(3243) <= not((inputs(160)) or (inputs(169)));
    layer0_outputs(3244) <= inputs(35);
    layer0_outputs(3245) <= not(inputs(238));
    layer0_outputs(3246) <= inputs(104);
    layer0_outputs(3247) <= not((inputs(137)) or (inputs(125)));
    layer0_outputs(3248) <= inputs(150);
    layer0_outputs(3249) <= not((inputs(240)) xor (inputs(207)));
    layer0_outputs(3250) <= not(inputs(133)) or (inputs(124));
    layer0_outputs(3251) <= not(inputs(18));
    layer0_outputs(3252) <= not((inputs(110)) and (inputs(32)));
    layer0_outputs(3253) <= not(inputs(41)) or (inputs(243));
    layer0_outputs(3254) <= inputs(100);
    layer0_outputs(3255) <= not(inputs(196));
    layer0_outputs(3256) <= not(inputs(148));
    layer0_outputs(3257) <= not((inputs(174)) or (inputs(65)));
    layer0_outputs(3258) <= not(inputs(251));
    layer0_outputs(3259) <= not((inputs(113)) or (inputs(49)));
    layer0_outputs(3260) <= (inputs(65)) or (inputs(217));
    layer0_outputs(3261) <= not(inputs(229)) or (inputs(225));
    layer0_outputs(3262) <= inputs(139);
    layer0_outputs(3263) <= (inputs(52)) or (inputs(60));
    layer0_outputs(3264) <= (inputs(184)) or (inputs(98));
    layer0_outputs(3265) <= (inputs(54)) and not (inputs(46));
    layer0_outputs(3266) <= (inputs(237)) or (inputs(97));
    layer0_outputs(3267) <= (inputs(244)) or (inputs(56));
    layer0_outputs(3268) <= '0';
    layer0_outputs(3269) <= inputs(115);
    layer0_outputs(3270) <= inputs(187);
    layer0_outputs(3271) <= (inputs(148)) and (inputs(70));
    layer0_outputs(3272) <= (inputs(52)) xor (inputs(235));
    layer0_outputs(3273) <= '1';
    layer0_outputs(3274) <= (inputs(170)) and not (inputs(51));
    layer0_outputs(3275) <= inputs(42);
    layer0_outputs(3276) <= not(inputs(193)) or (inputs(151));
    layer0_outputs(3277) <= not(inputs(118));
    layer0_outputs(3278) <= (inputs(135)) and not (inputs(235));
    layer0_outputs(3279) <= not(inputs(229));
    layer0_outputs(3280) <= inputs(214);
    layer0_outputs(3281) <= (inputs(219)) or (inputs(126));
    layer0_outputs(3282) <= not(inputs(14)) or (inputs(140));
    layer0_outputs(3283) <= (inputs(175)) or (inputs(142));
    layer0_outputs(3284) <= not(inputs(34)) or (inputs(92));
    layer0_outputs(3285) <= '1';
    layer0_outputs(3286) <= (inputs(178)) or (inputs(79));
    layer0_outputs(3287) <= not(inputs(25));
    layer0_outputs(3288) <= (inputs(93)) or (inputs(183));
    layer0_outputs(3289) <= '0';
    layer0_outputs(3290) <= not(inputs(58)) or (inputs(66));
    layer0_outputs(3291) <= (inputs(24)) or (inputs(177));
    layer0_outputs(3292) <= (inputs(236)) and not (inputs(125));
    layer0_outputs(3293) <= not((inputs(195)) or (inputs(185)));
    layer0_outputs(3294) <= not(inputs(24));
    layer0_outputs(3295) <= not(inputs(101));
    layer0_outputs(3296) <= (inputs(134)) and not (inputs(34));
    layer0_outputs(3297) <= (inputs(30)) and not (inputs(163));
    layer0_outputs(3298) <= (inputs(81)) or (inputs(98));
    layer0_outputs(3299) <= (inputs(86)) and not (inputs(240));
    layer0_outputs(3300) <= not(inputs(170));
    layer0_outputs(3301) <= (inputs(21)) and not (inputs(214));
    layer0_outputs(3302) <= not((inputs(252)) and (inputs(242)));
    layer0_outputs(3303) <= not(inputs(194));
    layer0_outputs(3304) <= inputs(235);
    layer0_outputs(3305) <= inputs(169);
    layer0_outputs(3306) <= inputs(187);
    layer0_outputs(3307) <= (inputs(221)) and not (inputs(49));
    layer0_outputs(3308) <= not(inputs(38));
    layer0_outputs(3309) <= (inputs(10)) and not (inputs(159));
    layer0_outputs(3310) <= (inputs(135)) or (inputs(207));
    layer0_outputs(3311) <= inputs(247);
    layer0_outputs(3312) <= inputs(26);
    layer0_outputs(3313) <= (inputs(7)) or (inputs(206));
    layer0_outputs(3314) <= not((inputs(228)) or (inputs(177)));
    layer0_outputs(3315) <= (inputs(147)) xor (inputs(63));
    layer0_outputs(3316) <= not((inputs(109)) or (inputs(85)));
    layer0_outputs(3317) <= (inputs(135)) and not (inputs(254));
    layer0_outputs(3318) <= (inputs(165)) or (inputs(200));
    layer0_outputs(3319) <= (inputs(10)) and not (inputs(194));
    layer0_outputs(3320) <= inputs(112);
    layer0_outputs(3321) <= '0';
    layer0_outputs(3322) <= not(inputs(248));
    layer0_outputs(3323) <= (inputs(246)) xor (inputs(250));
    layer0_outputs(3324) <= not(inputs(152)) or (inputs(50));
    layer0_outputs(3325) <= (inputs(104)) and not (inputs(80));
    layer0_outputs(3326) <= not(inputs(126));
    layer0_outputs(3327) <= not(inputs(210));
    layer0_outputs(3328) <= not((inputs(59)) xor (inputs(237)));
    layer0_outputs(3329) <= not(inputs(236)) or (inputs(44));
    layer0_outputs(3330) <= (inputs(216)) and not (inputs(140));
    layer0_outputs(3331) <= inputs(33);
    layer0_outputs(3332) <= (inputs(125)) and (inputs(93));
    layer0_outputs(3333) <= inputs(98);
    layer0_outputs(3334) <= inputs(88);
    layer0_outputs(3335) <= not((inputs(234)) xor (inputs(169)));
    layer0_outputs(3336) <= (inputs(174)) xor (inputs(43));
    layer0_outputs(3337) <= not(inputs(146));
    layer0_outputs(3338) <= not((inputs(219)) xor (inputs(67)));
    layer0_outputs(3339) <= not(inputs(135));
    layer0_outputs(3340) <= not((inputs(100)) and (inputs(78)));
    layer0_outputs(3341) <= '1';
    layer0_outputs(3342) <= not(inputs(9));
    layer0_outputs(3343) <= '0';
    layer0_outputs(3344) <= inputs(18);
    layer0_outputs(3345) <= not(inputs(45));
    layer0_outputs(3346) <= not((inputs(191)) or (inputs(137)));
    layer0_outputs(3347) <= not((inputs(207)) or (inputs(167)));
    layer0_outputs(3348) <= (inputs(97)) or (inputs(100));
    layer0_outputs(3349) <= (inputs(204)) and not (inputs(46));
    layer0_outputs(3350) <= (inputs(16)) or (inputs(225));
    layer0_outputs(3351) <= not((inputs(131)) xor (inputs(28)));
    layer0_outputs(3352) <= not((inputs(49)) or (inputs(68)));
    layer0_outputs(3353) <= (inputs(194)) or (inputs(201));
    layer0_outputs(3354) <= not(inputs(40)) or (inputs(120));
    layer0_outputs(3355) <= inputs(119);
    layer0_outputs(3356) <= not((inputs(181)) or (inputs(149)));
    layer0_outputs(3357) <= inputs(229);
    layer0_outputs(3358) <= not(inputs(131));
    layer0_outputs(3359) <= not(inputs(135));
    layer0_outputs(3360) <= (inputs(190)) and (inputs(5));
    layer0_outputs(3361) <= not((inputs(123)) or (inputs(217)));
    layer0_outputs(3362) <= not(inputs(231));
    layer0_outputs(3363) <= not((inputs(71)) or (inputs(177)));
    layer0_outputs(3364) <= not((inputs(224)) xor (inputs(32)));
    layer0_outputs(3365) <= (inputs(207)) and not (inputs(129));
    layer0_outputs(3366) <= (inputs(86)) xor (inputs(97));
    layer0_outputs(3367) <= '1';
    layer0_outputs(3368) <= not(inputs(111));
    layer0_outputs(3369) <= inputs(38);
    layer0_outputs(3370) <= (inputs(176)) or (inputs(42));
    layer0_outputs(3371) <= not(inputs(119));
    layer0_outputs(3372) <= not(inputs(182));
    layer0_outputs(3373) <= inputs(104);
    layer0_outputs(3374) <= not(inputs(13));
    layer0_outputs(3375) <= (inputs(198)) and not (inputs(96));
    layer0_outputs(3376) <= not((inputs(171)) xor (inputs(173)));
    layer0_outputs(3377) <= (inputs(213)) xor (inputs(195));
    layer0_outputs(3378) <= not(inputs(121)) or (inputs(194));
    layer0_outputs(3379) <= not(inputs(191));
    layer0_outputs(3380) <= inputs(60);
    layer0_outputs(3381) <= not((inputs(70)) xor (inputs(177)));
    layer0_outputs(3382) <= '1';
    layer0_outputs(3383) <= (inputs(61)) and (inputs(20));
    layer0_outputs(3384) <= not(inputs(205)) or (inputs(12));
    layer0_outputs(3385) <= inputs(87);
    layer0_outputs(3386) <= (inputs(27)) and (inputs(1));
    layer0_outputs(3387) <= inputs(21);
    layer0_outputs(3388) <= (inputs(119)) or (inputs(134));
    layer0_outputs(3389) <= not((inputs(87)) or (inputs(100)));
    layer0_outputs(3390) <= not(inputs(6)) or (inputs(15));
    layer0_outputs(3391) <= inputs(105);
    layer0_outputs(3392) <= not(inputs(233)) or (inputs(130));
    layer0_outputs(3393) <= (inputs(164)) or (inputs(104));
    layer0_outputs(3394) <= inputs(246);
    layer0_outputs(3395) <= (inputs(12)) or (inputs(134));
    layer0_outputs(3396) <= (inputs(188)) or (inputs(62));
    layer0_outputs(3397) <= (inputs(4)) and (inputs(144));
    layer0_outputs(3398) <= not(inputs(208)) or (inputs(161));
    layer0_outputs(3399) <= '0';
    layer0_outputs(3400) <= (inputs(138)) or (inputs(68));
    layer0_outputs(3401) <= not((inputs(44)) or (inputs(115)));
    layer0_outputs(3402) <= (inputs(188)) and (inputs(151));
    layer0_outputs(3403) <= not((inputs(237)) xor (inputs(179)));
    layer0_outputs(3404) <= inputs(232);
    layer0_outputs(3405) <= not(inputs(53));
    layer0_outputs(3406) <= not((inputs(243)) or (inputs(207)));
    layer0_outputs(3407) <= not(inputs(67));
    layer0_outputs(3408) <= inputs(131);
    layer0_outputs(3409) <= not(inputs(150)) or (inputs(232));
    layer0_outputs(3410) <= not(inputs(136)) or (inputs(209));
    layer0_outputs(3411) <= (inputs(127)) or (inputs(233));
    layer0_outputs(3412) <= (inputs(244)) and not (inputs(50));
    layer0_outputs(3413) <= not(inputs(86));
    layer0_outputs(3414) <= (inputs(61)) or (inputs(97));
    layer0_outputs(3415) <= (inputs(166)) and not (inputs(81));
    layer0_outputs(3416) <= (inputs(18)) and not (inputs(11));
    layer0_outputs(3417) <= inputs(203);
    layer0_outputs(3418) <= inputs(189);
    layer0_outputs(3419) <= not((inputs(114)) or (inputs(97)));
    layer0_outputs(3420) <= not((inputs(200)) and (inputs(200)));
    layer0_outputs(3421) <= (inputs(210)) and not (inputs(128));
    layer0_outputs(3422) <= (inputs(4)) xor (inputs(126));
    layer0_outputs(3423) <= not(inputs(10));
    layer0_outputs(3424) <= not((inputs(236)) xor (inputs(142)));
    layer0_outputs(3425) <= not(inputs(89));
    layer0_outputs(3426) <= (inputs(209)) or (inputs(24));
    layer0_outputs(3427) <= (inputs(190)) or (inputs(125));
    layer0_outputs(3428) <= (inputs(3)) and (inputs(253));
    layer0_outputs(3429) <= (inputs(102)) or (inputs(15));
    layer0_outputs(3430) <= inputs(163);
    layer0_outputs(3431) <= (inputs(38)) or (inputs(60));
    layer0_outputs(3432) <= not(inputs(21)) or (inputs(144));
    layer0_outputs(3433) <= (inputs(92)) and not (inputs(47));
    layer0_outputs(3434) <= not(inputs(10)) or (inputs(241));
    layer0_outputs(3435) <= not(inputs(238));
    layer0_outputs(3436) <= (inputs(74)) and not (inputs(196));
    layer0_outputs(3437) <= not(inputs(227));
    layer0_outputs(3438) <= not((inputs(174)) xor (inputs(116)));
    layer0_outputs(3439) <= not((inputs(177)) xor (inputs(236)));
    layer0_outputs(3440) <= '1';
    layer0_outputs(3441) <= not((inputs(60)) xor (inputs(20)));
    layer0_outputs(3442) <= not(inputs(200));
    layer0_outputs(3443) <= not(inputs(178));
    layer0_outputs(3444) <= (inputs(140)) and not (inputs(81));
    layer0_outputs(3445) <= '1';
    layer0_outputs(3446) <= (inputs(197)) xor (inputs(245));
    layer0_outputs(3447) <= inputs(99);
    layer0_outputs(3448) <= inputs(40);
    layer0_outputs(3449) <= not((inputs(104)) xor (inputs(127)));
    layer0_outputs(3450) <= (inputs(223)) or (inputs(139));
    layer0_outputs(3451) <= inputs(106);
    layer0_outputs(3452) <= inputs(138);
    layer0_outputs(3453) <= (inputs(35)) xor (inputs(77));
    layer0_outputs(3454) <= not(inputs(254)) or (inputs(62));
    layer0_outputs(3455) <= not(inputs(81));
    layer0_outputs(3456) <= not(inputs(161));
    layer0_outputs(3457) <= not(inputs(236)) or (inputs(204));
    layer0_outputs(3458) <= not((inputs(103)) or (inputs(255)));
    layer0_outputs(3459) <= not(inputs(26));
    layer0_outputs(3460) <= (inputs(138)) and not (inputs(132));
    layer0_outputs(3461) <= not(inputs(120)) or (inputs(85));
    layer0_outputs(3462) <= inputs(138);
    layer0_outputs(3463) <= not((inputs(184)) or (inputs(166)));
    layer0_outputs(3464) <= inputs(172);
    layer0_outputs(3465) <= not(inputs(168));
    layer0_outputs(3466) <= not(inputs(86));
    layer0_outputs(3467) <= inputs(138);
    layer0_outputs(3468) <= inputs(61);
    layer0_outputs(3469) <= not(inputs(138)) or (inputs(158));
    layer0_outputs(3470) <= not(inputs(157));
    layer0_outputs(3471) <= not(inputs(189)) or (inputs(41));
    layer0_outputs(3472) <= not((inputs(89)) or (inputs(105)));
    layer0_outputs(3473) <= not(inputs(148)) or (inputs(52));
    layer0_outputs(3474) <= inputs(201);
    layer0_outputs(3475) <= (inputs(5)) or (inputs(31));
    layer0_outputs(3476) <= not((inputs(243)) or (inputs(120)));
    layer0_outputs(3477) <= not(inputs(243));
    layer0_outputs(3478) <= not((inputs(220)) or (inputs(124)));
    layer0_outputs(3479) <= (inputs(132)) and not (inputs(170));
    layer0_outputs(3480) <= not(inputs(126));
    layer0_outputs(3481) <= (inputs(227)) and not (inputs(67));
    layer0_outputs(3482) <= inputs(87);
    layer0_outputs(3483) <= not(inputs(217)) or (inputs(91));
    layer0_outputs(3484) <= (inputs(221)) or (inputs(216));
    layer0_outputs(3485) <= not((inputs(93)) or (inputs(2)));
    layer0_outputs(3486) <= not((inputs(101)) and (inputs(169)));
    layer0_outputs(3487) <= (inputs(24)) and not (inputs(241));
    layer0_outputs(3488) <= not(inputs(249));
    layer0_outputs(3489) <= '1';
    layer0_outputs(3490) <= not(inputs(23)) or (inputs(113));
    layer0_outputs(3491) <= inputs(166);
    layer0_outputs(3492) <= (inputs(224)) or (inputs(19));
    layer0_outputs(3493) <= (inputs(234)) and not (inputs(17));
    layer0_outputs(3494) <= not(inputs(63));
    layer0_outputs(3495) <= inputs(158);
    layer0_outputs(3496) <= (inputs(5)) or (inputs(35));
    layer0_outputs(3497) <= (inputs(160)) xor (inputs(163));
    layer0_outputs(3498) <= not(inputs(152)) or (inputs(81));
    layer0_outputs(3499) <= '1';
    layer0_outputs(3500) <= inputs(160);
    layer0_outputs(3501) <= not((inputs(116)) or (inputs(137)));
    layer0_outputs(3502) <= not(inputs(234));
    layer0_outputs(3503) <= not(inputs(34)) or (inputs(78));
    layer0_outputs(3504) <= not((inputs(93)) and (inputs(12)));
    layer0_outputs(3505) <= not(inputs(105));
    layer0_outputs(3506) <= not(inputs(163)) or (inputs(151));
    layer0_outputs(3507) <= not(inputs(197)) or (inputs(15));
    layer0_outputs(3508) <= inputs(203);
    layer0_outputs(3509) <= '0';
    layer0_outputs(3510) <= not(inputs(234)) or (inputs(16));
    layer0_outputs(3511) <= (inputs(243)) and not (inputs(42));
    layer0_outputs(3512) <= not(inputs(166));
    layer0_outputs(3513) <= not(inputs(71)) or (inputs(151));
    layer0_outputs(3514) <= (inputs(156)) or (inputs(59));
    layer0_outputs(3515) <= not((inputs(0)) or (inputs(189)));
    layer0_outputs(3516) <= not(inputs(149));
    layer0_outputs(3517) <= not(inputs(189)) or (inputs(107));
    layer0_outputs(3518) <= (inputs(43)) and not (inputs(239));
    layer0_outputs(3519) <= not(inputs(158));
    layer0_outputs(3520) <= not((inputs(66)) or (inputs(20)));
    layer0_outputs(3521) <= '0';
    layer0_outputs(3522) <= not((inputs(190)) or (inputs(30)));
    layer0_outputs(3523) <= not(inputs(103));
    layer0_outputs(3524) <= (inputs(126)) or (inputs(182));
    layer0_outputs(3525) <= not(inputs(99)) or (inputs(208));
    layer0_outputs(3526) <= inputs(120);
    layer0_outputs(3527) <= (inputs(120)) or (inputs(34));
    layer0_outputs(3528) <= not(inputs(38)) or (inputs(255));
    layer0_outputs(3529) <= not(inputs(191));
    layer0_outputs(3530) <= not(inputs(254));
    layer0_outputs(3531) <= (inputs(125)) or (inputs(154));
    layer0_outputs(3532) <= not(inputs(219));
    layer0_outputs(3533) <= not(inputs(92));
    layer0_outputs(3534) <= not(inputs(10)) or (inputs(65));
    layer0_outputs(3535) <= '1';
    layer0_outputs(3536) <= inputs(16);
    layer0_outputs(3537) <= '0';
    layer0_outputs(3538) <= '1';
    layer0_outputs(3539) <= not((inputs(53)) xor (inputs(169)));
    layer0_outputs(3540) <= (inputs(8)) and not (inputs(199));
    layer0_outputs(3541) <= not(inputs(90)) or (inputs(249));
    layer0_outputs(3542) <= not((inputs(71)) xor (inputs(34)));
    layer0_outputs(3543) <= inputs(20);
    layer0_outputs(3544) <= inputs(27);
    layer0_outputs(3545) <= (inputs(174)) or (inputs(179));
    layer0_outputs(3546) <= not(inputs(54)) or (inputs(115));
    layer0_outputs(3547) <= not(inputs(134));
    layer0_outputs(3548) <= not((inputs(254)) or (inputs(253)));
    layer0_outputs(3549) <= not(inputs(40));
    layer0_outputs(3550) <= (inputs(166)) xor (inputs(132));
    layer0_outputs(3551) <= not((inputs(174)) or (inputs(40)));
    layer0_outputs(3552) <= not((inputs(105)) xor (inputs(124)));
    layer0_outputs(3553) <= not(inputs(14)) or (inputs(184));
    layer0_outputs(3554) <= not(inputs(79));
    layer0_outputs(3555) <= not(inputs(130));
    layer0_outputs(3556) <= not((inputs(129)) or (inputs(82)));
    layer0_outputs(3557) <= inputs(67);
    layer0_outputs(3558) <= inputs(242);
    layer0_outputs(3559) <= not((inputs(205)) or (inputs(255)));
    layer0_outputs(3560) <= inputs(126);
    layer0_outputs(3561) <= not(inputs(180));
    layer0_outputs(3562) <= (inputs(67)) and not (inputs(112));
    layer0_outputs(3563) <= not(inputs(58));
    layer0_outputs(3564) <= not((inputs(170)) or (inputs(177)));
    layer0_outputs(3565) <= (inputs(139)) or (inputs(202));
    layer0_outputs(3566) <= not(inputs(210));
    layer0_outputs(3567) <= not(inputs(85));
    layer0_outputs(3568) <= inputs(185);
    layer0_outputs(3569) <= not(inputs(232));
    layer0_outputs(3570) <= (inputs(150)) or (inputs(150));
    layer0_outputs(3571) <= '1';
    layer0_outputs(3572) <= not((inputs(218)) or (inputs(36)));
    layer0_outputs(3573) <= '1';
    layer0_outputs(3574) <= inputs(147);
    layer0_outputs(3575) <= not(inputs(206));
    layer0_outputs(3576) <= inputs(66);
    layer0_outputs(3577) <= not(inputs(132));
    layer0_outputs(3578) <= (inputs(115)) and not (inputs(210));
    layer0_outputs(3579) <= not(inputs(117));
    layer0_outputs(3580) <= '1';
    layer0_outputs(3581) <= (inputs(74)) or (inputs(188));
    layer0_outputs(3582) <= (inputs(142)) or (inputs(158));
    layer0_outputs(3583) <= inputs(202);
    layer0_outputs(3584) <= (inputs(198)) xor (inputs(253));
    layer0_outputs(3585) <= not(inputs(41));
    layer0_outputs(3586) <= inputs(219);
    layer0_outputs(3587) <= not((inputs(197)) or (inputs(191)));
    layer0_outputs(3588) <= inputs(192);
    layer0_outputs(3589) <= (inputs(245)) and not (inputs(162));
    layer0_outputs(3590) <= not(inputs(44)) or (inputs(73));
    layer0_outputs(3591) <= inputs(151);
    layer0_outputs(3592) <= '1';
    layer0_outputs(3593) <= (inputs(230)) xor (inputs(47));
    layer0_outputs(3594) <= (inputs(51)) or (inputs(193));
    layer0_outputs(3595) <= inputs(227);
    layer0_outputs(3596) <= (inputs(201)) and (inputs(55));
    layer0_outputs(3597) <= (inputs(235)) and not (inputs(234));
    layer0_outputs(3598) <= (inputs(151)) and not (inputs(249));
    layer0_outputs(3599) <= (inputs(139)) and not (inputs(45));
    layer0_outputs(3600) <= inputs(59);
    layer0_outputs(3601) <= (inputs(171)) xor (inputs(112));
    layer0_outputs(3602) <= (inputs(74)) and not (inputs(92));
    layer0_outputs(3603) <= (inputs(25)) or (inputs(2));
    layer0_outputs(3604) <= not((inputs(44)) and (inputs(120)));
    layer0_outputs(3605) <= not(inputs(163));
    layer0_outputs(3606) <= not((inputs(34)) xor (inputs(188)));
    layer0_outputs(3607) <= not(inputs(84));
    layer0_outputs(3608) <= not(inputs(221)) or (inputs(172));
    layer0_outputs(3609) <= (inputs(200)) xor (inputs(33));
    layer0_outputs(3610) <= not((inputs(65)) or (inputs(184)));
    layer0_outputs(3611) <= not((inputs(191)) or (inputs(106)));
    layer0_outputs(3612) <= (inputs(76)) or (inputs(61));
    layer0_outputs(3613) <= not(inputs(113));
    layer0_outputs(3614) <= '1';
    layer0_outputs(3615) <= not(inputs(55));
    layer0_outputs(3616) <= (inputs(76)) and not (inputs(157));
    layer0_outputs(3617) <= not((inputs(120)) or (inputs(94)));
    layer0_outputs(3618) <= (inputs(186)) or (inputs(49));
    layer0_outputs(3619) <= inputs(210);
    layer0_outputs(3620) <= (inputs(133)) or (inputs(85));
    layer0_outputs(3621) <= not((inputs(102)) or (inputs(44)));
    layer0_outputs(3622) <= not(inputs(215));
    layer0_outputs(3623) <= not((inputs(190)) or (inputs(164)));
    layer0_outputs(3624) <= not(inputs(117)) or (inputs(143));
    layer0_outputs(3625) <= '0';
    layer0_outputs(3626) <= not((inputs(24)) and (inputs(108)));
    layer0_outputs(3627) <= (inputs(34)) or (inputs(71));
    layer0_outputs(3628) <= inputs(73);
    layer0_outputs(3629) <= not((inputs(201)) or (inputs(209)));
    layer0_outputs(3630) <= (inputs(219)) and not (inputs(56));
    layer0_outputs(3631) <= (inputs(104)) or (inputs(22));
    layer0_outputs(3632) <= (inputs(5)) xor (inputs(161));
    layer0_outputs(3633) <= not((inputs(244)) or (inputs(222)));
    layer0_outputs(3634) <= (inputs(110)) xor (inputs(108));
    layer0_outputs(3635) <= (inputs(215)) or (inputs(223));
    layer0_outputs(3636) <= not(inputs(93)) or (inputs(174));
    layer0_outputs(3637) <= not(inputs(95));
    layer0_outputs(3638) <= inputs(252);
    layer0_outputs(3639) <= not(inputs(198)) or (inputs(122));
    layer0_outputs(3640) <= not((inputs(47)) xor (inputs(202)));
    layer0_outputs(3641) <= inputs(235);
    layer0_outputs(3642) <= not((inputs(205)) or (inputs(81)));
    layer0_outputs(3643) <= not(inputs(221));
    layer0_outputs(3644) <= not(inputs(14));
    layer0_outputs(3645) <= inputs(182);
    layer0_outputs(3646) <= (inputs(236)) and not (inputs(96));
    layer0_outputs(3647) <= not(inputs(153));
    layer0_outputs(3648) <= not(inputs(229));
    layer0_outputs(3649) <= not(inputs(82));
    layer0_outputs(3650) <= (inputs(138)) or (inputs(132));
    layer0_outputs(3651) <= not(inputs(202)) or (inputs(29));
    layer0_outputs(3652) <= (inputs(159)) or (inputs(59));
    layer0_outputs(3653) <= not((inputs(125)) or (inputs(49)));
    layer0_outputs(3654) <= '0';
    layer0_outputs(3655) <= (inputs(213)) or (inputs(173));
    layer0_outputs(3656) <= '1';
    layer0_outputs(3657) <= (inputs(195)) xor (inputs(146));
    layer0_outputs(3658) <= (inputs(125)) xor (inputs(181));
    layer0_outputs(3659) <= (inputs(43)) and not (inputs(204));
    layer0_outputs(3660) <= (inputs(2)) and (inputs(58));
    layer0_outputs(3661) <= (inputs(21)) and not (inputs(221));
    layer0_outputs(3662) <= (inputs(187)) or (inputs(155));
    layer0_outputs(3663) <= inputs(231);
    layer0_outputs(3664) <= inputs(208);
    layer0_outputs(3665) <= not(inputs(188));
    layer0_outputs(3666) <= (inputs(241)) and not (inputs(198));
    layer0_outputs(3667) <= '1';
    layer0_outputs(3668) <= (inputs(14)) and not (inputs(161));
    layer0_outputs(3669) <= not(inputs(21));
    layer0_outputs(3670) <= (inputs(181)) and not (inputs(97));
    layer0_outputs(3671) <= inputs(204);
    layer0_outputs(3672) <= not(inputs(158)) or (inputs(221));
    layer0_outputs(3673) <= (inputs(254)) xor (inputs(154));
    layer0_outputs(3674) <= not((inputs(220)) or (inputs(210)));
    layer0_outputs(3675) <= not(inputs(244)) or (inputs(198));
    layer0_outputs(3676) <= (inputs(140)) xor (inputs(244));
    layer0_outputs(3677) <= (inputs(10)) or (inputs(244));
    layer0_outputs(3678) <= (inputs(75)) and not (inputs(157));
    layer0_outputs(3679) <= not((inputs(227)) or (inputs(214)));
    layer0_outputs(3680) <= inputs(19);
    layer0_outputs(3681) <= (inputs(24)) and not (inputs(173));
    layer0_outputs(3682) <= (inputs(109)) and not (inputs(129));
    layer0_outputs(3683) <= inputs(140);
    layer0_outputs(3684) <= not((inputs(114)) or (inputs(57)));
    layer0_outputs(3685) <= not(inputs(158));
    layer0_outputs(3686) <= (inputs(46)) and not (inputs(1));
    layer0_outputs(3687) <= (inputs(70)) and (inputs(86));
    layer0_outputs(3688) <= inputs(64);
    layer0_outputs(3689) <= inputs(195);
    layer0_outputs(3690) <= (inputs(124)) and not (inputs(221));
    layer0_outputs(3691) <= '0';
    layer0_outputs(3692) <= not(inputs(32)) or (inputs(1));
    layer0_outputs(3693) <= (inputs(102)) and not (inputs(59));
    layer0_outputs(3694) <= (inputs(167)) or (inputs(166));
    layer0_outputs(3695) <= not((inputs(173)) xor (inputs(80)));
    layer0_outputs(3696) <= (inputs(224)) or (inputs(39));
    layer0_outputs(3697) <= '0';
    layer0_outputs(3698) <= (inputs(112)) xor (inputs(85));
    layer0_outputs(3699) <= (inputs(99)) or (inputs(176));
    layer0_outputs(3700) <= (inputs(69)) or (inputs(192));
    layer0_outputs(3701) <= not((inputs(205)) or (inputs(226)));
    layer0_outputs(3702) <= not((inputs(138)) or (inputs(166)));
    layer0_outputs(3703) <= (inputs(146)) and (inputs(173));
    layer0_outputs(3704) <= (inputs(55)) xor (inputs(23));
    layer0_outputs(3705) <= not(inputs(122));
    layer0_outputs(3706) <= not(inputs(3));
    layer0_outputs(3707) <= not(inputs(237)) or (inputs(200));
    layer0_outputs(3708) <= not(inputs(184));
    layer0_outputs(3709) <= (inputs(33)) or (inputs(206));
    layer0_outputs(3710) <= (inputs(125)) or (inputs(36));
    layer0_outputs(3711) <= (inputs(185)) or (inputs(210));
    layer0_outputs(3712) <= not((inputs(116)) xor (inputs(210)));
    layer0_outputs(3713) <= inputs(102);
    layer0_outputs(3714) <= inputs(17);
    layer0_outputs(3715) <= not(inputs(12));
    layer0_outputs(3716) <= not(inputs(73));
    layer0_outputs(3717) <= not(inputs(137));
    layer0_outputs(3718) <= not((inputs(0)) or (inputs(254)));
    layer0_outputs(3719) <= inputs(54);
    layer0_outputs(3720) <= (inputs(62)) and not (inputs(126));
    layer0_outputs(3721) <= not(inputs(236));
    layer0_outputs(3722) <= (inputs(169)) and not (inputs(22));
    layer0_outputs(3723) <= (inputs(40)) and not (inputs(252));
    layer0_outputs(3724) <= not(inputs(0)) or (inputs(14));
    layer0_outputs(3725) <= (inputs(72)) xor (inputs(17));
    layer0_outputs(3726) <= not((inputs(175)) or (inputs(221)));
    layer0_outputs(3727) <= inputs(212);
    layer0_outputs(3728) <= inputs(130);
    layer0_outputs(3729) <= not((inputs(186)) or (inputs(4)));
    layer0_outputs(3730) <= (inputs(171)) xor (inputs(150));
    layer0_outputs(3731) <= (inputs(223)) or (inputs(218));
    layer0_outputs(3732) <= (inputs(238)) or (inputs(18));
    layer0_outputs(3733) <= not((inputs(207)) or (inputs(237)));
    layer0_outputs(3734) <= (inputs(127)) or (inputs(114));
    layer0_outputs(3735) <= not(inputs(240));
    layer0_outputs(3736) <= '0';
    layer0_outputs(3737) <= (inputs(6)) or (inputs(110));
    layer0_outputs(3738) <= not(inputs(31));
    layer0_outputs(3739) <= (inputs(196)) and not (inputs(90));
    layer0_outputs(3740) <= (inputs(59)) or (inputs(194));
    layer0_outputs(3741) <= not(inputs(113));
    layer0_outputs(3742) <= (inputs(58)) and not (inputs(111));
    layer0_outputs(3743) <= (inputs(196)) or (inputs(127));
    layer0_outputs(3744) <= (inputs(255)) and not (inputs(164));
    layer0_outputs(3745) <= not(inputs(83)) or (inputs(238));
    layer0_outputs(3746) <= '0';
    layer0_outputs(3747) <= (inputs(36)) and (inputs(149));
    layer0_outputs(3748) <= not(inputs(211));
    layer0_outputs(3749) <= (inputs(184)) and not (inputs(122));
    layer0_outputs(3750) <= not(inputs(255)) or (inputs(138));
    layer0_outputs(3751) <= inputs(229);
    layer0_outputs(3752) <= (inputs(234)) xor (inputs(128));
    layer0_outputs(3753) <= not(inputs(181));
    layer0_outputs(3754) <= (inputs(90)) and not (inputs(86));
    layer0_outputs(3755) <= (inputs(145)) and not (inputs(147));
    layer0_outputs(3756) <= not(inputs(171));
    layer0_outputs(3757) <= not(inputs(157)) or (inputs(239));
    layer0_outputs(3758) <= not(inputs(99));
    layer0_outputs(3759) <= inputs(123);
    layer0_outputs(3760) <= (inputs(189)) or (inputs(190));
    layer0_outputs(3761) <= not(inputs(140)) or (inputs(41));
    layer0_outputs(3762) <= not(inputs(14));
    layer0_outputs(3763) <= inputs(248);
    layer0_outputs(3764) <= not((inputs(224)) or (inputs(35)));
    layer0_outputs(3765) <= not((inputs(35)) and (inputs(248)));
    layer0_outputs(3766) <= not((inputs(160)) or (inputs(143)));
    layer0_outputs(3767) <= not((inputs(17)) xor (inputs(111)));
    layer0_outputs(3768) <= not((inputs(171)) or (inputs(193)));
    layer0_outputs(3769) <= (inputs(247)) and not (inputs(240));
    layer0_outputs(3770) <= inputs(1);
    layer0_outputs(3771) <= '1';
    layer0_outputs(3772) <= inputs(170);
    layer0_outputs(3773) <= (inputs(236)) or (inputs(18));
    layer0_outputs(3774) <= not(inputs(67)) or (inputs(138));
    layer0_outputs(3775) <= inputs(193);
    layer0_outputs(3776) <= not(inputs(233)) or (inputs(251));
    layer0_outputs(3777) <= (inputs(227)) and not (inputs(91));
    layer0_outputs(3778) <= (inputs(119)) and not (inputs(156));
    layer0_outputs(3779) <= (inputs(253)) or (inputs(237));
    layer0_outputs(3780) <= not(inputs(2)) or (inputs(222));
    layer0_outputs(3781) <= not(inputs(164));
    layer0_outputs(3782) <= not(inputs(9)) or (inputs(205));
    layer0_outputs(3783) <= inputs(225);
    layer0_outputs(3784) <= not(inputs(104));
    layer0_outputs(3785) <= inputs(37);
    layer0_outputs(3786) <= not((inputs(174)) or (inputs(6)));
    layer0_outputs(3787) <= inputs(24);
    layer0_outputs(3788) <= not((inputs(29)) xor (inputs(65)));
    layer0_outputs(3789) <= inputs(17);
    layer0_outputs(3790) <= inputs(206);
    layer0_outputs(3791) <= not((inputs(243)) or (inputs(58)));
    layer0_outputs(3792) <= '1';
    layer0_outputs(3793) <= (inputs(216)) and not (inputs(0));
    layer0_outputs(3794) <= not(inputs(60));
    layer0_outputs(3795) <= (inputs(245)) or (inputs(199));
    layer0_outputs(3796) <= (inputs(116)) or (inputs(30));
    layer0_outputs(3797) <= '0';
    layer0_outputs(3798) <= '1';
    layer0_outputs(3799) <= '1';
    layer0_outputs(3800) <= not((inputs(132)) or (inputs(115)));
    layer0_outputs(3801) <= (inputs(100)) and not (inputs(78));
    layer0_outputs(3802) <= not((inputs(195)) or (inputs(143)));
    layer0_outputs(3803) <= not(inputs(121));
    layer0_outputs(3804) <= (inputs(132)) or (inputs(202));
    layer0_outputs(3805) <= (inputs(117)) and not (inputs(178));
    layer0_outputs(3806) <= (inputs(6)) and not (inputs(242));
    layer0_outputs(3807) <= '1';
    layer0_outputs(3808) <= (inputs(167)) and not (inputs(170));
    layer0_outputs(3809) <= (inputs(77)) or (inputs(132));
    layer0_outputs(3810) <= not((inputs(64)) or (inputs(218)));
    layer0_outputs(3811) <= (inputs(180)) and not (inputs(45));
    layer0_outputs(3812) <= (inputs(40)) or (inputs(69));
    layer0_outputs(3813) <= inputs(93);
    layer0_outputs(3814) <= (inputs(119)) xor (inputs(14));
    layer0_outputs(3815) <= not(inputs(54)) or (inputs(79));
    layer0_outputs(3816) <= (inputs(193)) or (inputs(156));
    layer0_outputs(3817) <= not(inputs(179)) or (inputs(149));
    layer0_outputs(3818) <= not((inputs(120)) or (inputs(252)));
    layer0_outputs(3819) <= (inputs(186)) or (inputs(205));
    layer0_outputs(3820) <= '1';
    layer0_outputs(3821) <= (inputs(39)) and not (inputs(175));
    layer0_outputs(3822) <= inputs(21);
    layer0_outputs(3823) <= inputs(73);
    layer0_outputs(3824) <= (inputs(47)) and (inputs(252));
    layer0_outputs(3825) <= inputs(210);
    layer0_outputs(3826) <= not((inputs(241)) or (inputs(174)));
    layer0_outputs(3827) <= (inputs(12)) and (inputs(41));
    layer0_outputs(3828) <= not(inputs(103));
    layer0_outputs(3829) <= not((inputs(64)) xor (inputs(34)));
    layer0_outputs(3830) <= inputs(97);
    layer0_outputs(3831) <= inputs(177);
    layer0_outputs(3832) <= not(inputs(204));
    layer0_outputs(3833) <= not(inputs(163));
    layer0_outputs(3834) <= not((inputs(40)) or (inputs(177)));
    layer0_outputs(3835) <= (inputs(101)) and (inputs(235));
    layer0_outputs(3836) <= inputs(136);
    layer0_outputs(3837) <= inputs(101);
    layer0_outputs(3838) <= (inputs(215)) xor (inputs(48));
    layer0_outputs(3839) <= inputs(92);
    layer0_outputs(3840) <= not((inputs(23)) xor (inputs(202)));
    layer0_outputs(3841) <= not((inputs(186)) or (inputs(68)));
    layer0_outputs(3842) <= inputs(176);
    layer0_outputs(3843) <= (inputs(161)) or (inputs(204));
    layer0_outputs(3844) <= not((inputs(133)) or (inputs(75)));
    layer0_outputs(3845) <= (inputs(49)) xor (inputs(65));
    layer0_outputs(3846) <= not((inputs(222)) xor (inputs(92)));
    layer0_outputs(3847) <= not(inputs(41));
    layer0_outputs(3848) <= (inputs(95)) or (inputs(228));
    layer0_outputs(3849) <= not((inputs(140)) or (inputs(129)));
    layer0_outputs(3850) <= (inputs(141)) or (inputs(186));
    layer0_outputs(3851) <= not((inputs(160)) xor (inputs(112)));
    layer0_outputs(3852) <= not(inputs(11));
    layer0_outputs(3853) <= (inputs(170)) and not (inputs(131));
    layer0_outputs(3854) <= not(inputs(255));
    layer0_outputs(3855) <= not(inputs(144)) or (inputs(45));
    layer0_outputs(3856) <= not((inputs(99)) xor (inputs(207)));
    layer0_outputs(3857) <= not((inputs(192)) xor (inputs(143)));
    layer0_outputs(3858) <= inputs(203);
    layer0_outputs(3859) <= inputs(118);
    layer0_outputs(3860) <= '1';
    layer0_outputs(3861) <= (inputs(118)) or (inputs(103));
    layer0_outputs(3862) <= inputs(199);
    layer0_outputs(3863) <= not((inputs(117)) or (inputs(124)));
    layer0_outputs(3864) <= '0';
    layer0_outputs(3865) <= inputs(199);
    layer0_outputs(3866) <= not(inputs(181)) or (inputs(158));
    layer0_outputs(3867) <= not((inputs(229)) and (inputs(93)));
    layer0_outputs(3868) <= inputs(172);
    layer0_outputs(3869) <= not(inputs(145));
    layer0_outputs(3870) <= not(inputs(54)) or (inputs(156));
    layer0_outputs(3871) <= inputs(211);
    layer0_outputs(3872) <= not((inputs(109)) or (inputs(155)));
    layer0_outputs(3873) <= (inputs(172)) and not (inputs(2));
    layer0_outputs(3874) <= '0';
    layer0_outputs(3875) <= (inputs(143)) or (inputs(79));
    layer0_outputs(3876) <= not(inputs(80));
    layer0_outputs(3877) <= not(inputs(102));
    layer0_outputs(3878) <= inputs(117);
    layer0_outputs(3879) <= (inputs(109)) xor (inputs(18));
    layer0_outputs(3880) <= (inputs(9)) and not (inputs(243));
    layer0_outputs(3881) <= not((inputs(121)) or (inputs(76)));
    layer0_outputs(3882) <= not(inputs(200));
    layer0_outputs(3883) <= inputs(153);
    layer0_outputs(3884) <= not((inputs(27)) and (inputs(112)));
    layer0_outputs(3885) <= '0';
    layer0_outputs(3886) <= inputs(59);
    layer0_outputs(3887) <= not((inputs(238)) or (inputs(218)));
    layer0_outputs(3888) <= (inputs(3)) and not (inputs(196));
    layer0_outputs(3889) <= not(inputs(199));
    layer0_outputs(3890) <= inputs(164);
    layer0_outputs(3891) <= not((inputs(210)) xor (inputs(176)));
    layer0_outputs(3892) <= (inputs(253)) and not (inputs(174));
    layer0_outputs(3893) <= not((inputs(250)) or (inputs(229)));
    layer0_outputs(3894) <= (inputs(23)) xor (inputs(130));
    layer0_outputs(3895) <= not((inputs(221)) or (inputs(7)));
    layer0_outputs(3896) <= inputs(51);
    layer0_outputs(3897) <= not((inputs(160)) or (inputs(33)));
    layer0_outputs(3898) <= (inputs(144)) and not (inputs(74));
    layer0_outputs(3899) <= '1';
    layer0_outputs(3900) <= not((inputs(60)) or (inputs(155)));
    layer0_outputs(3901) <= '0';
    layer0_outputs(3902) <= not((inputs(146)) or (inputs(9)));
    layer0_outputs(3903) <= inputs(131);
    layer0_outputs(3904) <= (inputs(189)) and not (inputs(15));
    layer0_outputs(3905) <= not(inputs(101)) or (inputs(239));
    layer0_outputs(3906) <= '0';
    layer0_outputs(3907) <= (inputs(255)) or (inputs(159));
    layer0_outputs(3908) <= not(inputs(238));
    layer0_outputs(3909) <= '0';
    layer0_outputs(3910) <= (inputs(142)) or (inputs(195));
    layer0_outputs(3911) <= inputs(24);
    layer0_outputs(3912) <= not(inputs(70));
    layer0_outputs(3913) <= not(inputs(32)) or (inputs(163));
    layer0_outputs(3914) <= not(inputs(26));
    layer0_outputs(3915) <= not(inputs(246)) or (inputs(15));
    layer0_outputs(3916) <= (inputs(60)) or (inputs(247));
    layer0_outputs(3917) <= (inputs(144)) and (inputs(46));
    layer0_outputs(3918) <= inputs(108);
    layer0_outputs(3919) <= not(inputs(73)) or (inputs(228));
    layer0_outputs(3920) <= not((inputs(135)) and (inputs(199)));
    layer0_outputs(3921) <= (inputs(140)) and not (inputs(250));
    layer0_outputs(3922) <= (inputs(216)) xor (inputs(7));
    layer0_outputs(3923) <= inputs(56);
    layer0_outputs(3924) <= not(inputs(101));
    layer0_outputs(3925) <= not((inputs(224)) or (inputs(210)));
    layer0_outputs(3926) <= (inputs(171)) or (inputs(128));
    layer0_outputs(3927) <= not(inputs(197));
    layer0_outputs(3928) <= not((inputs(254)) or (inputs(134)));
    layer0_outputs(3929) <= '0';
    layer0_outputs(3930) <= not((inputs(83)) or (inputs(220)));
    layer0_outputs(3931) <= inputs(173);
    layer0_outputs(3932) <= inputs(185);
    layer0_outputs(3933) <= not(inputs(131)) or (inputs(192));
    layer0_outputs(3934) <= (inputs(74)) and not (inputs(248));
    layer0_outputs(3935) <= not(inputs(248));
    layer0_outputs(3936) <= (inputs(230)) and not (inputs(3));
    layer0_outputs(3937) <= not(inputs(114));
    layer0_outputs(3938) <= (inputs(221)) or (inputs(130));
    layer0_outputs(3939) <= not((inputs(77)) or (inputs(129)));
    layer0_outputs(3940) <= not(inputs(61));
    layer0_outputs(3941) <= not(inputs(229));
    layer0_outputs(3942) <= (inputs(30)) or (inputs(209));
    layer0_outputs(3943) <= (inputs(151)) and not (inputs(247));
    layer0_outputs(3944) <= not(inputs(139)) or (inputs(97));
    layer0_outputs(3945) <= not(inputs(85));
    layer0_outputs(3946) <= not((inputs(202)) or (inputs(204)));
    layer0_outputs(3947) <= (inputs(72)) and not (inputs(48));
    layer0_outputs(3948) <= (inputs(52)) or (inputs(208));
    layer0_outputs(3949) <= not((inputs(111)) xor (inputs(166)));
    layer0_outputs(3950) <= not(inputs(41)) or (inputs(88));
    layer0_outputs(3951) <= not((inputs(141)) or (inputs(153)));
    layer0_outputs(3952) <= not(inputs(115));
    layer0_outputs(3953) <= (inputs(72)) and not (inputs(162));
    layer0_outputs(3954) <= '0';
    layer0_outputs(3955) <= inputs(57);
    layer0_outputs(3956) <= not((inputs(124)) or (inputs(42)));
    layer0_outputs(3957) <= not((inputs(97)) xor (inputs(49)));
    layer0_outputs(3958) <= not(inputs(88)) or (inputs(31));
    layer0_outputs(3959) <= (inputs(112)) or (inputs(196));
    layer0_outputs(3960) <= (inputs(211)) and not (inputs(17));
    layer0_outputs(3961) <= not(inputs(28)) or (inputs(12));
    layer0_outputs(3962) <= not(inputs(74)) or (inputs(143));
    layer0_outputs(3963) <= not(inputs(30));
    layer0_outputs(3964) <= not((inputs(53)) or (inputs(196)));
    layer0_outputs(3965) <= (inputs(43)) and not (inputs(236));
    layer0_outputs(3966) <= (inputs(198)) and not (inputs(234));
    layer0_outputs(3967) <= not(inputs(104)) or (inputs(53));
    layer0_outputs(3968) <= '0';
    layer0_outputs(3969) <= not((inputs(180)) and (inputs(46)));
    layer0_outputs(3970) <= not((inputs(206)) or (inputs(175)));
    layer0_outputs(3971) <= not(inputs(72));
    layer0_outputs(3972) <= not(inputs(162));
    layer0_outputs(3973) <= not((inputs(210)) or (inputs(76)));
    layer0_outputs(3974) <= not(inputs(115)) or (inputs(207));
    layer0_outputs(3975) <= not((inputs(164)) or (inputs(195)));
    layer0_outputs(3976) <= (inputs(167)) and (inputs(67));
    layer0_outputs(3977) <= (inputs(202)) and not (inputs(197));
    layer0_outputs(3978) <= not(inputs(87));
    layer0_outputs(3979) <= not((inputs(146)) or (inputs(111)));
    layer0_outputs(3980) <= not((inputs(143)) or (inputs(58)));
    layer0_outputs(3981) <= (inputs(200)) or (inputs(24));
    layer0_outputs(3982) <= not(inputs(229));
    layer0_outputs(3983) <= (inputs(72)) and not (inputs(176));
    layer0_outputs(3984) <= (inputs(59)) and not (inputs(160));
    layer0_outputs(3985) <= not((inputs(248)) and (inputs(4)));
    layer0_outputs(3986) <= not(inputs(58)) or (inputs(217));
    layer0_outputs(3987) <= not(inputs(77)) or (inputs(112));
    layer0_outputs(3988) <= not((inputs(138)) and (inputs(127)));
    layer0_outputs(3989) <= not(inputs(220));
    layer0_outputs(3990) <= (inputs(115)) and not (inputs(213));
    layer0_outputs(3991) <= (inputs(223)) or (inputs(21));
    layer0_outputs(3992) <= (inputs(37)) xor (inputs(7));
    layer0_outputs(3993) <= not((inputs(75)) and (inputs(106)));
    layer0_outputs(3994) <= (inputs(215)) or (inputs(24));
    layer0_outputs(3995) <= not((inputs(5)) and (inputs(249)));
    layer0_outputs(3996) <= not((inputs(228)) or (inputs(64)));
    layer0_outputs(3997) <= (inputs(75)) and (inputs(27));
    layer0_outputs(3998) <= not(inputs(174));
    layer0_outputs(3999) <= not(inputs(149));
    layer0_outputs(4000) <= not(inputs(212)) or (inputs(71));
    layer0_outputs(4001) <= not(inputs(115));
    layer0_outputs(4002) <= not(inputs(122));
    layer0_outputs(4003) <= '0';
    layer0_outputs(4004) <= inputs(228);
    layer0_outputs(4005) <= not((inputs(97)) or (inputs(249)));
    layer0_outputs(4006) <= not(inputs(145));
    layer0_outputs(4007) <= not((inputs(60)) or (inputs(5)));
    layer0_outputs(4008) <= not((inputs(146)) or (inputs(147)));
    layer0_outputs(4009) <= not((inputs(247)) or (inputs(230)));
    layer0_outputs(4010) <= inputs(61);
    layer0_outputs(4011) <= not((inputs(137)) or (inputs(15)));
    layer0_outputs(4012) <= (inputs(197)) or (inputs(187));
    layer0_outputs(4013) <= (inputs(121)) and not (inputs(160));
    layer0_outputs(4014) <= (inputs(52)) and not (inputs(112));
    layer0_outputs(4015) <= inputs(61);
    layer0_outputs(4016) <= not(inputs(134));
    layer0_outputs(4017) <= '1';
    layer0_outputs(4018) <= (inputs(155)) xor (inputs(107));
    layer0_outputs(4019) <= not(inputs(42)) or (inputs(74));
    layer0_outputs(4020) <= not((inputs(39)) or (inputs(247)));
    layer0_outputs(4021) <= (inputs(152)) and not (inputs(190));
    layer0_outputs(4022) <= not(inputs(181)) or (inputs(78));
    layer0_outputs(4023) <= not((inputs(109)) xor (inputs(121)));
    layer0_outputs(4024) <= not(inputs(124)) or (inputs(231));
    layer0_outputs(4025) <= not(inputs(213)) or (inputs(222));
    layer0_outputs(4026) <= (inputs(188)) and not (inputs(28));
    layer0_outputs(4027) <= not(inputs(246));
    layer0_outputs(4028) <= inputs(80);
    layer0_outputs(4029) <= (inputs(78)) and not (inputs(98));
    layer0_outputs(4030) <= not(inputs(92));
    layer0_outputs(4031) <= not((inputs(15)) or (inputs(164)));
    layer0_outputs(4032) <= not(inputs(152));
    layer0_outputs(4033) <= (inputs(96)) and not (inputs(65));
    layer0_outputs(4034) <= (inputs(198)) or (inputs(137));
    layer0_outputs(4035) <= not(inputs(162)) or (inputs(149));
    layer0_outputs(4036) <= not(inputs(59));
    layer0_outputs(4037) <= not((inputs(213)) and (inputs(37)));
    layer0_outputs(4038) <= '1';
    layer0_outputs(4039) <= '1';
    layer0_outputs(4040) <= (inputs(130)) and (inputs(73));
    layer0_outputs(4041) <= not((inputs(9)) or (inputs(37)));
    layer0_outputs(4042) <= inputs(255);
    layer0_outputs(4043) <= (inputs(236)) xor (inputs(192));
    layer0_outputs(4044) <= (inputs(246)) and not (inputs(220));
    layer0_outputs(4045) <= inputs(18);
    layer0_outputs(4046) <= not(inputs(90));
    layer0_outputs(4047) <= (inputs(57)) xor (inputs(118));
    layer0_outputs(4048) <= not(inputs(24));
    layer0_outputs(4049) <= not((inputs(113)) xor (inputs(39)));
    layer0_outputs(4050) <= not(inputs(62)) or (inputs(125));
    layer0_outputs(4051) <= not(inputs(88)) or (inputs(91));
    layer0_outputs(4052) <= '1';
    layer0_outputs(4053) <= '0';
    layer0_outputs(4054) <= inputs(128);
    layer0_outputs(4055) <= not(inputs(128)) or (inputs(214));
    layer0_outputs(4056) <= (inputs(240)) or (inputs(194));
    layer0_outputs(4057) <= not((inputs(44)) or (inputs(31)));
    layer0_outputs(4058) <= not((inputs(231)) or (inputs(237)));
    layer0_outputs(4059) <= not(inputs(37));
    layer0_outputs(4060) <= not((inputs(65)) and (inputs(138)));
    layer0_outputs(4061) <= not(inputs(69)) or (inputs(4));
    layer0_outputs(4062) <= (inputs(148)) or (inputs(145));
    layer0_outputs(4063) <= not((inputs(152)) xor (inputs(43)));
    layer0_outputs(4064) <= not((inputs(35)) and (inputs(240)));
    layer0_outputs(4065) <= inputs(210);
    layer0_outputs(4066) <= (inputs(24)) xor (inputs(71));
    layer0_outputs(4067) <= not(inputs(101));
    layer0_outputs(4068) <= not(inputs(84));
    layer0_outputs(4069) <= (inputs(104)) or (inputs(254));
    layer0_outputs(4070) <= inputs(71);
    layer0_outputs(4071) <= (inputs(177)) and not (inputs(52));
    layer0_outputs(4072) <= not(inputs(203));
    layer0_outputs(4073) <= not((inputs(91)) and (inputs(76)));
    layer0_outputs(4074) <= inputs(178);
    layer0_outputs(4075) <= (inputs(140)) xor (inputs(171));
    layer0_outputs(4076) <= not(inputs(39)) or (inputs(46));
    layer0_outputs(4077) <= (inputs(96)) xor (inputs(229));
    layer0_outputs(4078) <= not((inputs(30)) or (inputs(154)));
    layer0_outputs(4079) <= not(inputs(212));
    layer0_outputs(4080) <= not((inputs(124)) or (inputs(145)));
    layer0_outputs(4081) <= not(inputs(19)) or (inputs(241));
    layer0_outputs(4082) <= inputs(121);
    layer0_outputs(4083) <= (inputs(230)) and not (inputs(61));
    layer0_outputs(4084) <= not((inputs(101)) xor (inputs(81)));
    layer0_outputs(4085) <= not((inputs(221)) and (inputs(234)));
    layer0_outputs(4086) <= inputs(236);
    layer0_outputs(4087) <= '0';
    layer0_outputs(4088) <= (inputs(87)) and not (inputs(4));
    layer0_outputs(4089) <= (inputs(162)) or (inputs(214));
    layer0_outputs(4090) <= (inputs(146)) xor (inputs(217));
    layer0_outputs(4091) <= not((inputs(151)) or (inputs(222)));
    layer0_outputs(4092) <= (inputs(99)) and not (inputs(235));
    layer0_outputs(4093) <= not(inputs(55));
    layer0_outputs(4094) <= '0';
    layer0_outputs(4095) <= (inputs(32)) or (inputs(163));
    layer0_outputs(4096) <= (inputs(147)) or (inputs(0));
    layer0_outputs(4097) <= '0';
    layer0_outputs(4098) <= (inputs(74)) xor (inputs(57));
    layer0_outputs(4099) <= not(inputs(2));
    layer0_outputs(4100) <= (inputs(83)) and not (inputs(179));
    layer0_outputs(4101) <= inputs(41);
    layer0_outputs(4102) <= not((inputs(37)) xor (inputs(45)));
    layer0_outputs(4103) <= not((inputs(111)) or (inputs(122)));
    layer0_outputs(4104) <= not(inputs(149));
    layer0_outputs(4105) <= not((inputs(82)) or (inputs(86)));
    layer0_outputs(4106) <= (inputs(199)) and not (inputs(145));
    layer0_outputs(4107) <= not((inputs(3)) or (inputs(6)));
    layer0_outputs(4108) <= not(inputs(57));
    layer0_outputs(4109) <= inputs(66);
    layer0_outputs(4110) <= not(inputs(103));
    layer0_outputs(4111) <= not(inputs(44));
    layer0_outputs(4112) <= (inputs(254)) or (inputs(22));
    layer0_outputs(4113) <= (inputs(57)) and (inputs(109));
    layer0_outputs(4114) <= not((inputs(217)) or (inputs(236)));
    layer0_outputs(4115) <= not(inputs(225)) or (inputs(124));
    layer0_outputs(4116) <= '1';
    layer0_outputs(4117) <= not(inputs(69)) or (inputs(187));
    layer0_outputs(4118) <= not(inputs(74));
    layer0_outputs(4119) <= (inputs(253)) or (inputs(53));
    layer0_outputs(4120) <= (inputs(163)) or (inputs(173));
    layer0_outputs(4121) <= (inputs(111)) or (inputs(100));
    layer0_outputs(4122) <= inputs(45);
    layer0_outputs(4123) <= (inputs(224)) and (inputs(65));
    layer0_outputs(4124) <= inputs(233);
    layer0_outputs(4125) <= not((inputs(96)) or (inputs(62)));
    layer0_outputs(4126) <= not((inputs(159)) xor (inputs(208)));
    layer0_outputs(4127) <= (inputs(185)) and not (inputs(157));
    layer0_outputs(4128) <= inputs(88);
    layer0_outputs(4129) <= not(inputs(24)) or (inputs(100));
    layer0_outputs(4130) <= not((inputs(189)) xor (inputs(14)));
    layer0_outputs(4131) <= not(inputs(67)) or (inputs(158));
    layer0_outputs(4132) <= not((inputs(109)) or (inputs(27)));
    layer0_outputs(4133) <= '1';
    layer0_outputs(4134) <= (inputs(43)) and (inputs(113));
    layer0_outputs(4135) <= (inputs(202)) or (inputs(37));
    layer0_outputs(4136) <= inputs(41);
    layer0_outputs(4137) <= (inputs(163)) or (inputs(85));
    layer0_outputs(4138) <= (inputs(240)) or (inputs(25));
    layer0_outputs(4139) <= (inputs(67)) and not (inputs(58));
    layer0_outputs(4140) <= (inputs(10)) or (inputs(189));
    layer0_outputs(4141) <= (inputs(111)) or (inputs(68));
    layer0_outputs(4142) <= '1';
    layer0_outputs(4143) <= not(inputs(181));
    layer0_outputs(4144) <= inputs(152);
    layer0_outputs(4145) <= not(inputs(80));
    layer0_outputs(4146) <= (inputs(127)) or (inputs(67));
    layer0_outputs(4147) <= inputs(146);
    layer0_outputs(4148) <= not(inputs(89)) or (inputs(195));
    layer0_outputs(4149) <= inputs(4);
    layer0_outputs(4150) <= (inputs(47)) or (inputs(11));
    layer0_outputs(4151) <= not(inputs(204)) or (inputs(113));
    layer0_outputs(4152) <= not(inputs(172));
    layer0_outputs(4153) <= not(inputs(8)) or (inputs(10));
    layer0_outputs(4154) <= not(inputs(185));
    layer0_outputs(4155) <= inputs(55);
    layer0_outputs(4156) <= '1';
    layer0_outputs(4157) <= not(inputs(151));
    layer0_outputs(4158) <= (inputs(119)) and not (inputs(15));
    layer0_outputs(4159) <= not(inputs(202));
    layer0_outputs(4160) <= (inputs(132)) xor (inputs(36));
    layer0_outputs(4161) <= inputs(245);
    layer0_outputs(4162) <= (inputs(73)) and not (inputs(151));
    layer0_outputs(4163) <= (inputs(144)) xor (inputs(230));
    layer0_outputs(4164) <= not(inputs(139));
    layer0_outputs(4165) <= (inputs(7)) and not (inputs(160));
    layer0_outputs(4166) <= not((inputs(141)) and (inputs(94)));
    layer0_outputs(4167) <= not(inputs(28)) or (inputs(175));
    layer0_outputs(4168) <= not(inputs(210)) or (inputs(8));
    layer0_outputs(4169) <= not((inputs(87)) xor (inputs(186)));
    layer0_outputs(4170) <= (inputs(164)) or (inputs(129));
    layer0_outputs(4171) <= not((inputs(8)) or (inputs(106)));
    layer0_outputs(4172) <= not((inputs(53)) or (inputs(166)));
    layer0_outputs(4173) <= not(inputs(217));
    layer0_outputs(4174) <= '1';
    layer0_outputs(4175) <= not(inputs(8)) or (inputs(219));
    layer0_outputs(4176) <= not(inputs(120)) or (inputs(146));
    layer0_outputs(4177) <= not(inputs(253));
    layer0_outputs(4178) <= inputs(21);
    layer0_outputs(4179) <= (inputs(20)) xor (inputs(77));
    layer0_outputs(4180) <= (inputs(179)) or (inputs(185));
    layer0_outputs(4181) <= (inputs(180)) and not (inputs(75));
    layer0_outputs(4182) <= (inputs(85)) and not (inputs(221));
    layer0_outputs(4183) <= not((inputs(220)) or (inputs(196)));
    layer0_outputs(4184) <= not((inputs(81)) xor (inputs(252)));
    layer0_outputs(4185) <= (inputs(15)) xor (inputs(45));
    layer0_outputs(4186) <= (inputs(132)) and not (inputs(0));
    layer0_outputs(4187) <= (inputs(68)) or (inputs(116));
    layer0_outputs(4188) <= not(inputs(66)) or (inputs(107));
    layer0_outputs(4189) <= not((inputs(164)) xor (inputs(111)));
    layer0_outputs(4190) <= not(inputs(0));
    layer0_outputs(4191) <= (inputs(152)) and not (inputs(129));
    layer0_outputs(4192) <= inputs(218);
    layer0_outputs(4193) <= (inputs(80)) and (inputs(198));
    layer0_outputs(4194) <= inputs(191);
    layer0_outputs(4195) <= '1';
    layer0_outputs(4196) <= not((inputs(75)) xor (inputs(197)));
    layer0_outputs(4197) <= (inputs(51)) xor (inputs(97));
    layer0_outputs(4198) <= (inputs(88)) and not (inputs(196));
    layer0_outputs(4199) <= not(inputs(168));
    layer0_outputs(4200) <= (inputs(135)) and not (inputs(35));
    layer0_outputs(4201) <= '1';
    layer0_outputs(4202) <= (inputs(160)) and not (inputs(59));
    layer0_outputs(4203) <= inputs(82);
    layer0_outputs(4204) <= (inputs(214)) or (inputs(162));
    layer0_outputs(4205) <= '0';
    layer0_outputs(4206) <= inputs(108);
    layer0_outputs(4207) <= inputs(253);
    layer0_outputs(4208) <= inputs(145);
    layer0_outputs(4209) <= not(inputs(141));
    layer0_outputs(4210) <= not(inputs(170)) or (inputs(97));
    layer0_outputs(4211) <= not(inputs(107));
    layer0_outputs(4212) <= '1';
    layer0_outputs(4213) <= not((inputs(96)) or (inputs(50)));
    layer0_outputs(4214) <= not((inputs(227)) or (inputs(228)));
    layer0_outputs(4215) <= not((inputs(125)) or (inputs(139)));
    layer0_outputs(4216) <= (inputs(30)) and not (inputs(19));
    layer0_outputs(4217) <= '1';
    layer0_outputs(4218) <= (inputs(117)) and not (inputs(245));
    layer0_outputs(4219) <= not(inputs(78)) or (inputs(205));
    layer0_outputs(4220) <= not(inputs(233)) or (inputs(48));
    layer0_outputs(4221) <= (inputs(111)) or (inputs(23));
    layer0_outputs(4222) <= not(inputs(202));
    layer0_outputs(4223) <= inputs(225);
    layer0_outputs(4224) <= (inputs(226)) and not (inputs(1));
    layer0_outputs(4225) <= (inputs(192)) xor (inputs(11));
    layer0_outputs(4226) <= not(inputs(163)) or (inputs(62));
    layer0_outputs(4227) <= not((inputs(61)) xor (inputs(157)));
    layer0_outputs(4228) <= (inputs(201)) and (inputs(39));
    layer0_outputs(4229) <= not(inputs(248));
    layer0_outputs(4230) <= (inputs(102)) xor (inputs(132));
    layer0_outputs(4231) <= not(inputs(91)) or (inputs(235));
    layer0_outputs(4232) <= inputs(229);
    layer0_outputs(4233) <= inputs(154);
    layer0_outputs(4234) <= (inputs(202)) and not (inputs(79));
    layer0_outputs(4235) <= (inputs(120)) and not (inputs(47));
    layer0_outputs(4236) <= not(inputs(140)) or (inputs(214));
    layer0_outputs(4237) <= not(inputs(158));
    layer0_outputs(4238) <= '0';
    layer0_outputs(4239) <= not(inputs(130)) or (inputs(240));
    layer0_outputs(4240) <= (inputs(99)) and (inputs(131));
    layer0_outputs(4241) <= not(inputs(182));
    layer0_outputs(4242) <= not(inputs(137));
    layer0_outputs(4243) <= not((inputs(28)) xor (inputs(229)));
    layer0_outputs(4244) <= (inputs(175)) xor (inputs(167));
    layer0_outputs(4245) <= inputs(105);
    layer0_outputs(4246) <= not((inputs(174)) or (inputs(80)));
    layer0_outputs(4247) <= (inputs(40)) or (inputs(149));
    layer0_outputs(4248) <= inputs(193);
    layer0_outputs(4249) <= '0';
    layer0_outputs(4250) <= inputs(44);
    layer0_outputs(4251) <= not(inputs(106)) or (inputs(69));
    layer0_outputs(4252) <= not((inputs(76)) or (inputs(123)));
    layer0_outputs(4253) <= not(inputs(193));
    layer0_outputs(4254) <= (inputs(75)) and (inputs(15));
    layer0_outputs(4255) <= (inputs(40)) and not (inputs(146));
    layer0_outputs(4256) <= not(inputs(26)) or (inputs(114));
    layer0_outputs(4257) <= (inputs(157)) or (inputs(71));
    layer0_outputs(4258) <= not(inputs(165)) or (inputs(120));
    layer0_outputs(4259) <= (inputs(235)) and (inputs(6));
    layer0_outputs(4260) <= inputs(195);
    layer0_outputs(4261) <= inputs(122);
    layer0_outputs(4262) <= not(inputs(7)) or (inputs(144));
    layer0_outputs(4263) <= not(inputs(215)) or (inputs(44));
    layer0_outputs(4264) <= not(inputs(57));
    layer0_outputs(4265) <= not(inputs(97));
    layer0_outputs(4266) <= inputs(137);
    layer0_outputs(4267) <= (inputs(195)) xor (inputs(0));
    layer0_outputs(4268) <= not((inputs(176)) or (inputs(140)));
    layer0_outputs(4269) <= not(inputs(200)) or (inputs(159));
    layer0_outputs(4270) <= not(inputs(73));
    layer0_outputs(4271) <= not(inputs(235)) or (inputs(56));
    layer0_outputs(4272) <= (inputs(119)) and not (inputs(35));
    layer0_outputs(4273) <= (inputs(154)) and not (inputs(30));
    layer0_outputs(4274) <= not((inputs(86)) or (inputs(94)));
    layer0_outputs(4275) <= (inputs(234)) or (inputs(54));
    layer0_outputs(4276) <= not(inputs(217)) or (inputs(82));
    layer0_outputs(4277) <= not((inputs(113)) or (inputs(244)));
    layer0_outputs(4278) <= inputs(210);
    layer0_outputs(4279) <= (inputs(152)) or (inputs(84));
    layer0_outputs(4280) <= not(inputs(126)) or (inputs(17));
    layer0_outputs(4281) <= '0';
    layer0_outputs(4282) <= not((inputs(38)) or (inputs(49)));
    layer0_outputs(4283) <= not(inputs(198)) or (inputs(117));
    layer0_outputs(4284) <= (inputs(66)) and not (inputs(49));
    layer0_outputs(4285) <= (inputs(200)) or (inputs(180));
    layer0_outputs(4286) <= (inputs(142)) or (inputs(195));
    layer0_outputs(4287) <= not((inputs(24)) xor (inputs(177)));
    layer0_outputs(4288) <= not((inputs(199)) xor (inputs(152)));
    layer0_outputs(4289) <= not(inputs(35));
    layer0_outputs(4290) <= (inputs(131)) or (inputs(15));
    layer0_outputs(4291) <= (inputs(182)) and not (inputs(211));
    layer0_outputs(4292) <= (inputs(116)) xor (inputs(87));
    layer0_outputs(4293) <= not(inputs(136));
    layer0_outputs(4294) <= (inputs(198)) and not (inputs(3));
    layer0_outputs(4295) <= not(inputs(187)) or (inputs(30));
    layer0_outputs(4296) <= inputs(217);
    layer0_outputs(4297) <= (inputs(219)) and not (inputs(87));
    layer0_outputs(4298) <= not(inputs(56));
    layer0_outputs(4299) <= not(inputs(38)) or (inputs(141));
    layer0_outputs(4300) <= not(inputs(69));
    layer0_outputs(4301) <= not(inputs(221));
    layer0_outputs(4302) <= (inputs(141)) or (inputs(92));
    layer0_outputs(4303) <= (inputs(53)) and not (inputs(190));
    layer0_outputs(4304) <= inputs(219);
    layer0_outputs(4305) <= not(inputs(178));
    layer0_outputs(4306) <= not((inputs(226)) or (inputs(62)));
    layer0_outputs(4307) <= (inputs(136)) and (inputs(218));
    layer0_outputs(4308) <= not((inputs(45)) or (inputs(79)));
    layer0_outputs(4309) <= not((inputs(207)) or (inputs(244)));
    layer0_outputs(4310) <= (inputs(181)) or (inputs(66));
    layer0_outputs(4311) <= inputs(4);
    layer0_outputs(4312) <= not(inputs(165));
    layer0_outputs(4313) <= inputs(167);
    layer0_outputs(4314) <= '1';
    layer0_outputs(4315) <= not(inputs(153));
    layer0_outputs(4316) <= not(inputs(166)) or (inputs(158));
    layer0_outputs(4317) <= not(inputs(194));
    layer0_outputs(4318) <= not(inputs(91)) or (inputs(5));
    layer0_outputs(4319) <= not(inputs(43));
    layer0_outputs(4320) <= not(inputs(94));
    layer0_outputs(4321) <= not((inputs(42)) or (inputs(51)));
    layer0_outputs(4322) <= not((inputs(235)) or (inputs(116)));
    layer0_outputs(4323) <= (inputs(105)) xor (inputs(160));
    layer0_outputs(4324) <= (inputs(87)) xor (inputs(236));
    layer0_outputs(4325) <= (inputs(22)) and not (inputs(5));
    layer0_outputs(4326) <= (inputs(188)) and not (inputs(61));
    layer0_outputs(4327) <= not((inputs(10)) xor (inputs(6)));
    layer0_outputs(4328) <= not(inputs(86)) or (inputs(251));
    layer0_outputs(4329) <= inputs(56);
    layer0_outputs(4330) <= (inputs(242)) or (inputs(236));
    layer0_outputs(4331) <= inputs(142);
    layer0_outputs(4332) <= not((inputs(93)) xor (inputs(255)));
    layer0_outputs(4333) <= (inputs(57)) or (inputs(195));
    layer0_outputs(4334) <= (inputs(229)) and not (inputs(111));
    layer0_outputs(4335) <= not((inputs(31)) or (inputs(197)));
    layer0_outputs(4336) <= not((inputs(228)) and (inputs(228)));
    layer0_outputs(4337) <= not((inputs(210)) xor (inputs(181)));
    layer0_outputs(4338) <= inputs(232);
    layer0_outputs(4339) <= not(inputs(112));
    layer0_outputs(4340) <= (inputs(247)) and not (inputs(121));
    layer0_outputs(4341) <= '0';
    layer0_outputs(4342) <= inputs(26);
    layer0_outputs(4343) <= not((inputs(217)) xor (inputs(188)));
    layer0_outputs(4344) <= not(inputs(232)) or (inputs(208));
    layer0_outputs(4345) <= not(inputs(55));
    layer0_outputs(4346) <= (inputs(26)) xor (inputs(37));
    layer0_outputs(4347) <= not((inputs(209)) and (inputs(130)));
    layer0_outputs(4348) <= inputs(27);
    layer0_outputs(4349) <= (inputs(209)) and not (inputs(80));
    layer0_outputs(4350) <= (inputs(252)) and not (inputs(107));
    layer0_outputs(4351) <= not(inputs(42)) or (inputs(100));
    layer0_outputs(4352) <= not((inputs(40)) or (inputs(48)));
    layer0_outputs(4353) <= inputs(49);
    layer0_outputs(4354) <= not((inputs(61)) or (inputs(45)));
    layer0_outputs(4355) <= (inputs(209)) or (inputs(76));
    layer0_outputs(4356) <= not((inputs(99)) or (inputs(192)));
    layer0_outputs(4357) <= not((inputs(30)) or (inputs(117)));
    layer0_outputs(4358) <= not((inputs(4)) or (inputs(187)));
    layer0_outputs(4359) <= not(inputs(106));
    layer0_outputs(4360) <= not(inputs(8));
    layer0_outputs(4361) <= (inputs(254)) or (inputs(132));
    layer0_outputs(4362) <= (inputs(101)) and not (inputs(243));
    layer0_outputs(4363) <= not(inputs(195));
    layer0_outputs(4364) <= not((inputs(189)) or (inputs(55)));
    layer0_outputs(4365) <= not(inputs(146)) or (inputs(5));
    layer0_outputs(4366) <= not((inputs(197)) xor (inputs(228)));
    layer0_outputs(4367) <= (inputs(143)) or (inputs(44));
    layer0_outputs(4368) <= (inputs(85)) and (inputs(74));
    layer0_outputs(4369) <= not(inputs(76)) or (inputs(64));
    layer0_outputs(4370) <= inputs(175);
    layer0_outputs(4371) <= (inputs(113)) or (inputs(98));
    layer0_outputs(4372) <= (inputs(62)) or (inputs(96));
    layer0_outputs(4373) <= not((inputs(40)) or (inputs(236)));
    layer0_outputs(4374) <= not(inputs(164)) or (inputs(64));
    layer0_outputs(4375) <= (inputs(140)) and not (inputs(239));
    layer0_outputs(4376) <= not(inputs(203)) or (inputs(1));
    layer0_outputs(4377) <= not((inputs(17)) and (inputs(143)));
    layer0_outputs(4378) <= (inputs(221)) xor (inputs(61));
    layer0_outputs(4379) <= not(inputs(105));
    layer0_outputs(4380) <= not((inputs(141)) or (inputs(3)));
    layer0_outputs(4381) <= not((inputs(32)) or (inputs(214)));
    layer0_outputs(4382) <= (inputs(251)) and not (inputs(200));
    layer0_outputs(4383) <= (inputs(246)) or (inputs(138));
    layer0_outputs(4384) <= (inputs(33)) or (inputs(4));
    layer0_outputs(4385) <= inputs(180);
    layer0_outputs(4386) <= (inputs(109)) or (inputs(234));
    layer0_outputs(4387) <= not((inputs(225)) or (inputs(199)));
    layer0_outputs(4388) <= not(inputs(132)) or (inputs(14));
    layer0_outputs(4389) <= not((inputs(63)) or (inputs(55)));
    layer0_outputs(4390) <= (inputs(160)) or (inputs(57));
    layer0_outputs(4391) <= (inputs(129)) or (inputs(3));
    layer0_outputs(4392) <= not(inputs(228)) or (inputs(14));
    layer0_outputs(4393) <= inputs(15);
    layer0_outputs(4394) <= (inputs(160)) or (inputs(37));
    layer0_outputs(4395) <= inputs(61);
    layer0_outputs(4396) <= inputs(175);
    layer0_outputs(4397) <= (inputs(136)) or (inputs(107));
    layer0_outputs(4398) <= not(inputs(21)) or (inputs(221));
    layer0_outputs(4399) <= inputs(119);
    layer0_outputs(4400) <= '0';
    layer0_outputs(4401) <= not(inputs(58)) or (inputs(136));
    layer0_outputs(4402) <= not(inputs(90)) or (inputs(209));
    layer0_outputs(4403) <= not((inputs(179)) and (inputs(191)));
    layer0_outputs(4404) <= inputs(94);
    layer0_outputs(4405) <= not(inputs(218));
    layer0_outputs(4406) <= not((inputs(64)) or (inputs(206)));
    layer0_outputs(4407) <= not((inputs(84)) xor (inputs(92)));
    layer0_outputs(4408) <= inputs(165);
    layer0_outputs(4409) <= not(inputs(203));
    layer0_outputs(4410) <= (inputs(54)) and not (inputs(227));
    layer0_outputs(4411) <= not((inputs(36)) and (inputs(216)));
    layer0_outputs(4412) <= not(inputs(12));
    layer0_outputs(4413) <= not(inputs(214)) or (inputs(105));
    layer0_outputs(4414) <= (inputs(14)) or (inputs(83));
    layer0_outputs(4415) <= (inputs(212)) and not (inputs(11));
    layer0_outputs(4416) <= (inputs(19)) and not (inputs(20));
    layer0_outputs(4417) <= not(inputs(184)) or (inputs(118));
    layer0_outputs(4418) <= inputs(183);
    layer0_outputs(4419) <= not(inputs(67));
    layer0_outputs(4420) <= not((inputs(86)) or (inputs(42)));
    layer0_outputs(4421) <= '1';
    layer0_outputs(4422) <= not(inputs(121)) or (inputs(252));
    layer0_outputs(4423) <= not((inputs(157)) or (inputs(249)));
    layer0_outputs(4424) <= not((inputs(45)) or (inputs(80)));
    layer0_outputs(4425) <= (inputs(8)) and (inputs(64));
    layer0_outputs(4426) <= not(inputs(183)) or (inputs(17));
    layer0_outputs(4427) <= '1';
    layer0_outputs(4428) <= (inputs(25)) and (inputs(58));
    layer0_outputs(4429) <= inputs(164);
    layer0_outputs(4430) <= (inputs(98)) and not (inputs(222));
    layer0_outputs(4431) <= (inputs(189)) and (inputs(97));
    layer0_outputs(4432) <= (inputs(197)) xor (inputs(130));
    layer0_outputs(4433) <= not(inputs(79)) or (inputs(87));
    layer0_outputs(4434) <= not((inputs(72)) or (inputs(231)));
    layer0_outputs(4435) <= not(inputs(53));
    layer0_outputs(4436) <= inputs(113);
    layer0_outputs(4437) <= not(inputs(25)) or (inputs(232));
    layer0_outputs(4438) <= inputs(182);
    layer0_outputs(4439) <= not(inputs(24));
    layer0_outputs(4440) <= not((inputs(104)) or (inputs(4)));
    layer0_outputs(4441) <= not((inputs(223)) xor (inputs(162)));
    layer0_outputs(4442) <= inputs(47);
    layer0_outputs(4443) <= (inputs(185)) and not (inputs(177));
    layer0_outputs(4444) <= (inputs(103)) and (inputs(119));
    layer0_outputs(4445) <= not(inputs(108));
    layer0_outputs(4446) <= inputs(181);
    layer0_outputs(4447) <= not((inputs(247)) or (inputs(168)));
    layer0_outputs(4448) <= not(inputs(213));
    layer0_outputs(4449) <= not((inputs(242)) and (inputs(21)));
    layer0_outputs(4450) <= not((inputs(69)) or (inputs(115)));
    layer0_outputs(4451) <= (inputs(219)) and not (inputs(62));
    layer0_outputs(4452) <= inputs(142);
    layer0_outputs(4453) <= not(inputs(110));
    layer0_outputs(4454) <= inputs(102);
    layer0_outputs(4455) <= not(inputs(21));
    layer0_outputs(4456) <= not((inputs(177)) or (inputs(6)));
    layer0_outputs(4457) <= not(inputs(239));
    layer0_outputs(4458) <= (inputs(137)) and not (inputs(213));
    layer0_outputs(4459) <= not((inputs(76)) or (inputs(93)));
    layer0_outputs(4460) <= (inputs(104)) and (inputs(112));
    layer0_outputs(4461) <= not(inputs(123));
    layer0_outputs(4462) <= not((inputs(82)) xor (inputs(69)));
    layer0_outputs(4463) <= (inputs(221)) or (inputs(20));
    layer0_outputs(4464) <= not((inputs(130)) xor (inputs(148)));
    layer0_outputs(4465) <= not(inputs(234));
    layer0_outputs(4466) <= inputs(44);
    layer0_outputs(4467) <= '0';
    layer0_outputs(4468) <= (inputs(49)) and not (inputs(166));
    layer0_outputs(4469) <= not((inputs(51)) or (inputs(163)));
    layer0_outputs(4470) <= (inputs(179)) and not (inputs(243));
    layer0_outputs(4471) <= not((inputs(27)) or (inputs(184)));
    layer0_outputs(4472) <= not((inputs(232)) or (inputs(216)));
    layer0_outputs(4473) <= not(inputs(136));
    layer0_outputs(4474) <= '1';
    layer0_outputs(4475) <= (inputs(27)) and not (inputs(242));
    layer0_outputs(4476) <= inputs(128);
    layer0_outputs(4477) <= not(inputs(119)) or (inputs(85));
    layer0_outputs(4478) <= (inputs(95)) and not (inputs(241));
    layer0_outputs(4479) <= (inputs(129)) or (inputs(236));
    layer0_outputs(4480) <= not((inputs(4)) or (inputs(225)));
    layer0_outputs(4481) <= not((inputs(123)) and (inputs(222)));
    layer0_outputs(4482) <= (inputs(66)) xor (inputs(77));
    layer0_outputs(4483) <= not(inputs(147)) or (inputs(135));
    layer0_outputs(4484) <= inputs(71);
    layer0_outputs(4485) <= (inputs(161)) xor (inputs(131));
    layer0_outputs(4486) <= not(inputs(64)) or (inputs(63));
    layer0_outputs(4487) <= not((inputs(232)) or (inputs(162)));
    layer0_outputs(4488) <= inputs(154);
    layer0_outputs(4489) <= inputs(24);
    layer0_outputs(4490) <= not(inputs(211)) or (inputs(77));
    layer0_outputs(4491) <= not(inputs(96)) or (inputs(51));
    layer0_outputs(4492) <= not(inputs(110));
    layer0_outputs(4493) <= not(inputs(169));
    layer0_outputs(4494) <= (inputs(181)) or (inputs(42));
    layer0_outputs(4495) <= inputs(220);
    layer0_outputs(4496) <= inputs(74);
    layer0_outputs(4497) <= (inputs(100)) or (inputs(108));
    layer0_outputs(4498) <= not((inputs(201)) and (inputs(227)));
    layer0_outputs(4499) <= not(inputs(158));
    layer0_outputs(4500) <= not((inputs(153)) or (inputs(77)));
    layer0_outputs(4501) <= (inputs(134)) and not (inputs(140));
    layer0_outputs(4502) <= (inputs(145)) xor (inputs(131));
    layer0_outputs(4503) <= not((inputs(130)) and (inputs(236)));
    layer0_outputs(4504) <= not(inputs(253));
    layer0_outputs(4505) <= '0';
    layer0_outputs(4506) <= not(inputs(213));
    layer0_outputs(4507) <= inputs(166);
    layer0_outputs(4508) <= (inputs(138)) or (inputs(97));
    layer0_outputs(4509) <= not((inputs(13)) xor (inputs(46)));
    layer0_outputs(4510) <= not(inputs(23));
    layer0_outputs(4511) <= not(inputs(82));
    layer0_outputs(4512) <= '0';
    layer0_outputs(4513) <= (inputs(235)) and not (inputs(186));
    layer0_outputs(4514) <= not((inputs(112)) and (inputs(35)));
    layer0_outputs(4515) <= not((inputs(73)) or (inputs(19)));
    layer0_outputs(4516) <= (inputs(171)) and (inputs(20));
    layer0_outputs(4517) <= (inputs(184)) or (inputs(75));
    layer0_outputs(4518) <= not(inputs(9)) or (inputs(253));
    layer0_outputs(4519) <= inputs(65);
    layer0_outputs(4520) <= not(inputs(37));
    layer0_outputs(4521) <= (inputs(94)) and (inputs(150));
    layer0_outputs(4522) <= inputs(221);
    layer0_outputs(4523) <= (inputs(126)) xor (inputs(252));
    layer0_outputs(4524) <= (inputs(115)) and not (inputs(89));
    layer0_outputs(4525) <= (inputs(68)) and not (inputs(242));
    layer0_outputs(4526) <= not(inputs(228)) or (inputs(64));
    layer0_outputs(4527) <= (inputs(157)) and not (inputs(235));
    layer0_outputs(4528) <= not((inputs(161)) or (inputs(252)));
    layer0_outputs(4529) <= not(inputs(107));
    layer0_outputs(4530) <= not(inputs(167)) or (inputs(4));
    layer0_outputs(4531) <= not((inputs(210)) or (inputs(47)));
    layer0_outputs(4532) <= not((inputs(12)) or (inputs(154)));
    layer0_outputs(4533) <= (inputs(223)) xor (inputs(3));
    layer0_outputs(4534) <= '1';
    layer0_outputs(4535) <= not(inputs(119));
    layer0_outputs(4536) <= not((inputs(106)) or (inputs(5)));
    layer0_outputs(4537) <= (inputs(191)) and not (inputs(66));
    layer0_outputs(4538) <= not(inputs(227));
    layer0_outputs(4539) <= (inputs(196)) and not (inputs(118));
    layer0_outputs(4540) <= not((inputs(238)) xor (inputs(250)));
    layer0_outputs(4541) <= not(inputs(75)) or (inputs(142));
    layer0_outputs(4542) <= not(inputs(24));
    layer0_outputs(4543) <= not(inputs(25)) or (inputs(237));
    layer0_outputs(4544) <= inputs(53);
    layer0_outputs(4545) <= inputs(67);
    layer0_outputs(4546) <= not(inputs(153));
    layer0_outputs(4547) <= not((inputs(220)) or (inputs(27)));
    layer0_outputs(4548) <= not(inputs(213)) or (inputs(83));
    layer0_outputs(4549) <= not((inputs(154)) or (inputs(149)));
    layer0_outputs(4550) <= '0';
    layer0_outputs(4551) <= (inputs(77)) or (inputs(163));
    layer0_outputs(4552) <= not(inputs(39)) or (inputs(41));
    layer0_outputs(4553) <= '1';
    layer0_outputs(4554) <= (inputs(55)) and not (inputs(228));
    layer0_outputs(4555) <= not(inputs(8));
    layer0_outputs(4556) <= inputs(248);
    layer0_outputs(4557) <= inputs(109);
    layer0_outputs(4558) <= (inputs(114)) or (inputs(148));
    layer0_outputs(4559) <= not((inputs(136)) xor (inputs(146)));
    layer0_outputs(4560) <= (inputs(179)) or (inputs(151));
    layer0_outputs(4561) <= (inputs(178)) or (inputs(142));
    layer0_outputs(4562) <= (inputs(185)) and not (inputs(132));
    layer0_outputs(4563) <= not(inputs(124));
    layer0_outputs(4564) <= inputs(253);
    layer0_outputs(4565) <= not(inputs(151)) or (inputs(114));
    layer0_outputs(4566) <= (inputs(181)) xor (inputs(156));
    layer0_outputs(4567) <= inputs(28);
    layer0_outputs(4568) <= (inputs(167)) xor (inputs(109));
    layer0_outputs(4569) <= not(inputs(219));
    layer0_outputs(4570) <= not(inputs(24));
    layer0_outputs(4571) <= not((inputs(177)) and (inputs(93)));
    layer0_outputs(4572) <= not((inputs(4)) or (inputs(179)));
    layer0_outputs(4573) <= not(inputs(151)) or (inputs(86));
    layer0_outputs(4574) <= not((inputs(74)) and (inputs(138)));
    layer0_outputs(4575) <= inputs(108);
    layer0_outputs(4576) <= inputs(180);
    layer0_outputs(4577) <= not(inputs(126));
    layer0_outputs(4578) <= (inputs(107)) or (inputs(221));
    layer0_outputs(4579) <= inputs(83);
    layer0_outputs(4580) <= not(inputs(103));
    layer0_outputs(4581) <= not(inputs(79)) or (inputs(71));
    layer0_outputs(4582) <= not((inputs(3)) or (inputs(75)));
    layer0_outputs(4583) <= (inputs(173)) or (inputs(142));
    layer0_outputs(4584) <= not(inputs(117)) or (inputs(2));
    layer0_outputs(4585) <= not((inputs(3)) and (inputs(117)));
    layer0_outputs(4586) <= not((inputs(229)) or (inputs(211)));
    layer0_outputs(4587) <= not(inputs(224));
    layer0_outputs(4588) <= not((inputs(50)) and (inputs(217)));
    layer0_outputs(4589) <= not(inputs(29));
    layer0_outputs(4590) <= not((inputs(136)) xor (inputs(121)));
    layer0_outputs(4591) <= not((inputs(66)) or (inputs(227)));
    layer0_outputs(4592) <= not(inputs(145)) or (inputs(137));
    layer0_outputs(4593) <= not(inputs(112));
    layer0_outputs(4594) <= not(inputs(159)) or (inputs(11));
    layer0_outputs(4595) <= (inputs(99)) and not (inputs(158));
    layer0_outputs(4596) <= not((inputs(49)) or (inputs(88)));
    layer0_outputs(4597) <= not(inputs(162));
    layer0_outputs(4598) <= (inputs(134)) or (inputs(223));
    layer0_outputs(4599) <= inputs(90);
    layer0_outputs(4600) <= inputs(165);
    layer0_outputs(4601) <= (inputs(13)) and not (inputs(204));
    layer0_outputs(4602) <= inputs(118);
    layer0_outputs(4603) <= not(inputs(150));
    layer0_outputs(4604) <= not(inputs(199));
    layer0_outputs(4605) <= not((inputs(110)) or (inputs(130)));
    layer0_outputs(4606) <= inputs(168);
    layer0_outputs(4607) <= not((inputs(53)) or (inputs(116)));
    layer0_outputs(4608) <= not(inputs(139)) or (inputs(177));
    layer0_outputs(4609) <= inputs(85);
    layer0_outputs(4610) <= (inputs(133)) and not (inputs(210));
    layer0_outputs(4611) <= not(inputs(199)) or (inputs(36));
    layer0_outputs(4612) <= not(inputs(236));
    layer0_outputs(4613) <= (inputs(135)) and not (inputs(39));
    layer0_outputs(4614) <= not((inputs(53)) and (inputs(89)));
    layer0_outputs(4615) <= (inputs(249)) or (inputs(186));
    layer0_outputs(4616) <= inputs(231);
    layer0_outputs(4617) <= not(inputs(163));
    layer0_outputs(4618) <= not(inputs(167)) or (inputs(29));
    layer0_outputs(4619) <= (inputs(207)) or (inputs(254));
    layer0_outputs(4620) <= not(inputs(247));
    layer0_outputs(4621) <= inputs(69);
    layer0_outputs(4622) <= inputs(246);
    layer0_outputs(4623) <= not((inputs(125)) or (inputs(42)));
    layer0_outputs(4624) <= not((inputs(38)) or (inputs(50)));
    layer0_outputs(4625) <= inputs(53);
    layer0_outputs(4626) <= inputs(196);
    layer0_outputs(4627) <= not(inputs(177));
    layer0_outputs(4628) <= (inputs(7)) and not (inputs(38));
    layer0_outputs(4629) <= not(inputs(218));
    layer0_outputs(4630) <= not((inputs(192)) or (inputs(106)));
    layer0_outputs(4631) <= inputs(114);
    layer0_outputs(4632) <= '1';
    layer0_outputs(4633) <= (inputs(180)) and not (inputs(73));
    layer0_outputs(4634) <= (inputs(241)) and not (inputs(245));
    layer0_outputs(4635) <= not((inputs(17)) or (inputs(88)));
    layer0_outputs(4636) <= inputs(20);
    layer0_outputs(4637) <= not(inputs(106)) or (inputs(1));
    layer0_outputs(4638) <= inputs(97);
    layer0_outputs(4639) <= (inputs(109)) or (inputs(146));
    layer0_outputs(4640) <= not(inputs(184)) or (inputs(75));
    layer0_outputs(4641) <= inputs(202);
    layer0_outputs(4642) <= not(inputs(80)) or (inputs(60));
    layer0_outputs(4643) <= not(inputs(86)) or (inputs(139));
    layer0_outputs(4644) <= (inputs(65)) or (inputs(235));
    layer0_outputs(4645) <= inputs(147);
    layer0_outputs(4646) <= '0';
    layer0_outputs(4647) <= inputs(165);
    layer0_outputs(4648) <= not((inputs(100)) or (inputs(102)));
    layer0_outputs(4649) <= not(inputs(124)) or (inputs(132));
    layer0_outputs(4650) <= not((inputs(143)) or (inputs(226)));
    layer0_outputs(4651) <= inputs(178);
    layer0_outputs(4652) <= inputs(108);
    layer0_outputs(4653) <= not((inputs(96)) xor (inputs(70)));
    layer0_outputs(4654) <= (inputs(95)) or (inputs(182));
    layer0_outputs(4655) <= inputs(223);
    layer0_outputs(4656) <= not((inputs(140)) or (inputs(90)));
    layer0_outputs(4657) <= inputs(180);
    layer0_outputs(4658) <= inputs(147);
    layer0_outputs(4659) <= not((inputs(191)) or (inputs(209)));
    layer0_outputs(4660) <= (inputs(213)) and not (inputs(171));
    layer0_outputs(4661) <= not(inputs(114));
    layer0_outputs(4662) <= (inputs(68)) and not (inputs(225));
    layer0_outputs(4663) <= '0';
    layer0_outputs(4664) <= not((inputs(229)) or (inputs(237)));
    layer0_outputs(4665) <= (inputs(71)) and not (inputs(137));
    layer0_outputs(4666) <= (inputs(231)) or (inputs(207));
    layer0_outputs(4667) <= not(inputs(68));
    layer0_outputs(4668) <= (inputs(225)) and (inputs(189));
    layer0_outputs(4669) <= not(inputs(55));
    layer0_outputs(4670) <= inputs(197);
    layer0_outputs(4671) <= (inputs(93)) xor (inputs(62));
    layer0_outputs(4672) <= not(inputs(151));
    layer0_outputs(4673) <= inputs(165);
    layer0_outputs(4674) <= (inputs(209)) or (inputs(188));
    layer0_outputs(4675) <= not((inputs(6)) or (inputs(177)));
    layer0_outputs(4676) <= not(inputs(164)) or (inputs(112));
    layer0_outputs(4677) <= inputs(45);
    layer0_outputs(4678) <= inputs(64);
    layer0_outputs(4679) <= (inputs(121)) and not (inputs(147));
    layer0_outputs(4680) <= (inputs(46)) xor (inputs(149));
    layer0_outputs(4681) <= not((inputs(254)) or (inputs(54)));
    layer0_outputs(4682) <= not((inputs(226)) or (inputs(135)));
    layer0_outputs(4683) <= (inputs(64)) or (inputs(254));
    layer0_outputs(4684) <= (inputs(163)) xor (inputs(113));
    layer0_outputs(4685) <= not(inputs(99));
    layer0_outputs(4686) <= not(inputs(159));
    layer0_outputs(4687) <= not(inputs(19));
    layer0_outputs(4688) <= not(inputs(209));
    layer0_outputs(4689) <= not((inputs(35)) xor (inputs(46)));
    layer0_outputs(4690) <= not(inputs(41));
    layer0_outputs(4691) <= inputs(174);
    layer0_outputs(4692) <= (inputs(90)) or (inputs(18));
    layer0_outputs(4693) <= not(inputs(214));
    layer0_outputs(4694) <= (inputs(53)) or (inputs(48));
    layer0_outputs(4695) <= not((inputs(31)) xor (inputs(33)));
    layer0_outputs(4696) <= not((inputs(229)) and (inputs(20)));
    layer0_outputs(4697) <= '0';
    layer0_outputs(4698) <= not(inputs(211));
    layer0_outputs(4699) <= not((inputs(26)) or (inputs(59)));
    layer0_outputs(4700) <= not(inputs(140));
    layer0_outputs(4701) <= (inputs(46)) or (inputs(48));
    layer0_outputs(4702) <= inputs(45);
    layer0_outputs(4703) <= inputs(72);
    layer0_outputs(4704) <= not(inputs(55)) or (inputs(15));
    layer0_outputs(4705) <= inputs(227);
    layer0_outputs(4706) <= not(inputs(200));
    layer0_outputs(4707) <= (inputs(199)) or (inputs(254));
    layer0_outputs(4708) <= '0';
    layer0_outputs(4709) <= (inputs(202)) or (inputs(178));
    layer0_outputs(4710) <= (inputs(220)) and not (inputs(0));
    layer0_outputs(4711) <= inputs(4);
    layer0_outputs(4712) <= '1';
    layer0_outputs(4713) <= not(inputs(148));
    layer0_outputs(4714) <= (inputs(184)) and not (inputs(105));
    layer0_outputs(4715) <= not((inputs(101)) and (inputs(108)));
    layer0_outputs(4716) <= '0';
    layer0_outputs(4717) <= not(inputs(246));
    layer0_outputs(4718) <= not((inputs(4)) xor (inputs(186)));
    layer0_outputs(4719) <= not((inputs(169)) or (inputs(111)));
    layer0_outputs(4720) <= not(inputs(106)) or (inputs(97));
    layer0_outputs(4721) <= not((inputs(227)) or (inputs(175)));
    layer0_outputs(4722) <= inputs(11);
    layer0_outputs(4723) <= not(inputs(72));
    layer0_outputs(4724) <= not(inputs(252));
    layer0_outputs(4725) <= (inputs(140)) or (inputs(131));
    layer0_outputs(4726) <= not((inputs(228)) or (inputs(19)));
    layer0_outputs(4727) <= (inputs(146)) or (inputs(142));
    layer0_outputs(4728) <= not((inputs(167)) or (inputs(15)));
    layer0_outputs(4729) <= (inputs(0)) or (inputs(84));
    layer0_outputs(4730) <= inputs(147);
    layer0_outputs(4731) <= inputs(82);
    layer0_outputs(4732) <= (inputs(188)) and not (inputs(251));
    layer0_outputs(4733) <= not(inputs(141)) or (inputs(91));
    layer0_outputs(4734) <= not((inputs(71)) or (inputs(42)));
    layer0_outputs(4735) <= not(inputs(11)) or (inputs(246));
    layer0_outputs(4736) <= (inputs(230)) and not (inputs(22));
    layer0_outputs(4737) <= (inputs(112)) or (inputs(72));
    layer0_outputs(4738) <= (inputs(195)) and not (inputs(96));
    layer0_outputs(4739) <= not((inputs(217)) and (inputs(108)));
    layer0_outputs(4740) <= not((inputs(160)) or (inputs(231)));
    layer0_outputs(4741) <= (inputs(222)) and not (inputs(95));
    layer0_outputs(4742) <= not(inputs(210));
    layer0_outputs(4743) <= not(inputs(186)) or (inputs(251));
    layer0_outputs(4744) <= not((inputs(220)) or (inputs(223)));
    layer0_outputs(4745) <= not((inputs(215)) or (inputs(176)));
    layer0_outputs(4746) <= not((inputs(108)) xor (inputs(179)));
    layer0_outputs(4747) <= not((inputs(75)) or (inputs(108)));
    layer0_outputs(4748) <= inputs(175);
    layer0_outputs(4749) <= (inputs(92)) or (inputs(23));
    layer0_outputs(4750) <= inputs(30);
    layer0_outputs(4751) <= not(inputs(139));
    layer0_outputs(4752) <= not(inputs(153));
    layer0_outputs(4753) <= not(inputs(168)) or (inputs(202));
    layer0_outputs(4754) <= not(inputs(212)) or (inputs(237));
    layer0_outputs(4755) <= not(inputs(89));
    layer0_outputs(4756) <= (inputs(111)) or (inputs(212));
    layer0_outputs(4757) <= not((inputs(145)) xor (inputs(167)));
    layer0_outputs(4758) <= not(inputs(166));
    layer0_outputs(4759) <= not((inputs(19)) or (inputs(35)));
    layer0_outputs(4760) <= not(inputs(60));
    layer0_outputs(4761) <= (inputs(33)) or (inputs(2));
    layer0_outputs(4762) <= not(inputs(91)) or (inputs(63));
    layer0_outputs(4763) <= not(inputs(106)) or (inputs(128));
    layer0_outputs(4764) <= '0';
    layer0_outputs(4765) <= not(inputs(172));
    layer0_outputs(4766) <= (inputs(119)) or (inputs(190));
    layer0_outputs(4767) <= inputs(240);
    layer0_outputs(4768) <= '1';
    layer0_outputs(4769) <= inputs(57);
    layer0_outputs(4770) <= not(inputs(169));
    layer0_outputs(4771) <= not((inputs(206)) or (inputs(202)));
    layer0_outputs(4772) <= not(inputs(72)) or (inputs(186));
    layer0_outputs(4773) <= not((inputs(91)) and (inputs(104)));
    layer0_outputs(4774) <= not(inputs(152));
    layer0_outputs(4775) <= not(inputs(43));
    layer0_outputs(4776) <= not(inputs(185)) or (inputs(179));
    layer0_outputs(4777) <= inputs(213);
    layer0_outputs(4778) <= not((inputs(4)) or (inputs(133)));
    layer0_outputs(4779) <= (inputs(164)) xor (inputs(179));
    layer0_outputs(4780) <= inputs(88);
    layer0_outputs(4781) <= not((inputs(151)) xor (inputs(36)));
    layer0_outputs(4782) <= not((inputs(203)) xor (inputs(85)));
    layer0_outputs(4783) <= inputs(95);
    layer0_outputs(4784) <= not((inputs(22)) or (inputs(65)));
    layer0_outputs(4785) <= (inputs(131)) or (inputs(139));
    layer0_outputs(4786) <= (inputs(242)) and not (inputs(127));
    layer0_outputs(4787) <= (inputs(104)) or (inputs(122));
    layer0_outputs(4788) <= inputs(15);
    layer0_outputs(4789) <= not(inputs(223)) or (inputs(59));
    layer0_outputs(4790) <= not((inputs(77)) or (inputs(41)));
    layer0_outputs(4791) <= '0';
    layer0_outputs(4792) <= (inputs(44)) or (inputs(46));
    layer0_outputs(4793) <= (inputs(222)) and not (inputs(25));
    layer0_outputs(4794) <= not(inputs(216)) or (inputs(165));
    layer0_outputs(4795) <= (inputs(168)) and not (inputs(63));
    layer0_outputs(4796) <= not((inputs(11)) and (inputs(68)));
    layer0_outputs(4797) <= not(inputs(106));
    layer0_outputs(4798) <= (inputs(42)) or (inputs(17));
    layer0_outputs(4799) <= (inputs(214)) or (inputs(219));
    layer0_outputs(4800) <= (inputs(112)) or (inputs(247));
    layer0_outputs(4801) <= not(inputs(24));
    layer0_outputs(4802) <= (inputs(255)) and (inputs(33));
    layer0_outputs(4803) <= not(inputs(223));
    layer0_outputs(4804) <= not((inputs(86)) and (inputs(145)));
    layer0_outputs(4805) <= not(inputs(252));
    layer0_outputs(4806) <= (inputs(12)) and (inputs(57));
    layer0_outputs(4807) <= not(inputs(37));
    layer0_outputs(4808) <= not(inputs(180));
    layer0_outputs(4809) <= (inputs(114)) or (inputs(198));
    layer0_outputs(4810) <= inputs(82);
    layer0_outputs(4811) <= (inputs(180)) xor (inputs(8));
    layer0_outputs(4812) <= not(inputs(19));
    layer0_outputs(4813) <= not((inputs(139)) xor (inputs(206)));
    layer0_outputs(4814) <= '1';
    layer0_outputs(4815) <= not(inputs(73)) or (inputs(202));
    layer0_outputs(4816) <= (inputs(112)) or (inputs(75));
    layer0_outputs(4817) <= (inputs(198)) and (inputs(9));
    layer0_outputs(4818) <= not(inputs(249));
    layer0_outputs(4819) <= '1';
    layer0_outputs(4820) <= '0';
    layer0_outputs(4821) <= not((inputs(121)) and (inputs(230)));
    layer0_outputs(4822) <= not(inputs(182));
    layer0_outputs(4823) <= (inputs(191)) and not (inputs(229));
    layer0_outputs(4824) <= (inputs(147)) and (inputs(118));
    layer0_outputs(4825) <= not((inputs(183)) and (inputs(127)));
    layer0_outputs(4826) <= not(inputs(5)) or (inputs(106));
    layer0_outputs(4827) <= not(inputs(61));
    layer0_outputs(4828) <= (inputs(112)) and not (inputs(109));
    layer0_outputs(4829) <= not(inputs(170));
    layer0_outputs(4830) <= inputs(66);
    layer0_outputs(4831) <= (inputs(242)) or (inputs(187));
    layer0_outputs(4832) <= not(inputs(177)) or (inputs(252));
    layer0_outputs(4833) <= (inputs(70)) or (inputs(181));
    layer0_outputs(4834) <= not((inputs(172)) or (inputs(250)));
    layer0_outputs(4835) <= (inputs(99)) or (inputs(11));
    layer0_outputs(4836) <= not((inputs(207)) xor (inputs(210)));
    layer0_outputs(4837) <= (inputs(5)) or (inputs(31));
    layer0_outputs(4838) <= (inputs(84)) and not (inputs(215));
    layer0_outputs(4839) <= not((inputs(73)) and (inputs(180)));
    layer0_outputs(4840) <= not(inputs(135)) or (inputs(150));
    layer0_outputs(4841) <= (inputs(199)) and not (inputs(93));
    layer0_outputs(4842) <= (inputs(171)) and (inputs(210));
    layer0_outputs(4843) <= not(inputs(25)) or (inputs(113));
    layer0_outputs(4844) <= (inputs(103)) and not (inputs(33));
    layer0_outputs(4845) <= '0';
    layer0_outputs(4846) <= inputs(59);
    layer0_outputs(4847) <= (inputs(191)) and not (inputs(237));
    layer0_outputs(4848) <= (inputs(56)) or (inputs(161));
    layer0_outputs(4849) <= (inputs(187)) or (inputs(103));
    layer0_outputs(4850) <= not((inputs(235)) or (inputs(205)));
    layer0_outputs(4851) <= (inputs(238)) xor (inputs(213));
    layer0_outputs(4852) <= inputs(121);
    layer0_outputs(4853) <= inputs(201);
    layer0_outputs(4854) <= (inputs(100)) or (inputs(113));
    layer0_outputs(4855) <= inputs(8);
    layer0_outputs(4856) <= inputs(206);
    layer0_outputs(4857) <= inputs(136);
    layer0_outputs(4858) <= not(inputs(82));
    layer0_outputs(4859) <= (inputs(70)) or (inputs(20));
    layer0_outputs(4860) <= not(inputs(6)) or (inputs(33));
    layer0_outputs(4861) <= inputs(28);
    layer0_outputs(4862) <= inputs(99);
    layer0_outputs(4863) <= not(inputs(141));
    layer0_outputs(4864) <= not(inputs(246)) or (inputs(113));
    layer0_outputs(4865) <= (inputs(43)) xor (inputs(25));
    layer0_outputs(4866) <= inputs(54);
    layer0_outputs(4867) <= (inputs(114)) and not (inputs(160));
    layer0_outputs(4868) <= not(inputs(217));
    layer0_outputs(4869) <= not(inputs(148));
    layer0_outputs(4870) <= not((inputs(195)) xor (inputs(205)));
    layer0_outputs(4871) <= (inputs(20)) and not (inputs(171));
    layer0_outputs(4872) <= (inputs(229)) or (inputs(174));
    layer0_outputs(4873) <= (inputs(89)) and not (inputs(207));
    layer0_outputs(4874) <= not(inputs(92));
    layer0_outputs(4875) <= (inputs(189)) or (inputs(135));
    layer0_outputs(4876) <= not((inputs(108)) or (inputs(156)));
    layer0_outputs(4877) <= (inputs(218)) or (inputs(144));
    layer0_outputs(4878) <= not(inputs(12));
    layer0_outputs(4879) <= not((inputs(82)) or (inputs(115)));
    layer0_outputs(4880) <= inputs(115);
    layer0_outputs(4881) <= inputs(13);
    layer0_outputs(4882) <= inputs(29);
    layer0_outputs(4883) <= not((inputs(135)) or (inputs(175)));
    layer0_outputs(4884) <= not((inputs(116)) or (inputs(15)));
    layer0_outputs(4885) <= (inputs(2)) and not (inputs(90));
    layer0_outputs(4886) <= (inputs(27)) and not (inputs(203));
    layer0_outputs(4887) <= not(inputs(55));
    layer0_outputs(4888) <= not(inputs(175)) or (inputs(242));
    layer0_outputs(4889) <= not((inputs(131)) or (inputs(54)));
    layer0_outputs(4890) <= inputs(192);
    layer0_outputs(4891) <= (inputs(86)) and (inputs(37));
    layer0_outputs(4892) <= not((inputs(5)) xor (inputs(141)));
    layer0_outputs(4893) <= not(inputs(129));
    layer0_outputs(4894) <= not(inputs(83));
    layer0_outputs(4895) <= not(inputs(229)) or (inputs(119));
    layer0_outputs(4896) <= not(inputs(131)) or (inputs(242));
    layer0_outputs(4897) <= not((inputs(48)) or (inputs(60)));
    layer0_outputs(4898) <= (inputs(74)) and not (inputs(102));
    layer0_outputs(4899) <= inputs(69);
    layer0_outputs(4900) <= (inputs(241)) or (inputs(26));
    layer0_outputs(4901) <= not(inputs(116));
    layer0_outputs(4902) <= not((inputs(25)) xor (inputs(71)));
    layer0_outputs(4903) <= inputs(238);
    layer0_outputs(4904) <= not(inputs(143));
    layer0_outputs(4905) <= not(inputs(35)) or (inputs(250));
    layer0_outputs(4906) <= (inputs(233)) or (inputs(205));
    layer0_outputs(4907) <= '1';
    layer0_outputs(4908) <= not(inputs(165));
    layer0_outputs(4909) <= (inputs(184)) xor (inputs(232));
    layer0_outputs(4910) <= (inputs(184)) and not (inputs(103));
    layer0_outputs(4911) <= not((inputs(253)) and (inputs(193)));
    layer0_outputs(4912) <= not(inputs(22)) or (inputs(113));
    layer0_outputs(4913) <= (inputs(132)) or (inputs(148));
    layer0_outputs(4914) <= '1';
    layer0_outputs(4915) <= '1';
    layer0_outputs(4916) <= (inputs(68)) or (inputs(111));
    layer0_outputs(4917) <= not(inputs(248)) or (inputs(64));
    layer0_outputs(4918) <= not(inputs(195));
    layer0_outputs(4919) <= not(inputs(226)) or (inputs(89));
    layer0_outputs(4920) <= inputs(61);
    layer0_outputs(4921) <= '1';
    layer0_outputs(4922) <= not(inputs(95));
    layer0_outputs(4923) <= not(inputs(192));
    layer0_outputs(4924) <= (inputs(71)) and not (inputs(161));
    layer0_outputs(4925) <= inputs(212);
    layer0_outputs(4926) <= (inputs(221)) and (inputs(26));
    layer0_outputs(4927) <= (inputs(48)) and (inputs(200));
    layer0_outputs(4928) <= not(inputs(26));
    layer0_outputs(4929) <= not(inputs(32));
    layer0_outputs(4930) <= not((inputs(2)) or (inputs(228)));
    layer0_outputs(4931) <= (inputs(151)) and not (inputs(158));
    layer0_outputs(4932) <= not((inputs(95)) and (inputs(2)));
    layer0_outputs(4933) <= (inputs(253)) xor (inputs(156));
    layer0_outputs(4934) <= inputs(30);
    layer0_outputs(4935) <= (inputs(73)) or (inputs(94));
    layer0_outputs(4936) <= '1';
    layer0_outputs(4937) <= not(inputs(237));
    layer0_outputs(4938) <= not(inputs(138)) or (inputs(197));
    layer0_outputs(4939) <= not((inputs(91)) xor (inputs(19)));
    layer0_outputs(4940) <= (inputs(95)) and not (inputs(232));
    layer0_outputs(4941) <= (inputs(131)) and not (inputs(50));
    layer0_outputs(4942) <= (inputs(184)) and not (inputs(72));
    layer0_outputs(4943) <= not((inputs(203)) or (inputs(172)));
    layer0_outputs(4944) <= inputs(228);
    layer0_outputs(4945) <= not((inputs(8)) or (inputs(151)));
    layer0_outputs(4946) <= (inputs(132)) and not (inputs(19));
    layer0_outputs(4947) <= inputs(153);
    layer0_outputs(4948) <= inputs(1);
    layer0_outputs(4949) <= not(inputs(184));
    layer0_outputs(4950) <= (inputs(131)) or (inputs(193));
    layer0_outputs(4951) <= not(inputs(135)) or (inputs(226));
    layer0_outputs(4952) <= (inputs(4)) and not (inputs(170));
    layer0_outputs(4953) <= not((inputs(49)) xor (inputs(80)));
    layer0_outputs(4954) <= not((inputs(4)) or (inputs(59)));
    layer0_outputs(4955) <= not(inputs(137)) or (inputs(178));
    layer0_outputs(4956) <= '1';
    layer0_outputs(4957) <= not((inputs(166)) or (inputs(74)));
    layer0_outputs(4958) <= (inputs(174)) xor (inputs(71));
    layer0_outputs(4959) <= '0';
    layer0_outputs(4960) <= not(inputs(24)) or (inputs(253));
    layer0_outputs(4961) <= inputs(227);
    layer0_outputs(4962) <= not(inputs(135));
    layer0_outputs(4963) <= (inputs(166)) and not (inputs(125));
    layer0_outputs(4964) <= (inputs(102)) or (inputs(204));
    layer0_outputs(4965) <= not((inputs(181)) or (inputs(252)));
    layer0_outputs(4966) <= (inputs(152)) and (inputs(2));
    layer0_outputs(4967) <= inputs(47);
    layer0_outputs(4968) <= (inputs(147)) and not (inputs(254));
    layer0_outputs(4969) <= not(inputs(104));
    layer0_outputs(4970) <= not((inputs(153)) and (inputs(160)));
    layer0_outputs(4971) <= not(inputs(108)) or (inputs(132));
    layer0_outputs(4972) <= '0';
    layer0_outputs(4973) <= not((inputs(35)) xor (inputs(147)));
    layer0_outputs(4974) <= inputs(254);
    layer0_outputs(4975) <= (inputs(189)) or (inputs(38));
    layer0_outputs(4976) <= not(inputs(9)) or (inputs(128));
    layer0_outputs(4977) <= not((inputs(139)) and (inputs(24)));
    layer0_outputs(4978) <= '0';
    layer0_outputs(4979) <= not(inputs(219));
    layer0_outputs(4980) <= (inputs(75)) or (inputs(53));
    layer0_outputs(4981) <= not(inputs(202));
    layer0_outputs(4982) <= (inputs(241)) and not (inputs(209));
    layer0_outputs(4983) <= not((inputs(120)) or (inputs(223)));
    layer0_outputs(4984) <= (inputs(15)) and not (inputs(68));
    layer0_outputs(4985) <= (inputs(193)) or (inputs(214));
    layer0_outputs(4986) <= not((inputs(155)) or (inputs(229)));
    layer0_outputs(4987) <= not(inputs(90));
    layer0_outputs(4988) <= not(inputs(100)) or (inputs(36));
    layer0_outputs(4989) <= inputs(65);
    layer0_outputs(4990) <= (inputs(69)) and not (inputs(216));
    layer0_outputs(4991) <= not(inputs(162));
    layer0_outputs(4992) <= not((inputs(193)) or (inputs(221)));
    layer0_outputs(4993) <= not((inputs(24)) or (inputs(226)));
    layer0_outputs(4994) <= inputs(114);
    layer0_outputs(4995) <= (inputs(193)) and not (inputs(227));
    layer0_outputs(4996) <= (inputs(80)) or (inputs(16));
    layer0_outputs(4997) <= (inputs(140)) and not (inputs(224));
    layer0_outputs(4998) <= (inputs(255)) and not (inputs(41));
    layer0_outputs(4999) <= (inputs(78)) and (inputs(220));
    layer0_outputs(5000) <= (inputs(192)) or (inputs(235));
    layer0_outputs(5001) <= (inputs(125)) and not (inputs(41));
    layer0_outputs(5002) <= inputs(208);
    layer0_outputs(5003) <= (inputs(3)) or (inputs(148));
    layer0_outputs(5004) <= not((inputs(207)) xor (inputs(226)));
    layer0_outputs(5005) <= not((inputs(210)) or (inputs(91)));
    layer0_outputs(5006) <= not(inputs(119));
    layer0_outputs(5007) <= not((inputs(180)) or (inputs(9)));
    layer0_outputs(5008) <= inputs(25);
    layer0_outputs(5009) <= not(inputs(28)) or (inputs(252));
    layer0_outputs(5010) <= inputs(206);
    layer0_outputs(5011) <= (inputs(150)) and not (inputs(221));
    layer0_outputs(5012) <= inputs(92);
    layer0_outputs(5013) <= not(inputs(81)) or (inputs(85));
    layer0_outputs(5014) <= not(inputs(196)) or (inputs(45));
    layer0_outputs(5015) <= not(inputs(116)) or (inputs(147));
    layer0_outputs(5016) <= not(inputs(86));
    layer0_outputs(5017) <= '1';
    layer0_outputs(5018) <= not((inputs(110)) or (inputs(40)));
    layer0_outputs(5019) <= inputs(71);
    layer0_outputs(5020) <= (inputs(96)) and not (inputs(225));
    layer0_outputs(5021) <= (inputs(173)) and not (inputs(43));
    layer0_outputs(5022) <= inputs(57);
    layer0_outputs(5023) <= (inputs(66)) and not (inputs(119));
    layer0_outputs(5024) <= not(inputs(165));
    layer0_outputs(5025) <= inputs(234);
    layer0_outputs(5026) <= not(inputs(23)) or (inputs(223));
    layer0_outputs(5027) <= not(inputs(151)) or (inputs(117));
    layer0_outputs(5028) <= not(inputs(150));
    layer0_outputs(5029) <= not((inputs(240)) or (inputs(172)));
    layer0_outputs(5030) <= '0';
    layer0_outputs(5031) <= (inputs(182)) and not (inputs(26));
    layer0_outputs(5032) <= not((inputs(93)) or (inputs(147)));
    layer0_outputs(5033) <= inputs(179);
    layer0_outputs(5034) <= '0';
    layer0_outputs(5035) <= not(inputs(26)) or (inputs(170));
    layer0_outputs(5036) <= (inputs(146)) and not (inputs(66));
    layer0_outputs(5037) <= not(inputs(62));
    layer0_outputs(5038) <= not((inputs(168)) or (inputs(179)));
    layer0_outputs(5039) <= not((inputs(159)) xor (inputs(166)));
    layer0_outputs(5040) <= inputs(137);
    layer0_outputs(5041) <= not((inputs(7)) and (inputs(59)));
    layer0_outputs(5042) <= not(inputs(107));
    layer0_outputs(5043) <= (inputs(216)) and not (inputs(244));
    layer0_outputs(5044) <= not(inputs(179));
    layer0_outputs(5045) <= (inputs(59)) and not (inputs(11));
    layer0_outputs(5046) <= not(inputs(43));
    layer0_outputs(5047) <= not((inputs(155)) xor (inputs(14)));
    layer0_outputs(5048) <= (inputs(43)) and not (inputs(168));
    layer0_outputs(5049) <= not(inputs(47));
    layer0_outputs(5050) <= inputs(251);
    layer0_outputs(5051) <= not((inputs(24)) xor (inputs(54)));
    layer0_outputs(5052) <= not((inputs(23)) or (inputs(39)));
    layer0_outputs(5053) <= not(inputs(2));
    layer0_outputs(5054) <= not(inputs(109)) or (inputs(81));
    layer0_outputs(5055) <= inputs(62);
    layer0_outputs(5056) <= (inputs(245)) and not (inputs(93));
    layer0_outputs(5057) <= not(inputs(169)) or (inputs(78));
    layer0_outputs(5058) <= not((inputs(184)) or (inputs(1)));
    layer0_outputs(5059) <= not(inputs(22)) or (inputs(251));
    layer0_outputs(5060) <= (inputs(235)) or (inputs(16));
    layer0_outputs(5061) <= '1';
    layer0_outputs(5062) <= inputs(2);
    layer0_outputs(5063) <= '1';
    layer0_outputs(5064) <= not((inputs(250)) or (inputs(242)));
    layer0_outputs(5065) <= (inputs(204)) xor (inputs(169));
    layer0_outputs(5066) <= inputs(10);
    layer0_outputs(5067) <= (inputs(12)) and not (inputs(83));
    layer0_outputs(5068) <= not((inputs(146)) or (inputs(94)));
    layer0_outputs(5069) <= not(inputs(159));
    layer0_outputs(5070) <= (inputs(72)) and not (inputs(250));
    layer0_outputs(5071) <= (inputs(18)) or (inputs(141));
    layer0_outputs(5072) <= not(inputs(183)) or (inputs(91));
    layer0_outputs(5073) <= not(inputs(56)) or (inputs(29));
    layer0_outputs(5074) <= not(inputs(232));
    layer0_outputs(5075) <= (inputs(69)) xor (inputs(139));
    layer0_outputs(5076) <= (inputs(52)) or (inputs(243));
    layer0_outputs(5077) <= '0';
    layer0_outputs(5078) <= (inputs(133)) xor (inputs(209));
    layer0_outputs(5079) <= not(inputs(213));
    layer0_outputs(5080) <= not((inputs(70)) xor (inputs(251)));
    layer0_outputs(5081) <= (inputs(53)) and not (inputs(47));
    layer0_outputs(5082) <= not(inputs(85)) or (inputs(21));
    layer0_outputs(5083) <= '1';
    layer0_outputs(5084) <= inputs(180);
    layer0_outputs(5085) <= not((inputs(193)) or (inputs(223)));
    layer0_outputs(5086) <= '1';
    layer0_outputs(5087) <= inputs(109);
    layer0_outputs(5088) <= not((inputs(112)) or (inputs(89)));
    layer0_outputs(5089) <= (inputs(55)) and not (inputs(137));
    layer0_outputs(5090) <= not((inputs(160)) xor (inputs(231)));
    layer0_outputs(5091) <= not(inputs(51)) or (inputs(149));
    layer0_outputs(5092) <= not((inputs(223)) or (inputs(181)));
    layer0_outputs(5093) <= inputs(102);
    layer0_outputs(5094) <= not((inputs(104)) or (inputs(198)));
    layer0_outputs(5095) <= not((inputs(175)) xor (inputs(70)));
    layer0_outputs(5096) <= inputs(59);
    layer0_outputs(5097) <= not(inputs(220));
    layer0_outputs(5098) <= inputs(8);
    layer0_outputs(5099) <= inputs(179);
    layer0_outputs(5100) <= not((inputs(124)) and (inputs(136)));
    layer0_outputs(5101) <= not(inputs(116)) or (inputs(76));
    layer0_outputs(5102) <= not(inputs(55)) or (inputs(187));
    layer0_outputs(5103) <= not((inputs(44)) and (inputs(44)));
    layer0_outputs(5104) <= not((inputs(185)) and (inputs(179)));
    layer0_outputs(5105) <= inputs(231);
    layer0_outputs(5106) <= (inputs(160)) xor (inputs(172));
    layer0_outputs(5107) <= not(inputs(144));
    layer0_outputs(5108) <= not((inputs(230)) or (inputs(132)));
    layer0_outputs(5109) <= not((inputs(175)) and (inputs(107)));
    layer0_outputs(5110) <= not(inputs(94));
    layer0_outputs(5111) <= not(inputs(249)) or (inputs(56));
    layer0_outputs(5112) <= (inputs(144)) and not (inputs(85));
    layer0_outputs(5113) <= not(inputs(15));
    layer0_outputs(5114) <= (inputs(97)) or (inputs(153));
    layer0_outputs(5115) <= not(inputs(139));
    layer0_outputs(5116) <= not(inputs(59)) or (inputs(54));
    layer0_outputs(5117) <= (inputs(110)) and (inputs(225));
    layer0_outputs(5118) <= not(inputs(248));
    layer0_outputs(5119) <= (inputs(121)) and not (inputs(198));
    layer0_outputs(5120) <= not(inputs(114)) or (inputs(79));
    layer0_outputs(5121) <= (inputs(99)) or (inputs(173));
    layer0_outputs(5122) <= not((inputs(213)) and (inputs(184)));
    layer0_outputs(5123) <= (inputs(117)) and not (inputs(220));
    layer0_outputs(5124) <= not(inputs(183));
    layer0_outputs(5125) <= '0';
    layer0_outputs(5126) <= not(inputs(222));
    layer0_outputs(5127) <= not(inputs(118));
    layer0_outputs(5128) <= not(inputs(117));
    layer0_outputs(5129) <= (inputs(232)) or (inputs(202));
    layer0_outputs(5130) <= not(inputs(246));
    layer0_outputs(5131) <= not(inputs(172)) or (inputs(99));
    layer0_outputs(5132) <= inputs(92);
    layer0_outputs(5133) <= inputs(119);
    layer0_outputs(5134) <= not(inputs(114)) or (inputs(144));
    layer0_outputs(5135) <= (inputs(190)) and not (inputs(29));
    layer0_outputs(5136) <= not(inputs(24));
    layer0_outputs(5137) <= not((inputs(220)) or (inputs(7)));
    layer0_outputs(5138) <= not((inputs(74)) xor (inputs(241)));
    layer0_outputs(5139) <= inputs(110);
    layer0_outputs(5140) <= inputs(72);
    layer0_outputs(5141) <= not((inputs(93)) or (inputs(108)));
    layer0_outputs(5142) <= not(inputs(88));
    layer0_outputs(5143) <= inputs(219);
    layer0_outputs(5144) <= '1';
    layer0_outputs(5145) <= not(inputs(85));
    layer0_outputs(5146) <= not(inputs(179));
    layer0_outputs(5147) <= not((inputs(145)) or (inputs(83)));
    layer0_outputs(5148) <= not((inputs(111)) or (inputs(204)));
    layer0_outputs(5149) <= '1';
    layer0_outputs(5150) <= inputs(161);
    layer0_outputs(5151) <= inputs(131);
    layer0_outputs(5152) <= not((inputs(75)) or (inputs(0)));
    layer0_outputs(5153) <= inputs(202);
    layer0_outputs(5154) <= not(inputs(66));
    layer0_outputs(5155) <= inputs(27);
    layer0_outputs(5156) <= (inputs(237)) or (inputs(136));
    layer0_outputs(5157) <= inputs(5);
    layer0_outputs(5158) <= not(inputs(105));
    layer0_outputs(5159) <= (inputs(233)) or (inputs(167));
    layer0_outputs(5160) <= (inputs(56)) and (inputs(138));
    layer0_outputs(5161) <= not(inputs(211)) or (inputs(190));
    layer0_outputs(5162) <= (inputs(90)) and not (inputs(215));
    layer0_outputs(5163) <= (inputs(184)) or (inputs(195));
    layer0_outputs(5164) <= '1';
    layer0_outputs(5165) <= not((inputs(125)) and (inputs(67)));
    layer0_outputs(5166) <= (inputs(127)) and (inputs(41));
    layer0_outputs(5167) <= not(inputs(146));
    layer0_outputs(5168) <= not(inputs(141)) or (inputs(201));
    layer0_outputs(5169) <= not(inputs(122)) or (inputs(131));
    layer0_outputs(5170) <= not((inputs(243)) or (inputs(131)));
    layer0_outputs(5171) <= (inputs(159)) or (inputs(188));
    layer0_outputs(5172) <= inputs(132);
    layer0_outputs(5173) <= not(inputs(249));
    layer0_outputs(5174) <= (inputs(94)) or (inputs(37));
    layer0_outputs(5175) <= (inputs(5)) or (inputs(254));
    layer0_outputs(5176) <= not(inputs(222)) or (inputs(82));
    layer0_outputs(5177) <= not((inputs(228)) or (inputs(220)));
    layer0_outputs(5178) <= inputs(172);
    layer0_outputs(5179) <= (inputs(28)) or (inputs(130));
    layer0_outputs(5180) <= not((inputs(241)) or (inputs(242)));
    layer0_outputs(5181) <= (inputs(65)) and not (inputs(49));
    layer0_outputs(5182) <= (inputs(227)) and not (inputs(66));
    layer0_outputs(5183) <= not(inputs(40));
    layer0_outputs(5184) <= '1';
    layer0_outputs(5185) <= not(inputs(165));
    layer0_outputs(5186) <= not(inputs(12));
    layer0_outputs(5187) <= not(inputs(118));
    layer0_outputs(5188) <= (inputs(120)) and not (inputs(5));
    layer0_outputs(5189) <= not((inputs(28)) and (inputs(44)));
    layer0_outputs(5190) <= (inputs(69)) xor (inputs(13));
    layer0_outputs(5191) <= not(inputs(209));
    layer0_outputs(5192) <= not(inputs(180)) or (inputs(156));
    layer0_outputs(5193) <= inputs(231);
    layer0_outputs(5194) <= not(inputs(85));
    layer0_outputs(5195) <= (inputs(228)) and (inputs(114));
    layer0_outputs(5196) <= not((inputs(188)) or (inputs(4)));
    layer0_outputs(5197) <= not(inputs(234));
    layer0_outputs(5198) <= not(inputs(63));
    layer0_outputs(5199) <= not(inputs(119));
    layer0_outputs(5200) <= (inputs(34)) and not (inputs(251));
    layer0_outputs(5201) <= (inputs(252)) and not (inputs(2));
    layer0_outputs(5202) <= (inputs(223)) or (inputs(3));
    layer0_outputs(5203) <= not((inputs(60)) or (inputs(78)));
    layer0_outputs(5204) <= not(inputs(53)) or (inputs(44));
    layer0_outputs(5205) <= not((inputs(12)) or (inputs(18)));
    layer0_outputs(5206) <= inputs(7);
    layer0_outputs(5207) <= not(inputs(196)) or (inputs(1));
    layer0_outputs(5208) <= not(inputs(105));
    layer0_outputs(5209) <= not(inputs(141));
    layer0_outputs(5210) <= (inputs(76)) and (inputs(44));
    layer0_outputs(5211) <= not(inputs(149));
    layer0_outputs(5212) <= not(inputs(177)) or (inputs(158));
    layer0_outputs(5213) <= not(inputs(204));
    layer0_outputs(5214) <= not(inputs(201));
    layer0_outputs(5215) <= not((inputs(245)) xor (inputs(37)));
    layer0_outputs(5216) <= (inputs(168)) and (inputs(253));
    layer0_outputs(5217) <= inputs(212);
    layer0_outputs(5218) <= not(inputs(113));
    layer0_outputs(5219) <= (inputs(56)) and not (inputs(79));
    layer0_outputs(5220) <= not(inputs(21));
    layer0_outputs(5221) <= inputs(28);
    layer0_outputs(5222) <= not(inputs(212)) or (inputs(75));
    layer0_outputs(5223) <= not(inputs(83));
    layer0_outputs(5224) <= '1';
    layer0_outputs(5225) <= (inputs(62)) and (inputs(49));
    layer0_outputs(5226) <= inputs(87);
    layer0_outputs(5227) <= not(inputs(210));
    layer0_outputs(5228) <= not((inputs(77)) xor (inputs(43)));
    layer0_outputs(5229) <= not((inputs(99)) xor (inputs(182)));
    layer0_outputs(5230) <= not(inputs(46)) or (inputs(34));
    layer0_outputs(5231) <= not(inputs(192)) or (inputs(225));
    layer0_outputs(5232) <= not(inputs(4)) or (inputs(155));
    layer0_outputs(5233) <= not((inputs(218)) or (inputs(186)));
    layer0_outputs(5234) <= (inputs(22)) or (inputs(6));
    layer0_outputs(5235) <= inputs(120);
    layer0_outputs(5236) <= (inputs(2)) or (inputs(126));
    layer0_outputs(5237) <= not(inputs(37)) or (inputs(13));
    layer0_outputs(5238) <= not((inputs(50)) or (inputs(78)));
    layer0_outputs(5239) <= not(inputs(92));
    layer0_outputs(5240) <= (inputs(14)) or (inputs(96));
    layer0_outputs(5241) <= not(inputs(109));
    layer0_outputs(5242) <= (inputs(66)) xor (inputs(86));
    layer0_outputs(5243) <= not(inputs(50)) or (inputs(170));
    layer0_outputs(5244) <= not((inputs(246)) or (inputs(205)));
    layer0_outputs(5245) <= (inputs(33)) or (inputs(34));
    layer0_outputs(5246) <= (inputs(37)) and not (inputs(240));
    layer0_outputs(5247) <= '1';
    layer0_outputs(5248) <= (inputs(227)) or (inputs(0));
    layer0_outputs(5249) <= inputs(101);
    layer0_outputs(5250) <= (inputs(36)) and (inputs(60));
    layer0_outputs(5251) <= (inputs(10)) and not (inputs(60));
    layer0_outputs(5252) <= (inputs(194)) xor (inputs(38));
    layer0_outputs(5253) <= not((inputs(91)) xor (inputs(126)));
    layer0_outputs(5254) <= not((inputs(152)) and (inputs(156)));
    layer0_outputs(5255) <= not((inputs(193)) xor (inputs(5)));
    layer0_outputs(5256) <= inputs(52);
    layer0_outputs(5257) <= inputs(133);
    layer0_outputs(5258) <= '0';
    layer0_outputs(5259) <= (inputs(181)) and not (inputs(46));
    layer0_outputs(5260) <= not(inputs(21)) or (inputs(123));
    layer0_outputs(5261) <= (inputs(22)) and (inputs(63));
    layer0_outputs(5262) <= '1';
    layer0_outputs(5263) <= inputs(15);
    layer0_outputs(5264) <= (inputs(128)) or (inputs(156));
    layer0_outputs(5265) <= (inputs(244)) or (inputs(1));
    layer0_outputs(5266) <= (inputs(45)) xor (inputs(14));
    layer0_outputs(5267) <= (inputs(36)) and not (inputs(189));
    layer0_outputs(5268) <= not(inputs(72)) or (inputs(102));
    layer0_outputs(5269) <= inputs(138);
    layer0_outputs(5270) <= (inputs(92)) or (inputs(6));
    layer0_outputs(5271) <= not(inputs(19));
    layer0_outputs(5272) <= inputs(161);
    layer0_outputs(5273) <= not(inputs(9));
    layer0_outputs(5274) <= not(inputs(228)) or (inputs(35));
    layer0_outputs(5275) <= not(inputs(5)) or (inputs(221));
    layer0_outputs(5276) <= inputs(103);
    layer0_outputs(5277) <= (inputs(118)) and not (inputs(20));
    layer0_outputs(5278) <= inputs(180);
    layer0_outputs(5279) <= not((inputs(131)) or (inputs(82)));
    layer0_outputs(5280) <= inputs(89);
    layer0_outputs(5281) <= (inputs(72)) and (inputs(145));
    layer0_outputs(5282) <= not((inputs(157)) or (inputs(81)));
    layer0_outputs(5283) <= inputs(83);
    layer0_outputs(5284) <= (inputs(7)) and not (inputs(101));
    layer0_outputs(5285) <= '0';
    layer0_outputs(5286) <= '1';
    layer0_outputs(5287) <= not(inputs(104)) or (inputs(185));
    layer0_outputs(5288) <= not(inputs(209));
    layer0_outputs(5289) <= (inputs(63)) and not (inputs(19));
    layer0_outputs(5290) <= not(inputs(86));
    layer0_outputs(5291) <= not(inputs(175));
    layer0_outputs(5292) <= not(inputs(225));
    layer0_outputs(5293) <= (inputs(167)) or (inputs(223));
    layer0_outputs(5294) <= not(inputs(149)) or (inputs(26));
    layer0_outputs(5295) <= not((inputs(248)) and (inputs(83)));
    layer0_outputs(5296) <= (inputs(208)) or (inputs(237));
    layer0_outputs(5297) <= not((inputs(111)) or (inputs(190)));
    layer0_outputs(5298) <= (inputs(176)) and not (inputs(185));
    layer0_outputs(5299) <= (inputs(19)) or (inputs(153));
    layer0_outputs(5300) <= not((inputs(117)) or (inputs(93)));
    layer0_outputs(5301) <= not((inputs(23)) xor (inputs(246)));
    layer0_outputs(5302) <= (inputs(235)) or (inputs(237));
    layer0_outputs(5303) <= not((inputs(100)) or (inputs(149)));
    layer0_outputs(5304) <= (inputs(106)) and not (inputs(140));
    layer0_outputs(5305) <= not(inputs(65)) or (inputs(95));
    layer0_outputs(5306) <= (inputs(141)) and not (inputs(135));
    layer0_outputs(5307) <= not((inputs(185)) or (inputs(111)));
    layer0_outputs(5308) <= not((inputs(120)) xor (inputs(238)));
    layer0_outputs(5309) <= not(inputs(147));
    layer0_outputs(5310) <= (inputs(83)) xor (inputs(5));
    layer0_outputs(5311) <= not((inputs(94)) or (inputs(80)));
    layer0_outputs(5312) <= not((inputs(52)) or (inputs(45)));
    layer0_outputs(5313) <= not((inputs(151)) or (inputs(137)));
    layer0_outputs(5314) <= not((inputs(206)) or (inputs(158)));
    layer0_outputs(5315) <= not((inputs(195)) xor (inputs(16)));
    layer0_outputs(5316) <= (inputs(78)) and not (inputs(109));
    layer0_outputs(5317) <= (inputs(88)) and not (inputs(250));
    layer0_outputs(5318) <= (inputs(41)) and (inputs(58));
    layer0_outputs(5319) <= not(inputs(247)) or (inputs(64));
    layer0_outputs(5320) <= inputs(147);
    layer0_outputs(5321) <= (inputs(194)) xor (inputs(65));
    layer0_outputs(5322) <= not((inputs(248)) and (inputs(248)));
    layer0_outputs(5323) <= not(inputs(3));
    layer0_outputs(5324) <= not(inputs(8)) or (inputs(86));
    layer0_outputs(5325) <= not((inputs(112)) or (inputs(253)));
    layer0_outputs(5326) <= (inputs(185)) and not (inputs(128));
    layer0_outputs(5327) <= not(inputs(103)) or (inputs(222));
    layer0_outputs(5328) <= inputs(61);
    layer0_outputs(5329) <= inputs(114);
    layer0_outputs(5330) <= (inputs(209)) and not (inputs(214));
    layer0_outputs(5331) <= (inputs(24)) and not (inputs(145));
    layer0_outputs(5332) <= not(inputs(224)) or (inputs(143));
    layer0_outputs(5333) <= not((inputs(81)) or (inputs(212)));
    layer0_outputs(5334) <= (inputs(89)) xor (inputs(161));
    layer0_outputs(5335) <= not(inputs(182));
    layer0_outputs(5336) <= not(inputs(131)) or (inputs(44));
    layer0_outputs(5337) <= not(inputs(91)) or (inputs(182));
    layer0_outputs(5338) <= inputs(8);
    layer0_outputs(5339) <= not(inputs(98));
    layer0_outputs(5340) <= (inputs(94)) and not (inputs(122));
    layer0_outputs(5341) <= (inputs(56)) or (inputs(227));
    layer0_outputs(5342) <= not((inputs(107)) xor (inputs(172)));
    layer0_outputs(5343) <= (inputs(196)) xor (inputs(194));
    layer0_outputs(5344) <= not((inputs(90)) or (inputs(120)));
    layer0_outputs(5345) <= inputs(8);
    layer0_outputs(5346) <= (inputs(56)) and not (inputs(246));
    layer0_outputs(5347) <= not(inputs(114));
    layer0_outputs(5348) <= not(inputs(90));
    layer0_outputs(5349) <= inputs(200);
    layer0_outputs(5350) <= inputs(162);
    layer0_outputs(5351) <= not(inputs(213)) or (inputs(157));
    layer0_outputs(5352) <= not((inputs(109)) or (inputs(92)));
    layer0_outputs(5353) <= (inputs(222)) and not (inputs(241));
    layer0_outputs(5354) <= inputs(49);
    layer0_outputs(5355) <= inputs(94);
    layer0_outputs(5356) <= not((inputs(28)) and (inputs(26)));
    layer0_outputs(5357) <= not((inputs(51)) xor (inputs(69)));
    layer0_outputs(5358) <= inputs(212);
    layer0_outputs(5359) <= (inputs(19)) or (inputs(58));
    layer0_outputs(5360) <= not(inputs(249));
    layer0_outputs(5361) <= inputs(202);
    layer0_outputs(5362) <= (inputs(166)) and not (inputs(114));
    layer0_outputs(5363) <= not(inputs(181));
    layer0_outputs(5364) <= not(inputs(232));
    layer0_outputs(5365) <= not(inputs(115));
    layer0_outputs(5366) <= '1';
    layer0_outputs(5367) <= (inputs(1)) or (inputs(43));
    layer0_outputs(5368) <= not(inputs(202));
    layer0_outputs(5369) <= inputs(229);
    layer0_outputs(5370) <= (inputs(93)) and not (inputs(75));
    layer0_outputs(5371) <= not(inputs(92));
    layer0_outputs(5372) <= not((inputs(27)) or (inputs(140)));
    layer0_outputs(5373) <= not(inputs(201));
    layer0_outputs(5374) <= '1';
    layer0_outputs(5375) <= not(inputs(255)) or (inputs(129));
    layer0_outputs(5376) <= not(inputs(13)) or (inputs(106));
    layer0_outputs(5377) <= not((inputs(148)) or (inputs(180)));
    layer0_outputs(5378) <= (inputs(140)) or (inputs(129));
    layer0_outputs(5379) <= not(inputs(9));
    layer0_outputs(5380) <= not((inputs(105)) or (inputs(88)));
    layer0_outputs(5381) <= not((inputs(88)) or (inputs(247)));
    layer0_outputs(5382) <= not(inputs(26));
    layer0_outputs(5383) <= not((inputs(233)) or (inputs(79)));
    layer0_outputs(5384) <= not(inputs(247)) or (inputs(51));
    layer0_outputs(5385) <= (inputs(52)) xor (inputs(239));
    layer0_outputs(5386) <= not((inputs(227)) or (inputs(167)));
    layer0_outputs(5387) <= inputs(113);
    layer0_outputs(5388) <= not(inputs(37)) or (inputs(49));
    layer0_outputs(5389) <= (inputs(209)) and not (inputs(147));
    layer0_outputs(5390) <= '0';
    layer0_outputs(5391) <= not(inputs(83));
    layer0_outputs(5392) <= not((inputs(235)) or (inputs(147)));
    layer0_outputs(5393) <= inputs(141);
    layer0_outputs(5394) <= (inputs(9)) or (inputs(49));
    layer0_outputs(5395) <= not(inputs(85));
    layer0_outputs(5396) <= (inputs(33)) and not (inputs(77));
    layer0_outputs(5397) <= not(inputs(115));
    layer0_outputs(5398) <= (inputs(98)) or (inputs(100));
    layer0_outputs(5399) <= (inputs(56)) and not (inputs(116));
    layer0_outputs(5400) <= not(inputs(25));
    layer0_outputs(5401) <= (inputs(54)) and not (inputs(166));
    layer0_outputs(5402) <= not((inputs(46)) or (inputs(208)));
    layer0_outputs(5403) <= (inputs(27)) and not (inputs(157));
    layer0_outputs(5404) <= not(inputs(113)) or (inputs(221));
    layer0_outputs(5405) <= not(inputs(54)) or (inputs(253));
    layer0_outputs(5406) <= not((inputs(177)) and (inputs(249)));
    layer0_outputs(5407) <= not((inputs(81)) xor (inputs(186)));
    layer0_outputs(5408) <= not(inputs(121));
    layer0_outputs(5409) <= (inputs(97)) and (inputs(171));
    layer0_outputs(5410) <= (inputs(17)) or (inputs(157));
    layer0_outputs(5411) <= not((inputs(116)) or (inputs(14)));
    layer0_outputs(5412) <= (inputs(225)) and (inputs(250));
    layer0_outputs(5413) <= not(inputs(75));
    layer0_outputs(5414) <= inputs(229);
    layer0_outputs(5415) <= inputs(49);
    layer0_outputs(5416) <= not((inputs(70)) or (inputs(171)));
    layer0_outputs(5417) <= not((inputs(14)) or (inputs(61)));
    layer0_outputs(5418) <= not(inputs(34)) or (inputs(208));
    layer0_outputs(5419) <= not((inputs(115)) or (inputs(98)));
    layer0_outputs(5420) <= inputs(60);
    layer0_outputs(5421) <= not((inputs(197)) xor (inputs(115)));
    layer0_outputs(5422) <= (inputs(65)) xor (inputs(151));
    layer0_outputs(5423) <= not((inputs(167)) xor (inputs(50)));
    layer0_outputs(5424) <= not(inputs(189));
    layer0_outputs(5425) <= inputs(13);
    layer0_outputs(5426) <= inputs(191);
    layer0_outputs(5427) <= not(inputs(152)) or (inputs(11));
    layer0_outputs(5428) <= inputs(126);
    layer0_outputs(5429) <= inputs(131);
    layer0_outputs(5430) <= not(inputs(111)) or (inputs(244));
    layer0_outputs(5431) <= (inputs(62)) or (inputs(245));
    layer0_outputs(5432) <= not((inputs(209)) or (inputs(135)));
    layer0_outputs(5433) <= (inputs(93)) xor (inputs(243));
    layer0_outputs(5434) <= (inputs(238)) and not (inputs(105));
    layer0_outputs(5435) <= not(inputs(13)) or (inputs(177));
    layer0_outputs(5436) <= not((inputs(59)) and (inputs(56)));
    layer0_outputs(5437) <= inputs(229);
    layer0_outputs(5438) <= (inputs(81)) or (inputs(100));
    layer0_outputs(5439) <= (inputs(50)) or (inputs(128));
    layer0_outputs(5440) <= not((inputs(155)) and (inputs(169)));
    layer0_outputs(5441) <= not(inputs(235));
    layer0_outputs(5442) <= not((inputs(123)) xor (inputs(247)));
    layer0_outputs(5443) <= '1';
    layer0_outputs(5444) <= (inputs(88)) or (inputs(96));
    layer0_outputs(5445) <= inputs(128);
    layer0_outputs(5446) <= inputs(248);
    layer0_outputs(5447) <= inputs(63);
    layer0_outputs(5448) <= not(inputs(155));
    layer0_outputs(5449) <= not((inputs(152)) xor (inputs(116)));
    layer0_outputs(5450) <= (inputs(53)) and not (inputs(124));
    layer0_outputs(5451) <= (inputs(5)) or (inputs(31));
    layer0_outputs(5452) <= not((inputs(122)) or (inputs(106)));
    layer0_outputs(5453) <= not(inputs(214));
    layer0_outputs(5454) <= not(inputs(25)) or (inputs(204));
    layer0_outputs(5455) <= not((inputs(2)) or (inputs(201)));
    layer0_outputs(5456) <= (inputs(209)) and not (inputs(80));
    layer0_outputs(5457) <= inputs(184);
    layer0_outputs(5458) <= not(inputs(178));
    layer0_outputs(5459) <= not((inputs(223)) or (inputs(44)));
    layer0_outputs(5460) <= (inputs(184)) and (inputs(210));
    layer0_outputs(5461) <= inputs(209);
    layer0_outputs(5462) <= not(inputs(135)) or (inputs(114));
    layer0_outputs(5463) <= not(inputs(120));
    layer0_outputs(5464) <= (inputs(121)) and not (inputs(21));
    layer0_outputs(5465) <= not(inputs(106));
    layer0_outputs(5466) <= not(inputs(135)) or (inputs(110));
    layer0_outputs(5467) <= not((inputs(93)) or (inputs(44)));
    layer0_outputs(5468) <= not(inputs(35)) or (inputs(50));
    layer0_outputs(5469) <= not(inputs(248));
    layer0_outputs(5470) <= not(inputs(25)) or (inputs(9));
    layer0_outputs(5471) <= not(inputs(170));
    layer0_outputs(5472) <= (inputs(220)) and not (inputs(27));
    layer0_outputs(5473) <= not(inputs(7)) or (inputs(133));
    layer0_outputs(5474) <= not(inputs(73)) or (inputs(87));
    layer0_outputs(5475) <= (inputs(161)) and not (inputs(222));
    layer0_outputs(5476) <= not((inputs(118)) or (inputs(112)));
    layer0_outputs(5477) <= not((inputs(112)) or (inputs(15)));
    layer0_outputs(5478) <= not(inputs(21));
    layer0_outputs(5479) <= inputs(178);
    layer0_outputs(5480) <= (inputs(214)) and not (inputs(110));
    layer0_outputs(5481) <= not((inputs(152)) xor (inputs(211)));
    layer0_outputs(5482) <= not(inputs(228));
    layer0_outputs(5483) <= (inputs(221)) xor (inputs(26));
    layer0_outputs(5484) <= not((inputs(165)) or (inputs(67)));
    layer0_outputs(5485) <= not((inputs(161)) or (inputs(194)));
    layer0_outputs(5486) <= (inputs(90)) and not (inputs(81));
    layer0_outputs(5487) <= (inputs(118)) and not (inputs(15));
    layer0_outputs(5488) <= not((inputs(11)) xor (inputs(223)));
    layer0_outputs(5489) <= (inputs(73)) and not (inputs(153));
    layer0_outputs(5490) <= not(inputs(156));
    layer0_outputs(5491) <= not(inputs(158)) or (inputs(239));
    layer0_outputs(5492) <= (inputs(15)) xor (inputs(105));
    layer0_outputs(5493) <= not((inputs(135)) and (inputs(122)));
    layer0_outputs(5494) <= not((inputs(3)) or (inputs(65)));
    layer0_outputs(5495) <= (inputs(170)) or (inputs(205));
    layer0_outputs(5496) <= not((inputs(53)) xor (inputs(65)));
    layer0_outputs(5497) <= not((inputs(11)) or (inputs(75)));
    layer0_outputs(5498) <= (inputs(191)) or (inputs(226));
    layer0_outputs(5499) <= '0';
    layer0_outputs(5500) <= not(inputs(61)) or (inputs(221));
    layer0_outputs(5501) <= (inputs(226)) xor (inputs(23));
    layer0_outputs(5502) <= (inputs(109)) xor (inputs(190));
    layer0_outputs(5503) <= not((inputs(236)) or (inputs(126)));
    layer0_outputs(5504) <= not(inputs(216));
    layer0_outputs(5505) <= not(inputs(255));
    layer0_outputs(5506) <= (inputs(96)) xor (inputs(240));
    layer0_outputs(5507) <= not(inputs(126));
    layer0_outputs(5508) <= (inputs(163)) xor (inputs(165));
    layer0_outputs(5509) <= (inputs(254)) and not (inputs(220));
    layer0_outputs(5510) <= (inputs(194)) and not (inputs(128));
    layer0_outputs(5511) <= (inputs(196)) and not (inputs(94));
    layer0_outputs(5512) <= not(inputs(163));
    layer0_outputs(5513) <= inputs(142);
    layer0_outputs(5514) <= inputs(43);
    layer0_outputs(5515) <= not((inputs(125)) or (inputs(116)));
    layer0_outputs(5516) <= inputs(89);
    layer0_outputs(5517) <= not((inputs(148)) xor (inputs(128)));
    layer0_outputs(5518) <= not((inputs(1)) and (inputs(177)));
    layer0_outputs(5519) <= (inputs(218)) or (inputs(175));
    layer0_outputs(5520) <= '0';
    layer0_outputs(5521) <= not(inputs(203)) or (inputs(39));
    layer0_outputs(5522) <= not((inputs(61)) xor (inputs(74)));
    layer0_outputs(5523) <= not((inputs(135)) or (inputs(39)));
    layer0_outputs(5524) <= not(inputs(46)) or (inputs(203));
    layer0_outputs(5525) <= '0';
    layer0_outputs(5526) <= not(inputs(248));
    layer0_outputs(5527) <= not((inputs(113)) or (inputs(66)));
    layer0_outputs(5528) <= (inputs(23)) and not (inputs(144));
    layer0_outputs(5529) <= (inputs(45)) or (inputs(230));
    layer0_outputs(5530) <= (inputs(167)) and not (inputs(206));
    layer0_outputs(5531) <= '1';
    layer0_outputs(5532) <= not(inputs(186)) or (inputs(231));
    layer0_outputs(5533) <= not((inputs(44)) or (inputs(154)));
    layer0_outputs(5534) <= '0';
    layer0_outputs(5535) <= (inputs(70)) and not (inputs(163));
    layer0_outputs(5536) <= not(inputs(148));
    layer0_outputs(5537) <= not(inputs(207));
    layer0_outputs(5538) <= (inputs(184)) and not (inputs(130));
    layer0_outputs(5539) <= not(inputs(38));
    layer0_outputs(5540) <= (inputs(145)) and not (inputs(207));
    layer0_outputs(5541) <= not(inputs(209)) or (inputs(14));
    layer0_outputs(5542) <= not((inputs(74)) or (inputs(212)));
    layer0_outputs(5543) <= (inputs(221)) xor (inputs(126));
    layer0_outputs(5544) <= (inputs(143)) xor (inputs(92));
    layer0_outputs(5545) <= not((inputs(123)) or (inputs(176)));
    layer0_outputs(5546) <= inputs(71);
    layer0_outputs(5547) <= (inputs(168)) and not (inputs(177));
    layer0_outputs(5548) <= not((inputs(205)) or (inputs(246)));
    layer0_outputs(5549) <= (inputs(177)) xor (inputs(252));
    layer0_outputs(5550) <= inputs(233);
    layer0_outputs(5551) <= not(inputs(115)) or (inputs(207));
    layer0_outputs(5552) <= not(inputs(113));
    layer0_outputs(5553) <= not((inputs(197)) or (inputs(255)));
    layer0_outputs(5554) <= not(inputs(33)) or (inputs(111));
    layer0_outputs(5555) <= not((inputs(132)) or (inputs(240)));
    layer0_outputs(5556) <= not(inputs(215));
    layer0_outputs(5557) <= not(inputs(208));
    layer0_outputs(5558) <= inputs(138);
    layer0_outputs(5559) <= (inputs(14)) or (inputs(192));
    layer0_outputs(5560) <= inputs(167);
    layer0_outputs(5561) <= inputs(167);
    layer0_outputs(5562) <= (inputs(63)) and not (inputs(248));
    layer0_outputs(5563) <= not(inputs(51));
    layer0_outputs(5564) <= not((inputs(197)) and (inputs(153)));
    layer0_outputs(5565) <= not(inputs(118));
    layer0_outputs(5566) <= (inputs(62)) and not (inputs(36));
    layer0_outputs(5567) <= (inputs(208)) or (inputs(13));
    layer0_outputs(5568) <= inputs(178);
    layer0_outputs(5569) <= not(inputs(250)) or (inputs(10));
    layer0_outputs(5570) <= not((inputs(172)) and (inputs(12)));
    layer0_outputs(5571) <= not(inputs(241)) or (inputs(198));
    layer0_outputs(5572) <= (inputs(188)) or (inputs(87));
    layer0_outputs(5573) <= not(inputs(43));
    layer0_outputs(5574) <= not((inputs(235)) or (inputs(38)));
    layer0_outputs(5575) <= (inputs(59)) and not (inputs(91));
    layer0_outputs(5576) <= (inputs(254)) and not (inputs(47));
    layer0_outputs(5577) <= not((inputs(119)) or (inputs(47)));
    layer0_outputs(5578) <= not(inputs(88));
    layer0_outputs(5579) <= not(inputs(232));
    layer0_outputs(5580) <= not(inputs(45));
    layer0_outputs(5581) <= inputs(119);
    layer0_outputs(5582) <= not(inputs(111));
    layer0_outputs(5583) <= inputs(171);
    layer0_outputs(5584) <= not((inputs(69)) or (inputs(78)));
    layer0_outputs(5585) <= not((inputs(102)) or (inputs(248)));
    layer0_outputs(5586) <= not(inputs(109)) or (inputs(42));
    layer0_outputs(5587) <= not(inputs(122));
    layer0_outputs(5588) <= (inputs(118)) and not (inputs(109));
    layer0_outputs(5589) <= inputs(146);
    layer0_outputs(5590) <= not((inputs(138)) and (inputs(246)));
    layer0_outputs(5591) <= not((inputs(47)) xor (inputs(29)));
    layer0_outputs(5592) <= not(inputs(7));
    layer0_outputs(5593) <= (inputs(113)) and not (inputs(105));
    layer0_outputs(5594) <= not(inputs(183));
    layer0_outputs(5595) <= (inputs(237)) or (inputs(218));
    layer0_outputs(5596) <= (inputs(122)) and not (inputs(223));
    layer0_outputs(5597) <= not((inputs(217)) and (inputs(251)));
    layer0_outputs(5598) <= not((inputs(148)) xor (inputs(102)));
    layer0_outputs(5599) <= (inputs(182)) and (inputs(199));
    layer0_outputs(5600) <= (inputs(78)) or (inputs(7));
    layer0_outputs(5601) <= (inputs(81)) and not (inputs(150));
    layer0_outputs(5602) <= not((inputs(140)) or (inputs(172)));
    layer0_outputs(5603) <= (inputs(161)) and not (inputs(16));
    layer0_outputs(5604) <= inputs(53);
    layer0_outputs(5605) <= inputs(220);
    layer0_outputs(5606) <= inputs(163);
    layer0_outputs(5607) <= not((inputs(205)) xor (inputs(206)));
    layer0_outputs(5608) <= not(inputs(27)) or (inputs(54));
    layer0_outputs(5609) <= not(inputs(226));
    layer0_outputs(5610) <= inputs(97);
    layer0_outputs(5611) <= not(inputs(152)) or (inputs(85));
    layer0_outputs(5612) <= not((inputs(96)) or (inputs(80)));
    layer0_outputs(5613) <= not(inputs(242));
    layer0_outputs(5614) <= (inputs(18)) or (inputs(199));
    layer0_outputs(5615) <= not(inputs(157));
    layer0_outputs(5616) <= (inputs(4)) or (inputs(213));
    layer0_outputs(5617) <= (inputs(217)) and not (inputs(34));
    layer0_outputs(5618) <= not((inputs(94)) or (inputs(22)));
    layer0_outputs(5619) <= (inputs(239)) and (inputs(215));
    layer0_outputs(5620) <= (inputs(3)) xor (inputs(42));
    layer0_outputs(5621) <= not(inputs(174)) or (inputs(254));
    layer0_outputs(5622) <= not(inputs(203)) or (inputs(15));
    layer0_outputs(5623) <= not(inputs(131));
    layer0_outputs(5624) <= inputs(225);
    layer0_outputs(5625) <= not(inputs(100));
    layer0_outputs(5626) <= not((inputs(0)) xor (inputs(53)));
    layer0_outputs(5627) <= not(inputs(239));
    layer0_outputs(5628) <= not(inputs(68));
    layer0_outputs(5629) <= (inputs(168)) xor (inputs(217));
    layer0_outputs(5630) <= (inputs(122)) or (inputs(189));
    layer0_outputs(5631) <= inputs(206);
    layer0_outputs(5632) <= not(inputs(133)) or (inputs(79));
    layer0_outputs(5633) <= (inputs(134)) xor (inputs(92));
    layer0_outputs(5634) <= not(inputs(169)) or (inputs(145));
    layer0_outputs(5635) <= (inputs(79)) and not (inputs(225));
    layer0_outputs(5636) <= (inputs(44)) and not (inputs(239));
    layer0_outputs(5637) <= not((inputs(159)) xor (inputs(86)));
    layer0_outputs(5638) <= not(inputs(20)) or (inputs(52));
    layer0_outputs(5639) <= inputs(162);
    layer0_outputs(5640) <= not(inputs(64)) or (inputs(203));
    layer0_outputs(5641) <= (inputs(196)) and not (inputs(251));
    layer0_outputs(5642) <= (inputs(107)) and (inputs(96));
    layer0_outputs(5643) <= not((inputs(145)) xor (inputs(228)));
    layer0_outputs(5644) <= (inputs(117)) or (inputs(173));
    layer0_outputs(5645) <= not(inputs(197));
    layer0_outputs(5646) <= (inputs(133)) and not (inputs(225));
    layer0_outputs(5647) <= (inputs(178)) xor (inputs(135));
    layer0_outputs(5648) <= inputs(155);
    layer0_outputs(5649) <= not(inputs(147)) or (inputs(174));
    layer0_outputs(5650) <= (inputs(125)) and not (inputs(83));
    layer0_outputs(5651) <= (inputs(144)) and (inputs(72));
    layer0_outputs(5652) <= '1';
    layer0_outputs(5653) <= not(inputs(133)) or (inputs(172));
    layer0_outputs(5654) <= not(inputs(94));
    layer0_outputs(5655) <= (inputs(165)) and not (inputs(9));
    layer0_outputs(5656) <= not((inputs(122)) or (inputs(32)));
    layer0_outputs(5657) <= (inputs(188)) or (inputs(196));
    layer0_outputs(5658) <= not((inputs(67)) or (inputs(129)));
    layer0_outputs(5659) <= inputs(186);
    layer0_outputs(5660) <= not(inputs(52));
    layer0_outputs(5661) <= not(inputs(151));
    layer0_outputs(5662) <= (inputs(155)) and (inputs(2));
    layer0_outputs(5663) <= not(inputs(195));
    layer0_outputs(5664) <= (inputs(9)) or (inputs(212));
    layer0_outputs(5665) <= inputs(98);
    layer0_outputs(5666) <= not(inputs(155));
    layer0_outputs(5667) <= not(inputs(56));
    layer0_outputs(5668) <= inputs(213);
    layer0_outputs(5669) <= (inputs(112)) and not (inputs(206));
    layer0_outputs(5670) <= (inputs(152)) xor (inputs(17));
    layer0_outputs(5671) <= (inputs(0)) and not (inputs(166));
    layer0_outputs(5672) <= inputs(113);
    layer0_outputs(5673) <= not(inputs(212));
    layer0_outputs(5674) <= inputs(161);
    layer0_outputs(5675) <= '0';
    layer0_outputs(5676) <= inputs(129);
    layer0_outputs(5677) <= not(inputs(80));
    layer0_outputs(5678) <= inputs(30);
    layer0_outputs(5679) <= (inputs(130)) and not (inputs(59));
    layer0_outputs(5680) <= (inputs(207)) and not (inputs(5));
    layer0_outputs(5681) <= not((inputs(217)) xor (inputs(19)));
    layer0_outputs(5682) <= not(inputs(94));
    layer0_outputs(5683) <= '1';
    layer0_outputs(5684) <= not(inputs(37));
    layer0_outputs(5685) <= (inputs(29)) and (inputs(220));
    layer0_outputs(5686) <= '0';
    layer0_outputs(5687) <= not(inputs(101));
    layer0_outputs(5688) <= (inputs(87)) and not (inputs(158));
    layer0_outputs(5689) <= (inputs(161)) or (inputs(193));
    layer0_outputs(5690) <= '0';
    layer0_outputs(5691) <= (inputs(193)) and not (inputs(205));
    layer0_outputs(5692) <= '0';
    layer0_outputs(5693) <= (inputs(71)) or (inputs(236));
    layer0_outputs(5694) <= (inputs(31)) xor (inputs(119));
    layer0_outputs(5695) <= not(inputs(10));
    layer0_outputs(5696) <= (inputs(10)) xor (inputs(41));
    layer0_outputs(5697) <= not((inputs(26)) xor (inputs(64)));
    layer0_outputs(5698) <= (inputs(197)) xor (inputs(243));
    layer0_outputs(5699) <= (inputs(253)) or (inputs(132));
    layer0_outputs(5700) <= not((inputs(49)) xor (inputs(165)));
    layer0_outputs(5701) <= not((inputs(146)) or (inputs(136)));
    layer0_outputs(5702) <= (inputs(77)) xor (inputs(181));
    layer0_outputs(5703) <= (inputs(129)) or (inputs(62));
    layer0_outputs(5704) <= (inputs(8)) and not (inputs(66));
    layer0_outputs(5705) <= (inputs(90)) and not (inputs(229));
    layer0_outputs(5706) <= not(inputs(98)) or (inputs(55));
    layer0_outputs(5707) <= (inputs(126)) and not (inputs(40));
    layer0_outputs(5708) <= (inputs(107)) or (inputs(191));
    layer0_outputs(5709) <= not(inputs(206)) or (inputs(242));
    layer0_outputs(5710) <= not((inputs(7)) xor (inputs(254)));
    layer0_outputs(5711) <= (inputs(19)) or (inputs(195));
    layer0_outputs(5712) <= not((inputs(148)) or (inputs(126)));
    layer0_outputs(5713) <= inputs(62);
    layer0_outputs(5714) <= (inputs(72)) and not (inputs(0));
    layer0_outputs(5715) <= not(inputs(145));
    layer0_outputs(5716) <= not(inputs(77));
    layer0_outputs(5717) <= (inputs(169)) or (inputs(7));
    layer0_outputs(5718) <= not(inputs(105)) or (inputs(192));
    layer0_outputs(5719) <= not(inputs(107));
    layer0_outputs(5720) <= not(inputs(78));
    layer0_outputs(5721) <= inputs(206);
    layer0_outputs(5722) <= not(inputs(87));
    layer0_outputs(5723) <= (inputs(206)) or (inputs(116));
    layer0_outputs(5724) <= not((inputs(166)) xor (inputs(227)));
    layer0_outputs(5725) <= inputs(251);
    layer0_outputs(5726) <= not(inputs(125));
    layer0_outputs(5727) <= not(inputs(190));
    layer0_outputs(5728) <= not(inputs(218)) or (inputs(105));
    layer0_outputs(5729) <= not(inputs(230));
    layer0_outputs(5730) <= not(inputs(192));
    layer0_outputs(5731) <= (inputs(10)) or (inputs(26));
    layer0_outputs(5732) <= inputs(208);
    layer0_outputs(5733) <= inputs(210);
    layer0_outputs(5734) <= inputs(136);
    layer0_outputs(5735) <= inputs(52);
    layer0_outputs(5736) <= not(inputs(74)) or (inputs(248));
    layer0_outputs(5737) <= (inputs(33)) xor (inputs(154));
    layer0_outputs(5738) <= not((inputs(148)) or (inputs(112)));
    layer0_outputs(5739) <= (inputs(87)) xor (inputs(9));
    layer0_outputs(5740) <= (inputs(118)) xor (inputs(134));
    layer0_outputs(5741) <= (inputs(166)) and not (inputs(17));
    layer0_outputs(5742) <= not(inputs(113));
    layer0_outputs(5743) <= not(inputs(174));
    layer0_outputs(5744) <= (inputs(231)) and not (inputs(0));
    layer0_outputs(5745) <= inputs(118);
    layer0_outputs(5746) <= not((inputs(43)) xor (inputs(58)));
    layer0_outputs(5747) <= not((inputs(148)) or (inputs(191)));
    layer0_outputs(5748) <= (inputs(212)) and not (inputs(113));
    layer0_outputs(5749) <= (inputs(29)) and not (inputs(110));
    layer0_outputs(5750) <= not(inputs(120)) or (inputs(180));
    layer0_outputs(5751) <= '1';
    layer0_outputs(5752) <= (inputs(213)) and not (inputs(117));
    layer0_outputs(5753) <= not((inputs(5)) or (inputs(55)));
    layer0_outputs(5754) <= not((inputs(183)) or (inputs(230)));
    layer0_outputs(5755) <= inputs(75);
    layer0_outputs(5756) <= (inputs(71)) and not (inputs(134));
    layer0_outputs(5757) <= not(inputs(149));
    layer0_outputs(5758) <= (inputs(195)) and not (inputs(125));
    layer0_outputs(5759) <= not(inputs(196));
    layer0_outputs(5760) <= (inputs(221)) and not (inputs(113));
    layer0_outputs(5761) <= (inputs(134)) and not (inputs(239));
    layer0_outputs(5762) <= not(inputs(14)) or (inputs(58));
    layer0_outputs(5763) <= (inputs(164)) and not (inputs(220));
    layer0_outputs(5764) <= (inputs(7)) and not (inputs(97));
    layer0_outputs(5765) <= (inputs(86)) or (inputs(226));
    layer0_outputs(5766) <= not(inputs(51)) or (inputs(87));
    layer0_outputs(5767) <= not(inputs(71));
    layer0_outputs(5768) <= not(inputs(13));
    layer0_outputs(5769) <= not((inputs(53)) or (inputs(100)));
    layer0_outputs(5770) <= not(inputs(249));
    layer0_outputs(5771) <= (inputs(31)) or (inputs(166));
    layer0_outputs(5772) <= inputs(164);
    layer0_outputs(5773) <= not(inputs(133));
    layer0_outputs(5774) <= not(inputs(19)) or (inputs(63));
    layer0_outputs(5775) <= inputs(102);
    layer0_outputs(5776) <= not(inputs(250));
    layer0_outputs(5777) <= inputs(84);
    layer0_outputs(5778) <= inputs(187);
    layer0_outputs(5779) <= (inputs(190)) and not (inputs(254));
    layer0_outputs(5780) <= not((inputs(55)) and (inputs(75)));
    layer0_outputs(5781) <= (inputs(157)) and not (inputs(207));
    layer0_outputs(5782) <= not(inputs(120));
    layer0_outputs(5783) <= not((inputs(71)) xor (inputs(133)));
    layer0_outputs(5784) <= inputs(234);
    layer0_outputs(5785) <= not(inputs(23));
    layer0_outputs(5786) <= not((inputs(213)) and (inputs(81)));
    layer0_outputs(5787) <= '0';
    layer0_outputs(5788) <= inputs(212);
    layer0_outputs(5789) <= not((inputs(141)) or (inputs(129)));
    layer0_outputs(5790) <= '0';
    layer0_outputs(5791) <= not(inputs(246)) or (inputs(241));
    layer0_outputs(5792) <= (inputs(238)) or (inputs(166));
    layer0_outputs(5793) <= (inputs(48)) or (inputs(39));
    layer0_outputs(5794) <= (inputs(216)) and not (inputs(230));
    layer0_outputs(5795) <= inputs(189);
    layer0_outputs(5796) <= not(inputs(52));
    layer0_outputs(5797) <= '1';
    layer0_outputs(5798) <= not(inputs(8));
    layer0_outputs(5799) <= (inputs(245)) and not (inputs(25));
    layer0_outputs(5800) <= (inputs(198)) and not (inputs(186));
    layer0_outputs(5801) <= not(inputs(156));
    layer0_outputs(5802) <= (inputs(78)) or (inputs(59));
    layer0_outputs(5803) <= not((inputs(140)) and (inputs(86)));
    layer0_outputs(5804) <= not((inputs(194)) or (inputs(232)));
    layer0_outputs(5805) <= '1';
    layer0_outputs(5806) <= not(inputs(146));
    layer0_outputs(5807) <= not((inputs(142)) or (inputs(243)));
    layer0_outputs(5808) <= inputs(22);
    layer0_outputs(5809) <= (inputs(58)) and not (inputs(123));
    layer0_outputs(5810) <= not(inputs(122));
    layer0_outputs(5811) <= (inputs(77)) and (inputs(125));
    layer0_outputs(5812) <= (inputs(203)) xor (inputs(235));
    layer0_outputs(5813) <= '0';
    layer0_outputs(5814) <= (inputs(199)) and not (inputs(30));
    layer0_outputs(5815) <= (inputs(228)) and not (inputs(94));
    layer0_outputs(5816) <= not(inputs(61));
    layer0_outputs(5817) <= inputs(160);
    layer0_outputs(5818) <= (inputs(58)) xor (inputs(11));
    layer0_outputs(5819) <= not(inputs(203)) or (inputs(29));
    layer0_outputs(5820) <= not(inputs(114));
    layer0_outputs(5821) <= '1';
    layer0_outputs(5822) <= (inputs(2)) or (inputs(94));
    layer0_outputs(5823) <= not((inputs(180)) or (inputs(80)));
    layer0_outputs(5824) <= not((inputs(148)) xor (inputs(136)));
    layer0_outputs(5825) <= not(inputs(94));
    layer0_outputs(5826) <= inputs(72);
    layer0_outputs(5827) <= inputs(55);
    layer0_outputs(5828) <= inputs(229);
    layer0_outputs(5829) <= not(inputs(57));
    layer0_outputs(5830) <= (inputs(29)) or (inputs(113));
    layer0_outputs(5831) <= inputs(123);
    layer0_outputs(5832) <= not(inputs(155)) or (inputs(29));
    layer0_outputs(5833) <= (inputs(43)) or (inputs(185));
    layer0_outputs(5834) <= not((inputs(177)) or (inputs(127)));
    layer0_outputs(5835) <= not((inputs(164)) or (inputs(185)));
    layer0_outputs(5836) <= not(inputs(183));
    layer0_outputs(5837) <= (inputs(152)) and not (inputs(192));
    layer0_outputs(5838) <= not((inputs(21)) xor (inputs(177)));
    layer0_outputs(5839) <= (inputs(18)) xor (inputs(128));
    layer0_outputs(5840) <= (inputs(96)) or (inputs(99));
    layer0_outputs(5841) <= not(inputs(116));
    layer0_outputs(5842) <= '0';
    layer0_outputs(5843) <= not(inputs(183)) or (inputs(56));
    layer0_outputs(5844) <= not(inputs(119)) or (inputs(143));
    layer0_outputs(5845) <= (inputs(182)) and not (inputs(30));
    layer0_outputs(5846) <= (inputs(178)) and not (inputs(5));
    layer0_outputs(5847) <= not(inputs(221)) or (inputs(124));
    layer0_outputs(5848) <= not(inputs(60));
    layer0_outputs(5849) <= inputs(105);
    layer0_outputs(5850) <= not((inputs(180)) xor (inputs(228)));
    layer0_outputs(5851) <= not(inputs(142));
    layer0_outputs(5852) <= (inputs(107)) and not (inputs(116));
    layer0_outputs(5853) <= inputs(45);
    layer0_outputs(5854) <= (inputs(18)) or (inputs(106));
    layer0_outputs(5855) <= inputs(198);
    layer0_outputs(5856) <= inputs(115);
    layer0_outputs(5857) <= not(inputs(217)) or (inputs(140));
    layer0_outputs(5858) <= not(inputs(24)) or (inputs(243));
    layer0_outputs(5859) <= inputs(83);
    layer0_outputs(5860) <= not(inputs(226));
    layer0_outputs(5861) <= not((inputs(240)) or (inputs(168)));
    layer0_outputs(5862) <= (inputs(155)) and not (inputs(244));
    layer0_outputs(5863) <= (inputs(59)) or (inputs(75));
    layer0_outputs(5864) <= (inputs(37)) and (inputs(152));
    layer0_outputs(5865) <= not((inputs(94)) or (inputs(66)));
    layer0_outputs(5866) <= inputs(251);
    layer0_outputs(5867) <= not((inputs(240)) or (inputs(225)));
    layer0_outputs(5868) <= not((inputs(22)) or (inputs(49)));
    layer0_outputs(5869) <= not(inputs(20));
    layer0_outputs(5870) <= inputs(200);
    layer0_outputs(5871) <= not((inputs(142)) xor (inputs(3)));
    layer0_outputs(5872) <= (inputs(161)) and not (inputs(48));
    layer0_outputs(5873) <= not((inputs(30)) xor (inputs(110)));
    layer0_outputs(5874) <= not((inputs(254)) or (inputs(36)));
    layer0_outputs(5875) <= (inputs(139)) and not (inputs(241));
    layer0_outputs(5876) <= not((inputs(108)) and (inputs(57)));
    layer0_outputs(5877) <= not(inputs(70)) or (inputs(94));
    layer0_outputs(5878) <= not(inputs(231)) or (inputs(16));
    layer0_outputs(5879) <= (inputs(24)) and not (inputs(81));
    layer0_outputs(5880) <= not(inputs(246)) or (inputs(96));
    layer0_outputs(5881) <= (inputs(175)) or (inputs(164));
    layer0_outputs(5882) <= inputs(246);
    layer0_outputs(5883) <= inputs(70);
    layer0_outputs(5884) <= not(inputs(53)) or (inputs(72));
    layer0_outputs(5885) <= (inputs(35)) or (inputs(23));
    layer0_outputs(5886) <= inputs(135);
    layer0_outputs(5887) <= not((inputs(109)) or (inputs(193)));
    layer0_outputs(5888) <= not((inputs(99)) or (inputs(98)));
    layer0_outputs(5889) <= not((inputs(81)) xor (inputs(168)));
    layer0_outputs(5890) <= not(inputs(131)) or (inputs(58));
    layer0_outputs(5891) <= (inputs(235)) and not (inputs(185));
    layer0_outputs(5892) <= not((inputs(63)) or (inputs(135)));
    layer0_outputs(5893) <= (inputs(74)) or (inputs(78));
    layer0_outputs(5894) <= not(inputs(159)) or (inputs(250));
    layer0_outputs(5895) <= inputs(123);
    layer0_outputs(5896) <= not(inputs(164)) or (inputs(92));
    layer0_outputs(5897) <= not((inputs(93)) xor (inputs(17)));
    layer0_outputs(5898) <= not((inputs(214)) or (inputs(231)));
    layer0_outputs(5899) <= (inputs(35)) xor (inputs(52));
    layer0_outputs(5900) <= inputs(133);
    layer0_outputs(5901) <= '1';
    layer0_outputs(5902) <= not(inputs(168));
    layer0_outputs(5903) <= (inputs(226)) or (inputs(72));
    layer0_outputs(5904) <= (inputs(163)) and not (inputs(150));
    layer0_outputs(5905) <= not(inputs(159)) or (inputs(166));
    layer0_outputs(5906) <= not(inputs(226)) or (inputs(164));
    layer0_outputs(5907) <= not((inputs(218)) or (inputs(158)));
    layer0_outputs(5908) <= not(inputs(195));
    layer0_outputs(5909) <= (inputs(177)) or (inputs(208));
    layer0_outputs(5910) <= not(inputs(193)) or (inputs(120));
    layer0_outputs(5911) <= not((inputs(23)) xor (inputs(54)));
    layer0_outputs(5912) <= not((inputs(85)) or (inputs(140)));
    layer0_outputs(5913) <= (inputs(114)) or (inputs(101));
    layer0_outputs(5914) <= inputs(148);
    layer0_outputs(5915) <= inputs(164);
    layer0_outputs(5916) <= inputs(232);
    layer0_outputs(5917) <= inputs(92);
    layer0_outputs(5918) <= '1';
    layer0_outputs(5919) <= inputs(85);
    layer0_outputs(5920) <= not(inputs(139));
    layer0_outputs(5921) <= (inputs(158)) xor (inputs(90));
    layer0_outputs(5922) <= (inputs(178)) and not (inputs(61));
    layer0_outputs(5923) <= inputs(203);
    layer0_outputs(5924) <= not(inputs(94));
    layer0_outputs(5925) <= not(inputs(28)) or (inputs(239));
    layer0_outputs(5926) <= '0';
    layer0_outputs(5927) <= not(inputs(115));
    layer0_outputs(5928) <= inputs(232);
    layer0_outputs(5929) <= (inputs(233)) and (inputs(121));
    layer0_outputs(5930) <= (inputs(70)) and not (inputs(9));
    layer0_outputs(5931) <= (inputs(155)) and not (inputs(120));
    layer0_outputs(5932) <= not(inputs(129));
    layer0_outputs(5933) <= not(inputs(232));
    layer0_outputs(5934) <= inputs(226);
    layer0_outputs(5935) <= (inputs(49)) or (inputs(169));
    layer0_outputs(5936) <= not(inputs(169));
    layer0_outputs(5937) <= inputs(132);
    layer0_outputs(5938) <= (inputs(252)) and not (inputs(221));
    layer0_outputs(5939) <= (inputs(215)) and (inputs(252));
    layer0_outputs(5940) <= (inputs(187)) and not (inputs(62));
    layer0_outputs(5941) <= '0';
    layer0_outputs(5942) <= (inputs(87)) and not (inputs(167));
    layer0_outputs(5943) <= not(inputs(41));
    layer0_outputs(5944) <= (inputs(58)) or (inputs(34));
    layer0_outputs(5945) <= not(inputs(99));
    layer0_outputs(5946) <= (inputs(146)) and (inputs(254));
    layer0_outputs(5947) <= not((inputs(232)) or (inputs(226)));
    layer0_outputs(5948) <= not((inputs(242)) and (inputs(183)));
    layer0_outputs(5949) <= not(inputs(236)) or (inputs(41));
    layer0_outputs(5950) <= (inputs(223)) or (inputs(183));
    layer0_outputs(5951) <= (inputs(110)) xor (inputs(196));
    layer0_outputs(5952) <= (inputs(84)) and not (inputs(95));
    layer0_outputs(5953) <= inputs(106);
    layer0_outputs(5954) <= inputs(178);
    layer0_outputs(5955) <= (inputs(148)) and not (inputs(240));
    layer0_outputs(5956) <= (inputs(233)) and not (inputs(155));
    layer0_outputs(5957) <= '0';
    layer0_outputs(5958) <= (inputs(114)) and (inputs(228));
    layer0_outputs(5959) <= not(inputs(238));
    layer0_outputs(5960) <= (inputs(137)) xor (inputs(105));
    layer0_outputs(5961) <= not(inputs(43));
    layer0_outputs(5962) <= (inputs(249)) xor (inputs(0));
    layer0_outputs(5963) <= not(inputs(9));
    layer0_outputs(5964) <= inputs(7);
    layer0_outputs(5965) <= not((inputs(83)) and (inputs(90)));
    layer0_outputs(5966) <= not((inputs(59)) or (inputs(114)));
    layer0_outputs(5967) <= not((inputs(68)) xor (inputs(20)));
    layer0_outputs(5968) <= (inputs(132)) and not (inputs(7));
    layer0_outputs(5969) <= inputs(237);
    layer0_outputs(5970) <= (inputs(252)) and not (inputs(8));
    layer0_outputs(5971) <= not((inputs(134)) xor (inputs(255)));
    layer0_outputs(5972) <= (inputs(221)) xor (inputs(72));
    layer0_outputs(5973) <= (inputs(36)) or (inputs(62));
    layer0_outputs(5974) <= inputs(234);
    layer0_outputs(5975) <= not(inputs(245));
    layer0_outputs(5976) <= not(inputs(205));
    layer0_outputs(5977) <= inputs(212);
    layer0_outputs(5978) <= not(inputs(43)) or (inputs(181));
    layer0_outputs(5979) <= inputs(143);
    layer0_outputs(5980) <= (inputs(18)) and not (inputs(190));
    layer0_outputs(5981) <= not((inputs(170)) or (inputs(176)));
    layer0_outputs(5982) <= (inputs(219)) xor (inputs(120));
    layer0_outputs(5983) <= not(inputs(123)) or (inputs(83));
    layer0_outputs(5984) <= inputs(57);
    layer0_outputs(5985) <= not((inputs(250)) xor (inputs(46)));
    layer0_outputs(5986) <= (inputs(82)) and not (inputs(16));
    layer0_outputs(5987) <= (inputs(88)) or (inputs(205));
    layer0_outputs(5988) <= inputs(102);
    layer0_outputs(5989) <= '0';
    layer0_outputs(5990) <= (inputs(50)) xor (inputs(76));
    layer0_outputs(5991) <= not((inputs(168)) xor (inputs(253)));
    layer0_outputs(5992) <= (inputs(231)) and (inputs(203));
    layer0_outputs(5993) <= not(inputs(83));
    layer0_outputs(5994) <= not(inputs(233)) or (inputs(1));
    layer0_outputs(5995) <= not(inputs(3));
    layer0_outputs(5996) <= (inputs(130)) xor (inputs(189));
    layer0_outputs(5997) <= not(inputs(76)) or (inputs(176));
    layer0_outputs(5998) <= (inputs(24)) or (inputs(255));
    layer0_outputs(5999) <= (inputs(22)) and not (inputs(164));
    layer0_outputs(6000) <= (inputs(111)) or (inputs(59));
    layer0_outputs(6001) <= (inputs(43)) and not (inputs(233));
    layer0_outputs(6002) <= (inputs(103)) and not (inputs(2));
    layer0_outputs(6003) <= '1';
    layer0_outputs(6004) <= (inputs(106)) or (inputs(254));
    layer0_outputs(6005) <= not(inputs(215)) or (inputs(104));
    layer0_outputs(6006) <= not(inputs(245));
    layer0_outputs(6007) <= not(inputs(26)) or (inputs(167));
    layer0_outputs(6008) <= not((inputs(207)) xor (inputs(111)));
    layer0_outputs(6009) <= not((inputs(243)) or (inputs(111)));
    layer0_outputs(6010) <= not((inputs(60)) xor (inputs(4)));
    layer0_outputs(6011) <= (inputs(106)) and not (inputs(253));
    layer0_outputs(6012) <= inputs(89);
    layer0_outputs(6013) <= not(inputs(203));
    layer0_outputs(6014) <= inputs(145);
    layer0_outputs(6015) <= not(inputs(61));
    layer0_outputs(6016) <= inputs(98);
    layer0_outputs(6017) <= not(inputs(152)) or (inputs(146));
    layer0_outputs(6018) <= inputs(127);
    layer0_outputs(6019) <= (inputs(150)) and not (inputs(160));
    layer0_outputs(6020) <= (inputs(206)) and not (inputs(13));
    layer0_outputs(6021) <= '1';
    layer0_outputs(6022) <= inputs(189);
    layer0_outputs(6023) <= inputs(58);
    layer0_outputs(6024) <= (inputs(167)) or (inputs(222));
    layer0_outputs(6025) <= not(inputs(146)) or (inputs(1));
    layer0_outputs(6026) <= not(inputs(90)) or (inputs(149));
    layer0_outputs(6027) <= '1';
    layer0_outputs(6028) <= not((inputs(28)) or (inputs(84)));
    layer0_outputs(6029) <= not((inputs(112)) or (inputs(212)));
    layer0_outputs(6030) <= not(inputs(117));
    layer0_outputs(6031) <= (inputs(70)) and not (inputs(192));
    layer0_outputs(6032) <= inputs(45);
    layer0_outputs(6033) <= not((inputs(21)) or (inputs(77)));
    layer0_outputs(6034) <= not((inputs(35)) xor (inputs(66)));
    layer0_outputs(6035) <= (inputs(26)) and (inputs(84));
    layer0_outputs(6036) <= (inputs(124)) and not (inputs(220));
    layer0_outputs(6037) <= inputs(24);
    layer0_outputs(6038) <= not((inputs(131)) or (inputs(176)));
    layer0_outputs(6039) <= not((inputs(133)) xor (inputs(52)));
    layer0_outputs(6040) <= (inputs(99)) or (inputs(145));
    layer0_outputs(6041) <= (inputs(24)) xor (inputs(193));
    layer0_outputs(6042) <= (inputs(106)) and not (inputs(193));
    layer0_outputs(6043) <= not(inputs(27));
    layer0_outputs(6044) <= not(inputs(50));
    layer0_outputs(6045) <= not(inputs(28));
    layer0_outputs(6046) <= not(inputs(199)) or (inputs(220));
    layer0_outputs(6047) <= (inputs(171)) xor (inputs(138));
    layer0_outputs(6048) <= (inputs(155)) or (inputs(140));
    layer0_outputs(6049) <= inputs(74);
    layer0_outputs(6050) <= not((inputs(113)) and (inputs(65)));
    layer0_outputs(6051) <= inputs(73);
    layer0_outputs(6052) <= inputs(78);
    layer0_outputs(6053) <= '1';
    layer0_outputs(6054) <= inputs(40);
    layer0_outputs(6055) <= inputs(98);
    layer0_outputs(6056) <= not((inputs(139)) or (inputs(223)));
    layer0_outputs(6057) <= not((inputs(23)) xor (inputs(39)));
    layer0_outputs(6058) <= not(inputs(19)) or (inputs(253));
    layer0_outputs(6059) <= not(inputs(193));
    layer0_outputs(6060) <= not(inputs(119)) or (inputs(37));
    layer0_outputs(6061) <= inputs(165);
    layer0_outputs(6062) <= (inputs(188)) and (inputs(120));
    layer0_outputs(6063) <= (inputs(232)) or (inputs(161));
    layer0_outputs(6064) <= not(inputs(77));
    layer0_outputs(6065) <= '1';
    layer0_outputs(6066) <= not((inputs(149)) or (inputs(66)));
    layer0_outputs(6067) <= not(inputs(142)) or (inputs(230));
    layer0_outputs(6068) <= not((inputs(184)) or (inputs(216)));
    layer0_outputs(6069) <= not((inputs(73)) xor (inputs(252)));
    layer0_outputs(6070) <= not((inputs(1)) or (inputs(184)));
    layer0_outputs(6071) <= inputs(111);
    layer0_outputs(6072) <= '0';
    layer0_outputs(6073) <= (inputs(138)) or (inputs(251));
    layer0_outputs(6074) <= not((inputs(100)) or (inputs(155)));
    layer0_outputs(6075) <= not(inputs(243)) or (inputs(254));
    layer0_outputs(6076) <= not(inputs(131));
    layer0_outputs(6077) <= not((inputs(237)) or (inputs(149)));
    layer0_outputs(6078) <= not(inputs(102)) or (inputs(239));
    layer0_outputs(6079) <= not((inputs(133)) xor (inputs(103)));
    layer0_outputs(6080) <= '1';
    layer0_outputs(6081) <= not(inputs(235));
    layer0_outputs(6082) <= not((inputs(149)) or (inputs(90)));
    layer0_outputs(6083) <= inputs(113);
    layer0_outputs(6084) <= inputs(181);
    layer0_outputs(6085) <= not((inputs(42)) and (inputs(109)));
    layer0_outputs(6086) <= not(inputs(135));
    layer0_outputs(6087) <= not(inputs(129));
    layer0_outputs(6088) <= (inputs(100)) or (inputs(86));
    layer0_outputs(6089) <= (inputs(83)) and (inputs(89));
    layer0_outputs(6090) <= inputs(112);
    layer0_outputs(6091) <= not((inputs(157)) or (inputs(231)));
    layer0_outputs(6092) <= not((inputs(100)) and (inputs(212)));
    layer0_outputs(6093) <= '0';
    layer0_outputs(6094) <= (inputs(205)) and not (inputs(225));
    layer0_outputs(6095) <= not((inputs(171)) or (inputs(127)));
    layer0_outputs(6096) <= inputs(167);
    layer0_outputs(6097) <= (inputs(120)) and not (inputs(225));
    layer0_outputs(6098) <= not((inputs(217)) or (inputs(194)));
    layer0_outputs(6099) <= not(inputs(29)) or (inputs(147));
    layer0_outputs(6100) <= not((inputs(11)) and (inputs(24)));
    layer0_outputs(6101) <= not((inputs(164)) xor (inputs(146)));
    layer0_outputs(6102) <= not((inputs(213)) or (inputs(205)));
    layer0_outputs(6103) <= (inputs(163)) or (inputs(68));
    layer0_outputs(6104) <= inputs(59);
    layer0_outputs(6105) <= (inputs(85)) or (inputs(52));
    layer0_outputs(6106) <= not(inputs(135));
    layer0_outputs(6107) <= not((inputs(66)) and (inputs(55)));
    layer0_outputs(6108) <= '1';
    layer0_outputs(6109) <= inputs(229);
    layer0_outputs(6110) <= (inputs(76)) or (inputs(127));
    layer0_outputs(6111) <= '0';
    layer0_outputs(6112) <= (inputs(244)) or (inputs(126));
    layer0_outputs(6113) <= (inputs(179)) and not (inputs(222));
    layer0_outputs(6114) <= (inputs(30)) or (inputs(19));
    layer0_outputs(6115) <= (inputs(202)) xor (inputs(236));
    layer0_outputs(6116) <= '1';
    layer0_outputs(6117) <= not(inputs(15));
    layer0_outputs(6118) <= (inputs(216)) or (inputs(107));
    layer0_outputs(6119) <= (inputs(36)) or (inputs(246));
    layer0_outputs(6120) <= not((inputs(26)) or (inputs(174)));
    layer0_outputs(6121) <= not(inputs(215)) or (inputs(91));
    layer0_outputs(6122) <= '1';
    layer0_outputs(6123) <= not(inputs(151)) or (inputs(33));
    layer0_outputs(6124) <= (inputs(66)) and not (inputs(17));
    layer0_outputs(6125) <= '0';
    layer0_outputs(6126) <= not((inputs(197)) or (inputs(75)));
    layer0_outputs(6127) <= (inputs(21)) and not (inputs(97));
    layer0_outputs(6128) <= not(inputs(82));
    layer0_outputs(6129) <= not(inputs(117)) or (inputs(223));
    layer0_outputs(6130) <= (inputs(224)) and (inputs(46));
    layer0_outputs(6131) <= (inputs(4)) and not (inputs(12));
    layer0_outputs(6132) <= not(inputs(100)) or (inputs(74));
    layer0_outputs(6133) <= not((inputs(98)) and (inputs(181)));
    layer0_outputs(6134) <= (inputs(164)) and not (inputs(35));
    layer0_outputs(6135) <= (inputs(149)) or (inputs(57));
    layer0_outputs(6136) <= not((inputs(154)) or (inputs(218)));
    layer0_outputs(6137) <= (inputs(68)) and not (inputs(158));
    layer0_outputs(6138) <= not(inputs(215)) or (inputs(50));
    layer0_outputs(6139) <= inputs(118);
    layer0_outputs(6140) <= not(inputs(121));
    layer0_outputs(6141) <= (inputs(90)) xor (inputs(79));
    layer0_outputs(6142) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(6143) <= not((inputs(28)) and (inputs(42)));
    layer0_outputs(6144) <= inputs(181);
    layer0_outputs(6145) <= (inputs(122)) and not (inputs(32));
    layer0_outputs(6146) <= not(inputs(231));
    layer0_outputs(6147) <= not(inputs(226));
    layer0_outputs(6148) <= not(inputs(60));
    layer0_outputs(6149) <= (inputs(111)) or (inputs(118));
    layer0_outputs(6150) <= (inputs(245)) and not (inputs(51));
    layer0_outputs(6151) <= not(inputs(188)) or (inputs(159));
    layer0_outputs(6152) <= (inputs(58)) or (inputs(45));
    layer0_outputs(6153) <= (inputs(244)) and not (inputs(22));
    layer0_outputs(6154) <= (inputs(202)) or (inputs(96));
    layer0_outputs(6155) <= inputs(244);
    layer0_outputs(6156) <= inputs(105);
    layer0_outputs(6157) <= inputs(139);
    layer0_outputs(6158) <= not((inputs(253)) and (inputs(20)));
    layer0_outputs(6159) <= not((inputs(148)) xor (inputs(157)));
    layer0_outputs(6160) <= not((inputs(200)) or (inputs(118)));
    layer0_outputs(6161) <= (inputs(70)) xor (inputs(84));
    layer0_outputs(6162) <= (inputs(50)) and (inputs(31));
    layer0_outputs(6163) <= inputs(161);
    layer0_outputs(6164) <= inputs(213);
    layer0_outputs(6165) <= not(inputs(104));
    layer0_outputs(6166) <= not(inputs(21));
    layer0_outputs(6167) <= not(inputs(207));
    layer0_outputs(6168) <= not(inputs(227));
    layer0_outputs(6169) <= not(inputs(45)) or (inputs(60));
    layer0_outputs(6170) <= (inputs(178)) and (inputs(104));
    layer0_outputs(6171) <= (inputs(73)) and (inputs(153));
    layer0_outputs(6172) <= (inputs(67)) or (inputs(96));
    layer0_outputs(6173) <= (inputs(154)) or (inputs(202));
    layer0_outputs(6174) <= not(inputs(71));
    layer0_outputs(6175) <= not(inputs(229)) or (inputs(56));
    layer0_outputs(6176) <= not(inputs(104));
    layer0_outputs(6177) <= (inputs(74)) and not (inputs(112));
    layer0_outputs(6178) <= not((inputs(70)) or (inputs(185)));
    layer0_outputs(6179) <= inputs(121);
    layer0_outputs(6180) <= (inputs(133)) and not (inputs(181));
    layer0_outputs(6181) <= '1';
    layer0_outputs(6182) <= '1';
    layer0_outputs(6183) <= (inputs(223)) or (inputs(115));
    layer0_outputs(6184) <= not(inputs(83));
    layer0_outputs(6185) <= inputs(146);
    layer0_outputs(6186) <= not(inputs(133)) or (inputs(218));
    layer0_outputs(6187) <= not(inputs(194)) or (inputs(82));
    layer0_outputs(6188) <= not((inputs(163)) or (inputs(5)));
    layer0_outputs(6189) <= inputs(249);
    layer0_outputs(6190) <= (inputs(73)) or (inputs(43));
    layer0_outputs(6191) <= (inputs(155)) and not (inputs(171));
    layer0_outputs(6192) <= not(inputs(211)) or (inputs(89));
    layer0_outputs(6193) <= '1';
    layer0_outputs(6194) <= (inputs(156)) and (inputs(77));
    layer0_outputs(6195) <= inputs(165);
    layer0_outputs(6196) <= not(inputs(233));
    layer0_outputs(6197) <= not((inputs(255)) or (inputs(53)));
    layer0_outputs(6198) <= '1';
    layer0_outputs(6199) <= (inputs(141)) and not (inputs(154));
    layer0_outputs(6200) <= not(inputs(138));
    layer0_outputs(6201) <= not(inputs(104));
    layer0_outputs(6202) <= inputs(190);
    layer0_outputs(6203) <= (inputs(149)) xor (inputs(172));
    layer0_outputs(6204) <= (inputs(177)) or (inputs(182));
    layer0_outputs(6205) <= not((inputs(160)) or (inputs(249)));
    layer0_outputs(6206) <= not((inputs(156)) and (inputs(90)));
    layer0_outputs(6207) <= (inputs(89)) and not (inputs(249));
    layer0_outputs(6208) <= not((inputs(40)) or (inputs(121)));
    layer0_outputs(6209) <= (inputs(156)) and not (inputs(65));
    layer0_outputs(6210) <= '0';
    layer0_outputs(6211) <= not((inputs(183)) xor (inputs(242)));
    layer0_outputs(6212) <= not((inputs(77)) xor (inputs(37)));
    layer0_outputs(6213) <= not((inputs(37)) or (inputs(85)));
    layer0_outputs(6214) <= not((inputs(178)) xor (inputs(251)));
    layer0_outputs(6215) <= (inputs(39)) xor (inputs(42));
    layer0_outputs(6216) <= not((inputs(31)) xor (inputs(153)));
    layer0_outputs(6217) <= not((inputs(6)) or (inputs(41)));
    layer0_outputs(6218) <= not(inputs(209)) or (inputs(225));
    layer0_outputs(6219) <= not(inputs(46));
    layer0_outputs(6220) <= not((inputs(121)) or (inputs(253)));
    layer0_outputs(6221) <= not(inputs(45));
    layer0_outputs(6222) <= inputs(139);
    layer0_outputs(6223) <= not(inputs(235));
    layer0_outputs(6224) <= not((inputs(164)) or (inputs(38)));
    layer0_outputs(6225) <= not(inputs(123));
    layer0_outputs(6226) <= not(inputs(93)) or (inputs(33));
    layer0_outputs(6227) <= '1';
    layer0_outputs(6228) <= inputs(38);
    layer0_outputs(6229) <= not(inputs(147));
    layer0_outputs(6230) <= '1';
    layer0_outputs(6231) <= (inputs(178)) or (inputs(84));
    layer0_outputs(6232) <= inputs(77);
    layer0_outputs(6233) <= (inputs(228)) xor (inputs(213));
    layer0_outputs(6234) <= not((inputs(66)) or (inputs(97)));
    layer0_outputs(6235) <= not((inputs(178)) or (inputs(149)));
    layer0_outputs(6236) <= '0';
    layer0_outputs(6237) <= not((inputs(6)) or (inputs(44)));
    layer0_outputs(6238) <= (inputs(251)) and not (inputs(50));
    layer0_outputs(6239) <= not((inputs(108)) or (inputs(105)));
    layer0_outputs(6240) <= not((inputs(30)) or (inputs(82)));
    layer0_outputs(6241) <= (inputs(115)) xor (inputs(117));
    layer0_outputs(6242) <= inputs(169);
    layer0_outputs(6243) <= not((inputs(232)) or (inputs(1)));
    layer0_outputs(6244) <= (inputs(24)) or (inputs(216));
    layer0_outputs(6245) <= (inputs(9)) and not (inputs(65));
    layer0_outputs(6246) <= not(inputs(62));
    layer0_outputs(6247) <= inputs(51);
    layer0_outputs(6248) <= (inputs(157)) and not (inputs(240));
    layer0_outputs(6249) <= not(inputs(227)) or (inputs(243));
    layer0_outputs(6250) <= not((inputs(173)) and (inputs(154)));
    layer0_outputs(6251) <= inputs(223);
    layer0_outputs(6252) <= not(inputs(106));
    layer0_outputs(6253) <= (inputs(103)) and not (inputs(0));
    layer0_outputs(6254) <= not(inputs(91));
    layer0_outputs(6255) <= (inputs(106)) xor (inputs(141));
    layer0_outputs(6256) <= (inputs(152)) and not (inputs(176));
    layer0_outputs(6257) <= not(inputs(178));
    layer0_outputs(6258) <= not((inputs(26)) or (inputs(126)));
    layer0_outputs(6259) <= not(inputs(202));
    layer0_outputs(6260) <= (inputs(5)) xor (inputs(50));
    layer0_outputs(6261) <= '0';
    layer0_outputs(6262) <= not(inputs(87)) or (inputs(212));
    layer0_outputs(6263) <= (inputs(47)) and not (inputs(28));
    layer0_outputs(6264) <= not((inputs(8)) or (inputs(165)));
    layer0_outputs(6265) <= not(inputs(219));
    layer0_outputs(6266) <= not(inputs(208));
    layer0_outputs(6267) <= (inputs(135)) and (inputs(85));
    layer0_outputs(6268) <= not((inputs(79)) or (inputs(194)));
    layer0_outputs(6269) <= (inputs(36)) or (inputs(249));
    layer0_outputs(6270) <= not((inputs(217)) xor (inputs(222)));
    layer0_outputs(6271) <= not(inputs(162));
    layer0_outputs(6272) <= '1';
    layer0_outputs(6273) <= (inputs(189)) and not (inputs(254));
    layer0_outputs(6274) <= (inputs(226)) and not (inputs(81));
    layer0_outputs(6275) <= not(inputs(100)) or (inputs(125));
    layer0_outputs(6276) <= not(inputs(23));
    layer0_outputs(6277) <= not(inputs(73));
    layer0_outputs(6278) <= inputs(208);
    layer0_outputs(6279) <= (inputs(35)) or (inputs(239));
    layer0_outputs(6280) <= inputs(233);
    layer0_outputs(6281) <= not((inputs(223)) or (inputs(139)));
    layer0_outputs(6282) <= (inputs(56)) or (inputs(174));
    layer0_outputs(6283) <= not(inputs(35)) or (inputs(51));
    layer0_outputs(6284) <= (inputs(7)) or (inputs(194));
    layer0_outputs(6285) <= (inputs(229)) and not (inputs(58));
    layer0_outputs(6286) <= not(inputs(91));
    layer0_outputs(6287) <= not((inputs(74)) xor (inputs(242)));
    layer0_outputs(6288) <= not(inputs(96)) or (inputs(107));
    layer0_outputs(6289) <= (inputs(229)) and not (inputs(236));
    layer0_outputs(6290) <= (inputs(128)) xor (inputs(49));
    layer0_outputs(6291) <= not((inputs(53)) or (inputs(163)));
    layer0_outputs(6292) <= not((inputs(170)) and (inputs(54)));
    layer0_outputs(6293) <= (inputs(5)) or (inputs(144));
    layer0_outputs(6294) <= not(inputs(181));
    layer0_outputs(6295) <= inputs(28);
    layer0_outputs(6296) <= not((inputs(160)) or (inputs(230)));
    layer0_outputs(6297) <= (inputs(50)) and not (inputs(169));
    layer0_outputs(6298) <= (inputs(52)) and (inputs(97));
    layer0_outputs(6299) <= (inputs(110)) and not (inputs(222));
    layer0_outputs(6300) <= not(inputs(50)) or (inputs(234));
    layer0_outputs(6301) <= (inputs(247)) or (inputs(241));
    layer0_outputs(6302) <= not(inputs(206)) or (inputs(122));
    layer0_outputs(6303) <= inputs(198);
    layer0_outputs(6304) <= (inputs(147)) or (inputs(219));
    layer0_outputs(6305) <= inputs(148);
    layer0_outputs(6306) <= (inputs(198)) and not (inputs(154));
    layer0_outputs(6307) <= inputs(227);
    layer0_outputs(6308) <= '1';
    layer0_outputs(6309) <= (inputs(203)) and not (inputs(2));
    layer0_outputs(6310) <= inputs(244);
    layer0_outputs(6311) <= not((inputs(109)) or (inputs(65)));
    layer0_outputs(6312) <= (inputs(63)) or (inputs(64));
    layer0_outputs(6313) <= (inputs(93)) or (inputs(158));
    layer0_outputs(6314) <= not(inputs(51)) or (inputs(36));
    layer0_outputs(6315) <= not(inputs(89)) or (inputs(81));
    layer0_outputs(6316) <= (inputs(128)) xor (inputs(130));
    layer0_outputs(6317) <= (inputs(112)) or (inputs(29));
    layer0_outputs(6318) <= not(inputs(61));
    layer0_outputs(6319) <= (inputs(164)) and not (inputs(88));
    layer0_outputs(6320) <= not((inputs(253)) or (inputs(205)));
    layer0_outputs(6321) <= (inputs(243)) xor (inputs(97));
    layer0_outputs(6322) <= '0';
    layer0_outputs(6323) <= not(inputs(181));
    layer0_outputs(6324) <= not(inputs(72));
    layer0_outputs(6325) <= (inputs(126)) and not (inputs(169));
    layer0_outputs(6326) <= '1';
    layer0_outputs(6327) <= inputs(146);
    layer0_outputs(6328) <= not(inputs(201));
    layer0_outputs(6329) <= inputs(230);
    layer0_outputs(6330) <= not(inputs(182)) or (inputs(70));
    layer0_outputs(6331) <= (inputs(105)) xor (inputs(136));
    layer0_outputs(6332) <= inputs(22);
    layer0_outputs(6333) <= not(inputs(44)) or (inputs(23));
    layer0_outputs(6334) <= inputs(222);
    layer0_outputs(6335) <= not((inputs(100)) or (inputs(35)));
    layer0_outputs(6336) <= (inputs(249)) xor (inputs(56));
    layer0_outputs(6337) <= inputs(190);
    layer0_outputs(6338) <= '0';
    layer0_outputs(6339) <= inputs(86);
    layer0_outputs(6340) <= (inputs(120)) and not (inputs(125));
    layer0_outputs(6341) <= '0';
    layer0_outputs(6342) <= not(inputs(161)) or (inputs(217));
    layer0_outputs(6343) <= not((inputs(79)) or (inputs(22)));
    layer0_outputs(6344) <= '1';
    layer0_outputs(6345) <= (inputs(184)) xor (inputs(16));
    layer0_outputs(6346) <= (inputs(165)) or (inputs(188));
    layer0_outputs(6347) <= not((inputs(60)) xor (inputs(13)));
    layer0_outputs(6348) <= not(inputs(227)) or (inputs(3));
    layer0_outputs(6349) <= (inputs(24)) and not (inputs(103));
    layer0_outputs(6350) <= not(inputs(16)) or (inputs(46));
    layer0_outputs(6351) <= '1';
    layer0_outputs(6352) <= inputs(25);
    layer0_outputs(6353) <= not((inputs(230)) and (inputs(131)));
    layer0_outputs(6354) <= not(inputs(132)) or (inputs(33));
    layer0_outputs(6355) <= not(inputs(219)) or (inputs(182));
    layer0_outputs(6356) <= not(inputs(195));
    layer0_outputs(6357) <= (inputs(37)) and not (inputs(177));
    layer0_outputs(6358) <= inputs(193);
    layer0_outputs(6359) <= not(inputs(84));
    layer0_outputs(6360) <= not(inputs(67)) or (inputs(1));
    layer0_outputs(6361) <= not(inputs(22)) or (inputs(144));
    layer0_outputs(6362) <= not(inputs(184)) or (inputs(195));
    layer0_outputs(6363) <= not(inputs(41)) or (inputs(148));
    layer0_outputs(6364) <= inputs(130);
    layer0_outputs(6365) <= (inputs(222)) and not (inputs(128));
    layer0_outputs(6366) <= not(inputs(245)) or (inputs(139));
    layer0_outputs(6367) <= (inputs(2)) and not (inputs(192));
    layer0_outputs(6368) <= not(inputs(236));
    layer0_outputs(6369) <= (inputs(187)) xor (inputs(232));
    layer0_outputs(6370) <= not((inputs(172)) xor (inputs(137)));
    layer0_outputs(6371) <= not(inputs(226)) or (inputs(13));
    layer0_outputs(6372) <= not((inputs(228)) or (inputs(160)));
    layer0_outputs(6373) <= inputs(90);
    layer0_outputs(6374) <= not((inputs(184)) and (inputs(35)));
    layer0_outputs(6375) <= not(inputs(46));
    layer0_outputs(6376) <= inputs(63);
    layer0_outputs(6377) <= not((inputs(173)) or (inputs(97)));
    layer0_outputs(6378) <= inputs(232);
    layer0_outputs(6379) <= not(inputs(178)) or (inputs(31));
    layer0_outputs(6380) <= not((inputs(4)) or (inputs(92)));
    layer0_outputs(6381) <= not((inputs(195)) xor (inputs(78)));
    layer0_outputs(6382) <= not(inputs(234)) or (inputs(2));
    layer0_outputs(6383) <= (inputs(2)) and not (inputs(203));
    layer0_outputs(6384) <= inputs(197);
    layer0_outputs(6385) <= (inputs(50)) or (inputs(212));
    layer0_outputs(6386) <= (inputs(39)) or (inputs(4));
    layer0_outputs(6387) <= not(inputs(119)) or (inputs(255));
    layer0_outputs(6388) <= not(inputs(176)) or (inputs(169));
    layer0_outputs(6389) <= not((inputs(8)) xor (inputs(222)));
    layer0_outputs(6390) <= (inputs(237)) or (inputs(234));
    layer0_outputs(6391) <= (inputs(117)) and not (inputs(126));
    layer0_outputs(6392) <= inputs(81);
    layer0_outputs(6393) <= not((inputs(144)) or (inputs(7)));
    layer0_outputs(6394) <= '0';
    layer0_outputs(6395) <= not((inputs(22)) or (inputs(5)));
    layer0_outputs(6396) <= (inputs(242)) and not (inputs(244));
    layer0_outputs(6397) <= not(inputs(72)) or (inputs(16));
    layer0_outputs(6398) <= (inputs(229)) and (inputs(228));
    layer0_outputs(6399) <= not((inputs(253)) or (inputs(1)));
    layer0_outputs(6400) <= (inputs(103)) or (inputs(48));
    layer0_outputs(6401) <= not(inputs(201));
    layer0_outputs(6402) <= (inputs(224)) and (inputs(217));
    layer0_outputs(6403) <= not(inputs(245)) or (inputs(215));
    layer0_outputs(6404) <= (inputs(163)) or (inputs(151));
    layer0_outputs(6405) <= inputs(137);
    layer0_outputs(6406) <= not(inputs(22));
    layer0_outputs(6407) <= (inputs(49)) and not (inputs(67));
    layer0_outputs(6408) <= not(inputs(29));
    layer0_outputs(6409) <= (inputs(47)) and not (inputs(110));
    layer0_outputs(6410) <= (inputs(174)) and (inputs(214));
    layer0_outputs(6411) <= (inputs(104)) or (inputs(194));
    layer0_outputs(6412) <= not((inputs(131)) or (inputs(114)));
    layer0_outputs(6413) <= not(inputs(112));
    layer0_outputs(6414) <= not(inputs(101));
    layer0_outputs(6415) <= (inputs(54)) and not (inputs(168));
    layer0_outputs(6416) <= not(inputs(104));
    layer0_outputs(6417) <= not((inputs(146)) or (inputs(66)));
    layer0_outputs(6418) <= (inputs(164)) and (inputs(228));
    layer0_outputs(6419) <= not((inputs(136)) or (inputs(166)));
    layer0_outputs(6420) <= not((inputs(8)) or (inputs(250)));
    layer0_outputs(6421) <= not((inputs(8)) or (inputs(84)));
    layer0_outputs(6422) <= not((inputs(98)) or (inputs(170)));
    layer0_outputs(6423) <= not(inputs(80));
    layer0_outputs(6424) <= inputs(128);
    layer0_outputs(6425) <= not(inputs(79)) or (inputs(33));
    layer0_outputs(6426) <= (inputs(232)) xor (inputs(11));
    layer0_outputs(6427) <= not(inputs(125));
    layer0_outputs(6428) <= not((inputs(100)) or (inputs(52)));
    layer0_outputs(6429) <= not(inputs(2));
    layer0_outputs(6430) <= not(inputs(120));
    layer0_outputs(6431) <= not(inputs(43)) or (inputs(209));
    layer0_outputs(6432) <= '1';
    layer0_outputs(6433) <= (inputs(81)) and not (inputs(73));
    layer0_outputs(6434) <= not((inputs(3)) and (inputs(254)));
    layer0_outputs(6435) <= not(inputs(150)) or (inputs(142));
    layer0_outputs(6436) <= not(inputs(152));
    layer0_outputs(6437) <= not((inputs(179)) or (inputs(162)));
    layer0_outputs(6438) <= inputs(195);
    layer0_outputs(6439) <= not((inputs(208)) xor (inputs(238)));
    layer0_outputs(6440) <= not(inputs(43));
    layer0_outputs(6441) <= '0';
    layer0_outputs(6442) <= (inputs(169)) and not (inputs(102));
    layer0_outputs(6443) <= inputs(191);
    layer0_outputs(6444) <= not(inputs(223));
    layer0_outputs(6445) <= (inputs(52)) and not (inputs(125));
    layer0_outputs(6446) <= not((inputs(66)) or (inputs(117)));
    layer0_outputs(6447) <= not((inputs(245)) or (inputs(250)));
    layer0_outputs(6448) <= (inputs(91)) and not (inputs(194));
    layer0_outputs(6449) <= inputs(244);
    layer0_outputs(6450) <= not((inputs(52)) or (inputs(29)));
    layer0_outputs(6451) <= not(inputs(211));
    layer0_outputs(6452) <= (inputs(171)) xor (inputs(69));
    layer0_outputs(6453) <= not(inputs(122)) or (inputs(252));
    layer0_outputs(6454) <= inputs(17);
    layer0_outputs(6455) <= not(inputs(228)) or (inputs(89));
    layer0_outputs(6456) <= (inputs(231)) or (inputs(214));
    layer0_outputs(6457) <= inputs(137);
    layer0_outputs(6458) <= (inputs(145)) or (inputs(72));
    layer0_outputs(6459) <= not(inputs(236)) or (inputs(164));
    layer0_outputs(6460) <= not(inputs(110));
    layer0_outputs(6461) <= '0';
    layer0_outputs(6462) <= (inputs(163)) and (inputs(172));
    layer0_outputs(6463) <= (inputs(2)) or (inputs(105));
    layer0_outputs(6464) <= not((inputs(63)) or (inputs(106)));
    layer0_outputs(6465) <= inputs(181);
    layer0_outputs(6466) <= not((inputs(38)) or (inputs(83)));
    layer0_outputs(6467) <= inputs(229);
    layer0_outputs(6468) <= (inputs(99)) or (inputs(151));
    layer0_outputs(6469) <= not(inputs(75)) or (inputs(40));
    layer0_outputs(6470) <= not(inputs(73));
    layer0_outputs(6471) <= (inputs(237)) and not (inputs(105));
    layer0_outputs(6472) <= (inputs(139)) or (inputs(74));
    layer0_outputs(6473) <= (inputs(121)) and not (inputs(226));
    layer0_outputs(6474) <= inputs(136);
    layer0_outputs(6475) <= not((inputs(64)) or (inputs(166)));
    layer0_outputs(6476) <= not((inputs(87)) xor (inputs(89)));
    layer0_outputs(6477) <= inputs(71);
    layer0_outputs(6478) <= not(inputs(96));
    layer0_outputs(6479) <= inputs(75);
    layer0_outputs(6480) <= not(inputs(122)) or (inputs(182));
    layer0_outputs(6481) <= not(inputs(215));
    layer0_outputs(6482) <= (inputs(122)) or (inputs(148));
    layer0_outputs(6483) <= (inputs(91)) and (inputs(110));
    layer0_outputs(6484) <= inputs(248);
    layer0_outputs(6485) <= (inputs(22)) and not (inputs(144));
    layer0_outputs(6486) <= (inputs(83)) and not (inputs(234));
    layer0_outputs(6487) <= not((inputs(26)) or (inputs(110)));
    layer0_outputs(6488) <= not((inputs(14)) or (inputs(28)));
    layer0_outputs(6489) <= not(inputs(1)) or (inputs(81));
    layer0_outputs(6490) <= (inputs(162)) and not (inputs(248));
    layer0_outputs(6491) <= inputs(227);
    layer0_outputs(6492) <= not(inputs(111)) or (inputs(64));
    layer0_outputs(6493) <= not(inputs(248)) or (inputs(5));
    layer0_outputs(6494) <= not((inputs(221)) xor (inputs(74)));
    layer0_outputs(6495) <= not(inputs(82));
    layer0_outputs(6496) <= not(inputs(132));
    layer0_outputs(6497) <= not(inputs(102));
    layer0_outputs(6498) <= (inputs(25)) and not (inputs(197));
    layer0_outputs(6499) <= not(inputs(1));
    layer0_outputs(6500) <= inputs(13);
    layer0_outputs(6501) <= not(inputs(130));
    layer0_outputs(6502) <= not(inputs(144));
    layer0_outputs(6503) <= not(inputs(222)) or (inputs(206));
    layer0_outputs(6504) <= not(inputs(149));
    layer0_outputs(6505) <= not((inputs(141)) or (inputs(127)));
    layer0_outputs(6506) <= (inputs(164)) xor (inputs(114));
    layer0_outputs(6507) <= (inputs(163)) xor (inputs(53));
    layer0_outputs(6508) <= '0';
    layer0_outputs(6509) <= not(inputs(70));
    layer0_outputs(6510) <= '1';
    layer0_outputs(6511) <= (inputs(134)) and not (inputs(171));
    layer0_outputs(6512) <= not((inputs(203)) and (inputs(71)));
    layer0_outputs(6513) <= not((inputs(47)) or (inputs(62)));
    layer0_outputs(6514) <= not(inputs(89)) or (inputs(63));
    layer0_outputs(6515) <= not(inputs(94));
    layer0_outputs(6516) <= not(inputs(26));
    layer0_outputs(6517) <= '1';
    layer0_outputs(6518) <= '1';
    layer0_outputs(6519) <= (inputs(191)) and not (inputs(126));
    layer0_outputs(6520) <= not(inputs(169));
    layer0_outputs(6521) <= not(inputs(232));
    layer0_outputs(6522) <= not((inputs(115)) or (inputs(80)));
    layer0_outputs(6523) <= inputs(106);
    layer0_outputs(6524) <= not(inputs(211)) or (inputs(31));
    layer0_outputs(6525) <= not((inputs(208)) or (inputs(93)));
    layer0_outputs(6526) <= not(inputs(26)) or (inputs(192));
    layer0_outputs(6527) <= not(inputs(101)) or (inputs(244));
    layer0_outputs(6528) <= (inputs(233)) xor (inputs(245));
    layer0_outputs(6529) <= not(inputs(231));
    layer0_outputs(6530) <= not(inputs(43)) or (inputs(30));
    layer0_outputs(6531) <= not(inputs(71)) or (inputs(11));
    layer0_outputs(6532) <= '0';
    layer0_outputs(6533) <= not((inputs(106)) xor (inputs(221)));
    layer0_outputs(6534) <= (inputs(85)) and not (inputs(252));
    layer0_outputs(6535) <= not(inputs(151)) or (inputs(56));
    layer0_outputs(6536) <= (inputs(132)) and not (inputs(19));
    layer0_outputs(6537) <= inputs(153);
    layer0_outputs(6538) <= not((inputs(168)) or (inputs(142)));
    layer0_outputs(6539) <= (inputs(53)) xor (inputs(141));
    layer0_outputs(6540) <= inputs(237);
    layer0_outputs(6541) <= not((inputs(46)) or (inputs(18)));
    layer0_outputs(6542) <= not(inputs(25));
    layer0_outputs(6543) <= not(inputs(19));
    layer0_outputs(6544) <= (inputs(247)) xor (inputs(215));
    layer0_outputs(6545) <= not(inputs(106));
    layer0_outputs(6546) <= not(inputs(112));
    layer0_outputs(6547) <= inputs(23);
    layer0_outputs(6548) <= (inputs(161)) or (inputs(39));
    layer0_outputs(6549) <= (inputs(82)) and (inputs(137));
    layer0_outputs(6550) <= '0';
    layer0_outputs(6551) <= not((inputs(218)) or (inputs(222)));
    layer0_outputs(6552) <= not(inputs(90));
    layer0_outputs(6553) <= (inputs(227)) and (inputs(220));
    layer0_outputs(6554) <= not(inputs(94)) or (inputs(198));
    layer0_outputs(6555) <= (inputs(230)) and (inputs(90));
    layer0_outputs(6556) <= inputs(63);
    layer0_outputs(6557) <= not(inputs(155)) or (inputs(108));
    layer0_outputs(6558) <= inputs(190);
    layer0_outputs(6559) <= inputs(232);
    layer0_outputs(6560) <= (inputs(236)) xor (inputs(230));
    layer0_outputs(6561) <= (inputs(85)) and not (inputs(215));
    layer0_outputs(6562) <= not(inputs(132));
    layer0_outputs(6563) <= not((inputs(24)) and (inputs(26)));
    layer0_outputs(6564) <= inputs(103);
    layer0_outputs(6565) <= not(inputs(196));
    layer0_outputs(6566) <= (inputs(241)) or (inputs(137));
    layer0_outputs(6567) <= inputs(130);
    layer0_outputs(6568) <= (inputs(236)) and not (inputs(68));
    layer0_outputs(6569) <= not((inputs(54)) xor (inputs(29)));
    layer0_outputs(6570) <= not(inputs(14));
    layer0_outputs(6571) <= not(inputs(88)) or (inputs(211));
    layer0_outputs(6572) <= (inputs(156)) and not (inputs(3));
    layer0_outputs(6573) <= (inputs(145)) and not (inputs(103));
    layer0_outputs(6574) <= (inputs(155)) xor (inputs(137));
    layer0_outputs(6575) <= inputs(232);
    layer0_outputs(6576) <= (inputs(242)) xor (inputs(45));
    layer0_outputs(6577) <= (inputs(221)) or (inputs(201));
    layer0_outputs(6578) <= (inputs(41)) or (inputs(51));
    layer0_outputs(6579) <= '0';
    layer0_outputs(6580) <= not(inputs(36));
    layer0_outputs(6581) <= not(inputs(68)) or (inputs(239));
    layer0_outputs(6582) <= '0';
    layer0_outputs(6583) <= inputs(167);
    layer0_outputs(6584) <= not(inputs(219));
    layer0_outputs(6585) <= inputs(102);
    layer0_outputs(6586) <= (inputs(150)) and not (inputs(174));
    layer0_outputs(6587) <= (inputs(76)) and not (inputs(8));
    layer0_outputs(6588) <= inputs(22);
    layer0_outputs(6589) <= inputs(119);
    layer0_outputs(6590) <= not(inputs(57)) or (inputs(235));
    layer0_outputs(6591) <= inputs(169);
    layer0_outputs(6592) <= not((inputs(172)) or (inputs(67)));
    layer0_outputs(6593) <= (inputs(188)) or (inputs(39));
    layer0_outputs(6594) <= (inputs(232)) and not (inputs(52));
    layer0_outputs(6595) <= not(inputs(232)) or (inputs(128));
    layer0_outputs(6596) <= inputs(121);
    layer0_outputs(6597) <= (inputs(201)) and not (inputs(79));
    layer0_outputs(6598) <= inputs(66);
    layer0_outputs(6599) <= inputs(246);
    layer0_outputs(6600) <= not(inputs(143));
    layer0_outputs(6601) <= not(inputs(30));
    layer0_outputs(6602) <= not(inputs(196));
    layer0_outputs(6603) <= (inputs(93)) or (inputs(63));
    layer0_outputs(6604) <= not((inputs(141)) xor (inputs(106)));
    layer0_outputs(6605) <= (inputs(218)) and not (inputs(41));
    layer0_outputs(6606) <= '1';
    layer0_outputs(6607) <= inputs(57);
    layer0_outputs(6608) <= (inputs(243)) or (inputs(119));
    layer0_outputs(6609) <= (inputs(32)) or (inputs(20));
    layer0_outputs(6610) <= not(inputs(40));
    layer0_outputs(6611) <= not(inputs(212)) or (inputs(51));
    layer0_outputs(6612) <= (inputs(193)) or (inputs(63));
    layer0_outputs(6613) <= inputs(205);
    layer0_outputs(6614) <= '0';
    layer0_outputs(6615) <= (inputs(108)) and not (inputs(71));
    layer0_outputs(6616) <= not((inputs(97)) or (inputs(132)));
    layer0_outputs(6617) <= not(inputs(73));
    layer0_outputs(6618) <= not(inputs(104));
    layer0_outputs(6619) <= not((inputs(67)) or (inputs(154)));
    layer0_outputs(6620) <= not((inputs(29)) or (inputs(159)));
    layer0_outputs(6621) <= (inputs(250)) or (inputs(62));
    layer0_outputs(6622) <= (inputs(44)) or (inputs(127));
    layer0_outputs(6623) <= (inputs(157)) or (inputs(159));
    layer0_outputs(6624) <= not(inputs(88));
    layer0_outputs(6625) <= not(inputs(207));
    layer0_outputs(6626) <= not(inputs(26));
    layer0_outputs(6627) <= (inputs(81)) or (inputs(109));
    layer0_outputs(6628) <= inputs(46);
    layer0_outputs(6629) <= not((inputs(170)) xor (inputs(77)));
    layer0_outputs(6630) <= inputs(212);
    layer0_outputs(6631) <= (inputs(143)) or (inputs(113));
    layer0_outputs(6632) <= (inputs(223)) xor (inputs(127));
    layer0_outputs(6633) <= (inputs(74)) or (inputs(119));
    layer0_outputs(6634) <= not(inputs(131));
    layer0_outputs(6635) <= (inputs(84)) or (inputs(84));
    layer0_outputs(6636) <= (inputs(185)) xor (inputs(123));
    layer0_outputs(6637) <= not(inputs(27));
    layer0_outputs(6638) <= not(inputs(84));
    layer0_outputs(6639) <= not(inputs(205));
    layer0_outputs(6640) <= inputs(158);
    layer0_outputs(6641) <= not((inputs(157)) or (inputs(161)));
    layer0_outputs(6642) <= (inputs(105)) and not (inputs(79));
    layer0_outputs(6643) <= inputs(84);
    layer0_outputs(6644) <= not((inputs(68)) or (inputs(127)));
    layer0_outputs(6645) <= (inputs(178)) and not (inputs(20));
    layer0_outputs(6646) <= '1';
    layer0_outputs(6647) <= (inputs(69)) xor (inputs(104));
    layer0_outputs(6648) <= (inputs(194)) and not (inputs(128));
    layer0_outputs(6649) <= (inputs(196)) and not (inputs(80));
    layer0_outputs(6650) <= (inputs(126)) and not (inputs(47));
    layer0_outputs(6651) <= not(inputs(180)) or (inputs(81));
    layer0_outputs(6652) <= (inputs(69)) xor (inputs(63));
    layer0_outputs(6653) <= (inputs(7)) and not (inputs(190));
    layer0_outputs(6654) <= (inputs(232)) and not (inputs(107));
    layer0_outputs(6655) <= not((inputs(187)) xor (inputs(115)));
    layer0_outputs(6656) <= not((inputs(227)) or (inputs(141)));
    layer0_outputs(6657) <= (inputs(48)) xor (inputs(244));
    layer0_outputs(6658) <= inputs(150);
    layer0_outputs(6659) <= (inputs(217)) and (inputs(20));
    layer0_outputs(6660) <= inputs(128);
    layer0_outputs(6661) <= not((inputs(242)) or (inputs(248)));
    layer0_outputs(6662) <= inputs(57);
    layer0_outputs(6663) <= not(inputs(103)) or (inputs(7));
    layer0_outputs(6664) <= (inputs(189)) or (inputs(76));
    layer0_outputs(6665) <= (inputs(54)) xor (inputs(41));
    layer0_outputs(6666) <= not(inputs(99));
    layer0_outputs(6667) <= not(inputs(87)) or (inputs(145));
    layer0_outputs(6668) <= (inputs(153)) and (inputs(148));
    layer0_outputs(6669) <= inputs(82);
    layer0_outputs(6670) <= not((inputs(159)) or (inputs(181)));
    layer0_outputs(6671) <= not((inputs(124)) or (inputs(201)));
    layer0_outputs(6672) <= not(inputs(30)) or (inputs(222));
    layer0_outputs(6673) <= inputs(185);
    layer0_outputs(6674) <= (inputs(167)) and not (inputs(47));
    layer0_outputs(6675) <= not(inputs(133));
    layer0_outputs(6676) <= not((inputs(94)) or (inputs(175)));
    layer0_outputs(6677) <= not(inputs(233)) or (inputs(1));
    layer0_outputs(6678) <= not(inputs(133));
    layer0_outputs(6679) <= not(inputs(222));
    layer0_outputs(6680) <= not(inputs(219)) or (inputs(66));
    layer0_outputs(6681) <= not(inputs(36)) or (inputs(112));
    layer0_outputs(6682) <= not(inputs(162));
    layer0_outputs(6683) <= (inputs(212)) or (inputs(246));
    layer0_outputs(6684) <= not((inputs(91)) xor (inputs(162)));
    layer0_outputs(6685) <= not((inputs(190)) xor (inputs(176)));
    layer0_outputs(6686) <= inputs(127);
    layer0_outputs(6687) <= (inputs(124)) or (inputs(31));
    layer0_outputs(6688) <= not(inputs(120));
    layer0_outputs(6689) <= '0';
    layer0_outputs(6690) <= (inputs(67)) and not (inputs(231));
    layer0_outputs(6691) <= (inputs(193)) and not (inputs(33));
    layer0_outputs(6692) <= not((inputs(0)) or (inputs(245)));
    layer0_outputs(6693) <= not((inputs(177)) xor (inputs(133)));
    layer0_outputs(6694) <= inputs(237);
    layer0_outputs(6695) <= (inputs(175)) or (inputs(157));
    layer0_outputs(6696) <= not(inputs(53)) or (inputs(143));
    layer0_outputs(6697) <= not((inputs(147)) xor (inputs(94)));
    layer0_outputs(6698) <= (inputs(79)) or (inputs(163));
    layer0_outputs(6699) <= not((inputs(3)) or (inputs(153)));
    layer0_outputs(6700) <= not(inputs(161));
    layer0_outputs(6701) <= not((inputs(80)) xor (inputs(184)));
    layer0_outputs(6702) <= (inputs(155)) or (inputs(165));
    layer0_outputs(6703) <= inputs(191);
    layer0_outputs(6704) <= inputs(104);
    layer0_outputs(6705) <= not((inputs(2)) or (inputs(77)));
    layer0_outputs(6706) <= inputs(148);
    layer0_outputs(6707) <= not(inputs(210)) or (inputs(1));
    layer0_outputs(6708) <= '0';
    layer0_outputs(6709) <= not((inputs(100)) or (inputs(63)));
    layer0_outputs(6710) <= (inputs(34)) and (inputs(124));
    layer0_outputs(6711) <= not((inputs(180)) or (inputs(192)));
    layer0_outputs(6712) <= (inputs(215)) and (inputs(228));
    layer0_outputs(6713) <= not((inputs(23)) and (inputs(67)));
    layer0_outputs(6714) <= (inputs(124)) or (inputs(62));
    layer0_outputs(6715) <= not((inputs(92)) or (inputs(58)));
    layer0_outputs(6716) <= (inputs(22)) or (inputs(191));
    layer0_outputs(6717) <= not(inputs(76));
    layer0_outputs(6718) <= not(inputs(142)) or (inputs(223));
    layer0_outputs(6719) <= (inputs(14)) xor (inputs(145));
    layer0_outputs(6720) <= (inputs(235)) or (inputs(195));
    layer0_outputs(6721) <= '0';
    layer0_outputs(6722) <= not(inputs(124));
    layer0_outputs(6723) <= not(inputs(179));
    layer0_outputs(6724) <= inputs(100);
    layer0_outputs(6725) <= (inputs(109)) xor (inputs(38));
    layer0_outputs(6726) <= not((inputs(58)) or (inputs(165)));
    layer0_outputs(6727) <= inputs(166);
    layer0_outputs(6728) <= not((inputs(65)) and (inputs(97)));
    layer0_outputs(6729) <= not((inputs(249)) or (inputs(18)));
    layer0_outputs(6730) <= not((inputs(219)) xor (inputs(188)));
    layer0_outputs(6731) <= (inputs(229)) xor (inputs(251));
    layer0_outputs(6732) <= not((inputs(164)) or (inputs(174)));
    layer0_outputs(6733) <= (inputs(86)) and (inputs(103));
    layer0_outputs(6734) <= not((inputs(199)) or (inputs(96)));
    layer0_outputs(6735) <= (inputs(55)) and not (inputs(252));
    layer0_outputs(6736) <= not(inputs(226));
    layer0_outputs(6737) <= (inputs(87)) and not (inputs(174));
    layer0_outputs(6738) <= (inputs(19)) xor (inputs(231));
    layer0_outputs(6739) <= not((inputs(59)) or (inputs(111)));
    layer0_outputs(6740) <= not(inputs(55));
    layer0_outputs(6741) <= (inputs(38)) or (inputs(70));
    layer0_outputs(6742) <= '0';
    layer0_outputs(6743) <= (inputs(132)) xor (inputs(189));
    layer0_outputs(6744) <= inputs(234);
    layer0_outputs(6745) <= (inputs(111)) or (inputs(132));
    layer0_outputs(6746) <= inputs(75);
    layer0_outputs(6747) <= (inputs(209)) and not (inputs(174));
    layer0_outputs(6748) <= not((inputs(151)) or (inputs(206)));
    layer0_outputs(6749) <= '0';
    layer0_outputs(6750) <= not((inputs(241)) and (inputs(237)));
    layer0_outputs(6751) <= not(inputs(232));
    layer0_outputs(6752) <= '1';
    layer0_outputs(6753) <= (inputs(116)) and not (inputs(251));
    layer0_outputs(6754) <= '1';
    layer0_outputs(6755) <= not(inputs(229)) or (inputs(49));
    layer0_outputs(6756) <= not(inputs(6));
    layer0_outputs(6757) <= not(inputs(149)) or (inputs(215));
    layer0_outputs(6758) <= not((inputs(42)) and (inputs(62)));
    layer0_outputs(6759) <= not(inputs(8)) or (inputs(118));
    layer0_outputs(6760) <= not(inputs(86)) or (inputs(159));
    layer0_outputs(6761) <= not((inputs(96)) or (inputs(85)));
    layer0_outputs(6762) <= inputs(106);
    layer0_outputs(6763) <= (inputs(162)) or (inputs(85));
    layer0_outputs(6764) <= (inputs(99)) and not (inputs(127));
    layer0_outputs(6765) <= (inputs(20)) or (inputs(18));
    layer0_outputs(6766) <= inputs(27);
    layer0_outputs(6767) <= (inputs(54)) or (inputs(146));
    layer0_outputs(6768) <= (inputs(168)) and not (inputs(78));
    layer0_outputs(6769) <= not(inputs(155)) or (inputs(82));
    layer0_outputs(6770) <= (inputs(223)) or (inputs(5));
    layer0_outputs(6771) <= inputs(36);
    layer0_outputs(6772) <= inputs(18);
    layer0_outputs(6773) <= not((inputs(79)) or (inputs(12)));
    layer0_outputs(6774) <= not((inputs(146)) xor (inputs(228)));
    layer0_outputs(6775) <= (inputs(150)) xor (inputs(149));
    layer0_outputs(6776) <= (inputs(104)) and not (inputs(145));
    layer0_outputs(6777) <= inputs(70);
    layer0_outputs(6778) <= not((inputs(73)) or (inputs(6)));
    layer0_outputs(6779) <= (inputs(31)) or (inputs(28));
    layer0_outputs(6780) <= not((inputs(128)) xor (inputs(100)));
    layer0_outputs(6781) <= (inputs(192)) and not (inputs(95));
    layer0_outputs(6782) <= not(inputs(58));
    layer0_outputs(6783) <= not(inputs(26)) or (inputs(145));
    layer0_outputs(6784) <= not(inputs(198));
    layer0_outputs(6785) <= not(inputs(57));
    layer0_outputs(6786) <= not(inputs(53)) or (inputs(190));
    layer0_outputs(6787) <= not(inputs(189));
    layer0_outputs(6788) <= not((inputs(180)) xor (inputs(6)));
    layer0_outputs(6789) <= '0';
    layer0_outputs(6790) <= inputs(102);
    layer0_outputs(6791) <= (inputs(218)) or (inputs(198));
    layer0_outputs(6792) <= (inputs(37)) and not (inputs(129));
    layer0_outputs(6793) <= (inputs(92)) or (inputs(111));
    layer0_outputs(6794) <= not((inputs(47)) or (inputs(228)));
    layer0_outputs(6795) <= inputs(187);
    layer0_outputs(6796) <= inputs(115);
    layer0_outputs(6797) <= (inputs(244)) xor (inputs(115));
    layer0_outputs(6798) <= not(inputs(124));
    layer0_outputs(6799) <= '0';
    layer0_outputs(6800) <= inputs(87);
    layer0_outputs(6801) <= (inputs(180)) and not (inputs(29));
    layer0_outputs(6802) <= '1';
    layer0_outputs(6803) <= '0';
    layer0_outputs(6804) <= (inputs(135)) or (inputs(118));
    layer0_outputs(6805) <= not((inputs(144)) xor (inputs(102)));
    layer0_outputs(6806) <= (inputs(6)) xor (inputs(110));
    layer0_outputs(6807) <= (inputs(203)) and not (inputs(97));
    layer0_outputs(6808) <= not(inputs(115)) or (inputs(58));
    layer0_outputs(6809) <= not(inputs(52)) or (inputs(181));
    layer0_outputs(6810) <= not((inputs(19)) and (inputs(232)));
    layer0_outputs(6811) <= not(inputs(42)) or (inputs(144));
    layer0_outputs(6812) <= not(inputs(226)) or (inputs(239));
    layer0_outputs(6813) <= not(inputs(133));
    layer0_outputs(6814) <= (inputs(50)) and not (inputs(142));
    layer0_outputs(6815) <= not(inputs(124));
    layer0_outputs(6816) <= not(inputs(80)) or (inputs(66));
    layer0_outputs(6817) <= not((inputs(70)) xor (inputs(117)));
    layer0_outputs(6818) <= not(inputs(91));
    layer0_outputs(6819) <= not((inputs(68)) xor (inputs(189)));
    layer0_outputs(6820) <= (inputs(231)) and not (inputs(9));
    layer0_outputs(6821) <= not((inputs(2)) or (inputs(22)));
    layer0_outputs(6822) <= '1';
    layer0_outputs(6823) <= not(inputs(246)) or (inputs(55));
    layer0_outputs(6824) <= inputs(27);
    layer0_outputs(6825) <= (inputs(28)) xor (inputs(94));
    layer0_outputs(6826) <= not(inputs(166)) or (inputs(116));
    layer0_outputs(6827) <= not(inputs(127));
    layer0_outputs(6828) <= not(inputs(83)) or (inputs(235));
    layer0_outputs(6829) <= not(inputs(117));
    layer0_outputs(6830) <= '0';
    layer0_outputs(6831) <= (inputs(24)) and not (inputs(225));
    layer0_outputs(6832) <= inputs(135);
    layer0_outputs(6833) <= '1';
    layer0_outputs(6834) <= not((inputs(242)) or (inputs(240)));
    layer0_outputs(6835) <= (inputs(8)) xor (inputs(170));
    layer0_outputs(6836) <= not((inputs(108)) or (inputs(113)));
    layer0_outputs(6837) <= not(inputs(194));
    layer0_outputs(6838) <= not((inputs(2)) or (inputs(239)));
    layer0_outputs(6839) <= not(inputs(218)) or (inputs(72));
    layer0_outputs(6840) <= not((inputs(15)) or (inputs(62)));
    layer0_outputs(6841) <= (inputs(205)) or (inputs(210));
    layer0_outputs(6842) <= not((inputs(9)) or (inputs(130)));
    layer0_outputs(6843) <= inputs(148);
    layer0_outputs(6844) <= (inputs(189)) or (inputs(225));
    layer0_outputs(6845) <= not((inputs(137)) xor (inputs(237)));
    layer0_outputs(6846) <= not(inputs(18));
    layer0_outputs(6847) <= not(inputs(164));
    layer0_outputs(6848) <= not((inputs(38)) xor (inputs(225)));
    layer0_outputs(6849) <= inputs(102);
    layer0_outputs(6850) <= not((inputs(14)) or (inputs(197)));
    layer0_outputs(6851) <= not(inputs(79)) or (inputs(222));
    layer0_outputs(6852) <= inputs(42);
    layer0_outputs(6853) <= inputs(207);
    layer0_outputs(6854) <= inputs(228);
    layer0_outputs(6855) <= (inputs(243)) and (inputs(93));
    layer0_outputs(6856) <= inputs(132);
    layer0_outputs(6857) <= (inputs(221)) xor (inputs(142));
    layer0_outputs(6858) <= (inputs(118)) or (inputs(198));
    layer0_outputs(6859) <= not(inputs(54));
    layer0_outputs(6860) <= (inputs(180)) xor (inputs(177));
    layer0_outputs(6861) <= not(inputs(218)) or (inputs(98));
    layer0_outputs(6862) <= not((inputs(63)) xor (inputs(132)));
    layer0_outputs(6863) <= inputs(202);
    layer0_outputs(6864) <= not(inputs(172)) or (inputs(98));
    layer0_outputs(6865) <= not(inputs(121)) or (inputs(39));
    layer0_outputs(6866) <= '1';
    layer0_outputs(6867) <= not(inputs(138));
    layer0_outputs(6868) <= (inputs(38)) and not (inputs(217));
    layer0_outputs(6869) <= (inputs(109)) or (inputs(144));
    layer0_outputs(6870) <= (inputs(72)) and not (inputs(253));
    layer0_outputs(6871) <= (inputs(68)) xor (inputs(67));
    layer0_outputs(6872) <= not(inputs(37)) or (inputs(211));
    layer0_outputs(6873) <= (inputs(34)) or (inputs(240));
    layer0_outputs(6874) <= not((inputs(3)) xor (inputs(153)));
    layer0_outputs(6875) <= not((inputs(53)) or (inputs(203)));
    layer0_outputs(6876) <= '0';
    layer0_outputs(6877) <= not((inputs(38)) or (inputs(206)));
    layer0_outputs(6878) <= '1';
    layer0_outputs(6879) <= '1';
    layer0_outputs(6880) <= inputs(81);
    layer0_outputs(6881) <= inputs(147);
    layer0_outputs(6882) <= not((inputs(164)) or (inputs(158)));
    layer0_outputs(6883) <= not(inputs(83));
    layer0_outputs(6884) <= (inputs(147)) and not (inputs(72));
    layer0_outputs(6885) <= (inputs(253)) or (inputs(117));
    layer0_outputs(6886) <= '1';
    layer0_outputs(6887) <= not(inputs(122));
    layer0_outputs(6888) <= not(inputs(72)) or (inputs(123));
    layer0_outputs(6889) <= not((inputs(89)) or (inputs(214)));
    layer0_outputs(6890) <= (inputs(120)) or (inputs(80));
    layer0_outputs(6891) <= not((inputs(117)) or (inputs(231)));
    layer0_outputs(6892) <= not(inputs(97));
    layer0_outputs(6893) <= not((inputs(31)) or (inputs(247)));
    layer0_outputs(6894) <= (inputs(181)) or (inputs(251));
    layer0_outputs(6895) <= inputs(160);
    layer0_outputs(6896) <= not((inputs(182)) or (inputs(99)));
    layer0_outputs(6897) <= (inputs(210)) and (inputs(117));
    layer0_outputs(6898) <= not((inputs(134)) xor (inputs(148)));
    layer0_outputs(6899) <= (inputs(158)) and (inputs(186));
    layer0_outputs(6900) <= not((inputs(53)) xor (inputs(206)));
    layer0_outputs(6901) <= not((inputs(105)) and (inputs(154)));
    layer0_outputs(6902) <= inputs(174);
    layer0_outputs(6903) <= not((inputs(39)) or (inputs(9)));
    layer0_outputs(6904) <= (inputs(203)) and not (inputs(20));
    layer0_outputs(6905) <= not((inputs(16)) or (inputs(22)));
    layer0_outputs(6906) <= (inputs(218)) and not (inputs(173));
    layer0_outputs(6907) <= not((inputs(6)) or (inputs(57)));
    layer0_outputs(6908) <= inputs(188);
    layer0_outputs(6909) <= inputs(161);
    layer0_outputs(6910) <= inputs(25);
    layer0_outputs(6911) <= not((inputs(211)) or (inputs(14)));
    layer0_outputs(6912) <= inputs(12);
    layer0_outputs(6913) <= (inputs(109)) and (inputs(153));
    layer0_outputs(6914) <= not((inputs(244)) or (inputs(3)));
    layer0_outputs(6915) <= not((inputs(79)) or (inputs(192)));
    layer0_outputs(6916) <= not(inputs(81));
    layer0_outputs(6917) <= not((inputs(222)) or (inputs(168)));
    layer0_outputs(6918) <= not(inputs(182));
    layer0_outputs(6919) <= not((inputs(210)) or (inputs(202)));
    layer0_outputs(6920) <= inputs(120);
    layer0_outputs(6921) <= inputs(70);
    layer0_outputs(6922) <= not((inputs(53)) or (inputs(16)));
    layer0_outputs(6923) <= inputs(72);
    layer0_outputs(6924) <= (inputs(27)) or (inputs(223));
    layer0_outputs(6925) <= not(inputs(184)) or (inputs(142));
    layer0_outputs(6926) <= not(inputs(115));
    layer0_outputs(6927) <= inputs(190);
    layer0_outputs(6928) <= not((inputs(119)) or (inputs(73)));
    layer0_outputs(6929) <= not(inputs(233));
    layer0_outputs(6930) <= not((inputs(134)) xor (inputs(227)));
    layer0_outputs(6931) <= (inputs(34)) or (inputs(193));
    layer0_outputs(6932) <= not((inputs(109)) or (inputs(255)));
    layer0_outputs(6933) <= (inputs(124)) and (inputs(182));
    layer0_outputs(6934) <= inputs(176);
    layer0_outputs(6935) <= not(inputs(107)) or (inputs(97));
    layer0_outputs(6936) <= (inputs(36)) or (inputs(186));
    layer0_outputs(6937) <= not((inputs(153)) or (inputs(110)));
    layer0_outputs(6938) <= not((inputs(131)) xor (inputs(103)));
    layer0_outputs(6939) <= (inputs(250)) and not (inputs(80));
    layer0_outputs(6940) <= (inputs(143)) or (inputs(95));
    layer0_outputs(6941) <= (inputs(207)) or (inputs(188));
    layer0_outputs(6942) <= not((inputs(250)) or (inputs(0)));
    layer0_outputs(6943) <= (inputs(56)) and not (inputs(103));
    layer0_outputs(6944) <= inputs(230);
    layer0_outputs(6945) <= not(inputs(218)) or (inputs(12));
    layer0_outputs(6946) <= not(inputs(34));
    layer0_outputs(6947) <= inputs(189);
    layer0_outputs(6948) <= not(inputs(63)) or (inputs(17));
    layer0_outputs(6949) <= (inputs(165)) or (inputs(48));
    layer0_outputs(6950) <= (inputs(119)) and not (inputs(19));
    layer0_outputs(6951) <= (inputs(118)) and not (inputs(253));
    layer0_outputs(6952) <= not(inputs(101)) or (inputs(241));
    layer0_outputs(6953) <= inputs(181);
    layer0_outputs(6954) <= (inputs(229)) or (inputs(207));
    layer0_outputs(6955) <= inputs(205);
    layer0_outputs(6956) <= '0';
    layer0_outputs(6957) <= not((inputs(210)) or (inputs(54)));
    layer0_outputs(6958) <= not(inputs(186));
    layer0_outputs(6959) <= not(inputs(195));
    layer0_outputs(6960) <= '0';
    layer0_outputs(6961) <= '0';
    layer0_outputs(6962) <= not((inputs(26)) or (inputs(187)));
    layer0_outputs(6963) <= not(inputs(35));
    layer0_outputs(6964) <= (inputs(72)) and not (inputs(138));
    layer0_outputs(6965) <= (inputs(115)) and not (inputs(162));
    layer0_outputs(6966) <= (inputs(60)) and not (inputs(28));
    layer0_outputs(6967) <= not(inputs(154)) or (inputs(41));
    layer0_outputs(6968) <= inputs(204);
    layer0_outputs(6969) <= not(inputs(111));
    layer0_outputs(6970) <= not(inputs(156)) or (inputs(64));
    layer0_outputs(6971) <= not(inputs(3)) or (inputs(238));
    layer0_outputs(6972) <= (inputs(187)) xor (inputs(105));
    layer0_outputs(6973) <= not((inputs(80)) xor (inputs(69)));
    layer0_outputs(6974) <= inputs(122);
    layer0_outputs(6975) <= not((inputs(56)) or (inputs(255)));
    layer0_outputs(6976) <= not(inputs(233)) or (inputs(225));
    layer0_outputs(6977) <= (inputs(240)) and (inputs(119));
    layer0_outputs(6978) <= not(inputs(213));
    layer0_outputs(6979) <= not((inputs(26)) and (inputs(32)));
    layer0_outputs(6980) <= not(inputs(16));
    layer0_outputs(6981) <= (inputs(117)) xor (inputs(4));
    layer0_outputs(6982) <= not((inputs(179)) or (inputs(119)));
    layer0_outputs(6983) <= not((inputs(204)) or (inputs(93)));
    layer0_outputs(6984) <= inputs(60);
    layer0_outputs(6985) <= not(inputs(101));
    layer0_outputs(6986) <= not(inputs(149));
    layer0_outputs(6987) <= not((inputs(114)) or (inputs(121)));
    layer0_outputs(6988) <= not((inputs(105)) or (inputs(159)));
    layer0_outputs(6989) <= (inputs(206)) or (inputs(202));
    layer0_outputs(6990) <= inputs(157);
    layer0_outputs(6991) <= not((inputs(33)) xor (inputs(209)));
    layer0_outputs(6992) <= (inputs(121)) and not (inputs(207));
    layer0_outputs(6993) <= not((inputs(23)) or (inputs(174)));
    layer0_outputs(6994) <= not((inputs(181)) or (inputs(34)));
    layer0_outputs(6995) <= not(inputs(85));
    layer0_outputs(6996) <= (inputs(158)) or (inputs(214));
    layer0_outputs(6997) <= (inputs(32)) and not (inputs(122));
    layer0_outputs(6998) <= not((inputs(195)) or (inputs(173)));
    layer0_outputs(6999) <= '0';
    layer0_outputs(7000) <= inputs(219);
    layer0_outputs(7001) <= (inputs(125)) and not (inputs(221));
    layer0_outputs(7002) <= inputs(136);
    layer0_outputs(7003) <= '1';
    layer0_outputs(7004) <= not(inputs(180)) or (inputs(247));
    layer0_outputs(7005) <= not((inputs(46)) and (inputs(188)));
    layer0_outputs(7006) <= not(inputs(76));
    layer0_outputs(7007) <= (inputs(240)) and not (inputs(90));
    layer0_outputs(7008) <= (inputs(58)) xor (inputs(89));
    layer0_outputs(7009) <= not(inputs(139)) or (inputs(93));
    layer0_outputs(7010) <= inputs(185);
    layer0_outputs(7011) <= (inputs(204)) or (inputs(3));
    layer0_outputs(7012) <= (inputs(38)) and not (inputs(67));
    layer0_outputs(7013) <= not(inputs(41));
    layer0_outputs(7014) <= not(inputs(189));
    layer0_outputs(7015) <= inputs(225);
    layer0_outputs(7016) <= not(inputs(138)) or (inputs(6));
    layer0_outputs(7017) <= inputs(233);
    layer0_outputs(7018) <= (inputs(129)) xor (inputs(101));
    layer0_outputs(7019) <= not((inputs(37)) and (inputs(167)));
    layer0_outputs(7020) <= not(inputs(10));
    layer0_outputs(7021) <= (inputs(157)) or (inputs(68));
    layer0_outputs(7022) <= not(inputs(125)) or (inputs(63));
    layer0_outputs(7023) <= not((inputs(204)) or (inputs(244)));
    layer0_outputs(7024) <= inputs(237);
    layer0_outputs(7025) <= not(inputs(101));
    layer0_outputs(7026) <= not((inputs(135)) or (inputs(15)));
    layer0_outputs(7027) <= (inputs(171)) or (inputs(201));
    layer0_outputs(7028) <= (inputs(124)) and (inputs(169));
    layer0_outputs(7029) <= not(inputs(73)) or (inputs(127));
    layer0_outputs(7030) <= not(inputs(61)) or (inputs(138));
    layer0_outputs(7031) <= not(inputs(134));
    layer0_outputs(7032) <= (inputs(64)) xor (inputs(212));
    layer0_outputs(7033) <= not(inputs(2));
    layer0_outputs(7034) <= inputs(118);
    layer0_outputs(7035) <= not(inputs(82)) or (inputs(17));
    layer0_outputs(7036) <= '1';
    layer0_outputs(7037) <= (inputs(49)) and not (inputs(143));
    layer0_outputs(7038) <= inputs(147);
    layer0_outputs(7039) <= not(inputs(119));
    layer0_outputs(7040) <= not(inputs(163));
    layer0_outputs(7041) <= not(inputs(238));
    layer0_outputs(7042) <= not(inputs(184)) or (inputs(227));
    layer0_outputs(7043) <= (inputs(115)) and not (inputs(176));
    layer0_outputs(7044) <= not((inputs(156)) or (inputs(223)));
    layer0_outputs(7045) <= not(inputs(123));
    layer0_outputs(7046) <= not(inputs(201));
    layer0_outputs(7047) <= not(inputs(25)) or (inputs(31));
    layer0_outputs(7048) <= inputs(197);
    layer0_outputs(7049) <= inputs(90);
    layer0_outputs(7050) <= (inputs(20)) and not (inputs(174));
    layer0_outputs(7051) <= inputs(211);
    layer0_outputs(7052) <= (inputs(61)) or (inputs(31));
    layer0_outputs(7053) <= (inputs(201)) and (inputs(36));
    layer0_outputs(7054) <= not((inputs(32)) or (inputs(38)));
    layer0_outputs(7055) <= inputs(25);
    layer0_outputs(7056) <= not(inputs(210)) or (inputs(97));
    layer0_outputs(7057) <= (inputs(227)) or (inputs(231));
    layer0_outputs(7058) <= (inputs(71)) and not (inputs(247));
    layer0_outputs(7059) <= not(inputs(116));
    layer0_outputs(7060) <= not(inputs(178)) or (inputs(181));
    layer0_outputs(7061) <= not(inputs(175)) or (inputs(178));
    layer0_outputs(7062) <= inputs(183);
    layer0_outputs(7063) <= not((inputs(254)) xor (inputs(160)));
    layer0_outputs(7064) <= not(inputs(114));
    layer0_outputs(7065) <= not(inputs(194));
    layer0_outputs(7066) <= (inputs(101)) or (inputs(255));
    layer0_outputs(7067) <= inputs(194);
    layer0_outputs(7068) <= not((inputs(43)) or (inputs(131)));
    layer0_outputs(7069) <= not(inputs(227));
    layer0_outputs(7070) <= not((inputs(53)) or (inputs(176)));
    layer0_outputs(7071) <= not(inputs(229)) or (inputs(119));
    layer0_outputs(7072) <= inputs(102);
    layer0_outputs(7073) <= inputs(135);
    layer0_outputs(7074) <= not(inputs(121));
    layer0_outputs(7075) <= (inputs(231)) and not (inputs(199));
    layer0_outputs(7076) <= not((inputs(83)) or (inputs(110)));
    layer0_outputs(7077) <= not((inputs(27)) xor (inputs(200)));
    layer0_outputs(7078) <= inputs(43);
    layer0_outputs(7079) <= '1';
    layer0_outputs(7080) <= not((inputs(122)) or (inputs(82)));
    layer0_outputs(7081) <= not((inputs(243)) or (inputs(62)));
    layer0_outputs(7082) <= '1';
    layer0_outputs(7083) <= not((inputs(224)) xor (inputs(3)));
    layer0_outputs(7084) <= inputs(46);
    layer0_outputs(7085) <= inputs(187);
    layer0_outputs(7086) <= inputs(138);
    layer0_outputs(7087) <= (inputs(168)) or (inputs(223));
    layer0_outputs(7088) <= inputs(195);
    layer0_outputs(7089) <= inputs(30);
    layer0_outputs(7090) <= (inputs(115)) xor (inputs(147));
    layer0_outputs(7091) <= not((inputs(55)) or (inputs(32)));
    layer0_outputs(7092) <= (inputs(0)) and not (inputs(156));
    layer0_outputs(7093) <= not((inputs(0)) or (inputs(125)));
    layer0_outputs(7094) <= not((inputs(207)) xor (inputs(156)));
    layer0_outputs(7095) <= not(inputs(178));
    layer0_outputs(7096) <= (inputs(149)) or (inputs(68));
    layer0_outputs(7097) <= inputs(26);
    layer0_outputs(7098) <= not(inputs(48)) or (inputs(251));
    layer0_outputs(7099) <= not((inputs(145)) xor (inputs(186)));
    layer0_outputs(7100) <= not((inputs(162)) xor (inputs(248)));
    layer0_outputs(7101) <= (inputs(156)) or (inputs(118));
    layer0_outputs(7102) <= not(inputs(56)) or (inputs(252));
    layer0_outputs(7103) <= not(inputs(44));
    layer0_outputs(7104) <= (inputs(46)) and not (inputs(145));
    layer0_outputs(7105) <= not(inputs(75));
    layer0_outputs(7106) <= (inputs(148)) and (inputs(137));
    layer0_outputs(7107) <= (inputs(34)) or (inputs(207));
    layer0_outputs(7108) <= (inputs(218)) xor (inputs(79));
    layer0_outputs(7109) <= (inputs(87)) and (inputs(108));
    layer0_outputs(7110) <= not(inputs(221)) or (inputs(50));
    layer0_outputs(7111) <= not((inputs(208)) xor (inputs(153)));
    layer0_outputs(7112) <= inputs(177);
    layer0_outputs(7113) <= (inputs(2)) or (inputs(227));
    layer0_outputs(7114) <= not(inputs(185));
    layer0_outputs(7115) <= inputs(161);
    layer0_outputs(7116) <= not((inputs(204)) or (inputs(98)));
    layer0_outputs(7117) <= inputs(194);
    layer0_outputs(7118) <= not(inputs(218));
    layer0_outputs(7119) <= (inputs(226)) or (inputs(43));
    layer0_outputs(7120) <= inputs(39);
    layer0_outputs(7121) <= (inputs(133)) and (inputs(37));
    layer0_outputs(7122) <= '1';
    layer0_outputs(7123) <= not(inputs(76));
    layer0_outputs(7124) <= (inputs(179)) and not (inputs(251));
    layer0_outputs(7125) <= inputs(166);
    layer0_outputs(7126) <= inputs(230);
    layer0_outputs(7127) <= not(inputs(56));
    layer0_outputs(7128) <= (inputs(118)) and not (inputs(27));
    layer0_outputs(7129) <= inputs(82);
    layer0_outputs(7130) <= (inputs(38)) xor (inputs(246));
    layer0_outputs(7131) <= not(inputs(36)) or (inputs(206));
    layer0_outputs(7132) <= not(inputs(136)) or (inputs(41));
    layer0_outputs(7133) <= not(inputs(146)) or (inputs(131));
    layer0_outputs(7134) <= inputs(136);
    layer0_outputs(7135) <= (inputs(250)) and not (inputs(142));
    layer0_outputs(7136) <= (inputs(184)) or (inputs(32));
    layer0_outputs(7137) <= not((inputs(152)) xor (inputs(78)));
    layer0_outputs(7138) <= not(inputs(127)) or (inputs(34));
    layer0_outputs(7139) <= (inputs(23)) or (inputs(216));
    layer0_outputs(7140) <= not(inputs(103)) or (inputs(176));
    layer0_outputs(7141) <= not(inputs(156)) or (inputs(239));
    layer0_outputs(7142) <= (inputs(41)) or (inputs(34));
    layer0_outputs(7143) <= not(inputs(52));
    layer0_outputs(7144) <= (inputs(208)) or (inputs(165));
    layer0_outputs(7145) <= (inputs(108)) or (inputs(110));
    layer0_outputs(7146) <= inputs(140);
    layer0_outputs(7147) <= not((inputs(99)) xor (inputs(87)));
    layer0_outputs(7148) <= not(inputs(75)) or (inputs(46));
    layer0_outputs(7149) <= (inputs(111)) xor (inputs(91));
    layer0_outputs(7150) <= not(inputs(230));
    layer0_outputs(7151) <= not((inputs(143)) and (inputs(217)));
    layer0_outputs(7152) <= not(inputs(137));
    layer0_outputs(7153) <= (inputs(200)) and (inputs(20));
    layer0_outputs(7154) <= not((inputs(139)) or (inputs(14)));
    layer0_outputs(7155) <= '1';
    layer0_outputs(7156) <= not((inputs(49)) xor (inputs(25)));
    layer0_outputs(7157) <= (inputs(235)) and (inputs(248));
    layer0_outputs(7158) <= inputs(174);
    layer0_outputs(7159) <= not(inputs(191));
    layer0_outputs(7160) <= not(inputs(47));
    layer0_outputs(7161) <= not(inputs(230));
    layer0_outputs(7162) <= not((inputs(127)) xor (inputs(90)));
    layer0_outputs(7163) <= (inputs(255)) and not (inputs(95));
    layer0_outputs(7164) <= not(inputs(200));
    layer0_outputs(7165) <= not((inputs(13)) and (inputs(251)));
    layer0_outputs(7166) <= (inputs(174)) or (inputs(73));
    layer0_outputs(7167) <= (inputs(165)) or (inputs(133));
    layer0_outputs(7168) <= not((inputs(29)) xor (inputs(145)));
    layer0_outputs(7169) <= not((inputs(217)) or (inputs(237)));
    layer0_outputs(7170) <= (inputs(189)) or (inputs(108));
    layer0_outputs(7171) <= inputs(167);
    layer0_outputs(7172) <= not((inputs(85)) or (inputs(44)));
    layer0_outputs(7173) <= (inputs(229)) xor (inputs(64));
    layer0_outputs(7174) <= (inputs(120)) or (inputs(252));
    layer0_outputs(7175) <= not((inputs(209)) xor (inputs(202)));
    layer0_outputs(7176) <= not(inputs(66)) or (inputs(159));
    layer0_outputs(7177) <= (inputs(136)) and not (inputs(176));
    layer0_outputs(7178) <= (inputs(195)) and not (inputs(122));
    layer0_outputs(7179) <= not(inputs(210));
    layer0_outputs(7180) <= not((inputs(115)) xor (inputs(101)));
    layer0_outputs(7181) <= not(inputs(75)) or (inputs(113));
    layer0_outputs(7182) <= (inputs(136)) or (inputs(184));
    layer0_outputs(7183) <= not(inputs(75));
    layer0_outputs(7184) <= '1';
    layer0_outputs(7185) <= not((inputs(63)) xor (inputs(23)));
    layer0_outputs(7186) <= '1';
    layer0_outputs(7187) <= inputs(35);
    layer0_outputs(7188) <= (inputs(181)) or (inputs(167));
    layer0_outputs(7189) <= not(inputs(166));
    layer0_outputs(7190) <= not(inputs(210));
    layer0_outputs(7191) <= not(inputs(198));
    layer0_outputs(7192) <= (inputs(87)) and not (inputs(130));
    layer0_outputs(7193) <= (inputs(158)) and not (inputs(14));
    layer0_outputs(7194) <= inputs(167);
    layer0_outputs(7195) <= not(inputs(85)) or (inputs(226));
    layer0_outputs(7196) <= not(inputs(146));
    layer0_outputs(7197) <= '1';
    layer0_outputs(7198) <= not(inputs(82));
    layer0_outputs(7199) <= (inputs(117)) and not (inputs(45));
    layer0_outputs(7200) <= not((inputs(58)) xor (inputs(176)));
    layer0_outputs(7201) <= (inputs(179)) and not (inputs(60));
    layer0_outputs(7202) <= (inputs(29)) xor (inputs(197));
    layer0_outputs(7203) <= not((inputs(8)) or (inputs(122)));
    layer0_outputs(7204) <= (inputs(41)) or (inputs(225));
    layer0_outputs(7205) <= not((inputs(136)) and (inputs(107)));
    layer0_outputs(7206) <= not(inputs(227));
    layer0_outputs(7207) <= inputs(46);
    layer0_outputs(7208) <= inputs(244);
    layer0_outputs(7209) <= inputs(22);
    layer0_outputs(7210) <= (inputs(202)) or (inputs(175));
    layer0_outputs(7211) <= not((inputs(137)) xor (inputs(199)));
    layer0_outputs(7212) <= not((inputs(189)) and (inputs(112)));
    layer0_outputs(7213) <= inputs(98);
    layer0_outputs(7214) <= (inputs(91)) xor (inputs(94));
    layer0_outputs(7215) <= inputs(70);
    layer0_outputs(7216) <= inputs(98);
    layer0_outputs(7217) <= inputs(77);
    layer0_outputs(7218) <= not(inputs(213)) or (inputs(48));
    layer0_outputs(7219) <= not(inputs(25)) or (inputs(208));
    layer0_outputs(7220) <= not(inputs(145));
    layer0_outputs(7221) <= not((inputs(239)) and (inputs(107)));
    layer0_outputs(7222) <= not(inputs(92));
    layer0_outputs(7223) <= not(inputs(176));
    layer0_outputs(7224) <= inputs(73);
    layer0_outputs(7225) <= '0';
    layer0_outputs(7226) <= not(inputs(207)) or (inputs(143));
    layer0_outputs(7227) <= not(inputs(243)) or (inputs(145));
    layer0_outputs(7228) <= (inputs(149)) or (inputs(167));
    layer0_outputs(7229) <= inputs(85);
    layer0_outputs(7230) <= (inputs(71)) or (inputs(41));
    layer0_outputs(7231) <= (inputs(22)) or (inputs(49));
    layer0_outputs(7232) <= '0';
    layer0_outputs(7233) <= (inputs(90)) or (inputs(208));
    layer0_outputs(7234) <= not((inputs(22)) or (inputs(192)));
    layer0_outputs(7235) <= not(inputs(231)) or (inputs(29));
    layer0_outputs(7236) <= (inputs(16)) and (inputs(36));
    layer0_outputs(7237) <= '0';
    layer0_outputs(7238) <= not(inputs(165));
    layer0_outputs(7239) <= (inputs(122)) and (inputs(91));
    layer0_outputs(7240) <= not((inputs(138)) or (inputs(219)));
    layer0_outputs(7241) <= not(inputs(189));
    layer0_outputs(7242) <= (inputs(140)) or (inputs(252));
    layer0_outputs(7243) <= '1';
    layer0_outputs(7244) <= not((inputs(21)) or (inputs(55)));
    layer0_outputs(7245) <= not(inputs(101)) or (inputs(93));
    layer0_outputs(7246) <= not((inputs(29)) or (inputs(209)));
    layer0_outputs(7247) <= (inputs(11)) and not (inputs(204));
    layer0_outputs(7248) <= (inputs(222)) or (inputs(86));
    layer0_outputs(7249) <= not((inputs(142)) or (inputs(214)));
    layer0_outputs(7250) <= (inputs(93)) and not (inputs(127));
    layer0_outputs(7251) <= not(inputs(156)) or (inputs(6));
    layer0_outputs(7252) <= not((inputs(186)) and (inputs(214)));
    layer0_outputs(7253) <= inputs(69);
    layer0_outputs(7254) <= (inputs(185)) or (inputs(51));
    layer0_outputs(7255) <= inputs(110);
    layer0_outputs(7256) <= not(inputs(252)) or (inputs(157));
    layer0_outputs(7257) <= (inputs(166)) and not (inputs(15));
    layer0_outputs(7258) <= (inputs(69)) and not (inputs(176));
    layer0_outputs(7259) <= (inputs(138)) or (inputs(239));
    layer0_outputs(7260) <= not(inputs(53)) or (inputs(61));
    layer0_outputs(7261) <= not(inputs(71));
    layer0_outputs(7262) <= not(inputs(147));
    layer0_outputs(7263) <= inputs(158);
    layer0_outputs(7264) <= '1';
    layer0_outputs(7265) <= '0';
    layer0_outputs(7266) <= (inputs(5)) and (inputs(217));
    layer0_outputs(7267) <= inputs(67);
    layer0_outputs(7268) <= not(inputs(90));
    layer0_outputs(7269) <= not(inputs(218)) or (inputs(70));
    layer0_outputs(7270) <= not(inputs(66)) or (inputs(180));
    layer0_outputs(7271) <= not((inputs(254)) xor (inputs(205)));
    layer0_outputs(7272) <= not((inputs(244)) or (inputs(57)));
    layer0_outputs(7273) <= not(inputs(105)) or (inputs(15));
    layer0_outputs(7274) <= (inputs(84)) or (inputs(84));
    layer0_outputs(7275) <= not((inputs(150)) xor (inputs(6)));
    layer0_outputs(7276) <= '1';
    layer0_outputs(7277) <= inputs(189);
    layer0_outputs(7278) <= not(inputs(188));
    layer0_outputs(7279) <= (inputs(137)) or (inputs(32));
    layer0_outputs(7280) <= (inputs(18)) and not (inputs(196));
    layer0_outputs(7281) <= (inputs(183)) or (inputs(186));
    layer0_outputs(7282) <= (inputs(77)) and not (inputs(205));
    layer0_outputs(7283) <= (inputs(164)) and not (inputs(30));
    layer0_outputs(7284) <= inputs(211);
    layer0_outputs(7285) <= inputs(176);
    layer0_outputs(7286) <= not(inputs(217));
    layer0_outputs(7287) <= (inputs(161)) or (inputs(1));
    layer0_outputs(7288) <= (inputs(19)) xor (inputs(147));
    layer0_outputs(7289) <= (inputs(3)) xor (inputs(174));
    layer0_outputs(7290) <= inputs(33);
    layer0_outputs(7291) <= not((inputs(138)) xor (inputs(168)));
    layer0_outputs(7292) <= not(inputs(84)) or (inputs(222));
    layer0_outputs(7293) <= (inputs(223)) or (inputs(28));
    layer0_outputs(7294) <= (inputs(124)) or (inputs(154));
    layer0_outputs(7295) <= not((inputs(211)) and (inputs(43)));
    layer0_outputs(7296) <= (inputs(192)) and not (inputs(129));
    layer0_outputs(7297) <= (inputs(142)) xor (inputs(68));
    layer0_outputs(7298) <= not((inputs(81)) and (inputs(239)));
    layer0_outputs(7299) <= (inputs(255)) or (inputs(89));
    layer0_outputs(7300) <= inputs(103);
    layer0_outputs(7301) <= (inputs(119)) and not (inputs(134));
    layer0_outputs(7302) <= not(inputs(178));
    layer0_outputs(7303) <= (inputs(226)) or (inputs(78));
    layer0_outputs(7304) <= inputs(97);
    layer0_outputs(7305) <= not(inputs(13));
    layer0_outputs(7306) <= (inputs(249)) xor (inputs(152));
    layer0_outputs(7307) <= inputs(188);
    layer0_outputs(7308) <= inputs(219);
    layer0_outputs(7309) <= not(inputs(194));
    layer0_outputs(7310) <= not((inputs(65)) or (inputs(104)));
    layer0_outputs(7311) <= (inputs(176)) or (inputs(79));
    layer0_outputs(7312) <= (inputs(38)) and not (inputs(130));
    layer0_outputs(7313) <= not(inputs(217));
    layer0_outputs(7314) <= not((inputs(90)) and (inputs(28)));
    layer0_outputs(7315) <= (inputs(215)) and not (inputs(46));
    layer0_outputs(7316) <= (inputs(0)) or (inputs(35));
    layer0_outputs(7317) <= (inputs(187)) xor (inputs(76));
    layer0_outputs(7318) <= '0';
    layer0_outputs(7319) <= not(inputs(195));
    layer0_outputs(7320) <= (inputs(143)) or (inputs(247));
    layer0_outputs(7321) <= not(inputs(163));
    layer0_outputs(7322) <= not(inputs(117));
    layer0_outputs(7323) <= not((inputs(129)) or (inputs(69)));
    layer0_outputs(7324) <= not(inputs(187));
    layer0_outputs(7325) <= not((inputs(151)) and (inputs(57)));
    layer0_outputs(7326) <= '0';
    layer0_outputs(7327) <= inputs(53);
    layer0_outputs(7328) <= '0';
    layer0_outputs(7329) <= not(inputs(227)) or (inputs(13));
    layer0_outputs(7330) <= not(inputs(179));
    layer0_outputs(7331) <= not((inputs(8)) or (inputs(111)));
    layer0_outputs(7332) <= '1';
    layer0_outputs(7333) <= (inputs(203)) xor (inputs(234));
    layer0_outputs(7334) <= not(inputs(209)) or (inputs(210));
    layer0_outputs(7335) <= inputs(122);
    layer0_outputs(7336) <= inputs(0);
    layer0_outputs(7337) <= inputs(26);
    layer0_outputs(7338) <= not((inputs(228)) xor (inputs(61)));
    layer0_outputs(7339) <= inputs(44);
    layer0_outputs(7340) <= not(inputs(98));
    layer0_outputs(7341) <= not(inputs(247)) or (inputs(54));
    layer0_outputs(7342) <= '1';
    layer0_outputs(7343) <= (inputs(184)) and not (inputs(67));
    layer0_outputs(7344) <= (inputs(55)) and not (inputs(164));
    layer0_outputs(7345) <= (inputs(123)) or (inputs(22));
    layer0_outputs(7346) <= '0';
    layer0_outputs(7347) <= not(inputs(142)) or (inputs(104));
    layer0_outputs(7348) <= not((inputs(129)) or (inputs(78)));
    layer0_outputs(7349) <= (inputs(35)) and not (inputs(244));
    layer0_outputs(7350) <= (inputs(20)) and not (inputs(201));
    layer0_outputs(7351) <= (inputs(52)) and not (inputs(235));
    layer0_outputs(7352) <= (inputs(166)) and not (inputs(86));
    layer0_outputs(7353) <= not(inputs(193)) or (inputs(252));
    layer0_outputs(7354) <= not((inputs(110)) and (inputs(159)));
    layer0_outputs(7355) <= (inputs(233)) and not (inputs(110));
    layer0_outputs(7356) <= not((inputs(37)) and (inputs(226)));
    layer0_outputs(7357) <= not(inputs(151));
    layer0_outputs(7358) <= (inputs(60)) and not (inputs(182));
    layer0_outputs(7359) <= inputs(58);
    layer0_outputs(7360) <= inputs(255);
    layer0_outputs(7361) <= (inputs(127)) xor (inputs(107));
    layer0_outputs(7362) <= not((inputs(156)) xor (inputs(234)));
    layer0_outputs(7363) <= (inputs(33)) or (inputs(29));
    layer0_outputs(7364) <= (inputs(247)) and not (inputs(105));
    layer0_outputs(7365) <= inputs(70);
    layer0_outputs(7366) <= (inputs(245)) or (inputs(86));
    layer0_outputs(7367) <= not(inputs(211));
    layer0_outputs(7368) <= not(inputs(214));
    layer0_outputs(7369) <= (inputs(186)) and not (inputs(41));
    layer0_outputs(7370) <= inputs(194);
    layer0_outputs(7371) <= (inputs(78)) or (inputs(155));
    layer0_outputs(7372) <= not(inputs(150));
    layer0_outputs(7373) <= not(inputs(93));
    layer0_outputs(7374) <= not(inputs(122)) or (inputs(212));
    layer0_outputs(7375) <= inputs(176);
    layer0_outputs(7376) <= not(inputs(164)) or (inputs(155));
    layer0_outputs(7377) <= not(inputs(82)) or (inputs(192));
    layer0_outputs(7378) <= not(inputs(18)) or (inputs(219));
    layer0_outputs(7379) <= not((inputs(245)) and (inputs(218)));
    layer0_outputs(7380) <= not(inputs(254));
    layer0_outputs(7381) <= (inputs(75)) and not (inputs(101));
    layer0_outputs(7382) <= not((inputs(134)) xor (inputs(151)));
    layer0_outputs(7383) <= '0';
    layer0_outputs(7384) <= not(inputs(155)) or (inputs(34));
    layer0_outputs(7385) <= inputs(253);
    layer0_outputs(7386) <= inputs(70);
    layer0_outputs(7387) <= not((inputs(126)) xor (inputs(107)));
    layer0_outputs(7388) <= (inputs(74)) or (inputs(185));
    layer0_outputs(7389) <= not(inputs(242)) or (inputs(170));
    layer0_outputs(7390) <= not((inputs(218)) xor (inputs(186)));
    layer0_outputs(7391) <= (inputs(176)) or (inputs(228));
    layer0_outputs(7392) <= not(inputs(193));
    layer0_outputs(7393) <= not((inputs(101)) xor (inputs(116)));
    layer0_outputs(7394) <= inputs(12);
    layer0_outputs(7395) <= not((inputs(242)) or (inputs(13)));
    layer0_outputs(7396) <= not((inputs(247)) and (inputs(171)));
    layer0_outputs(7397) <= not(inputs(63));
    layer0_outputs(7398) <= inputs(52);
    layer0_outputs(7399) <= (inputs(49)) and not (inputs(160));
    layer0_outputs(7400) <= (inputs(215)) and (inputs(235));
    layer0_outputs(7401) <= '0';
    layer0_outputs(7402) <= inputs(51);
    layer0_outputs(7403) <= not((inputs(133)) and (inputs(137)));
    layer0_outputs(7404) <= not(inputs(211));
    layer0_outputs(7405) <= not(inputs(96)) or (inputs(125));
    layer0_outputs(7406) <= not(inputs(40));
    layer0_outputs(7407) <= inputs(21);
    layer0_outputs(7408) <= not(inputs(166)) or (inputs(193));
    layer0_outputs(7409) <= inputs(130);
    layer0_outputs(7410) <= not(inputs(240));
    layer0_outputs(7411) <= (inputs(133)) and not (inputs(138));
    layer0_outputs(7412) <= (inputs(98)) or (inputs(84));
    layer0_outputs(7413) <= '0';
    layer0_outputs(7414) <= inputs(35);
    layer0_outputs(7415) <= not(inputs(137));
    layer0_outputs(7416) <= not((inputs(252)) or (inputs(51)));
    layer0_outputs(7417) <= not((inputs(65)) or (inputs(96)));
    layer0_outputs(7418) <= '0';
    layer0_outputs(7419) <= not(inputs(156)) or (inputs(51));
    layer0_outputs(7420) <= not((inputs(8)) or (inputs(239)));
    layer0_outputs(7421) <= not((inputs(25)) xor (inputs(87)));
    layer0_outputs(7422) <= not((inputs(52)) or (inputs(78)));
    layer0_outputs(7423) <= not((inputs(201)) and (inputs(155)));
    layer0_outputs(7424) <= (inputs(8)) and (inputs(42));
    layer0_outputs(7425) <= not(inputs(137)) or (inputs(250));
    layer0_outputs(7426) <= '1';
    layer0_outputs(7427) <= (inputs(102)) and not (inputs(67));
    layer0_outputs(7428) <= not((inputs(33)) or (inputs(155)));
    layer0_outputs(7429) <= not(inputs(104));
    layer0_outputs(7430) <= (inputs(72)) xor (inputs(65));
    layer0_outputs(7431) <= not(inputs(20));
    layer0_outputs(7432) <= (inputs(81)) xor (inputs(114));
    layer0_outputs(7433) <= (inputs(219)) and not (inputs(240));
    layer0_outputs(7434) <= not(inputs(246));
    layer0_outputs(7435) <= (inputs(75)) or (inputs(143));
    layer0_outputs(7436) <= (inputs(91)) or (inputs(126));
    layer0_outputs(7437) <= (inputs(195)) or (inputs(215));
    layer0_outputs(7438) <= not(inputs(141));
    layer0_outputs(7439) <= (inputs(133)) and not (inputs(226));
    layer0_outputs(7440) <= '0';
    layer0_outputs(7441) <= (inputs(209)) and not (inputs(124));
    layer0_outputs(7442) <= not(inputs(105));
    layer0_outputs(7443) <= '0';
    layer0_outputs(7444) <= inputs(129);
    layer0_outputs(7445) <= not((inputs(21)) or (inputs(183)));
    layer0_outputs(7446) <= (inputs(0)) and not (inputs(30));
    layer0_outputs(7447) <= not((inputs(255)) xor (inputs(98)));
    layer0_outputs(7448) <= inputs(237);
    layer0_outputs(7449) <= inputs(35);
    layer0_outputs(7450) <= not(inputs(40)) or (inputs(251));
    layer0_outputs(7451) <= (inputs(83)) and (inputs(250));
    layer0_outputs(7452) <= not(inputs(102));
    layer0_outputs(7453) <= not(inputs(255));
    layer0_outputs(7454) <= (inputs(196)) xor (inputs(225));
    layer0_outputs(7455) <= (inputs(163)) or (inputs(236));
    layer0_outputs(7456) <= not(inputs(232));
    layer0_outputs(7457) <= inputs(213);
    layer0_outputs(7458) <= (inputs(89)) and (inputs(38));
    layer0_outputs(7459) <= not(inputs(237));
    layer0_outputs(7460) <= not((inputs(27)) or (inputs(4)));
    layer0_outputs(7461) <= not((inputs(189)) xor (inputs(187)));
    layer0_outputs(7462) <= (inputs(35)) and not (inputs(57));
    layer0_outputs(7463) <= (inputs(231)) or (inputs(221));
    layer0_outputs(7464) <= (inputs(165)) or (inputs(182));
    layer0_outputs(7465) <= (inputs(234)) or (inputs(251));
    layer0_outputs(7466) <= (inputs(128)) or (inputs(174));
    layer0_outputs(7467) <= (inputs(24)) and (inputs(42));
    layer0_outputs(7468) <= inputs(228);
    layer0_outputs(7469) <= not((inputs(245)) or (inputs(145)));
    layer0_outputs(7470) <= not(inputs(85)) or (inputs(140));
    layer0_outputs(7471) <= inputs(24);
    layer0_outputs(7472) <= (inputs(88)) and not (inputs(142));
    layer0_outputs(7473) <= (inputs(95)) xor (inputs(11));
    layer0_outputs(7474) <= not((inputs(187)) or (inputs(5)));
    layer0_outputs(7475) <= (inputs(172)) and not (inputs(216));
    layer0_outputs(7476) <= inputs(67);
    layer0_outputs(7477) <= '1';
    layer0_outputs(7478) <= (inputs(95)) or (inputs(161));
    layer0_outputs(7479) <= not((inputs(216)) or (inputs(84)));
    layer0_outputs(7480) <= not(inputs(121)) or (inputs(195));
    layer0_outputs(7481) <= not((inputs(180)) xor (inputs(250)));
    layer0_outputs(7482) <= '1';
    layer0_outputs(7483) <= (inputs(231)) and not (inputs(142));
    layer0_outputs(7484) <= '0';
    layer0_outputs(7485) <= (inputs(117)) or (inputs(190));
    layer0_outputs(7486) <= not(inputs(125));
    layer0_outputs(7487) <= inputs(247);
    layer0_outputs(7488) <= (inputs(196)) or (inputs(95));
    layer0_outputs(7489) <= not(inputs(104)) or (inputs(33));
    layer0_outputs(7490) <= not((inputs(184)) xor (inputs(150)));
    layer0_outputs(7491) <= not((inputs(156)) or (inputs(189)));
    layer0_outputs(7492) <= (inputs(32)) or (inputs(41));
    layer0_outputs(7493) <= not(inputs(192)) or (inputs(229));
    layer0_outputs(7494) <= inputs(46);
    layer0_outputs(7495) <= (inputs(212)) and (inputs(191));
    layer0_outputs(7496) <= not(inputs(12));
    layer0_outputs(7497) <= (inputs(23)) or (inputs(244));
    layer0_outputs(7498) <= (inputs(162)) and not (inputs(143));
    layer0_outputs(7499) <= '0';
    layer0_outputs(7500) <= (inputs(129)) and not (inputs(118));
    layer0_outputs(7501) <= not(inputs(248)) or (inputs(238));
    layer0_outputs(7502) <= (inputs(151)) and not (inputs(76));
    layer0_outputs(7503) <= not(inputs(235));
    layer0_outputs(7504) <= not((inputs(191)) or (inputs(27)));
    layer0_outputs(7505) <= not(inputs(222));
    layer0_outputs(7506) <= (inputs(132)) and not (inputs(134));
    layer0_outputs(7507) <= (inputs(59)) and not (inputs(136));
    layer0_outputs(7508) <= not((inputs(238)) or (inputs(95)));
    layer0_outputs(7509) <= not(inputs(69));
    layer0_outputs(7510) <= '0';
    layer0_outputs(7511) <= not(inputs(242));
    layer0_outputs(7512) <= not((inputs(19)) xor (inputs(142)));
    layer0_outputs(7513) <= (inputs(53)) and (inputs(13));
    layer0_outputs(7514) <= (inputs(239)) and not (inputs(46));
    layer0_outputs(7515) <= (inputs(54)) and not (inputs(249));
    layer0_outputs(7516) <= inputs(43);
    layer0_outputs(7517) <= (inputs(204)) xor (inputs(127));
    layer0_outputs(7518) <= not(inputs(24)) or (inputs(161));
    layer0_outputs(7519) <= (inputs(170)) xor (inputs(107));
    layer0_outputs(7520) <= (inputs(219)) and (inputs(214));
    layer0_outputs(7521) <= not(inputs(137));
    layer0_outputs(7522) <= not(inputs(227)) or (inputs(78));
    layer0_outputs(7523) <= (inputs(238)) and not (inputs(157));
    layer0_outputs(7524) <= (inputs(156)) and (inputs(245));
    layer0_outputs(7525) <= not(inputs(46));
    layer0_outputs(7526) <= not((inputs(238)) xor (inputs(61)));
    layer0_outputs(7527) <= not(inputs(36)) or (inputs(36));
    layer0_outputs(7528) <= not(inputs(39)) or (inputs(162));
    layer0_outputs(7529) <= inputs(14);
    layer0_outputs(7530) <= not(inputs(56));
    layer0_outputs(7531) <= not(inputs(2));
    layer0_outputs(7532) <= not(inputs(72));
    layer0_outputs(7533) <= inputs(49);
    layer0_outputs(7534) <= not((inputs(114)) or (inputs(220)));
    layer0_outputs(7535) <= not((inputs(163)) xor (inputs(171)));
    layer0_outputs(7536) <= not(inputs(138)) or (inputs(248));
    layer0_outputs(7537) <= (inputs(118)) or (inputs(117));
    layer0_outputs(7538) <= '0';
    layer0_outputs(7539) <= (inputs(200)) and not (inputs(10));
    layer0_outputs(7540) <= (inputs(239)) or (inputs(74));
    layer0_outputs(7541) <= not(inputs(34));
    layer0_outputs(7542) <= not(inputs(12));
    layer0_outputs(7543) <= (inputs(206)) and not (inputs(222));
    layer0_outputs(7544) <= not(inputs(138));
    layer0_outputs(7545) <= not(inputs(246));
    layer0_outputs(7546) <= (inputs(172)) and not (inputs(35));
    layer0_outputs(7547) <= not((inputs(42)) or (inputs(127)));
    layer0_outputs(7548) <= inputs(56);
    layer0_outputs(7549) <= (inputs(26)) and not (inputs(40));
    layer0_outputs(7550) <= (inputs(88)) and not (inputs(129));
    layer0_outputs(7551) <= (inputs(28)) or (inputs(153));
    layer0_outputs(7552) <= (inputs(240)) and not (inputs(206));
    layer0_outputs(7553) <= not(inputs(169));
    layer0_outputs(7554) <= not(inputs(94));
    layer0_outputs(7555) <= not(inputs(70));
    layer0_outputs(7556) <= not(inputs(154)) or (inputs(48));
    layer0_outputs(7557) <= (inputs(176)) xor (inputs(215));
    layer0_outputs(7558) <= '1';
    layer0_outputs(7559) <= not(inputs(58)) or (inputs(33));
    layer0_outputs(7560) <= not(inputs(234)) or (inputs(4));
    layer0_outputs(7561) <= inputs(163);
    layer0_outputs(7562) <= inputs(147);
    layer0_outputs(7563) <= not(inputs(246));
    layer0_outputs(7564) <= inputs(105);
    layer0_outputs(7565) <= inputs(196);
    layer0_outputs(7566) <= inputs(254);
    layer0_outputs(7567) <= not((inputs(93)) or (inputs(123)));
    layer0_outputs(7568) <= inputs(142);
    layer0_outputs(7569) <= not(inputs(9)) or (inputs(226));
    layer0_outputs(7570) <= not(inputs(136)) or (inputs(194));
    layer0_outputs(7571) <= '0';
    layer0_outputs(7572) <= not(inputs(130));
    layer0_outputs(7573) <= (inputs(4)) and (inputs(186));
    layer0_outputs(7574) <= not(inputs(53)) or (inputs(175));
    layer0_outputs(7575) <= '0';
    layer0_outputs(7576) <= not(inputs(94));
    layer0_outputs(7577) <= (inputs(169)) or (inputs(143));
    layer0_outputs(7578) <= (inputs(78)) or (inputs(161));
    layer0_outputs(7579) <= (inputs(100)) and not (inputs(119));
    layer0_outputs(7580) <= (inputs(32)) or (inputs(29));
    layer0_outputs(7581) <= inputs(162);
    layer0_outputs(7582) <= (inputs(31)) or (inputs(118));
    layer0_outputs(7583) <= inputs(142);
    layer0_outputs(7584) <= not(inputs(247));
    layer0_outputs(7585) <= (inputs(223)) and not (inputs(33));
    layer0_outputs(7586) <= not(inputs(125));
    layer0_outputs(7587) <= not(inputs(217));
    layer0_outputs(7588) <= not(inputs(196)) or (inputs(86));
    layer0_outputs(7589) <= not((inputs(29)) and (inputs(128)));
    layer0_outputs(7590) <= inputs(170);
    layer0_outputs(7591) <= not(inputs(99));
    layer0_outputs(7592) <= (inputs(172)) or (inputs(159));
    layer0_outputs(7593) <= not(inputs(116)) or (inputs(35));
    layer0_outputs(7594) <= not((inputs(194)) xor (inputs(141)));
    layer0_outputs(7595) <= (inputs(209)) and not (inputs(129));
    layer0_outputs(7596) <= not((inputs(241)) or (inputs(101)));
    layer0_outputs(7597) <= not(inputs(182)) or (inputs(63));
    layer0_outputs(7598) <= not(inputs(184));
    layer0_outputs(7599) <= not(inputs(60)) or (inputs(251));
    layer0_outputs(7600) <= not(inputs(203));
    layer0_outputs(7601) <= not(inputs(217)) or (inputs(246));
    layer0_outputs(7602) <= (inputs(136)) and not (inputs(241));
    layer0_outputs(7603) <= not(inputs(160));
    layer0_outputs(7604) <= not(inputs(222)) or (inputs(208));
    layer0_outputs(7605) <= (inputs(84)) and not (inputs(48));
    layer0_outputs(7606) <= not(inputs(118)) or (inputs(142));
    layer0_outputs(7607) <= not(inputs(146)) or (inputs(104));
    layer0_outputs(7608) <= not(inputs(219)) or (inputs(170));
    layer0_outputs(7609) <= (inputs(160)) or (inputs(157));
    layer0_outputs(7610) <= (inputs(118)) and not (inputs(175));
    layer0_outputs(7611) <= '0';
    layer0_outputs(7612) <= not(inputs(89)) or (inputs(4));
    layer0_outputs(7613) <= (inputs(191)) and not (inputs(32));
    layer0_outputs(7614) <= '1';
    layer0_outputs(7615) <= not(inputs(161)) or (inputs(70));
    layer0_outputs(7616) <= '0';
    layer0_outputs(7617) <= (inputs(198)) or (inputs(73));
    layer0_outputs(7618) <= (inputs(248)) and not (inputs(35));
    layer0_outputs(7619) <= (inputs(232)) and not (inputs(33));
    layer0_outputs(7620) <= not(inputs(204));
    layer0_outputs(7621) <= not(inputs(40)) or (inputs(100));
    layer0_outputs(7622) <= '0';
    layer0_outputs(7623) <= not((inputs(76)) xor (inputs(0)));
    layer0_outputs(7624) <= (inputs(45)) and not (inputs(242));
    layer0_outputs(7625) <= (inputs(91)) or (inputs(63));
    layer0_outputs(7626) <= not((inputs(237)) or (inputs(253)));
    layer0_outputs(7627) <= not(inputs(83));
    layer0_outputs(7628) <= not(inputs(231));
    layer0_outputs(7629) <= inputs(13);
    layer0_outputs(7630) <= '0';
    layer0_outputs(7631) <= not(inputs(59));
    layer0_outputs(7632) <= not((inputs(74)) xor (inputs(173)));
    layer0_outputs(7633) <= (inputs(161)) xor (inputs(230));
    layer0_outputs(7634) <= (inputs(225)) and not (inputs(14));
    layer0_outputs(7635) <= not((inputs(201)) xor (inputs(71)));
    layer0_outputs(7636) <= not(inputs(158));
    layer0_outputs(7637) <= inputs(191);
    layer0_outputs(7638) <= not((inputs(24)) and (inputs(30)));
    layer0_outputs(7639) <= not((inputs(17)) or (inputs(238)));
    layer0_outputs(7640) <= (inputs(235)) or (inputs(110));
    layer0_outputs(7641) <= '1';
    layer0_outputs(7642) <= (inputs(94)) and not (inputs(32));
    layer0_outputs(7643) <= inputs(149);
    layer0_outputs(7644) <= (inputs(156)) or (inputs(65));
    layer0_outputs(7645) <= (inputs(89)) or (inputs(228));
    layer0_outputs(7646) <= inputs(210);
    layer0_outputs(7647) <= (inputs(80)) xor (inputs(103));
    layer0_outputs(7648) <= not(inputs(189));
    layer0_outputs(7649) <= not((inputs(218)) or (inputs(93)));
    layer0_outputs(7650) <= (inputs(76)) and (inputs(9));
    layer0_outputs(7651) <= inputs(109);
    layer0_outputs(7652) <= not(inputs(150)) or (inputs(13));
    layer0_outputs(7653) <= not(inputs(247)) or (inputs(79));
    layer0_outputs(7654) <= not((inputs(94)) or (inputs(238)));
    layer0_outputs(7655) <= inputs(92);
    layer0_outputs(7656) <= not((inputs(104)) or (inputs(60)));
    layer0_outputs(7657) <= inputs(130);
    layer0_outputs(7658) <= (inputs(71)) and not (inputs(76));
    layer0_outputs(7659) <= inputs(164);
    layer0_outputs(7660) <= '1';
    layer0_outputs(7661) <= inputs(118);
    layer0_outputs(7662) <= not((inputs(7)) xor (inputs(78)));
    layer0_outputs(7663) <= not(inputs(234));
    layer0_outputs(7664) <= inputs(101);
    layer0_outputs(7665) <= (inputs(174)) xor (inputs(106));
    layer0_outputs(7666) <= inputs(248);
    layer0_outputs(7667) <= not((inputs(83)) or (inputs(239)));
    layer0_outputs(7668) <= inputs(254);
    layer0_outputs(7669) <= '0';
    layer0_outputs(7670) <= (inputs(76)) and not (inputs(56));
    layer0_outputs(7671) <= (inputs(147)) and not (inputs(51));
    layer0_outputs(7672) <= inputs(183);
    layer0_outputs(7673) <= inputs(134);
    layer0_outputs(7674) <= not(inputs(126));
    layer0_outputs(7675) <= not((inputs(75)) and (inputs(100)));
    layer0_outputs(7676) <= not((inputs(228)) and (inputs(101)));
    layer0_outputs(7677) <= not(inputs(163)) or (inputs(251));
    layer0_outputs(7678) <= inputs(201);
    layer0_outputs(7679) <= not((inputs(118)) or (inputs(173)));
    layer0_outputs(7680) <= not((inputs(180)) or (inputs(62)));
    layer0_outputs(7681) <= inputs(230);
    layer0_outputs(7682) <= not((inputs(134)) or (inputs(29)));
    layer0_outputs(7683) <= inputs(19);
    layer0_outputs(7684) <= not(inputs(183));
    layer0_outputs(7685) <= '1';
    layer0_outputs(7686) <= not(inputs(229));
    layer0_outputs(7687) <= not((inputs(234)) or (inputs(215)));
    layer0_outputs(7688) <= not(inputs(69)) or (inputs(134));
    layer0_outputs(7689) <= not((inputs(135)) and (inputs(227)));
    layer0_outputs(7690) <= (inputs(50)) xor (inputs(6));
    layer0_outputs(7691) <= (inputs(243)) or (inputs(74));
    layer0_outputs(7692) <= (inputs(236)) and (inputs(217));
    layer0_outputs(7693) <= (inputs(145)) or (inputs(247));
    layer0_outputs(7694) <= not(inputs(24)) or (inputs(163));
    layer0_outputs(7695) <= not(inputs(24));
    layer0_outputs(7696) <= '0';
    layer0_outputs(7697) <= (inputs(27)) or (inputs(1));
    layer0_outputs(7698) <= not(inputs(155));
    layer0_outputs(7699) <= not(inputs(196));
    layer0_outputs(7700) <= '1';
    layer0_outputs(7701) <= (inputs(81)) and not (inputs(105));
    layer0_outputs(7702) <= not((inputs(43)) xor (inputs(110)));
    layer0_outputs(7703) <= not(inputs(245));
    layer0_outputs(7704) <= not((inputs(18)) or (inputs(211)));
    layer0_outputs(7705) <= not(inputs(103)) or (inputs(109));
    layer0_outputs(7706) <= '0';
    layer0_outputs(7707) <= (inputs(218)) or (inputs(61));
    layer0_outputs(7708) <= (inputs(201)) or (inputs(239));
    layer0_outputs(7709) <= (inputs(238)) or (inputs(32));
    layer0_outputs(7710) <= not((inputs(154)) or (inputs(190)));
    layer0_outputs(7711) <= (inputs(68)) and not (inputs(172));
    layer0_outputs(7712) <= '1';
    layer0_outputs(7713) <= not(inputs(213));
    layer0_outputs(7714) <= not((inputs(28)) or (inputs(178)));
    layer0_outputs(7715) <= not(inputs(77)) or (inputs(209));
    layer0_outputs(7716) <= not(inputs(54));
    layer0_outputs(7717) <= not(inputs(85)) or (inputs(61));
    layer0_outputs(7718) <= not((inputs(213)) or (inputs(144)));
    layer0_outputs(7719) <= (inputs(135)) and not (inputs(155));
    layer0_outputs(7720) <= not(inputs(102));
    layer0_outputs(7721) <= inputs(180);
    layer0_outputs(7722) <= (inputs(137)) and (inputs(58));
    layer0_outputs(7723) <= not(inputs(188)) or (inputs(66));
    layer0_outputs(7724) <= inputs(106);
    layer0_outputs(7725) <= (inputs(55)) and not (inputs(123));
    layer0_outputs(7726) <= (inputs(141)) or (inputs(156));
    layer0_outputs(7727) <= not((inputs(180)) xor (inputs(129)));
    layer0_outputs(7728) <= (inputs(160)) xor (inputs(162));
    layer0_outputs(7729) <= inputs(234);
    layer0_outputs(7730) <= (inputs(71)) xor (inputs(51));
    layer0_outputs(7731) <= (inputs(33)) and not (inputs(56));
    layer0_outputs(7732) <= not((inputs(150)) or (inputs(31)));
    layer0_outputs(7733) <= (inputs(136)) or (inputs(242));
    layer0_outputs(7734) <= (inputs(63)) or (inputs(201));
    layer0_outputs(7735) <= not((inputs(17)) or (inputs(59)));
    layer0_outputs(7736) <= not(inputs(178));
    layer0_outputs(7737) <= not(inputs(52));
    layer0_outputs(7738) <= inputs(163);
    layer0_outputs(7739) <= inputs(152);
    layer0_outputs(7740) <= not(inputs(106)) or (inputs(194));
    layer0_outputs(7741) <= (inputs(211)) and not (inputs(151));
    layer0_outputs(7742) <= (inputs(187)) and not (inputs(26));
    layer0_outputs(7743) <= not((inputs(129)) or (inputs(170)));
    layer0_outputs(7744) <= inputs(49);
    layer0_outputs(7745) <= not(inputs(51)) or (inputs(173));
    layer0_outputs(7746) <= not((inputs(206)) or (inputs(115)));
    layer0_outputs(7747) <= not((inputs(204)) xor (inputs(80)));
    layer0_outputs(7748) <= (inputs(18)) or (inputs(120));
    layer0_outputs(7749) <= (inputs(19)) and not (inputs(28));
    layer0_outputs(7750) <= (inputs(178)) and not (inputs(14));
    layer0_outputs(7751) <= inputs(164);
    layer0_outputs(7752) <= not((inputs(74)) xor (inputs(146)));
    layer0_outputs(7753) <= (inputs(158)) and not (inputs(62));
    layer0_outputs(7754) <= not((inputs(181)) or (inputs(197)));
    layer0_outputs(7755) <= (inputs(140)) or (inputs(154));
    layer0_outputs(7756) <= inputs(68);
    layer0_outputs(7757) <= not((inputs(66)) or (inputs(43)));
    layer0_outputs(7758) <= (inputs(184)) and not (inputs(227));
    layer0_outputs(7759) <= not((inputs(131)) or (inputs(78)));
    layer0_outputs(7760) <= inputs(79);
    layer0_outputs(7761) <= not(inputs(182));
    layer0_outputs(7762) <= not(inputs(51));
    layer0_outputs(7763) <= not(inputs(72));
    layer0_outputs(7764) <= not((inputs(188)) or (inputs(176)));
    layer0_outputs(7765) <= not(inputs(104));
    layer0_outputs(7766) <= (inputs(167)) and not (inputs(127));
    layer0_outputs(7767) <= inputs(121);
    layer0_outputs(7768) <= not((inputs(211)) or (inputs(210)));
    layer0_outputs(7769) <= not((inputs(122)) or (inputs(42)));
    layer0_outputs(7770) <= not(inputs(72));
    layer0_outputs(7771) <= not(inputs(187));
    layer0_outputs(7772) <= (inputs(27)) and (inputs(119));
    layer0_outputs(7773) <= not((inputs(171)) xor (inputs(142)));
    layer0_outputs(7774) <= not(inputs(225));
    layer0_outputs(7775) <= not((inputs(114)) and (inputs(183)));
    layer0_outputs(7776) <= (inputs(22)) and not (inputs(176));
    layer0_outputs(7777) <= (inputs(147)) and not (inputs(236));
    layer0_outputs(7778) <= not(inputs(150)) or (inputs(29));
    layer0_outputs(7779) <= (inputs(90)) and (inputs(37));
    layer0_outputs(7780) <= (inputs(150)) and not (inputs(232));
    layer0_outputs(7781) <= inputs(85);
    layer0_outputs(7782) <= not((inputs(32)) xor (inputs(157)));
    layer0_outputs(7783) <= not((inputs(235)) xor (inputs(219)));
    layer0_outputs(7784) <= not((inputs(85)) and (inputs(27)));
    layer0_outputs(7785) <= (inputs(11)) or (inputs(112));
    layer0_outputs(7786) <= not((inputs(107)) and (inputs(195)));
    layer0_outputs(7787) <= (inputs(104)) and (inputs(132));
    layer0_outputs(7788) <= '0';
    layer0_outputs(7789) <= '1';
    layer0_outputs(7790) <= not((inputs(236)) xor (inputs(228)));
    layer0_outputs(7791) <= (inputs(33)) and not (inputs(145));
    layer0_outputs(7792) <= inputs(19);
    layer0_outputs(7793) <= not(inputs(179)) or (inputs(121));
    layer0_outputs(7794) <= (inputs(222)) and not (inputs(234));
    layer0_outputs(7795) <= not((inputs(112)) or (inputs(162)));
    layer0_outputs(7796) <= inputs(207);
    layer0_outputs(7797) <= inputs(86);
    layer0_outputs(7798) <= not((inputs(23)) or (inputs(49)));
    layer0_outputs(7799) <= (inputs(175)) or (inputs(248));
    layer0_outputs(7800) <= inputs(169);
    layer0_outputs(7801) <= inputs(24);
    layer0_outputs(7802) <= not((inputs(238)) or (inputs(67)));
    layer0_outputs(7803) <= (inputs(157)) and not (inputs(255));
    layer0_outputs(7804) <= (inputs(255)) xor (inputs(33));
    layer0_outputs(7805) <= not((inputs(21)) or (inputs(65)));
    layer0_outputs(7806) <= not((inputs(203)) xor (inputs(18)));
    layer0_outputs(7807) <= (inputs(65)) xor (inputs(84));
    layer0_outputs(7808) <= not((inputs(135)) and (inputs(242)));
    layer0_outputs(7809) <= (inputs(90)) and not (inputs(187));
    layer0_outputs(7810) <= (inputs(189)) xor (inputs(219));
    layer0_outputs(7811) <= (inputs(144)) and not (inputs(12));
    layer0_outputs(7812) <= inputs(236);
    layer0_outputs(7813) <= not((inputs(77)) xor (inputs(80)));
    layer0_outputs(7814) <= not((inputs(220)) or (inputs(33)));
    layer0_outputs(7815) <= '1';
    layer0_outputs(7816) <= '0';
    layer0_outputs(7817) <= not(inputs(21));
    layer0_outputs(7818) <= not((inputs(104)) or (inputs(38)));
    layer0_outputs(7819) <= inputs(138);
    layer0_outputs(7820) <= not(inputs(179));
    layer0_outputs(7821) <= inputs(51);
    layer0_outputs(7822) <= not(inputs(236));
    layer0_outputs(7823) <= not((inputs(24)) and (inputs(73)));
    layer0_outputs(7824) <= not(inputs(111));
    layer0_outputs(7825) <= inputs(213);
    layer0_outputs(7826) <= (inputs(245)) or (inputs(63));
    layer0_outputs(7827) <= (inputs(230)) and (inputs(162));
    layer0_outputs(7828) <= (inputs(143)) xor (inputs(95));
    layer0_outputs(7829) <= not((inputs(78)) or (inputs(186)));
    layer0_outputs(7830) <= not((inputs(214)) or (inputs(229)));
    layer0_outputs(7831) <= (inputs(182)) or (inputs(68));
    layer0_outputs(7832) <= not((inputs(117)) xor (inputs(196)));
    layer0_outputs(7833) <= not((inputs(162)) or (inputs(187)));
    layer0_outputs(7834) <= (inputs(136)) or (inputs(255));
    layer0_outputs(7835) <= not(inputs(130));
    layer0_outputs(7836) <= not((inputs(230)) xor (inputs(235)));
    layer0_outputs(7837) <= (inputs(242)) xor (inputs(134));
    layer0_outputs(7838) <= not(inputs(8));
    layer0_outputs(7839) <= not(inputs(25));
    layer0_outputs(7840) <= inputs(150);
    layer0_outputs(7841) <= not((inputs(185)) xor (inputs(87)));
    layer0_outputs(7842) <= not(inputs(52));
    layer0_outputs(7843) <= not(inputs(246)) or (inputs(223));
    layer0_outputs(7844) <= not((inputs(22)) or (inputs(136)));
    layer0_outputs(7845) <= not(inputs(101));
    layer0_outputs(7846) <= not((inputs(131)) and (inputs(190)));
    layer0_outputs(7847) <= not(inputs(194)) or (inputs(107));
    layer0_outputs(7848) <= not(inputs(89)) or (inputs(100));
    layer0_outputs(7849) <= not((inputs(168)) and (inputs(144)));
    layer0_outputs(7850) <= inputs(247);
    layer0_outputs(7851) <= not((inputs(29)) or (inputs(220)));
    layer0_outputs(7852) <= (inputs(251)) xor (inputs(44));
    layer0_outputs(7853) <= (inputs(179)) xor (inputs(0));
    layer0_outputs(7854) <= inputs(30);
    layer0_outputs(7855) <= (inputs(28)) xor (inputs(198));
    layer0_outputs(7856) <= not((inputs(233)) or (inputs(81)));
    layer0_outputs(7857) <= inputs(185);
    layer0_outputs(7858) <= inputs(146);
    layer0_outputs(7859) <= inputs(89);
    layer0_outputs(7860) <= inputs(231);
    layer0_outputs(7861) <= not(inputs(101)) or (inputs(224));
    layer0_outputs(7862) <= inputs(93);
    layer0_outputs(7863) <= (inputs(119)) and not (inputs(58));
    layer0_outputs(7864) <= '0';
    layer0_outputs(7865) <= inputs(75);
    layer0_outputs(7866) <= not(inputs(92));
    layer0_outputs(7867) <= not(inputs(155));
    layer0_outputs(7868) <= (inputs(114)) or (inputs(145));
    layer0_outputs(7869) <= not(inputs(117));
    layer0_outputs(7870) <= inputs(34);
    layer0_outputs(7871) <= not(inputs(39));
    layer0_outputs(7872) <= not(inputs(247));
    layer0_outputs(7873) <= not((inputs(27)) or (inputs(26)));
    layer0_outputs(7874) <= inputs(98);
    layer0_outputs(7875) <= not(inputs(76));
    layer0_outputs(7876) <= (inputs(231)) and not (inputs(34));
    layer0_outputs(7877) <= (inputs(19)) and not (inputs(128));
    layer0_outputs(7878) <= not(inputs(245)) or (inputs(84));
    layer0_outputs(7879) <= inputs(95);
    layer0_outputs(7880) <= not(inputs(25));
    layer0_outputs(7881) <= (inputs(86)) or (inputs(51));
    layer0_outputs(7882) <= not(inputs(231));
    layer0_outputs(7883) <= not(inputs(228)) or (inputs(97));
    layer0_outputs(7884) <= '1';
    layer0_outputs(7885) <= inputs(7);
    layer0_outputs(7886) <= not(inputs(93)) or (inputs(116));
    layer0_outputs(7887) <= '0';
    layer0_outputs(7888) <= not((inputs(114)) xor (inputs(6)));
    layer0_outputs(7889) <= not(inputs(228));
    layer0_outputs(7890) <= inputs(189);
    layer0_outputs(7891) <= (inputs(98)) and not (inputs(144));
    layer0_outputs(7892) <= not((inputs(181)) or (inputs(70)));
    layer0_outputs(7893) <= not((inputs(64)) and (inputs(82)));
    layer0_outputs(7894) <= not(inputs(73));
    layer0_outputs(7895) <= not(inputs(91));
    layer0_outputs(7896) <= not((inputs(217)) or (inputs(17)));
    layer0_outputs(7897) <= (inputs(215)) and not (inputs(154));
    layer0_outputs(7898) <= (inputs(198)) and (inputs(61));
    layer0_outputs(7899) <= not((inputs(197)) xor (inputs(100)));
    layer0_outputs(7900) <= (inputs(52)) or (inputs(125));
    layer0_outputs(7901) <= not(inputs(217));
    layer0_outputs(7902) <= not(inputs(164));
    layer0_outputs(7903) <= inputs(112);
    layer0_outputs(7904) <= not((inputs(203)) or (inputs(185)));
    layer0_outputs(7905) <= not((inputs(177)) xor (inputs(225)));
    layer0_outputs(7906) <= (inputs(135)) and not (inputs(197));
    layer0_outputs(7907) <= not(inputs(202));
    layer0_outputs(7908) <= not((inputs(26)) and (inputs(217)));
    layer0_outputs(7909) <= (inputs(244)) xor (inputs(77));
    layer0_outputs(7910) <= not((inputs(116)) xor (inputs(145)));
    layer0_outputs(7911) <= (inputs(213)) and not (inputs(71));
    layer0_outputs(7912) <= not(inputs(83)) or (inputs(176));
    layer0_outputs(7913) <= not(inputs(121)) or (inputs(224));
    layer0_outputs(7914) <= not(inputs(213)) or (inputs(115));
    layer0_outputs(7915) <= (inputs(237)) or (inputs(238));
    layer0_outputs(7916) <= (inputs(37)) and (inputs(39));
    layer0_outputs(7917) <= (inputs(25)) and not (inputs(254));
    layer0_outputs(7918) <= (inputs(155)) xor (inputs(3));
    layer0_outputs(7919) <= not((inputs(214)) or (inputs(88)));
    layer0_outputs(7920) <= inputs(148);
    layer0_outputs(7921) <= not(inputs(33));
    layer0_outputs(7922) <= not(inputs(43)) or (inputs(123));
    layer0_outputs(7923) <= (inputs(103)) xor (inputs(108));
    layer0_outputs(7924) <= inputs(100);
    layer0_outputs(7925) <= not((inputs(197)) or (inputs(12)));
    layer0_outputs(7926) <= not(inputs(48)) or (inputs(170));
    layer0_outputs(7927) <= not(inputs(63)) or (inputs(128));
    layer0_outputs(7928) <= not((inputs(245)) and (inputs(76)));
    layer0_outputs(7929) <= not(inputs(91)) or (inputs(176));
    layer0_outputs(7930) <= inputs(53);
    layer0_outputs(7931) <= '0';
    layer0_outputs(7932) <= inputs(139);
    layer0_outputs(7933) <= not((inputs(168)) xor (inputs(230)));
    layer0_outputs(7934) <= not((inputs(2)) or (inputs(23)));
    layer0_outputs(7935) <= (inputs(186)) and not (inputs(139));
    layer0_outputs(7936) <= inputs(234);
    layer0_outputs(7937) <= not((inputs(176)) or (inputs(5)));
    layer0_outputs(7938) <= not((inputs(79)) or (inputs(160)));
    layer0_outputs(7939) <= not(inputs(37)) or (inputs(101));
    layer0_outputs(7940) <= not((inputs(79)) xor (inputs(110)));
    layer0_outputs(7941) <= not(inputs(117)) or (inputs(221));
    layer0_outputs(7942) <= not(inputs(194)) or (inputs(8));
    layer0_outputs(7943) <= not((inputs(172)) xor (inputs(251)));
    layer0_outputs(7944) <= not(inputs(60)) or (inputs(191));
    layer0_outputs(7945) <= inputs(94);
    layer0_outputs(7946) <= inputs(104);
    layer0_outputs(7947) <= '1';
    layer0_outputs(7948) <= (inputs(255)) or (inputs(154));
    layer0_outputs(7949) <= (inputs(102)) or (inputs(193));
    layer0_outputs(7950) <= not(inputs(75));
    layer0_outputs(7951) <= inputs(13);
    layer0_outputs(7952) <= not(inputs(89)) or (inputs(100));
    layer0_outputs(7953) <= not((inputs(104)) or (inputs(151)));
    layer0_outputs(7954) <= (inputs(114)) and not (inputs(107));
    layer0_outputs(7955) <= not((inputs(85)) or (inputs(206)));
    layer0_outputs(7956) <= not((inputs(173)) xor (inputs(254)));
    layer0_outputs(7957) <= (inputs(175)) xor (inputs(145));
    layer0_outputs(7958) <= not((inputs(47)) or (inputs(44)));
    layer0_outputs(7959) <= inputs(95);
    layer0_outputs(7960) <= '1';
    layer0_outputs(7961) <= not(inputs(121));
    layer0_outputs(7962) <= not(inputs(219));
    layer0_outputs(7963) <= (inputs(6)) or (inputs(44));
    layer0_outputs(7964) <= not(inputs(4)) or (inputs(44));
    layer0_outputs(7965) <= (inputs(139)) and (inputs(129));
    layer0_outputs(7966) <= not((inputs(158)) or (inputs(214)));
    layer0_outputs(7967) <= (inputs(158)) and not (inputs(49));
    layer0_outputs(7968) <= (inputs(239)) or (inputs(20));
    layer0_outputs(7969) <= not(inputs(145));
    layer0_outputs(7970) <= not(inputs(145));
    layer0_outputs(7971) <= (inputs(38)) or (inputs(31));
    layer0_outputs(7972) <= not(inputs(20)) or (inputs(247));
    layer0_outputs(7973) <= not((inputs(26)) and (inputs(13)));
    layer0_outputs(7974) <= not(inputs(218));
    layer0_outputs(7975) <= not((inputs(207)) xor (inputs(251)));
    layer0_outputs(7976) <= (inputs(239)) or (inputs(165));
    layer0_outputs(7977) <= not(inputs(33));
    layer0_outputs(7978) <= (inputs(69)) or (inputs(147));
    layer0_outputs(7979) <= inputs(93);
    layer0_outputs(7980) <= not(inputs(101));
    layer0_outputs(7981) <= not(inputs(88));
    layer0_outputs(7982) <= not(inputs(146));
    layer0_outputs(7983) <= not(inputs(136));
    layer0_outputs(7984) <= inputs(133);
    layer0_outputs(7985) <= inputs(68);
    layer0_outputs(7986) <= (inputs(136)) and (inputs(83));
    layer0_outputs(7987) <= inputs(161);
    layer0_outputs(7988) <= inputs(188);
    layer0_outputs(7989) <= inputs(108);
    layer0_outputs(7990) <= not((inputs(147)) or (inputs(130)));
    layer0_outputs(7991) <= not(inputs(69)) or (inputs(173));
    layer0_outputs(7992) <= not(inputs(23));
    layer0_outputs(7993) <= not(inputs(27)) or (inputs(144));
    layer0_outputs(7994) <= (inputs(181)) and not (inputs(114));
    layer0_outputs(7995) <= not((inputs(216)) and (inputs(155)));
    layer0_outputs(7996) <= not(inputs(153));
    layer0_outputs(7997) <= (inputs(229)) and not (inputs(47));
    layer0_outputs(7998) <= not((inputs(238)) or (inputs(121)));
    layer0_outputs(7999) <= not(inputs(108));
    layer0_outputs(8000) <= not(inputs(78)) or (inputs(238));
    layer0_outputs(8001) <= not((inputs(175)) or (inputs(228)));
    layer0_outputs(8002) <= (inputs(195)) and not (inputs(63));
    layer0_outputs(8003) <= (inputs(21)) or (inputs(124));
    layer0_outputs(8004) <= not(inputs(207)) or (inputs(138));
    layer0_outputs(8005) <= (inputs(102)) xor (inputs(97));
    layer0_outputs(8006) <= inputs(67);
    layer0_outputs(8007) <= not(inputs(168));
    layer0_outputs(8008) <= not((inputs(118)) or (inputs(181)));
    layer0_outputs(8009) <= (inputs(106)) and not (inputs(234));
    layer0_outputs(8010) <= not((inputs(211)) or (inputs(195)));
    layer0_outputs(8011) <= inputs(32);
    layer0_outputs(8012) <= not(inputs(72)) or (inputs(224));
    layer0_outputs(8013) <= not((inputs(158)) and (inputs(121)));
    layer0_outputs(8014) <= '1';
    layer0_outputs(8015) <= not((inputs(32)) or (inputs(224)));
    layer0_outputs(8016) <= not((inputs(221)) xor (inputs(122)));
    layer0_outputs(8017) <= not((inputs(21)) or (inputs(195)));
    layer0_outputs(8018) <= not((inputs(158)) or (inputs(210)));
    layer0_outputs(8019) <= inputs(250);
    layer0_outputs(8020) <= not(inputs(113));
    layer0_outputs(8021) <= inputs(105);
    layer0_outputs(8022) <= not(inputs(11));
    layer0_outputs(8023) <= not(inputs(42)) or (inputs(25));
    layer0_outputs(8024) <= not((inputs(1)) or (inputs(142)));
    layer0_outputs(8025) <= (inputs(8)) or (inputs(65));
    layer0_outputs(8026) <= inputs(194);
    layer0_outputs(8027) <= not((inputs(243)) or (inputs(191)));
    layer0_outputs(8028) <= not(inputs(4)) or (inputs(66));
    layer0_outputs(8029) <= inputs(46);
    layer0_outputs(8030) <= (inputs(135)) and (inputs(109));
    layer0_outputs(8031) <= not(inputs(226)) or (inputs(29));
    layer0_outputs(8032) <= inputs(174);
    layer0_outputs(8033) <= not((inputs(150)) or (inputs(166)));
    layer0_outputs(8034) <= (inputs(42)) and not (inputs(252));
    layer0_outputs(8035) <= not(inputs(222)) or (inputs(47));
    layer0_outputs(8036) <= not(inputs(66));
    layer0_outputs(8037) <= not((inputs(23)) xor (inputs(79)));
    layer0_outputs(8038) <= '0';
    layer0_outputs(8039) <= inputs(70);
    layer0_outputs(8040) <= not(inputs(190)) or (inputs(89));
    layer0_outputs(8041) <= (inputs(179)) and not (inputs(30));
    layer0_outputs(8042) <= not((inputs(186)) xor (inputs(121)));
    layer0_outputs(8043) <= not(inputs(9)) or (inputs(182));
    layer0_outputs(8044) <= (inputs(124)) and (inputs(88));
    layer0_outputs(8045) <= '1';
    layer0_outputs(8046) <= (inputs(116)) xor (inputs(235));
    layer0_outputs(8047) <= not((inputs(233)) and (inputs(220)));
    layer0_outputs(8048) <= (inputs(18)) xor (inputs(43));
    layer0_outputs(8049) <= (inputs(204)) and not (inputs(92));
    layer0_outputs(8050) <= (inputs(17)) and not (inputs(254));
    layer0_outputs(8051) <= not((inputs(6)) xor (inputs(70)));
    layer0_outputs(8052) <= not((inputs(2)) xor (inputs(91)));
    layer0_outputs(8053) <= not(inputs(122)) or (inputs(112));
    layer0_outputs(8054) <= not(inputs(193)) or (inputs(11));
    layer0_outputs(8055) <= not(inputs(101));
    layer0_outputs(8056) <= not(inputs(116)) or (inputs(33));
    layer0_outputs(8057) <= '0';
    layer0_outputs(8058) <= not((inputs(89)) or (inputs(177)));
    layer0_outputs(8059) <= '1';
    layer0_outputs(8060) <= not((inputs(226)) or (inputs(254)));
    layer0_outputs(8061) <= (inputs(163)) or (inputs(235));
    layer0_outputs(8062) <= '0';
    layer0_outputs(8063) <= not(inputs(170)) or (inputs(40));
    layer0_outputs(8064) <= not(inputs(118));
    layer0_outputs(8065) <= not((inputs(177)) xor (inputs(139)));
    layer0_outputs(8066) <= '0';
    layer0_outputs(8067) <= not((inputs(170)) and (inputs(47)));
    layer0_outputs(8068) <= not((inputs(116)) or (inputs(193)));
    layer0_outputs(8069) <= not((inputs(111)) or (inputs(21)));
    layer0_outputs(8070) <= not(inputs(201)) or (inputs(242));
    layer0_outputs(8071) <= '1';
    layer0_outputs(8072) <= inputs(120);
    layer0_outputs(8073) <= not(inputs(230));
    layer0_outputs(8074) <= (inputs(173)) or (inputs(175));
    layer0_outputs(8075) <= not((inputs(22)) or (inputs(32)));
    layer0_outputs(8076) <= not((inputs(68)) xor (inputs(81)));
    layer0_outputs(8077) <= not((inputs(173)) xor (inputs(122)));
    layer0_outputs(8078) <= not((inputs(207)) or (inputs(188)));
    layer0_outputs(8079) <= '1';
    layer0_outputs(8080) <= not(inputs(126));
    layer0_outputs(8081) <= not(inputs(37)) or (inputs(235));
    layer0_outputs(8082) <= not(inputs(163)) or (inputs(15));
    layer0_outputs(8083) <= not(inputs(154));
    layer0_outputs(8084) <= inputs(100);
    layer0_outputs(8085) <= (inputs(221)) and not (inputs(111));
    layer0_outputs(8086) <= inputs(195);
    layer0_outputs(8087) <= '0';
    layer0_outputs(8088) <= not((inputs(236)) xor (inputs(225)));
    layer0_outputs(8089) <= (inputs(226)) or (inputs(21));
    layer0_outputs(8090) <= (inputs(21)) and not (inputs(142));
    layer0_outputs(8091) <= (inputs(72)) or (inputs(182));
    layer0_outputs(8092) <= not(inputs(93)) or (inputs(63));
    layer0_outputs(8093) <= not(inputs(200));
    layer0_outputs(8094) <= not(inputs(208));
    layer0_outputs(8095) <= not((inputs(23)) or (inputs(246)));
    layer0_outputs(8096) <= (inputs(19)) and not (inputs(144));
    layer0_outputs(8097) <= not((inputs(91)) or (inputs(49)));
    layer0_outputs(8098) <= inputs(147);
    layer0_outputs(8099) <= inputs(77);
    layer0_outputs(8100) <= not(inputs(129));
    layer0_outputs(8101) <= (inputs(129)) and not (inputs(254));
    layer0_outputs(8102) <= inputs(75);
    layer0_outputs(8103) <= not(inputs(236)) or (inputs(124));
    layer0_outputs(8104) <= not(inputs(40));
    layer0_outputs(8105) <= not(inputs(7));
    layer0_outputs(8106) <= not(inputs(243)) or (inputs(74));
    layer0_outputs(8107) <= not(inputs(60)) or (inputs(16));
    layer0_outputs(8108) <= not((inputs(64)) or (inputs(205)));
    layer0_outputs(8109) <= not(inputs(210));
    layer0_outputs(8110) <= not(inputs(136)) or (inputs(232));
    layer0_outputs(8111) <= not(inputs(99));
    layer0_outputs(8112) <= not(inputs(255)) or (inputs(163));
    layer0_outputs(8113) <= (inputs(155)) xor (inputs(188));
    layer0_outputs(8114) <= not(inputs(24));
    layer0_outputs(8115) <= not(inputs(154));
    layer0_outputs(8116) <= not(inputs(168)) or (inputs(103));
    layer0_outputs(8117) <= (inputs(237)) xor (inputs(82));
    layer0_outputs(8118) <= (inputs(236)) or (inputs(48));
    layer0_outputs(8119) <= inputs(52);
    layer0_outputs(8120) <= (inputs(1)) and (inputs(134));
    layer0_outputs(8121) <= (inputs(224)) or (inputs(4));
    layer0_outputs(8122) <= (inputs(154)) or (inputs(54));
    layer0_outputs(8123) <= inputs(25);
    layer0_outputs(8124) <= not((inputs(46)) or (inputs(96)));
    layer0_outputs(8125) <= '0';
    layer0_outputs(8126) <= (inputs(242)) and not (inputs(234));
    layer0_outputs(8127) <= inputs(169);
    layer0_outputs(8128) <= inputs(180);
    layer0_outputs(8129) <= not(inputs(166));
    layer0_outputs(8130) <= not((inputs(239)) xor (inputs(52)));
    layer0_outputs(8131) <= inputs(66);
    layer0_outputs(8132) <= (inputs(234)) and (inputs(166));
    layer0_outputs(8133) <= (inputs(38)) and (inputs(38));
    layer0_outputs(8134) <= not((inputs(12)) or (inputs(36)));
    layer0_outputs(8135) <= inputs(19);
    layer0_outputs(8136) <= (inputs(171)) xor (inputs(76));
    layer0_outputs(8137) <= inputs(39);
    layer0_outputs(8138) <= not(inputs(15)) or (inputs(119));
    layer0_outputs(8139) <= not(inputs(60));
    layer0_outputs(8140) <= '0';
    layer0_outputs(8141) <= not(inputs(183)) or (inputs(94));
    layer0_outputs(8142) <= not((inputs(76)) or (inputs(23)));
    layer0_outputs(8143) <= not(inputs(145));
    layer0_outputs(8144) <= (inputs(95)) or (inputs(58));
    layer0_outputs(8145) <= not(inputs(59)) or (inputs(191));
    layer0_outputs(8146) <= inputs(86);
    layer0_outputs(8147) <= (inputs(184)) and (inputs(3));
    layer0_outputs(8148) <= (inputs(29)) xor (inputs(17));
    layer0_outputs(8149) <= not((inputs(82)) or (inputs(246)));
    layer0_outputs(8150) <= not((inputs(52)) or (inputs(211)));
    layer0_outputs(8151) <= (inputs(204)) and not (inputs(145));
    layer0_outputs(8152) <= not(inputs(246)) or (inputs(93));
    layer0_outputs(8153) <= not(inputs(187));
    layer0_outputs(8154) <= (inputs(137)) and not (inputs(236));
    layer0_outputs(8155) <= not((inputs(234)) or (inputs(225)));
    layer0_outputs(8156) <= not((inputs(255)) or (inputs(245)));
    layer0_outputs(8157) <= not(inputs(143));
    layer0_outputs(8158) <= inputs(198);
    layer0_outputs(8159) <= not((inputs(235)) or (inputs(242)));
    layer0_outputs(8160) <= '1';
    layer0_outputs(8161) <= not(inputs(112)) or (inputs(236));
    layer0_outputs(8162) <= not(inputs(6));
    layer0_outputs(8163) <= not(inputs(172));
    layer0_outputs(8164) <= '1';
    layer0_outputs(8165) <= not(inputs(166));
    layer0_outputs(8166) <= (inputs(152)) and not (inputs(78));
    layer0_outputs(8167) <= not((inputs(194)) xor (inputs(164)));
    layer0_outputs(8168) <= inputs(1);
    layer0_outputs(8169) <= (inputs(244)) or (inputs(47));
    layer0_outputs(8170) <= not((inputs(168)) or (inputs(199)));
    layer0_outputs(8171) <= (inputs(85)) or (inputs(130));
    layer0_outputs(8172) <= not(inputs(198));
    layer0_outputs(8173) <= not((inputs(214)) or (inputs(230)));
    layer0_outputs(8174) <= (inputs(224)) xor (inputs(248));
    layer0_outputs(8175) <= inputs(195);
    layer0_outputs(8176) <= not((inputs(167)) xor (inputs(237)));
    layer0_outputs(8177) <= not(inputs(30)) or (inputs(255));
    layer0_outputs(8178) <= not((inputs(108)) or (inputs(100)));
    layer0_outputs(8179) <= not(inputs(99));
    layer0_outputs(8180) <= '0';
    layer0_outputs(8181) <= (inputs(195)) and not (inputs(129));
    layer0_outputs(8182) <= not((inputs(191)) or (inputs(146)));
    layer0_outputs(8183) <= (inputs(150)) and (inputs(203));
    layer0_outputs(8184) <= not(inputs(163));
    layer0_outputs(8185) <= inputs(90);
    layer0_outputs(8186) <= not(inputs(89)) or (inputs(16));
    layer0_outputs(8187) <= not(inputs(23)) or (inputs(176));
    layer0_outputs(8188) <= '0';
    layer0_outputs(8189) <= inputs(217);
    layer0_outputs(8190) <= (inputs(165)) or (inputs(165));
    layer0_outputs(8191) <= (inputs(136)) or (inputs(30));
    layer0_outputs(8192) <= inputs(163);
    layer0_outputs(8193) <= (inputs(250)) and not (inputs(208));
    layer0_outputs(8194) <= (inputs(169)) xor (inputs(236));
    layer0_outputs(8195) <= not(inputs(65)) or (inputs(159));
    layer0_outputs(8196) <= inputs(215);
    layer0_outputs(8197) <= not((inputs(236)) and (inputs(249)));
    layer0_outputs(8198) <= not((inputs(23)) or (inputs(96)));
    layer0_outputs(8199) <= (inputs(195)) and not (inputs(111));
    layer0_outputs(8200) <= not(inputs(29));
    layer0_outputs(8201) <= (inputs(227)) or (inputs(72));
    layer0_outputs(8202) <= not(inputs(103)) or (inputs(254));
    layer0_outputs(8203) <= not((inputs(229)) or (inputs(253)));
    layer0_outputs(8204) <= inputs(233);
    layer0_outputs(8205) <= not((inputs(17)) xor (inputs(135)));
    layer0_outputs(8206) <= not((inputs(35)) xor (inputs(154)));
    layer0_outputs(8207) <= (inputs(37)) and not (inputs(252));
    layer0_outputs(8208) <= '0';
    layer0_outputs(8209) <= (inputs(235)) or (inputs(141));
    layer0_outputs(8210) <= inputs(129);
    layer0_outputs(8211) <= (inputs(207)) xor (inputs(121));
    layer0_outputs(8212) <= not(inputs(157));
    layer0_outputs(8213) <= (inputs(184)) xor (inputs(154));
    layer0_outputs(8214) <= (inputs(222)) xor (inputs(249));
    layer0_outputs(8215) <= not((inputs(138)) and (inputs(153)));
    layer0_outputs(8216) <= inputs(72);
    layer0_outputs(8217) <= not((inputs(199)) or (inputs(125)));
    layer0_outputs(8218) <= inputs(180);
    layer0_outputs(8219) <= (inputs(38)) and not (inputs(220));
    layer0_outputs(8220) <= inputs(51);
    layer0_outputs(8221) <= (inputs(47)) or (inputs(92));
    layer0_outputs(8222) <= not(inputs(45)) or (inputs(83));
    layer0_outputs(8223) <= (inputs(85)) and not (inputs(212));
    layer0_outputs(8224) <= inputs(37);
    layer0_outputs(8225) <= (inputs(81)) or (inputs(16));
    layer0_outputs(8226) <= not(inputs(102));
    layer0_outputs(8227) <= not((inputs(21)) xor (inputs(51)));
    layer0_outputs(8228) <= not((inputs(100)) or (inputs(211)));
    layer0_outputs(8229) <= not(inputs(231)) or (inputs(93));
    layer0_outputs(8230) <= (inputs(194)) and not (inputs(236));
    layer0_outputs(8231) <= inputs(30);
    layer0_outputs(8232) <= inputs(129);
    layer0_outputs(8233) <= (inputs(181)) and not (inputs(24));
    layer0_outputs(8234) <= (inputs(170)) and not (inputs(134));
    layer0_outputs(8235) <= inputs(210);
    layer0_outputs(8236) <= not(inputs(40)) or (inputs(212));
    layer0_outputs(8237) <= (inputs(119)) and not (inputs(164));
    layer0_outputs(8238) <= not(inputs(4)) or (inputs(35));
    layer0_outputs(8239) <= (inputs(150)) and not (inputs(56));
    layer0_outputs(8240) <= not(inputs(194));
    layer0_outputs(8241) <= inputs(215);
    layer0_outputs(8242) <= (inputs(52)) and not (inputs(26));
    layer0_outputs(8243) <= not((inputs(55)) xor (inputs(8)));
    layer0_outputs(8244) <= (inputs(134)) and not (inputs(111));
    layer0_outputs(8245) <= inputs(9);
    layer0_outputs(8246) <= not(inputs(23));
    layer0_outputs(8247) <= (inputs(188)) xor (inputs(192));
    layer0_outputs(8248) <= not(inputs(92)) or (inputs(248));
    layer0_outputs(8249) <= (inputs(211)) and not (inputs(13));
    layer0_outputs(8250) <= not(inputs(56));
    layer0_outputs(8251) <= (inputs(84)) and not (inputs(239));
    layer0_outputs(8252) <= '1';
    layer0_outputs(8253) <= not((inputs(129)) or (inputs(84)));
    layer0_outputs(8254) <= not(inputs(85)) or (inputs(78));
    layer0_outputs(8255) <= (inputs(251)) and not (inputs(250));
    layer0_outputs(8256) <= (inputs(107)) or (inputs(52));
    layer0_outputs(8257) <= (inputs(81)) xor (inputs(189));
    layer0_outputs(8258) <= not((inputs(26)) and (inputs(64)));
    layer0_outputs(8259) <= not((inputs(175)) and (inputs(81)));
    layer0_outputs(8260) <= (inputs(144)) or (inputs(112));
    layer0_outputs(8261) <= not((inputs(30)) and (inputs(11)));
    layer0_outputs(8262) <= not((inputs(59)) or (inputs(75)));
    layer0_outputs(8263) <= not(inputs(82));
    layer0_outputs(8264) <= not(inputs(112));
    layer0_outputs(8265) <= not(inputs(104)) or (inputs(113));
    layer0_outputs(8266) <= '1';
    layer0_outputs(8267) <= not((inputs(78)) or (inputs(59)));
    layer0_outputs(8268) <= not(inputs(44)) or (inputs(187));
    layer0_outputs(8269) <= inputs(195);
    layer0_outputs(8270) <= inputs(169);
    layer0_outputs(8271) <= not((inputs(108)) and (inputs(231)));
    layer0_outputs(8272) <= (inputs(13)) or (inputs(15));
    layer0_outputs(8273) <= not(inputs(168));
    layer0_outputs(8274) <= '1';
    layer0_outputs(8275) <= '0';
    layer0_outputs(8276) <= not((inputs(221)) xor (inputs(237)));
    layer0_outputs(8277) <= not(inputs(122)) or (inputs(57));
    layer0_outputs(8278) <= (inputs(147)) or (inputs(238));
    layer0_outputs(8279) <= not(inputs(193));
    layer0_outputs(8280) <= (inputs(255)) or (inputs(237));
    layer0_outputs(8281) <= not((inputs(23)) or (inputs(33)));
    layer0_outputs(8282) <= not(inputs(171)) or (inputs(131));
    layer0_outputs(8283) <= (inputs(71)) xor (inputs(197));
    layer0_outputs(8284) <= inputs(20);
    layer0_outputs(8285) <= not(inputs(139));
    layer0_outputs(8286) <= not(inputs(168)) or (inputs(186));
    layer0_outputs(8287) <= not((inputs(229)) xor (inputs(96)));
    layer0_outputs(8288) <= not((inputs(32)) or (inputs(199)));
    layer0_outputs(8289) <= not(inputs(167)) or (inputs(101));
    layer0_outputs(8290) <= not((inputs(218)) or (inputs(190)));
    layer0_outputs(8291) <= (inputs(133)) and (inputs(153));
    layer0_outputs(8292) <= (inputs(150)) or (inputs(134));
    layer0_outputs(8293) <= (inputs(76)) or (inputs(160));
    layer0_outputs(8294) <= (inputs(60)) and not (inputs(238));
    layer0_outputs(8295) <= not(inputs(245)) or (inputs(48));
    layer0_outputs(8296) <= '1';
    layer0_outputs(8297) <= not((inputs(142)) or (inputs(205)));
    layer0_outputs(8298) <= inputs(83);
    layer0_outputs(8299) <= (inputs(105)) xor (inputs(73));
    layer0_outputs(8300) <= (inputs(34)) xor (inputs(97));
    layer0_outputs(8301) <= not(inputs(105));
    layer0_outputs(8302) <= (inputs(180)) and not (inputs(37));
    layer0_outputs(8303) <= (inputs(52)) or (inputs(207));
    layer0_outputs(8304) <= inputs(49);
    layer0_outputs(8305) <= inputs(137);
    layer0_outputs(8306) <= (inputs(110)) and not (inputs(96));
    layer0_outputs(8307) <= not(inputs(196));
    layer0_outputs(8308) <= not(inputs(137)) or (inputs(22));
    layer0_outputs(8309) <= (inputs(0)) and (inputs(131));
    layer0_outputs(8310) <= not((inputs(204)) or (inputs(207)));
    layer0_outputs(8311) <= not(inputs(108)) or (inputs(37));
    layer0_outputs(8312) <= (inputs(37)) and not (inputs(224));
    layer0_outputs(8313) <= (inputs(70)) or (inputs(32));
    layer0_outputs(8314) <= (inputs(212)) or (inputs(177));
    layer0_outputs(8315) <= (inputs(107)) xor (inputs(111));
    layer0_outputs(8316) <= inputs(90);
    layer0_outputs(8317) <= not(inputs(183)) or (inputs(114));
    layer0_outputs(8318) <= not((inputs(80)) xor (inputs(77)));
    layer0_outputs(8319) <= not((inputs(241)) or (inputs(94)));
    layer0_outputs(8320) <= inputs(234);
    layer0_outputs(8321) <= not((inputs(243)) and (inputs(202)));
    layer0_outputs(8322) <= not(inputs(10));
    layer0_outputs(8323) <= not(inputs(51));
    layer0_outputs(8324) <= not(inputs(119));
    layer0_outputs(8325) <= (inputs(238)) and (inputs(64));
    layer0_outputs(8326) <= (inputs(47)) and (inputs(212));
    layer0_outputs(8327) <= not(inputs(95));
    layer0_outputs(8328) <= not(inputs(105)) or (inputs(113));
    layer0_outputs(8329) <= not((inputs(62)) and (inputs(211)));
    layer0_outputs(8330) <= (inputs(50)) or (inputs(158));
    layer0_outputs(8331) <= (inputs(1)) and (inputs(81));
    layer0_outputs(8332) <= not((inputs(64)) xor (inputs(52)));
    layer0_outputs(8333) <= not(inputs(156)) or (inputs(194));
    layer0_outputs(8334) <= (inputs(52)) or (inputs(190));
    layer0_outputs(8335) <= not((inputs(129)) xor (inputs(147)));
    layer0_outputs(8336) <= (inputs(135)) and not (inputs(65));
    layer0_outputs(8337) <= not((inputs(208)) and (inputs(185)));
    layer0_outputs(8338) <= not(inputs(139));
    layer0_outputs(8339) <= inputs(239);
    layer0_outputs(8340) <= (inputs(137)) and (inputs(155));
    layer0_outputs(8341) <= '0';
    layer0_outputs(8342) <= not((inputs(76)) and (inputs(103)));
    layer0_outputs(8343) <= (inputs(126)) xor (inputs(11));
    layer0_outputs(8344) <= inputs(212);
    layer0_outputs(8345) <= not((inputs(179)) or (inputs(144)));
    layer0_outputs(8346) <= '1';
    layer0_outputs(8347) <= not(inputs(105));
    layer0_outputs(8348) <= (inputs(152)) xor (inputs(138));
    layer0_outputs(8349) <= inputs(150);
    layer0_outputs(8350) <= inputs(230);
    layer0_outputs(8351) <= (inputs(242)) or (inputs(97));
    layer0_outputs(8352) <= (inputs(98)) or (inputs(110));
    layer0_outputs(8353) <= (inputs(117)) xor (inputs(131));
    layer0_outputs(8354) <= (inputs(135)) and not (inputs(84));
    layer0_outputs(8355) <= '0';
    layer0_outputs(8356) <= not((inputs(148)) or (inputs(165)));
    layer0_outputs(8357) <= '1';
    layer0_outputs(8358) <= not((inputs(225)) xor (inputs(151)));
    layer0_outputs(8359) <= (inputs(8)) or (inputs(28));
    layer0_outputs(8360) <= (inputs(2)) or (inputs(139));
    layer0_outputs(8361) <= not((inputs(3)) and (inputs(127)));
    layer0_outputs(8362) <= not(inputs(216)) or (inputs(135));
    layer0_outputs(8363) <= not((inputs(90)) xor (inputs(110)));
    layer0_outputs(8364) <= not(inputs(230));
    layer0_outputs(8365) <= not(inputs(10)) or (inputs(74));
    layer0_outputs(8366) <= not((inputs(252)) xor (inputs(253)));
    layer0_outputs(8367) <= (inputs(42)) and not (inputs(147));
    layer0_outputs(8368) <= '1';
    layer0_outputs(8369) <= not(inputs(35));
    layer0_outputs(8370) <= '1';
    layer0_outputs(8371) <= not(inputs(83));
    layer0_outputs(8372) <= not(inputs(40)) or (inputs(19));
    layer0_outputs(8373) <= not(inputs(126)) or (inputs(212));
    layer0_outputs(8374) <= not((inputs(108)) or (inputs(128)));
    layer0_outputs(8375) <= (inputs(68)) and not (inputs(8));
    layer0_outputs(8376) <= inputs(159);
    layer0_outputs(8377) <= not(inputs(149)) or (inputs(80));
    layer0_outputs(8378) <= not(inputs(134)) or (inputs(155));
    layer0_outputs(8379) <= inputs(234);
    layer0_outputs(8380) <= inputs(147);
    layer0_outputs(8381) <= not(inputs(25));
    layer0_outputs(8382) <= not((inputs(235)) or (inputs(11)));
    layer0_outputs(8383) <= (inputs(10)) or (inputs(171));
    layer0_outputs(8384) <= not(inputs(6)) or (inputs(197));
    layer0_outputs(8385) <= not(inputs(15)) or (inputs(63));
    layer0_outputs(8386) <= '1';
    layer0_outputs(8387) <= (inputs(31)) or (inputs(20));
    layer0_outputs(8388) <= (inputs(230)) or (inputs(248));
    layer0_outputs(8389) <= not(inputs(98));
    layer0_outputs(8390) <= (inputs(73)) and not (inputs(165));
    layer0_outputs(8391) <= (inputs(138)) and not (inputs(24));
    layer0_outputs(8392) <= inputs(74);
    layer0_outputs(8393) <= not((inputs(192)) xor (inputs(10)));
    layer0_outputs(8394) <= not((inputs(205)) or (inputs(82)));
    layer0_outputs(8395) <= not(inputs(32));
    layer0_outputs(8396) <= (inputs(19)) xor (inputs(194));
    layer0_outputs(8397) <= (inputs(172)) and not (inputs(10));
    layer0_outputs(8398) <= (inputs(210)) and not (inputs(167));
    layer0_outputs(8399) <= (inputs(55)) and (inputs(39));
    layer0_outputs(8400) <= not((inputs(169)) or (inputs(64)));
    layer0_outputs(8401) <= not(inputs(22)) or (inputs(220));
    layer0_outputs(8402) <= (inputs(113)) or (inputs(6));
    layer0_outputs(8403) <= (inputs(92)) and not (inputs(24));
    layer0_outputs(8404) <= not(inputs(69));
    layer0_outputs(8405) <= not(inputs(57));
    layer0_outputs(8406) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(8407) <= not((inputs(164)) and (inputs(106)));
    layer0_outputs(8408) <= not((inputs(68)) or (inputs(195)));
    layer0_outputs(8409) <= (inputs(72)) and not (inputs(183));
    layer0_outputs(8410) <= (inputs(85)) and not (inputs(191));
    layer0_outputs(8411) <= inputs(209);
    layer0_outputs(8412) <= inputs(128);
    layer0_outputs(8413) <= inputs(197);
    layer0_outputs(8414) <= (inputs(79)) or (inputs(160));
    layer0_outputs(8415) <= (inputs(31)) xor (inputs(109));
    layer0_outputs(8416) <= not(inputs(24));
    layer0_outputs(8417) <= (inputs(255)) or (inputs(175));
    layer0_outputs(8418) <= not((inputs(79)) or (inputs(22)));
    layer0_outputs(8419) <= not(inputs(131)) or (inputs(89));
    layer0_outputs(8420) <= (inputs(144)) and not (inputs(120));
    layer0_outputs(8421) <= '1';
    layer0_outputs(8422) <= inputs(151);
    layer0_outputs(8423) <= (inputs(103)) and not (inputs(174));
    layer0_outputs(8424) <= not(inputs(136)) or (inputs(98));
    layer0_outputs(8425) <= not((inputs(242)) xor (inputs(108)));
    layer0_outputs(8426) <= not((inputs(169)) xor (inputs(231)));
    layer0_outputs(8427) <= (inputs(233)) and not (inputs(238));
    layer0_outputs(8428) <= (inputs(55)) or (inputs(121));
    layer0_outputs(8429) <= not(inputs(78)) or (inputs(118));
    layer0_outputs(8430) <= (inputs(12)) or (inputs(19));
    layer0_outputs(8431) <= not((inputs(36)) or (inputs(148)));
    layer0_outputs(8432) <= inputs(178);
    layer0_outputs(8433) <= inputs(184);
    layer0_outputs(8434) <= not(inputs(161));
    layer0_outputs(8435) <= not(inputs(218)) or (inputs(11));
    layer0_outputs(8436) <= not(inputs(186)) or (inputs(131));
    layer0_outputs(8437) <= not((inputs(86)) or (inputs(172)));
    layer0_outputs(8438) <= inputs(94);
    layer0_outputs(8439) <= (inputs(33)) xor (inputs(237));
    layer0_outputs(8440) <= inputs(31);
    layer0_outputs(8441) <= (inputs(218)) or (inputs(124));
    layer0_outputs(8442) <= (inputs(4)) or (inputs(55));
    layer0_outputs(8443) <= (inputs(67)) and not (inputs(133));
    layer0_outputs(8444) <= inputs(163);
    layer0_outputs(8445) <= inputs(45);
    layer0_outputs(8446) <= '0';
    layer0_outputs(8447) <= (inputs(113)) or (inputs(96));
    layer0_outputs(8448) <= not((inputs(177)) or (inputs(229)));
    layer0_outputs(8449) <= inputs(228);
    layer0_outputs(8450) <= not(inputs(231)) or (inputs(108));
    layer0_outputs(8451) <= not(inputs(112));
    layer0_outputs(8452) <= not(inputs(70)) or (inputs(239));
    layer0_outputs(8453) <= inputs(12);
    layer0_outputs(8454) <= (inputs(250)) or (inputs(113));
    layer0_outputs(8455) <= (inputs(163)) or (inputs(224));
    layer0_outputs(8456) <= not(inputs(130));
    layer0_outputs(8457) <= (inputs(161)) xor (inputs(49));
    layer0_outputs(8458) <= not(inputs(70)) or (inputs(221));
    layer0_outputs(8459) <= inputs(140);
    layer0_outputs(8460) <= not(inputs(213));
    layer0_outputs(8461) <= not(inputs(89));
    layer0_outputs(8462) <= not((inputs(206)) xor (inputs(69)));
    layer0_outputs(8463) <= not((inputs(154)) or (inputs(156)));
    layer0_outputs(8464) <= inputs(211);
    layer0_outputs(8465) <= not(inputs(85));
    layer0_outputs(8466) <= not(inputs(143));
    layer0_outputs(8467) <= '0';
    layer0_outputs(8468) <= not((inputs(234)) or (inputs(17)));
    layer0_outputs(8469) <= (inputs(76)) and not (inputs(191));
    layer0_outputs(8470) <= (inputs(133)) and not (inputs(95));
    layer0_outputs(8471) <= '1';
    layer0_outputs(8472) <= not((inputs(38)) or (inputs(235)));
    layer0_outputs(8473) <= not(inputs(13));
    layer0_outputs(8474) <= not(inputs(128));
    layer0_outputs(8475) <= inputs(228);
    layer0_outputs(8476) <= not((inputs(245)) and (inputs(217)));
    layer0_outputs(8477) <= not(inputs(16));
    layer0_outputs(8478) <= (inputs(204)) or (inputs(31));
    layer0_outputs(8479) <= (inputs(47)) xor (inputs(124));
    layer0_outputs(8480) <= (inputs(236)) or (inputs(92));
    layer0_outputs(8481) <= not(inputs(143)) or (inputs(1));
    layer0_outputs(8482) <= (inputs(183)) and not (inputs(113));
    layer0_outputs(8483) <= (inputs(249)) or (inputs(230));
    layer0_outputs(8484) <= (inputs(248)) and (inputs(197));
    layer0_outputs(8485) <= not(inputs(4)) or (inputs(20));
    layer0_outputs(8486) <= not((inputs(26)) or (inputs(188)));
    layer0_outputs(8487) <= (inputs(184)) and not (inputs(109));
    layer0_outputs(8488) <= inputs(170);
    layer0_outputs(8489) <= inputs(234);
    layer0_outputs(8490) <= not(inputs(190));
    layer0_outputs(8491) <= not(inputs(169));
    layer0_outputs(8492) <= not(inputs(212)) or (inputs(243));
    layer0_outputs(8493) <= (inputs(27)) and not (inputs(109));
    layer0_outputs(8494) <= not((inputs(89)) and (inputs(21)));
    layer0_outputs(8495) <= not((inputs(38)) or (inputs(211)));
    layer0_outputs(8496) <= inputs(186);
    layer0_outputs(8497) <= not(inputs(245)) or (inputs(116));
    layer0_outputs(8498) <= (inputs(216)) and not (inputs(128));
    layer0_outputs(8499) <= (inputs(168)) and not (inputs(83));
    layer0_outputs(8500) <= '1';
    layer0_outputs(8501) <= inputs(189);
    layer0_outputs(8502) <= (inputs(42)) or (inputs(64));
    layer0_outputs(8503) <= inputs(88);
    layer0_outputs(8504) <= not((inputs(232)) xor (inputs(244)));
    layer0_outputs(8505) <= (inputs(169)) and not (inputs(47));
    layer0_outputs(8506) <= not(inputs(229));
    layer0_outputs(8507) <= (inputs(89)) and not (inputs(38));
    layer0_outputs(8508) <= inputs(166);
    layer0_outputs(8509) <= inputs(96);
    layer0_outputs(8510) <= not(inputs(105));
    layer0_outputs(8511) <= not((inputs(166)) xor (inputs(104)));
    layer0_outputs(8512) <= inputs(45);
    layer0_outputs(8513) <= not(inputs(198)) or (inputs(88));
    layer0_outputs(8514) <= not(inputs(3)) or (inputs(14));
    layer0_outputs(8515) <= inputs(68);
    layer0_outputs(8516) <= not((inputs(240)) xor (inputs(194)));
    layer0_outputs(8517) <= not(inputs(210));
    layer0_outputs(8518) <= not((inputs(49)) or (inputs(187)));
    layer0_outputs(8519) <= not((inputs(153)) or (inputs(12)));
    layer0_outputs(8520) <= not(inputs(21));
    layer0_outputs(8521) <= not(inputs(140)) or (inputs(253));
    layer0_outputs(8522) <= not((inputs(155)) and (inputs(247)));
    layer0_outputs(8523) <= (inputs(117)) and not (inputs(254));
    layer0_outputs(8524) <= not(inputs(28));
    layer0_outputs(8525) <= (inputs(147)) and not (inputs(47));
    layer0_outputs(8526) <= not(inputs(227)) or (inputs(62));
    layer0_outputs(8527) <= (inputs(40)) or (inputs(181));
    layer0_outputs(8528) <= not((inputs(246)) and (inputs(217)));
    layer0_outputs(8529) <= inputs(193);
    layer0_outputs(8530) <= not(inputs(53)) or (inputs(241));
    layer0_outputs(8531) <= not((inputs(87)) or (inputs(147)));
    layer0_outputs(8532) <= inputs(234);
    layer0_outputs(8533) <= not((inputs(206)) or (inputs(42)));
    layer0_outputs(8534) <= (inputs(172)) or (inputs(146));
    layer0_outputs(8535) <= inputs(113);
    layer0_outputs(8536) <= not(inputs(0)) or (inputs(234));
    layer0_outputs(8537) <= inputs(165);
    layer0_outputs(8538) <= not(inputs(103));
    layer0_outputs(8539) <= inputs(235);
    layer0_outputs(8540) <= not((inputs(124)) or (inputs(188)));
    layer0_outputs(8541) <= (inputs(142)) or (inputs(59));
    layer0_outputs(8542) <= '1';
    layer0_outputs(8543) <= not(inputs(58));
    layer0_outputs(8544) <= (inputs(46)) and not (inputs(109));
    layer0_outputs(8545) <= not(inputs(180));
    layer0_outputs(8546) <= not((inputs(105)) or (inputs(212)));
    layer0_outputs(8547) <= not(inputs(46));
    layer0_outputs(8548) <= not((inputs(69)) xor (inputs(174)));
    layer0_outputs(8549) <= not(inputs(1));
    layer0_outputs(8550) <= inputs(43);
    layer0_outputs(8551) <= (inputs(106)) and not (inputs(152));
    layer0_outputs(8552) <= inputs(161);
    layer0_outputs(8553) <= inputs(30);
    layer0_outputs(8554) <= '1';
    layer0_outputs(8555) <= (inputs(78)) and not (inputs(131));
    layer0_outputs(8556) <= not(inputs(247));
    layer0_outputs(8557) <= (inputs(105)) or (inputs(224));
    layer0_outputs(8558) <= not(inputs(183));
    layer0_outputs(8559) <= (inputs(152)) and not (inputs(158));
    layer0_outputs(8560) <= not((inputs(167)) or (inputs(238)));
    layer0_outputs(8561) <= not(inputs(165)) or (inputs(155));
    layer0_outputs(8562) <= not(inputs(227)) or (inputs(10));
    layer0_outputs(8563) <= inputs(221);
    layer0_outputs(8564) <= not(inputs(173));
    layer0_outputs(8565) <= not(inputs(254));
    layer0_outputs(8566) <= not(inputs(239)) or (inputs(47));
    layer0_outputs(8567) <= not((inputs(215)) xor (inputs(96)));
    layer0_outputs(8568) <= not((inputs(6)) or (inputs(61)));
    layer0_outputs(8569) <= (inputs(168)) or (inputs(163));
    layer0_outputs(8570) <= (inputs(223)) and not (inputs(232));
    layer0_outputs(8571) <= inputs(83);
    layer0_outputs(8572) <= not((inputs(250)) xor (inputs(118)));
    layer0_outputs(8573) <= (inputs(188)) or (inputs(105));
    layer0_outputs(8574) <= not(inputs(195)) or (inputs(130));
    layer0_outputs(8575) <= (inputs(254)) or (inputs(159));
    layer0_outputs(8576) <= not((inputs(146)) and (inputs(72)));
    layer0_outputs(8577) <= not((inputs(140)) xor (inputs(247)));
    layer0_outputs(8578) <= inputs(77);
    layer0_outputs(8579) <= inputs(46);
    layer0_outputs(8580) <= inputs(55);
    layer0_outputs(8581) <= (inputs(170)) or (inputs(216));
    layer0_outputs(8582) <= not(inputs(99)) or (inputs(82));
    layer0_outputs(8583) <= not(inputs(244)) or (inputs(219));
    layer0_outputs(8584) <= '1';
    layer0_outputs(8585) <= not(inputs(78));
    layer0_outputs(8586) <= (inputs(151)) or (inputs(171));
    layer0_outputs(8587) <= (inputs(235)) and not (inputs(127));
    layer0_outputs(8588) <= (inputs(143)) or (inputs(180));
    layer0_outputs(8589) <= (inputs(17)) or (inputs(209));
    layer0_outputs(8590) <= not(inputs(209));
    layer0_outputs(8591) <= not(inputs(130)) or (inputs(230));
    layer0_outputs(8592) <= not(inputs(126));
    layer0_outputs(8593) <= (inputs(240)) and (inputs(185));
    layer0_outputs(8594) <= (inputs(65)) and not (inputs(12));
    layer0_outputs(8595) <= (inputs(183)) xor (inputs(122));
    layer0_outputs(8596) <= not(inputs(87));
    layer0_outputs(8597) <= inputs(74);
    layer0_outputs(8598) <= not(inputs(158)) or (inputs(187));
    layer0_outputs(8599) <= not(inputs(79));
    layer0_outputs(8600) <= not((inputs(244)) xor (inputs(248)));
    layer0_outputs(8601) <= (inputs(133)) and (inputs(84));
    layer0_outputs(8602) <= not(inputs(44)) or (inputs(144));
    layer0_outputs(8603) <= '1';
    layer0_outputs(8604) <= (inputs(61)) or (inputs(172));
    layer0_outputs(8605) <= inputs(90);
    layer0_outputs(8606) <= not((inputs(146)) or (inputs(150)));
    layer0_outputs(8607) <= (inputs(52)) and not (inputs(190));
    layer0_outputs(8608) <= (inputs(216)) xor (inputs(17));
    layer0_outputs(8609) <= not(inputs(230)) or (inputs(235));
    layer0_outputs(8610) <= not((inputs(95)) or (inputs(234)));
    layer0_outputs(8611) <= not(inputs(241));
    layer0_outputs(8612) <= inputs(150);
    layer0_outputs(8613) <= not(inputs(201)) or (inputs(71));
    layer0_outputs(8614) <= inputs(129);
    layer0_outputs(8615) <= (inputs(250)) and (inputs(10));
    layer0_outputs(8616) <= not(inputs(157));
    layer0_outputs(8617) <= not((inputs(189)) and (inputs(124)));
    layer0_outputs(8618) <= (inputs(153)) or (inputs(138));
    layer0_outputs(8619) <= not((inputs(212)) or (inputs(193)));
    layer0_outputs(8620) <= (inputs(3)) or (inputs(16));
    layer0_outputs(8621) <= not(inputs(102)) or (inputs(207));
    layer0_outputs(8622) <= (inputs(104)) and (inputs(40));
    layer0_outputs(8623) <= not(inputs(146));
    layer0_outputs(8624) <= (inputs(121)) and not (inputs(186));
    layer0_outputs(8625) <= not(inputs(208));
    layer0_outputs(8626) <= '1';
    layer0_outputs(8627) <= not(inputs(59)) or (inputs(109));
    layer0_outputs(8628) <= inputs(91);
    layer0_outputs(8629) <= '0';
    layer0_outputs(8630) <= not(inputs(222));
    layer0_outputs(8631) <= (inputs(225)) xor (inputs(174));
    layer0_outputs(8632) <= (inputs(23)) and not (inputs(191));
    layer0_outputs(8633) <= not(inputs(203));
    layer0_outputs(8634) <= (inputs(126)) or (inputs(32));
    layer0_outputs(8635) <= not(inputs(76));
    layer0_outputs(8636) <= inputs(61);
    layer0_outputs(8637) <= (inputs(91)) or (inputs(108));
    layer0_outputs(8638) <= not((inputs(218)) or (inputs(54)));
    layer0_outputs(8639) <= not(inputs(39));
    layer0_outputs(8640) <= (inputs(51)) or (inputs(17));
    layer0_outputs(8641) <= not((inputs(150)) and (inputs(181)));
    layer0_outputs(8642) <= not((inputs(181)) or (inputs(212)));
    layer0_outputs(8643) <= not(inputs(214)) or (inputs(155));
    layer0_outputs(8644) <= inputs(148);
    layer0_outputs(8645) <= not(inputs(149)) or (inputs(79));
    layer0_outputs(8646) <= (inputs(188)) xor (inputs(124));
    layer0_outputs(8647) <= (inputs(191)) or (inputs(219));
    layer0_outputs(8648) <= (inputs(99)) and not (inputs(209));
    layer0_outputs(8649) <= not(inputs(8));
    layer0_outputs(8650) <= (inputs(98)) xor (inputs(68));
    layer0_outputs(8651) <= inputs(224);
    layer0_outputs(8652) <= not(inputs(36));
    layer0_outputs(8653) <= not(inputs(123));
    layer0_outputs(8654) <= (inputs(213)) and not (inputs(116));
    layer0_outputs(8655) <= not((inputs(255)) or (inputs(133)));
    layer0_outputs(8656) <= (inputs(160)) or (inputs(202));
    layer0_outputs(8657) <= inputs(21);
    layer0_outputs(8658) <= not(inputs(29)) or (inputs(162));
    layer0_outputs(8659) <= inputs(197);
    layer0_outputs(8660) <= not(inputs(119)) or (inputs(96));
    layer0_outputs(8661) <= not((inputs(176)) or (inputs(204)));
    layer0_outputs(8662) <= (inputs(137)) and not (inputs(134));
    layer0_outputs(8663) <= inputs(166);
    layer0_outputs(8664) <= not((inputs(33)) and (inputs(182)));
    layer0_outputs(8665) <= (inputs(177)) or (inputs(10));
    layer0_outputs(8666) <= (inputs(229)) or (inputs(177));
    layer0_outputs(8667) <= not((inputs(99)) or (inputs(215)));
    layer0_outputs(8668) <= not(inputs(88)) or (inputs(250));
    layer0_outputs(8669) <= inputs(183);
    layer0_outputs(8670) <= (inputs(216)) or (inputs(111));
    layer0_outputs(8671) <= inputs(156);
    layer0_outputs(8672) <= not((inputs(210)) or (inputs(197)));
    layer0_outputs(8673) <= not(inputs(52)) or (inputs(17));
    layer0_outputs(8674) <= not((inputs(219)) and (inputs(58)));
    layer0_outputs(8675) <= (inputs(146)) and not (inputs(17));
    layer0_outputs(8676) <= not(inputs(15));
    layer0_outputs(8677) <= not((inputs(159)) or (inputs(233)));
    layer0_outputs(8678) <= (inputs(102)) and (inputs(229));
    layer0_outputs(8679) <= (inputs(55)) xor (inputs(197));
    layer0_outputs(8680) <= inputs(226);
    layer0_outputs(8681) <= not(inputs(199)) or (inputs(162));
    layer0_outputs(8682) <= (inputs(223)) and not (inputs(233));
    layer0_outputs(8683) <= not(inputs(245));
    layer0_outputs(8684) <= not((inputs(151)) or (inputs(2)));
    layer0_outputs(8685) <= not(inputs(220));
    layer0_outputs(8686) <= not((inputs(89)) or (inputs(50)));
    layer0_outputs(8687) <= (inputs(171)) or (inputs(191));
    layer0_outputs(8688) <= (inputs(12)) or (inputs(111));
    layer0_outputs(8689) <= not((inputs(80)) or (inputs(194)));
    layer0_outputs(8690) <= not(inputs(109));
    layer0_outputs(8691) <= not((inputs(234)) xor (inputs(186)));
    layer0_outputs(8692) <= not(inputs(104)) or (inputs(189));
    layer0_outputs(8693) <= not((inputs(179)) xor (inputs(0)));
    layer0_outputs(8694) <= not(inputs(88)) or (inputs(193));
    layer0_outputs(8695) <= not(inputs(209));
    layer0_outputs(8696) <= inputs(167);
    layer0_outputs(8697) <= not(inputs(85));
    layer0_outputs(8698) <= inputs(124);
    layer0_outputs(8699) <= '1';
    layer0_outputs(8700) <= inputs(183);
    layer0_outputs(8701) <= (inputs(108)) xor (inputs(63));
    layer0_outputs(8702) <= '1';
    layer0_outputs(8703) <= (inputs(6)) and not (inputs(29));
    layer0_outputs(8704) <= inputs(99);
    layer0_outputs(8705) <= not(inputs(67)) or (inputs(216));
    layer0_outputs(8706) <= not(inputs(249));
    layer0_outputs(8707) <= not(inputs(210));
    layer0_outputs(8708) <= not((inputs(4)) or (inputs(45)));
    layer0_outputs(8709) <= inputs(2);
    layer0_outputs(8710) <= inputs(190);
    layer0_outputs(8711) <= (inputs(201)) and not (inputs(47));
    layer0_outputs(8712) <= not((inputs(8)) and (inputs(192)));
    layer0_outputs(8713) <= not((inputs(16)) xor (inputs(41)));
    layer0_outputs(8714) <= (inputs(239)) or (inputs(184));
    layer0_outputs(8715) <= (inputs(18)) xor (inputs(240));
    layer0_outputs(8716) <= '0';
    layer0_outputs(8717) <= not((inputs(6)) or (inputs(163)));
    layer0_outputs(8718) <= not(inputs(76));
    layer0_outputs(8719) <= '1';
    layer0_outputs(8720) <= not((inputs(34)) or (inputs(196)));
    layer0_outputs(8721) <= inputs(85);
    layer0_outputs(8722) <= not(inputs(181));
    layer0_outputs(8723) <= not(inputs(193));
    layer0_outputs(8724) <= (inputs(39)) and not (inputs(147));
    layer0_outputs(8725) <= not(inputs(33)) or (inputs(144));
    layer0_outputs(8726) <= (inputs(151)) or (inputs(31));
    layer0_outputs(8727) <= inputs(167);
    layer0_outputs(8728) <= not(inputs(2));
    layer0_outputs(8729) <= inputs(63);
    layer0_outputs(8730) <= inputs(207);
    layer0_outputs(8731) <= inputs(92);
    layer0_outputs(8732) <= '1';
    layer0_outputs(8733) <= (inputs(69)) and not (inputs(142));
    layer0_outputs(8734) <= not((inputs(114)) or (inputs(117)));
    layer0_outputs(8735) <= '0';
    layer0_outputs(8736) <= not(inputs(19)) or (inputs(233));
    layer0_outputs(8737) <= (inputs(244)) and not (inputs(196));
    layer0_outputs(8738) <= inputs(160);
    layer0_outputs(8739) <= (inputs(250)) xor (inputs(133));
    layer0_outputs(8740) <= inputs(182);
    layer0_outputs(8741) <= not(inputs(235));
    layer0_outputs(8742) <= '1';
    layer0_outputs(8743) <= not(inputs(25));
    layer0_outputs(8744) <= '0';
    layer0_outputs(8745) <= not((inputs(118)) xor (inputs(185)));
    layer0_outputs(8746) <= (inputs(94)) or (inputs(193));
    layer0_outputs(8747) <= (inputs(168)) or (inputs(98));
    layer0_outputs(8748) <= inputs(126);
    layer0_outputs(8749) <= not((inputs(49)) or (inputs(106)));
    layer0_outputs(8750) <= not((inputs(112)) or (inputs(29)));
    layer0_outputs(8751) <= (inputs(107)) xor (inputs(64));
    layer0_outputs(8752) <= inputs(136);
    layer0_outputs(8753) <= not((inputs(189)) xor (inputs(38)));
    layer0_outputs(8754) <= (inputs(153)) or (inputs(188));
    layer0_outputs(8755) <= not(inputs(187));
    layer0_outputs(8756) <= '1';
    layer0_outputs(8757) <= (inputs(37)) xor (inputs(38));
    layer0_outputs(8758) <= (inputs(143)) and not (inputs(102));
    layer0_outputs(8759) <= not(inputs(120)) or (inputs(2));
    layer0_outputs(8760) <= not((inputs(100)) or (inputs(145)));
    layer0_outputs(8761) <= inputs(76);
    layer0_outputs(8762) <= inputs(72);
    layer0_outputs(8763) <= not(inputs(213));
    layer0_outputs(8764) <= not((inputs(8)) or (inputs(35)));
    layer0_outputs(8765) <= (inputs(41)) and (inputs(205));
    layer0_outputs(8766) <= (inputs(202)) and not (inputs(113));
    layer0_outputs(8767) <= inputs(61);
    layer0_outputs(8768) <= (inputs(159)) and not (inputs(250));
    layer0_outputs(8769) <= not((inputs(76)) and (inputs(167)));
    layer0_outputs(8770) <= (inputs(32)) and not (inputs(39));
    layer0_outputs(8771) <= not((inputs(184)) xor (inputs(182)));
    layer0_outputs(8772) <= (inputs(75)) or (inputs(166));
    layer0_outputs(8773) <= not(inputs(233));
    layer0_outputs(8774) <= (inputs(103)) and not (inputs(91));
    layer0_outputs(8775) <= (inputs(152)) and not (inputs(46));
    layer0_outputs(8776) <= (inputs(99)) or (inputs(69));
    layer0_outputs(8777) <= not(inputs(131));
    layer0_outputs(8778) <= not(inputs(106)) or (inputs(112));
    layer0_outputs(8779) <= inputs(94);
    layer0_outputs(8780) <= not(inputs(58));
    layer0_outputs(8781) <= (inputs(9)) and (inputs(60));
    layer0_outputs(8782) <= (inputs(173)) or (inputs(192));
    layer0_outputs(8783) <= not((inputs(45)) or (inputs(65)));
    layer0_outputs(8784) <= (inputs(126)) xor (inputs(13));
    layer0_outputs(8785) <= (inputs(116)) and not (inputs(243));
    layer0_outputs(8786) <= not((inputs(15)) and (inputs(124)));
    layer0_outputs(8787) <= (inputs(216)) and (inputs(159));
    layer0_outputs(8788) <= inputs(116);
    layer0_outputs(8789) <= not(inputs(35)) or (inputs(240));
    layer0_outputs(8790) <= (inputs(70)) and not (inputs(104));
    layer0_outputs(8791) <= (inputs(101)) and not (inputs(16));
    layer0_outputs(8792) <= not(inputs(29));
    layer0_outputs(8793) <= inputs(176);
    layer0_outputs(8794) <= not((inputs(97)) and (inputs(191)));
    layer0_outputs(8795) <= not(inputs(216)) or (inputs(95));
    layer0_outputs(8796) <= not(inputs(155)) or (inputs(145));
    layer0_outputs(8797) <= not(inputs(76));
    layer0_outputs(8798) <= (inputs(79)) xor (inputs(198));
    layer0_outputs(8799) <= inputs(125);
    layer0_outputs(8800) <= not((inputs(248)) or (inputs(194)));
    layer0_outputs(8801) <= not((inputs(1)) or (inputs(25)));
    layer0_outputs(8802) <= (inputs(219)) xor (inputs(233));
    layer0_outputs(8803) <= not(inputs(87)) or (inputs(12));
    layer0_outputs(8804) <= inputs(29);
    layer0_outputs(8805) <= (inputs(209)) xor (inputs(175));
    layer0_outputs(8806) <= not(inputs(212));
    layer0_outputs(8807) <= inputs(145);
    layer0_outputs(8808) <= (inputs(42)) or (inputs(73));
    layer0_outputs(8809) <= not((inputs(91)) or (inputs(131)));
    layer0_outputs(8810) <= inputs(152);
    layer0_outputs(8811) <= inputs(128);
    layer0_outputs(8812) <= inputs(86);
    layer0_outputs(8813) <= not(inputs(71)) or (inputs(254));
    layer0_outputs(8814) <= not((inputs(252)) or (inputs(218)));
    layer0_outputs(8815) <= (inputs(223)) and (inputs(160));
    layer0_outputs(8816) <= not((inputs(164)) xor (inputs(117)));
    layer0_outputs(8817) <= '0';
    layer0_outputs(8818) <= (inputs(115)) or (inputs(164));
    layer0_outputs(8819) <= not(inputs(152));
    layer0_outputs(8820) <= inputs(8);
    layer0_outputs(8821) <= (inputs(52)) or (inputs(1));
    layer0_outputs(8822) <= not((inputs(199)) xor (inputs(241)));
    layer0_outputs(8823) <= not(inputs(60));
    layer0_outputs(8824) <= not(inputs(73));
    layer0_outputs(8825) <= (inputs(132)) xor (inputs(21));
    layer0_outputs(8826) <= not(inputs(195)) or (inputs(79));
    layer0_outputs(8827) <= inputs(103);
    layer0_outputs(8828) <= not(inputs(98));
    layer0_outputs(8829) <= not(inputs(130)) or (inputs(87));
    layer0_outputs(8830) <= not((inputs(45)) or (inputs(232)));
    layer0_outputs(8831) <= not(inputs(187)) or (inputs(248));
    layer0_outputs(8832) <= not(inputs(37)) or (inputs(213));
    layer0_outputs(8833) <= (inputs(145)) xor (inputs(179));
    layer0_outputs(8834) <= not((inputs(134)) or (inputs(77)));
    layer0_outputs(8835) <= (inputs(45)) and not (inputs(107));
    layer0_outputs(8836) <= not(inputs(44));
    layer0_outputs(8837) <= not(inputs(165));
    layer0_outputs(8838) <= (inputs(45)) and not (inputs(224));
    layer0_outputs(8839) <= not((inputs(220)) xor (inputs(192)));
    layer0_outputs(8840) <= not((inputs(70)) xor (inputs(126)));
    layer0_outputs(8841) <= not(inputs(152)) or (inputs(47));
    layer0_outputs(8842) <= (inputs(230)) xor (inputs(105));
    layer0_outputs(8843) <= not(inputs(164)) or (inputs(94));
    layer0_outputs(8844) <= '1';
    layer0_outputs(8845) <= not((inputs(33)) or (inputs(149)));
    layer0_outputs(8846) <= (inputs(99)) or (inputs(82));
    layer0_outputs(8847) <= inputs(20);
    layer0_outputs(8848) <= (inputs(146)) or (inputs(96));
    layer0_outputs(8849) <= inputs(150);
    layer0_outputs(8850) <= not(inputs(151)) or (inputs(55));
    layer0_outputs(8851) <= not(inputs(73));
    layer0_outputs(8852) <= not((inputs(47)) xor (inputs(67)));
    layer0_outputs(8853) <= not(inputs(230));
    layer0_outputs(8854) <= not(inputs(214)) or (inputs(15));
    layer0_outputs(8855) <= '1';
    layer0_outputs(8856) <= not((inputs(109)) or (inputs(41)));
    layer0_outputs(8857) <= (inputs(141)) or (inputs(155));
    layer0_outputs(8858) <= (inputs(56)) and not (inputs(30));
    layer0_outputs(8859) <= not((inputs(205)) and (inputs(253)));
    layer0_outputs(8860) <= (inputs(144)) or (inputs(179));
    layer0_outputs(8861) <= not(inputs(118)) or (inputs(38));
    layer0_outputs(8862) <= not(inputs(201)) or (inputs(228));
    layer0_outputs(8863) <= not(inputs(195)) or (inputs(94));
    layer0_outputs(8864) <= (inputs(247)) and not (inputs(62));
    layer0_outputs(8865) <= not(inputs(182));
    layer0_outputs(8866) <= (inputs(139)) xor (inputs(203));
    layer0_outputs(8867) <= inputs(27);
    layer0_outputs(8868) <= not(inputs(123)) or (inputs(129));
    layer0_outputs(8869) <= (inputs(246)) and not (inputs(148));
    layer0_outputs(8870) <= inputs(43);
    layer0_outputs(8871) <= (inputs(200)) and not (inputs(203));
    layer0_outputs(8872) <= (inputs(57)) and not (inputs(206));
    layer0_outputs(8873) <= inputs(146);
    layer0_outputs(8874) <= inputs(146);
    layer0_outputs(8875) <= (inputs(0)) and (inputs(32));
    layer0_outputs(8876) <= (inputs(201)) or (inputs(173));
    layer0_outputs(8877) <= not(inputs(130));
    layer0_outputs(8878) <= not(inputs(211));
    layer0_outputs(8879) <= inputs(229);
    layer0_outputs(8880) <= (inputs(34)) and not (inputs(63));
    layer0_outputs(8881) <= (inputs(156)) or (inputs(141));
    layer0_outputs(8882) <= (inputs(12)) or (inputs(141));
    layer0_outputs(8883) <= not(inputs(31));
    layer0_outputs(8884) <= inputs(92);
    layer0_outputs(8885) <= not(inputs(114));
    layer0_outputs(8886) <= not((inputs(239)) or (inputs(28)));
    layer0_outputs(8887) <= '1';
    layer0_outputs(8888) <= not(inputs(94));
    layer0_outputs(8889) <= not((inputs(54)) or (inputs(96)));
    layer0_outputs(8890) <= not((inputs(212)) and (inputs(246)));
    layer0_outputs(8891) <= not((inputs(189)) xor (inputs(221)));
    layer0_outputs(8892) <= not(inputs(94)) or (inputs(121));
    layer0_outputs(8893) <= not(inputs(74));
    layer0_outputs(8894) <= not(inputs(117)) or (inputs(175));
    layer0_outputs(8895) <= not((inputs(19)) or (inputs(68)));
    layer0_outputs(8896) <= (inputs(127)) or (inputs(232));
    layer0_outputs(8897) <= not((inputs(179)) or (inputs(210)));
    layer0_outputs(8898) <= not(inputs(196)) or (inputs(140));
    layer0_outputs(8899) <= not(inputs(111)) or (inputs(7));
    layer0_outputs(8900) <= not(inputs(233));
    layer0_outputs(8901) <= not(inputs(27));
    layer0_outputs(8902) <= not((inputs(177)) or (inputs(60)));
    layer0_outputs(8903) <= not((inputs(179)) xor (inputs(52)));
    layer0_outputs(8904) <= not(inputs(5)) or (inputs(37));
    layer0_outputs(8905) <= not(inputs(117)) or (inputs(171));
    layer0_outputs(8906) <= inputs(34);
    layer0_outputs(8907) <= (inputs(7)) or (inputs(139));
    layer0_outputs(8908) <= (inputs(57)) and not (inputs(82));
    layer0_outputs(8909) <= not(inputs(25));
    layer0_outputs(8910) <= not(inputs(189));
    layer0_outputs(8911) <= (inputs(192)) or (inputs(214));
    layer0_outputs(8912) <= inputs(120);
    layer0_outputs(8913) <= not(inputs(198)) or (inputs(191));
    layer0_outputs(8914) <= (inputs(75)) and not (inputs(192));
    layer0_outputs(8915) <= (inputs(128)) and not (inputs(10));
    layer0_outputs(8916) <= not(inputs(226));
    layer0_outputs(8917) <= (inputs(178)) xor (inputs(160));
    layer0_outputs(8918) <= '0';
    layer0_outputs(8919) <= not((inputs(163)) xor (inputs(69)));
    layer0_outputs(8920) <= not((inputs(240)) or (inputs(18)));
    layer0_outputs(8921) <= not(inputs(233)) or (inputs(50));
    layer0_outputs(8922) <= '1';
    layer0_outputs(8923) <= not((inputs(0)) and (inputs(16)));
    layer0_outputs(8924) <= '1';
    layer0_outputs(8925) <= not(inputs(152));
    layer0_outputs(8926) <= not(inputs(211));
    layer0_outputs(8927) <= (inputs(184)) and not (inputs(31));
    layer0_outputs(8928) <= (inputs(98)) or (inputs(60));
    layer0_outputs(8929) <= (inputs(144)) or (inputs(32));
    layer0_outputs(8930) <= not((inputs(66)) and (inputs(140)));
    layer0_outputs(8931) <= (inputs(22)) xor (inputs(67));
    layer0_outputs(8932) <= inputs(69);
    layer0_outputs(8933) <= not((inputs(39)) and (inputs(171)));
    layer0_outputs(8934) <= not((inputs(159)) or (inputs(3)));
    layer0_outputs(8935) <= (inputs(88)) xor (inputs(139));
    layer0_outputs(8936) <= (inputs(245)) and not (inputs(148));
    layer0_outputs(8937) <= '1';
    layer0_outputs(8938) <= inputs(19);
    layer0_outputs(8939) <= not(inputs(39));
    layer0_outputs(8940) <= inputs(249);
    layer0_outputs(8941) <= (inputs(143)) and not (inputs(39));
    layer0_outputs(8942) <= inputs(97);
    layer0_outputs(8943) <= not((inputs(138)) and (inputs(202)));
    layer0_outputs(8944) <= not(inputs(173));
    layer0_outputs(8945) <= not(inputs(108)) or (inputs(228));
    layer0_outputs(8946) <= (inputs(233)) and (inputs(90));
    layer0_outputs(8947) <= (inputs(137)) and not (inputs(171));
    layer0_outputs(8948) <= not(inputs(22));
    layer0_outputs(8949) <= not((inputs(154)) and (inputs(101)));
    layer0_outputs(8950) <= inputs(140);
    layer0_outputs(8951) <= not(inputs(228));
    layer0_outputs(8952) <= not(inputs(229)) or (inputs(114));
    layer0_outputs(8953) <= not((inputs(178)) or (inputs(84)));
    layer0_outputs(8954) <= '0';
    layer0_outputs(8955) <= not(inputs(183)) or (inputs(239));
    layer0_outputs(8956) <= (inputs(180)) and (inputs(246));
    layer0_outputs(8957) <= not((inputs(241)) xor (inputs(224)));
    layer0_outputs(8958) <= not(inputs(104));
    layer0_outputs(8959) <= (inputs(193)) or (inputs(48));
    layer0_outputs(8960) <= not((inputs(1)) xor (inputs(110)));
    layer0_outputs(8961) <= not(inputs(230));
    layer0_outputs(8962) <= '0';
    layer0_outputs(8963) <= (inputs(125)) or (inputs(2));
    layer0_outputs(8964) <= (inputs(87)) xor (inputs(128));
    layer0_outputs(8965) <= (inputs(93)) or (inputs(58));
    layer0_outputs(8966) <= not(inputs(255)) or (inputs(152));
    layer0_outputs(8967) <= (inputs(212)) and not (inputs(3));
    layer0_outputs(8968) <= (inputs(94)) or (inputs(6));
    layer0_outputs(8969) <= (inputs(22)) or (inputs(9));
    layer0_outputs(8970) <= not((inputs(57)) xor (inputs(102)));
    layer0_outputs(8971) <= not(inputs(161)) or (inputs(247));
    layer0_outputs(8972) <= (inputs(160)) and not (inputs(82));
    layer0_outputs(8973) <= not(inputs(57));
    layer0_outputs(8974) <= not(inputs(164));
    layer0_outputs(8975) <= inputs(164);
    layer0_outputs(8976) <= inputs(75);
    layer0_outputs(8977) <= not((inputs(155)) or (inputs(188)));
    layer0_outputs(8978) <= inputs(25);
    layer0_outputs(8979) <= (inputs(122)) and not (inputs(209));
    layer0_outputs(8980) <= not((inputs(238)) xor (inputs(100)));
    layer0_outputs(8981) <= not(inputs(21));
    layer0_outputs(8982) <= not(inputs(0)) or (inputs(80));
    layer0_outputs(8983) <= (inputs(34)) and not (inputs(132));
    layer0_outputs(8984) <= (inputs(5)) and not (inputs(38));
    layer0_outputs(8985) <= (inputs(195)) and not (inputs(13));
    layer0_outputs(8986) <= (inputs(51)) or (inputs(153));
    layer0_outputs(8987) <= '0';
    layer0_outputs(8988) <= not((inputs(66)) or (inputs(101)));
    layer0_outputs(8989) <= not(inputs(163));
    layer0_outputs(8990) <= not((inputs(227)) or (inputs(150)));
    layer0_outputs(8991) <= (inputs(76)) and (inputs(181));
    layer0_outputs(8992) <= not(inputs(116));
    layer0_outputs(8993) <= not(inputs(90));
    layer0_outputs(8994) <= not(inputs(187));
    layer0_outputs(8995) <= not((inputs(192)) or (inputs(196)));
    layer0_outputs(8996) <= not((inputs(225)) xor (inputs(148)));
    layer0_outputs(8997) <= not(inputs(37)) or (inputs(39));
    layer0_outputs(8998) <= not(inputs(239)) or (inputs(39));
    layer0_outputs(8999) <= (inputs(221)) xor (inputs(72));
    layer0_outputs(9000) <= not(inputs(45));
    layer0_outputs(9001) <= not(inputs(90));
    layer0_outputs(9002) <= (inputs(70)) xor (inputs(83));
    layer0_outputs(9003) <= not(inputs(21));
    layer0_outputs(9004) <= not((inputs(22)) or (inputs(8)));
    layer0_outputs(9005) <= not(inputs(255));
    layer0_outputs(9006) <= inputs(164);
    layer0_outputs(9007) <= (inputs(20)) and not (inputs(113));
    layer0_outputs(9008) <= not((inputs(227)) or (inputs(81)));
    layer0_outputs(9009) <= inputs(220);
    layer0_outputs(9010) <= (inputs(37)) and not (inputs(164));
    layer0_outputs(9011) <= not(inputs(218)) or (inputs(48));
    layer0_outputs(9012) <= not((inputs(154)) and (inputs(221)));
    layer0_outputs(9013) <= not(inputs(2)) or (inputs(112));
    layer0_outputs(9014) <= not(inputs(203));
    layer0_outputs(9015) <= not(inputs(184));
    layer0_outputs(9016) <= not((inputs(126)) or (inputs(57)));
    layer0_outputs(9017) <= not((inputs(98)) xor (inputs(132)));
    layer0_outputs(9018) <= not(inputs(148)) or (inputs(30));
    layer0_outputs(9019) <= inputs(114);
    layer0_outputs(9020) <= (inputs(141)) and not (inputs(35));
    layer0_outputs(9021) <= inputs(238);
    layer0_outputs(9022) <= not((inputs(83)) or (inputs(252)));
    layer0_outputs(9023) <= not((inputs(167)) or (inputs(36)));
    layer0_outputs(9024) <= (inputs(55)) or (inputs(17));
    layer0_outputs(9025) <= (inputs(172)) or (inputs(171));
    layer0_outputs(9026) <= inputs(147);
    layer0_outputs(9027) <= not(inputs(37)) or (inputs(130));
    layer0_outputs(9028) <= (inputs(108)) and not (inputs(250));
    layer0_outputs(9029) <= (inputs(20)) and not (inputs(223));
    layer0_outputs(9030) <= not((inputs(118)) xor (inputs(149)));
    layer0_outputs(9031) <= not(inputs(185)) or (inputs(224));
    layer0_outputs(9032) <= (inputs(233)) and not (inputs(226));
    layer0_outputs(9033) <= inputs(125);
    layer0_outputs(9034) <= inputs(3);
    layer0_outputs(9035) <= (inputs(180)) and (inputs(232));
    layer0_outputs(9036) <= not(inputs(148));
    layer0_outputs(9037) <= not(inputs(129));
    layer0_outputs(9038) <= (inputs(14)) xor (inputs(103));
    layer0_outputs(9039) <= inputs(229);
    layer0_outputs(9040) <= inputs(154);
    layer0_outputs(9041) <= (inputs(31)) and not (inputs(154));
    layer0_outputs(9042) <= (inputs(0)) or (inputs(144));
    layer0_outputs(9043) <= not(inputs(19));
    layer0_outputs(9044) <= (inputs(138)) xor (inputs(63));
    layer0_outputs(9045) <= not((inputs(220)) or (inputs(199)));
    layer0_outputs(9046) <= inputs(159);
    layer0_outputs(9047) <= (inputs(107)) or (inputs(162));
    layer0_outputs(9048) <= not(inputs(159)) or (inputs(17));
    layer0_outputs(9049) <= not(inputs(99));
    layer0_outputs(9050) <= '0';
    layer0_outputs(9051) <= not(inputs(248)) or (inputs(14));
    layer0_outputs(9052) <= (inputs(211)) and (inputs(188));
    layer0_outputs(9053) <= (inputs(106)) and not (inputs(255));
    layer0_outputs(9054) <= (inputs(141)) and not (inputs(122));
    layer0_outputs(9055) <= inputs(108);
    layer0_outputs(9056) <= (inputs(118)) or (inputs(173));
    layer0_outputs(9057) <= not((inputs(126)) or (inputs(191)));
    layer0_outputs(9058) <= (inputs(121)) and (inputs(21));
    layer0_outputs(9059) <= (inputs(228)) and not (inputs(48));
    layer0_outputs(9060) <= not((inputs(177)) xor (inputs(216)));
    layer0_outputs(9061) <= not((inputs(75)) and (inputs(29)));
    layer0_outputs(9062) <= not(inputs(166));
    layer0_outputs(9063) <= not((inputs(142)) or (inputs(86)));
    layer0_outputs(9064) <= inputs(109);
    layer0_outputs(9065) <= (inputs(105)) and not (inputs(1));
    layer0_outputs(9066) <= (inputs(2)) and not (inputs(96));
    layer0_outputs(9067) <= not(inputs(142)) or (inputs(208));
    layer0_outputs(9068) <= (inputs(237)) and not (inputs(154));
    layer0_outputs(9069) <= not(inputs(228));
    layer0_outputs(9070) <= not(inputs(186));
    layer0_outputs(9071) <= not(inputs(80)) or (inputs(232));
    layer0_outputs(9072) <= not((inputs(6)) or (inputs(205)));
    layer0_outputs(9073) <= (inputs(204)) or (inputs(201));
    layer0_outputs(9074) <= inputs(118);
    layer0_outputs(9075) <= not((inputs(203)) xor (inputs(30)));
    layer0_outputs(9076) <= (inputs(119)) or (inputs(14));
    layer0_outputs(9077) <= not(inputs(103)) or (inputs(1));
    layer0_outputs(9078) <= not(inputs(4));
    layer0_outputs(9079) <= not(inputs(167));
    layer0_outputs(9080) <= not(inputs(144));
    layer0_outputs(9081) <= not(inputs(234));
    layer0_outputs(9082) <= not(inputs(114));
    layer0_outputs(9083) <= (inputs(177)) xor (inputs(227));
    layer0_outputs(9084) <= (inputs(233)) and not (inputs(44));
    layer0_outputs(9085) <= not(inputs(152));
    layer0_outputs(9086) <= not((inputs(54)) or (inputs(178)));
    layer0_outputs(9087) <= (inputs(80)) and (inputs(189));
    layer0_outputs(9088) <= (inputs(75)) or (inputs(35));
    layer0_outputs(9089) <= not(inputs(61));
    layer0_outputs(9090) <= not((inputs(220)) and (inputs(78)));
    layer0_outputs(9091) <= (inputs(168)) xor (inputs(36));
    layer0_outputs(9092) <= not((inputs(67)) xor (inputs(21)));
    layer0_outputs(9093) <= (inputs(2)) and not (inputs(244));
    layer0_outputs(9094) <= not(inputs(211));
    layer0_outputs(9095) <= not(inputs(114));
    layer0_outputs(9096) <= inputs(20);
    layer0_outputs(9097) <= (inputs(37)) and not (inputs(128));
    layer0_outputs(9098) <= inputs(239);
    layer0_outputs(9099) <= (inputs(90)) and not (inputs(247));
    layer0_outputs(9100) <= (inputs(81)) and not (inputs(162));
    layer0_outputs(9101) <= not(inputs(154));
    layer0_outputs(9102) <= (inputs(217)) and not (inputs(109));
    layer0_outputs(9103) <= inputs(108);
    layer0_outputs(9104) <= (inputs(55)) or (inputs(112));
    layer0_outputs(9105) <= not(inputs(203));
    layer0_outputs(9106) <= not(inputs(245));
    layer0_outputs(9107) <= not(inputs(177));
    layer0_outputs(9108) <= '1';
    layer0_outputs(9109) <= not(inputs(107)) or (inputs(253));
    layer0_outputs(9110) <= '1';
    layer0_outputs(9111) <= (inputs(235)) xor (inputs(64));
    layer0_outputs(9112) <= not(inputs(95));
    layer0_outputs(9113) <= (inputs(77)) and (inputs(70));
    layer0_outputs(9114) <= '1';
    layer0_outputs(9115) <= (inputs(188)) or (inputs(146));
    layer0_outputs(9116) <= (inputs(246)) and (inputs(170));
    layer0_outputs(9117) <= not((inputs(61)) or (inputs(177)));
    layer0_outputs(9118) <= (inputs(179)) xor (inputs(165));
    layer0_outputs(9119) <= inputs(218);
    layer0_outputs(9120) <= not((inputs(96)) xor (inputs(85)));
    layer0_outputs(9121) <= not(inputs(231)) or (inputs(89));
    layer0_outputs(9122) <= (inputs(165)) or (inputs(101));
    layer0_outputs(9123) <= inputs(88);
    layer0_outputs(9124) <= (inputs(188)) or (inputs(103));
    layer0_outputs(9125) <= not((inputs(127)) or (inputs(69)));
    layer0_outputs(9126) <= not(inputs(68)) or (inputs(223));
    layer0_outputs(9127) <= inputs(127);
    layer0_outputs(9128) <= inputs(199);
    layer0_outputs(9129) <= not(inputs(215));
    layer0_outputs(9130) <= not(inputs(197)) or (inputs(67));
    layer0_outputs(9131) <= (inputs(0)) xor (inputs(151));
    layer0_outputs(9132) <= not((inputs(228)) or (inputs(108)));
    layer0_outputs(9133) <= inputs(107);
    layer0_outputs(9134) <= (inputs(50)) xor (inputs(81));
    layer0_outputs(9135) <= not(inputs(82));
    layer0_outputs(9136) <= (inputs(111)) or (inputs(223));
    layer0_outputs(9137) <= not((inputs(153)) or (inputs(238)));
    layer0_outputs(9138) <= not(inputs(95));
    layer0_outputs(9139) <= (inputs(167)) and not (inputs(45));
    layer0_outputs(9140) <= (inputs(204)) or (inputs(197));
    layer0_outputs(9141) <= (inputs(250)) or (inputs(28));
    layer0_outputs(9142) <= not(inputs(3));
    layer0_outputs(9143) <= not(inputs(51));
    layer0_outputs(9144) <= not(inputs(149));
    layer0_outputs(9145) <= (inputs(6)) and (inputs(222));
    layer0_outputs(9146) <= (inputs(11)) or (inputs(97));
    layer0_outputs(9147) <= (inputs(215)) and not (inputs(51));
    layer0_outputs(9148) <= (inputs(79)) or (inputs(180));
    layer0_outputs(9149) <= not(inputs(140));
    layer0_outputs(9150) <= not(inputs(115));
    layer0_outputs(9151) <= not((inputs(52)) xor (inputs(143)));
    layer0_outputs(9152) <= not((inputs(133)) or (inputs(82)));
    layer0_outputs(9153) <= (inputs(116)) or (inputs(183));
    layer0_outputs(9154) <= inputs(160);
    layer0_outputs(9155) <= not(inputs(99)) or (inputs(18));
    layer0_outputs(9156) <= not(inputs(120)) or (inputs(96));
    layer0_outputs(9157) <= '1';
    layer0_outputs(9158) <= inputs(243);
    layer0_outputs(9159) <= inputs(42);
    layer0_outputs(9160) <= not(inputs(92));
    layer0_outputs(9161) <= not(inputs(31)) or (inputs(91));
    layer0_outputs(9162) <= (inputs(52)) or (inputs(78));
    layer0_outputs(9163) <= not(inputs(121));
    layer0_outputs(9164) <= not((inputs(76)) and (inputs(66)));
    layer0_outputs(9165) <= inputs(183);
    layer0_outputs(9166) <= (inputs(202)) and not (inputs(6));
    layer0_outputs(9167) <= not(inputs(157)) or (inputs(188));
    layer0_outputs(9168) <= not(inputs(167));
    layer0_outputs(9169) <= not(inputs(170));
    layer0_outputs(9170) <= (inputs(15)) and not (inputs(156));
    layer0_outputs(9171) <= inputs(129);
    layer0_outputs(9172) <= (inputs(167)) and not (inputs(159));
    layer0_outputs(9173) <= not(inputs(63));
    layer0_outputs(9174) <= '1';
    layer0_outputs(9175) <= not(inputs(180)) or (inputs(46));
    layer0_outputs(9176) <= not(inputs(66));
    layer0_outputs(9177) <= not((inputs(165)) or (inputs(130)));
    layer0_outputs(9178) <= not(inputs(186));
    layer0_outputs(9179) <= '1';
    layer0_outputs(9180) <= not(inputs(168));
    layer0_outputs(9181) <= (inputs(115)) and not (inputs(122));
    layer0_outputs(9182) <= not((inputs(107)) or (inputs(16)));
    layer0_outputs(9183) <= not(inputs(117));
    layer0_outputs(9184) <= not((inputs(79)) and (inputs(191)));
    layer0_outputs(9185) <= (inputs(115)) or (inputs(21));
    layer0_outputs(9186) <= not(inputs(24)) or (inputs(216));
    layer0_outputs(9187) <= (inputs(157)) and not (inputs(49));
    layer0_outputs(9188) <= not(inputs(23));
    layer0_outputs(9189) <= (inputs(1)) and (inputs(254));
    layer0_outputs(9190) <= '0';
    layer0_outputs(9191) <= not((inputs(139)) and (inputs(189)));
    layer0_outputs(9192) <= (inputs(213)) and not (inputs(121));
    layer0_outputs(9193) <= (inputs(2)) or (inputs(194));
    layer0_outputs(9194) <= not(inputs(241));
    layer0_outputs(9195) <= not((inputs(136)) and (inputs(15)));
    layer0_outputs(9196) <= (inputs(182)) and not (inputs(76));
    layer0_outputs(9197) <= (inputs(255)) and not (inputs(18));
    layer0_outputs(9198) <= inputs(19);
    layer0_outputs(9199) <= not((inputs(66)) xor (inputs(5)));
    layer0_outputs(9200) <= not(inputs(252));
    layer0_outputs(9201) <= (inputs(218)) or (inputs(222));
    layer0_outputs(9202) <= (inputs(86)) and (inputs(6));
    layer0_outputs(9203) <= (inputs(236)) and not (inputs(176));
    layer0_outputs(9204) <= not(inputs(101)) or (inputs(18));
    layer0_outputs(9205) <= inputs(67);
    layer0_outputs(9206) <= not((inputs(144)) xor (inputs(103)));
    layer0_outputs(9207) <= not(inputs(6));
    layer0_outputs(9208) <= inputs(168);
    layer0_outputs(9209) <= (inputs(240)) or (inputs(204));
    layer0_outputs(9210) <= inputs(149);
    layer0_outputs(9211) <= inputs(140);
    layer0_outputs(9212) <= (inputs(9)) or (inputs(127));
    layer0_outputs(9213) <= inputs(40);
    layer0_outputs(9214) <= not((inputs(240)) xor (inputs(247)));
    layer0_outputs(9215) <= (inputs(89)) xor (inputs(157));
    layer0_outputs(9216) <= not((inputs(193)) xor (inputs(235)));
    layer0_outputs(9217) <= (inputs(244)) and not (inputs(127));
    layer0_outputs(9218) <= (inputs(61)) and not (inputs(190));
    layer0_outputs(9219) <= (inputs(76)) or (inputs(162));
    layer0_outputs(9220) <= not(inputs(252)) or (inputs(64));
    layer0_outputs(9221) <= inputs(123);
    layer0_outputs(9222) <= '0';
    layer0_outputs(9223) <= '1';
    layer0_outputs(9224) <= not(inputs(132)) or (inputs(238));
    layer0_outputs(9225) <= (inputs(0)) or (inputs(73));
    layer0_outputs(9226) <= not((inputs(29)) xor (inputs(62)));
    layer0_outputs(9227) <= (inputs(1)) or (inputs(12));
    layer0_outputs(9228) <= not(inputs(153));
    layer0_outputs(9229) <= not(inputs(140)) or (inputs(253));
    layer0_outputs(9230) <= (inputs(148)) and not (inputs(246));
    layer0_outputs(9231) <= (inputs(50)) or (inputs(151));
    layer0_outputs(9232) <= not((inputs(110)) or (inputs(25)));
    layer0_outputs(9233) <= not(inputs(155)) or (inputs(75));
    layer0_outputs(9234) <= inputs(47);
    layer0_outputs(9235) <= inputs(33);
    layer0_outputs(9236) <= not(inputs(88)) or (inputs(27));
    layer0_outputs(9237) <= (inputs(77)) or (inputs(110));
    layer0_outputs(9238) <= (inputs(99)) or (inputs(23));
    layer0_outputs(9239) <= not((inputs(237)) or (inputs(226)));
    layer0_outputs(9240) <= (inputs(86)) xor (inputs(127));
    layer0_outputs(9241) <= (inputs(129)) xor (inputs(116));
    layer0_outputs(9242) <= not((inputs(177)) or (inputs(217)));
    layer0_outputs(9243) <= not((inputs(205)) xor (inputs(162)));
    layer0_outputs(9244) <= not((inputs(64)) xor (inputs(133)));
    layer0_outputs(9245) <= (inputs(86)) and not (inputs(48));
    layer0_outputs(9246) <= not((inputs(32)) or (inputs(226)));
    layer0_outputs(9247) <= inputs(190);
    layer0_outputs(9248) <= (inputs(196)) and not (inputs(174));
    layer0_outputs(9249) <= not(inputs(142));
    layer0_outputs(9250) <= inputs(104);
    layer0_outputs(9251) <= not(inputs(187)) or (inputs(59));
    layer0_outputs(9252) <= not(inputs(143)) or (inputs(225));
    layer0_outputs(9253) <= not((inputs(10)) or (inputs(50)));
    layer0_outputs(9254) <= '0';
    layer0_outputs(9255) <= '0';
    layer0_outputs(9256) <= inputs(169);
    layer0_outputs(9257) <= (inputs(233)) or (inputs(142));
    layer0_outputs(9258) <= not(inputs(145));
    layer0_outputs(9259) <= inputs(8);
    layer0_outputs(9260) <= inputs(161);
    layer0_outputs(9261) <= not(inputs(38)) or (inputs(176));
    layer0_outputs(9262) <= inputs(146);
    layer0_outputs(9263) <= not(inputs(204));
    layer0_outputs(9264) <= inputs(122);
    layer0_outputs(9265) <= not((inputs(210)) or (inputs(180)));
    layer0_outputs(9266) <= (inputs(134)) and (inputs(67));
    layer0_outputs(9267) <= not(inputs(13)) or (inputs(206));
    layer0_outputs(9268) <= not(inputs(130));
    layer0_outputs(9269) <= not((inputs(179)) xor (inputs(95)));
    layer0_outputs(9270) <= not((inputs(126)) xor (inputs(156)));
    layer0_outputs(9271) <= not((inputs(201)) xor (inputs(185)));
    layer0_outputs(9272) <= (inputs(114)) or (inputs(14));
    layer0_outputs(9273) <= not(inputs(226));
    layer0_outputs(9274) <= not(inputs(8)) or (inputs(159));
    layer0_outputs(9275) <= not(inputs(248));
    layer0_outputs(9276) <= '1';
    layer0_outputs(9277) <= (inputs(127)) and not (inputs(209));
    layer0_outputs(9278) <= not(inputs(64)) or (inputs(102));
    layer0_outputs(9279) <= not(inputs(19));
    layer0_outputs(9280) <= (inputs(224)) xor (inputs(157));
    layer0_outputs(9281) <= inputs(220);
    layer0_outputs(9282) <= (inputs(22)) and not (inputs(183));
    layer0_outputs(9283) <= (inputs(196)) or (inputs(98));
    layer0_outputs(9284) <= (inputs(55)) and not (inputs(255));
    layer0_outputs(9285) <= inputs(103);
    layer0_outputs(9286) <= inputs(23);
    layer0_outputs(9287) <= (inputs(84)) and not (inputs(248));
    layer0_outputs(9288) <= (inputs(172)) or (inputs(188));
    layer0_outputs(9289) <= inputs(201);
    layer0_outputs(9290) <= (inputs(151)) and not (inputs(215));
    layer0_outputs(9291) <= not((inputs(159)) or (inputs(120)));
    layer0_outputs(9292) <= inputs(3);
    layer0_outputs(9293) <= not((inputs(107)) xor (inputs(181)));
    layer0_outputs(9294) <= inputs(43);
    layer0_outputs(9295) <= (inputs(228)) and not (inputs(179));
    layer0_outputs(9296) <= inputs(152);
    layer0_outputs(9297) <= (inputs(219)) or (inputs(223));
    layer0_outputs(9298) <= (inputs(231)) or (inputs(27));
    layer0_outputs(9299) <= not((inputs(230)) or (inputs(206)));
    layer0_outputs(9300) <= not((inputs(34)) or (inputs(122)));
    layer0_outputs(9301) <= inputs(242);
    layer0_outputs(9302) <= not(inputs(55)) or (inputs(46));
    layer0_outputs(9303) <= not((inputs(90)) xor (inputs(190)));
    layer0_outputs(9304) <= not(inputs(1));
    layer0_outputs(9305) <= not(inputs(186)) or (inputs(109));
    layer0_outputs(9306) <= not((inputs(12)) xor (inputs(46)));
    layer0_outputs(9307) <= not(inputs(219)) or (inputs(44));
    layer0_outputs(9308) <= (inputs(47)) and not (inputs(253));
    layer0_outputs(9309) <= (inputs(246)) and not (inputs(233));
    layer0_outputs(9310) <= not(inputs(216)) or (inputs(165));
    layer0_outputs(9311) <= (inputs(176)) or (inputs(189));
    layer0_outputs(9312) <= not(inputs(136)) or (inputs(14));
    layer0_outputs(9313) <= not((inputs(123)) xor (inputs(130)));
    layer0_outputs(9314) <= not(inputs(101)) or (inputs(123));
    layer0_outputs(9315) <= (inputs(20)) and not (inputs(252));
    layer0_outputs(9316) <= (inputs(177)) and not (inputs(223));
    layer0_outputs(9317) <= (inputs(229)) and not (inputs(220));
    layer0_outputs(9318) <= (inputs(57)) and (inputs(231));
    layer0_outputs(9319) <= not((inputs(206)) or (inputs(28)));
    layer0_outputs(9320) <= (inputs(38)) and not (inputs(252));
    layer0_outputs(9321) <= (inputs(232)) and (inputs(67));
    layer0_outputs(9322) <= not((inputs(203)) or (inputs(58)));
    layer0_outputs(9323) <= (inputs(30)) and (inputs(18));
    layer0_outputs(9324) <= not(inputs(100));
    layer0_outputs(9325) <= (inputs(60)) xor (inputs(231));
    layer0_outputs(9326) <= (inputs(13)) xor (inputs(74));
    layer0_outputs(9327) <= not(inputs(49));
    layer0_outputs(9328) <= not((inputs(115)) xor (inputs(227)));
    layer0_outputs(9329) <= (inputs(195)) or (inputs(129));
    layer0_outputs(9330) <= inputs(140);
    layer0_outputs(9331) <= not(inputs(19)) or (inputs(241));
    layer0_outputs(9332) <= (inputs(99)) or (inputs(248));
    layer0_outputs(9333) <= (inputs(62)) and not (inputs(109));
    layer0_outputs(9334) <= inputs(165);
    layer0_outputs(9335) <= '1';
    layer0_outputs(9336) <= (inputs(227)) and not (inputs(98));
    layer0_outputs(9337) <= inputs(4);
    layer0_outputs(9338) <= not((inputs(16)) and (inputs(115)));
    layer0_outputs(9339) <= '1';
    layer0_outputs(9340) <= (inputs(154)) or (inputs(85));
    layer0_outputs(9341) <= inputs(165);
    layer0_outputs(9342) <= not(inputs(197));
    layer0_outputs(9343) <= not((inputs(120)) xor (inputs(163)));
    layer0_outputs(9344) <= (inputs(126)) or (inputs(101));
    layer0_outputs(9345) <= (inputs(54)) and (inputs(161));
    layer0_outputs(9346) <= not((inputs(147)) or (inputs(93)));
    layer0_outputs(9347) <= inputs(138);
    layer0_outputs(9348) <= inputs(241);
    layer0_outputs(9349) <= inputs(101);
    layer0_outputs(9350) <= (inputs(218)) and (inputs(234));
    layer0_outputs(9351) <= not((inputs(44)) or (inputs(47)));
    layer0_outputs(9352) <= not(inputs(23));
    layer0_outputs(9353) <= (inputs(77)) xor (inputs(13));
    layer0_outputs(9354) <= inputs(163);
    layer0_outputs(9355) <= not((inputs(61)) or (inputs(209)));
    layer0_outputs(9356) <= (inputs(238)) and not (inputs(50));
    layer0_outputs(9357) <= not(inputs(14)) or (inputs(59));
    layer0_outputs(9358) <= inputs(200);
    layer0_outputs(9359) <= '0';
    layer0_outputs(9360) <= not(inputs(8)) or (inputs(159));
    layer0_outputs(9361) <= not(inputs(196));
    layer0_outputs(9362) <= inputs(21);
    layer0_outputs(9363) <= not((inputs(94)) xor (inputs(123)));
    layer0_outputs(9364) <= inputs(39);
    layer0_outputs(9365) <= not(inputs(123));
    layer0_outputs(9366) <= not(inputs(161)) or (inputs(160));
    layer0_outputs(9367) <= not(inputs(13));
    layer0_outputs(9368) <= (inputs(176)) and (inputs(17));
    layer0_outputs(9369) <= inputs(110);
    layer0_outputs(9370) <= '0';
    layer0_outputs(9371) <= not((inputs(140)) xor (inputs(186)));
    layer0_outputs(9372) <= (inputs(56)) and not (inputs(8));
    layer0_outputs(9373) <= (inputs(105)) and not (inputs(205));
    layer0_outputs(9374) <= not((inputs(179)) or (inputs(175)));
    layer0_outputs(9375) <= inputs(215);
    layer0_outputs(9376) <= (inputs(135)) xor (inputs(144));
    layer0_outputs(9377) <= not((inputs(135)) or (inputs(32)));
    layer0_outputs(9378) <= (inputs(1)) and not (inputs(216));
    layer0_outputs(9379) <= inputs(158);
    layer0_outputs(9380) <= inputs(222);
    layer0_outputs(9381) <= (inputs(123)) or (inputs(237));
    layer0_outputs(9382) <= not(inputs(144));
    layer0_outputs(9383) <= not(inputs(229));
    layer0_outputs(9384) <= inputs(108);
    layer0_outputs(9385) <= not(inputs(198)) or (inputs(247));
    layer0_outputs(9386) <= (inputs(64)) and not (inputs(2));
    layer0_outputs(9387) <= not(inputs(153));
    layer0_outputs(9388) <= not(inputs(49));
    layer0_outputs(9389) <= not(inputs(198)) or (inputs(48));
    layer0_outputs(9390) <= inputs(14);
    layer0_outputs(9391) <= not(inputs(142));
    layer0_outputs(9392) <= (inputs(228)) and not (inputs(215));
    layer0_outputs(9393) <= (inputs(21)) or (inputs(36));
    layer0_outputs(9394) <= not(inputs(123)) or (inputs(74));
    layer0_outputs(9395) <= inputs(178);
    layer0_outputs(9396) <= (inputs(92)) or (inputs(92));
    layer0_outputs(9397) <= (inputs(185)) or (inputs(115));
    layer0_outputs(9398) <= not((inputs(224)) or (inputs(34)));
    layer0_outputs(9399) <= not(inputs(37));
    layer0_outputs(9400) <= inputs(152);
    layer0_outputs(9401) <= not(inputs(20)) or (inputs(140));
    layer0_outputs(9402) <= inputs(114);
    layer0_outputs(9403) <= (inputs(69)) or (inputs(160));
    layer0_outputs(9404) <= '1';
    layer0_outputs(9405) <= (inputs(168)) xor (inputs(33));
    layer0_outputs(9406) <= not(inputs(109)) or (inputs(175));
    layer0_outputs(9407) <= '1';
    layer0_outputs(9408) <= (inputs(9)) and (inputs(111));
    layer0_outputs(9409) <= inputs(112);
    layer0_outputs(9410) <= not((inputs(15)) and (inputs(0)));
    layer0_outputs(9411) <= not((inputs(209)) or (inputs(210)));
    layer0_outputs(9412) <= not(inputs(127));
    layer0_outputs(9413) <= (inputs(190)) or (inputs(78));
    layer0_outputs(9414) <= (inputs(238)) or (inputs(243));
    layer0_outputs(9415) <= not((inputs(180)) xor (inputs(174)));
    layer0_outputs(9416) <= not(inputs(88));
    layer0_outputs(9417) <= not((inputs(3)) and (inputs(96)));
    layer0_outputs(9418) <= inputs(121);
    layer0_outputs(9419) <= '0';
    layer0_outputs(9420) <= (inputs(103)) and (inputs(124));
    layer0_outputs(9421) <= inputs(140);
    layer0_outputs(9422) <= not(inputs(109));
    layer0_outputs(9423) <= not((inputs(179)) xor (inputs(157)));
    layer0_outputs(9424) <= (inputs(1)) or (inputs(150));
    layer0_outputs(9425) <= (inputs(118)) and not (inputs(177));
    layer0_outputs(9426) <= inputs(164);
    layer0_outputs(9427) <= '0';
    layer0_outputs(9428) <= inputs(102);
    layer0_outputs(9429) <= not((inputs(123)) or (inputs(50)));
    layer0_outputs(9430) <= not(inputs(148));
    layer0_outputs(9431) <= not((inputs(129)) or (inputs(146)));
    layer0_outputs(9432) <= inputs(106);
    layer0_outputs(9433) <= not(inputs(232));
    layer0_outputs(9434) <= (inputs(146)) xor (inputs(113));
    layer0_outputs(9435) <= not((inputs(112)) or (inputs(39)));
    layer0_outputs(9436) <= inputs(251);
    layer0_outputs(9437) <= not((inputs(22)) or (inputs(4)));
    layer0_outputs(9438) <= (inputs(239)) or (inputs(115));
    layer0_outputs(9439) <= not((inputs(155)) or (inputs(189)));
    layer0_outputs(9440) <= not(inputs(210)) or (inputs(29));
    layer0_outputs(9441) <= not(inputs(105));
    layer0_outputs(9442) <= not((inputs(131)) xor (inputs(165)));
    layer0_outputs(9443) <= not(inputs(137));
    layer0_outputs(9444) <= not((inputs(187)) xor (inputs(90)));
    layer0_outputs(9445) <= inputs(206);
    layer0_outputs(9446) <= inputs(169);
    layer0_outputs(9447) <= inputs(223);
    layer0_outputs(9448) <= inputs(202);
    layer0_outputs(9449) <= (inputs(252)) or (inputs(165));
    layer0_outputs(9450) <= inputs(230);
    layer0_outputs(9451) <= (inputs(243)) and not (inputs(234));
    layer0_outputs(9452) <= (inputs(27)) and not (inputs(161));
    layer0_outputs(9453) <= not((inputs(206)) and (inputs(53)));
    layer0_outputs(9454) <= inputs(4);
    layer0_outputs(9455) <= (inputs(94)) and not (inputs(137));
    layer0_outputs(9456) <= not(inputs(185));
    layer0_outputs(9457) <= (inputs(32)) xor (inputs(184));
    layer0_outputs(9458) <= not(inputs(196));
    layer0_outputs(9459) <= not(inputs(65));
    layer0_outputs(9460) <= not((inputs(167)) and (inputs(250)));
    layer0_outputs(9461) <= inputs(41);
    layer0_outputs(9462) <= not((inputs(13)) xor (inputs(138)));
    layer0_outputs(9463) <= not((inputs(83)) and (inputs(54)));
    layer0_outputs(9464) <= not(inputs(159));
    layer0_outputs(9465) <= not(inputs(220)) or (inputs(143));
    layer0_outputs(9466) <= not((inputs(152)) or (inputs(253)));
    layer0_outputs(9467) <= not((inputs(16)) xor (inputs(116)));
    layer0_outputs(9468) <= not(inputs(67)) or (inputs(175));
    layer0_outputs(9469) <= inputs(39);
    layer0_outputs(9470) <= not((inputs(87)) or (inputs(161)));
    layer0_outputs(9471) <= (inputs(254)) and not (inputs(241));
    layer0_outputs(9472) <= (inputs(90)) and (inputs(43));
    layer0_outputs(9473) <= '1';
    layer0_outputs(9474) <= '0';
    layer0_outputs(9475) <= (inputs(41)) and not (inputs(131));
    layer0_outputs(9476) <= not((inputs(173)) xor (inputs(118)));
    layer0_outputs(9477) <= (inputs(188)) and (inputs(226));
    layer0_outputs(9478) <= (inputs(53)) or (inputs(38));
    layer0_outputs(9479) <= not((inputs(34)) xor (inputs(106)));
    layer0_outputs(9480) <= (inputs(132)) and not (inputs(172));
    layer0_outputs(9481) <= '1';
    layer0_outputs(9482) <= not(inputs(74)) or (inputs(71));
    layer0_outputs(9483) <= inputs(44);
    layer0_outputs(9484) <= '1';
    layer0_outputs(9485) <= inputs(182);
    layer0_outputs(9486) <= (inputs(206)) or (inputs(105));
    layer0_outputs(9487) <= not((inputs(72)) and (inputs(118)));
    layer0_outputs(9488) <= (inputs(223)) or (inputs(198));
    layer0_outputs(9489) <= (inputs(97)) or (inputs(233));
    layer0_outputs(9490) <= not(inputs(39));
    layer0_outputs(9491) <= not((inputs(48)) or (inputs(74)));
    layer0_outputs(9492) <= not(inputs(110));
    layer0_outputs(9493) <= not(inputs(231));
    layer0_outputs(9494) <= not(inputs(27)) or (inputs(169));
    layer0_outputs(9495) <= '1';
    layer0_outputs(9496) <= (inputs(13)) and not (inputs(224));
    layer0_outputs(9497) <= (inputs(199)) xor (inputs(79));
    layer0_outputs(9498) <= not(inputs(58));
    layer0_outputs(9499) <= (inputs(20)) xor (inputs(130));
    layer0_outputs(9500) <= (inputs(24)) or (inputs(160));
    layer0_outputs(9501) <= (inputs(74)) and not (inputs(250));
    layer0_outputs(9502) <= not(inputs(148)) or (inputs(107));
    layer0_outputs(9503) <= (inputs(38)) and not (inputs(157));
    layer0_outputs(9504) <= (inputs(220)) and (inputs(22));
    layer0_outputs(9505) <= (inputs(117)) or (inputs(219));
    layer0_outputs(9506) <= (inputs(230)) xor (inputs(63));
    layer0_outputs(9507) <= not(inputs(203)) or (inputs(75));
    layer0_outputs(9508) <= (inputs(22)) and not (inputs(202));
    layer0_outputs(9509) <= '0';
    layer0_outputs(9510) <= not(inputs(206));
    layer0_outputs(9511) <= (inputs(6)) and (inputs(213));
    layer0_outputs(9512) <= not((inputs(56)) xor (inputs(3)));
    layer0_outputs(9513) <= not(inputs(13));
    layer0_outputs(9514) <= not(inputs(105));
    layer0_outputs(9515) <= not(inputs(178)) or (inputs(184));
    layer0_outputs(9516) <= inputs(234);
    layer0_outputs(9517) <= not(inputs(42));
    layer0_outputs(9518) <= not(inputs(233)) or (inputs(19));
    layer0_outputs(9519) <= (inputs(129)) or (inputs(10));
    layer0_outputs(9520) <= not((inputs(153)) or (inputs(113)));
    layer0_outputs(9521) <= (inputs(89)) xor (inputs(18));
    layer0_outputs(9522) <= (inputs(53)) and not (inputs(197));
    layer0_outputs(9523) <= not((inputs(185)) or (inputs(187)));
    layer0_outputs(9524) <= not(inputs(248)) or (inputs(199));
    layer0_outputs(9525) <= not(inputs(137)) or (inputs(12));
    layer0_outputs(9526) <= not(inputs(89));
    layer0_outputs(9527) <= not(inputs(58));
    layer0_outputs(9528) <= inputs(99);
    layer0_outputs(9529) <= not(inputs(149)) or (inputs(48));
    layer0_outputs(9530) <= inputs(80);
    layer0_outputs(9531) <= not((inputs(64)) or (inputs(68)));
    layer0_outputs(9532) <= not((inputs(239)) and (inputs(139)));
    layer0_outputs(9533) <= (inputs(153)) xor (inputs(105));
    layer0_outputs(9534) <= not(inputs(143));
    layer0_outputs(9535) <= (inputs(33)) xor (inputs(240));
    layer0_outputs(9536) <= not((inputs(229)) or (inputs(182)));
    layer0_outputs(9537) <= (inputs(124)) and not (inputs(40));
    layer0_outputs(9538) <= inputs(204);
    layer0_outputs(9539) <= not((inputs(241)) or (inputs(84)));
    layer0_outputs(9540) <= not(inputs(167)) or (inputs(224));
    layer0_outputs(9541) <= (inputs(237)) or (inputs(85));
    layer0_outputs(9542) <= not(inputs(193)) or (inputs(112));
    layer0_outputs(9543) <= (inputs(188)) and not (inputs(12));
    layer0_outputs(9544) <= (inputs(176)) and not (inputs(173));
    layer0_outputs(9545) <= inputs(90);
    layer0_outputs(9546) <= not((inputs(207)) xor (inputs(2)));
    layer0_outputs(9547) <= inputs(25);
    layer0_outputs(9548) <= '1';
    layer0_outputs(9549) <= not(inputs(128));
    layer0_outputs(9550) <= inputs(180);
    layer0_outputs(9551) <= not(inputs(42)) or (inputs(159));
    layer0_outputs(9552) <= inputs(109);
    layer0_outputs(9553) <= (inputs(28)) xor (inputs(159));
    layer0_outputs(9554) <= (inputs(71)) and not (inputs(58));
    layer0_outputs(9555) <= inputs(102);
    layer0_outputs(9556) <= (inputs(178)) xor (inputs(23));
    layer0_outputs(9557) <= not(inputs(198)) or (inputs(27));
    layer0_outputs(9558) <= inputs(179);
    layer0_outputs(9559) <= (inputs(10)) or (inputs(101));
    layer0_outputs(9560) <= not(inputs(55));
    layer0_outputs(9561) <= not(inputs(222));
    layer0_outputs(9562) <= not(inputs(239));
    layer0_outputs(9563) <= (inputs(27)) or (inputs(95));
    layer0_outputs(9564) <= not(inputs(120)) or (inputs(201));
    layer0_outputs(9565) <= (inputs(168)) or (inputs(219));
    layer0_outputs(9566) <= not(inputs(130)) or (inputs(143));
    layer0_outputs(9567) <= inputs(202);
    layer0_outputs(9568) <= (inputs(240)) xor (inputs(16));
    layer0_outputs(9569) <= not(inputs(11));
    layer0_outputs(9570) <= not((inputs(83)) xor (inputs(216)));
    layer0_outputs(9571) <= (inputs(216)) or (inputs(199));
    layer0_outputs(9572) <= not(inputs(125));
    layer0_outputs(9573) <= (inputs(214)) and not (inputs(254));
    layer0_outputs(9574) <= (inputs(130)) and (inputs(155));
    layer0_outputs(9575) <= inputs(198);
    layer0_outputs(9576) <= not((inputs(245)) xor (inputs(120)));
    layer0_outputs(9577) <= not(inputs(214)) or (inputs(0));
    layer0_outputs(9578) <= (inputs(201)) or (inputs(122));
    layer0_outputs(9579) <= not(inputs(238));
    layer0_outputs(9580) <= not((inputs(140)) or (inputs(207)));
    layer0_outputs(9581) <= (inputs(181)) xor (inputs(2));
    layer0_outputs(9582) <= not(inputs(62));
    layer0_outputs(9583) <= not(inputs(168));
    layer0_outputs(9584) <= not(inputs(61)) or (inputs(210));
    layer0_outputs(9585) <= (inputs(37)) and not (inputs(247));
    layer0_outputs(9586) <= (inputs(149)) and (inputs(56));
    layer0_outputs(9587) <= not(inputs(114));
    layer0_outputs(9588) <= not(inputs(247)) or (inputs(32));
    layer0_outputs(9589) <= not(inputs(18)) or (inputs(51));
    layer0_outputs(9590) <= not(inputs(181));
    layer0_outputs(9591) <= inputs(214);
    layer0_outputs(9592) <= (inputs(139)) or (inputs(120));
    layer0_outputs(9593) <= not((inputs(92)) and (inputs(199)));
    layer0_outputs(9594) <= '0';
    layer0_outputs(9595) <= not(inputs(2));
    layer0_outputs(9596) <= (inputs(4)) or (inputs(123));
    layer0_outputs(9597) <= (inputs(57)) or (inputs(227));
    layer0_outputs(9598) <= not(inputs(154));
    layer0_outputs(9599) <= not((inputs(248)) xor (inputs(9)));
    layer0_outputs(9600) <= not(inputs(183)) or (inputs(198));
    layer0_outputs(9601) <= not(inputs(117));
    layer0_outputs(9602) <= not(inputs(25));
    layer0_outputs(9603) <= not(inputs(186));
    layer0_outputs(9604) <= inputs(164);
    layer0_outputs(9605) <= '0';
    layer0_outputs(9606) <= inputs(136);
    layer0_outputs(9607) <= not(inputs(115));
    layer0_outputs(9608) <= (inputs(154)) or (inputs(92));
    layer0_outputs(9609) <= not(inputs(10)) or (inputs(119));
    layer0_outputs(9610) <= not(inputs(206));
    layer0_outputs(9611) <= not(inputs(131));
    layer0_outputs(9612) <= (inputs(21)) or (inputs(16));
    layer0_outputs(9613) <= not(inputs(93));
    layer0_outputs(9614) <= (inputs(153)) and (inputs(228));
    layer0_outputs(9615) <= inputs(167);
    layer0_outputs(9616) <= inputs(225);
    layer0_outputs(9617) <= (inputs(24)) and not (inputs(153));
    layer0_outputs(9618) <= not(inputs(59));
    layer0_outputs(9619) <= '1';
    layer0_outputs(9620) <= (inputs(31)) and not (inputs(163));
    layer0_outputs(9621) <= not(inputs(51)) or (inputs(146));
    layer0_outputs(9622) <= not(inputs(152)) or (inputs(208));
    layer0_outputs(9623) <= '1';
    layer0_outputs(9624) <= not((inputs(62)) or (inputs(150)));
    layer0_outputs(9625) <= not(inputs(97)) or (inputs(208));
    layer0_outputs(9626) <= (inputs(139)) or (inputs(192));
    layer0_outputs(9627) <= not((inputs(252)) or (inputs(133)));
    layer0_outputs(9628) <= not((inputs(144)) or (inputs(142)));
    layer0_outputs(9629) <= not((inputs(246)) or (inputs(7)));
    layer0_outputs(9630) <= not(inputs(46));
    layer0_outputs(9631) <= (inputs(170)) and not (inputs(97));
    layer0_outputs(9632) <= not(inputs(160));
    layer0_outputs(9633) <= (inputs(240)) and not (inputs(87));
    layer0_outputs(9634) <= (inputs(106)) and not (inputs(43));
    layer0_outputs(9635) <= '0';
    layer0_outputs(9636) <= (inputs(203)) and not (inputs(31));
    layer0_outputs(9637) <= (inputs(139)) or (inputs(93));
    layer0_outputs(9638) <= inputs(98);
    layer0_outputs(9639) <= (inputs(230)) and not (inputs(142));
    layer0_outputs(9640) <= not(inputs(253));
    layer0_outputs(9641) <= not(inputs(118));
    layer0_outputs(9642) <= (inputs(51)) and not (inputs(176));
    layer0_outputs(9643) <= not((inputs(221)) xor (inputs(139)));
    layer0_outputs(9644) <= (inputs(132)) and not (inputs(26));
    layer0_outputs(9645) <= inputs(30);
    layer0_outputs(9646) <= (inputs(214)) and not (inputs(110));
    layer0_outputs(9647) <= (inputs(236)) xor (inputs(159));
    layer0_outputs(9648) <= (inputs(207)) and not (inputs(63));
    layer0_outputs(9649) <= not((inputs(161)) or (inputs(187)));
    layer0_outputs(9650) <= '1';
    layer0_outputs(9651) <= (inputs(13)) or (inputs(144));
    layer0_outputs(9652) <= (inputs(60)) or (inputs(251));
    layer0_outputs(9653) <= (inputs(80)) and not (inputs(26));
    layer0_outputs(9654) <= not(inputs(74));
    layer0_outputs(9655) <= (inputs(77)) or (inputs(9));
    layer0_outputs(9656) <= not(inputs(123)) or (inputs(22));
    layer0_outputs(9657) <= (inputs(17)) or (inputs(182));
    layer0_outputs(9658) <= not(inputs(131));
    layer0_outputs(9659) <= (inputs(4)) or (inputs(228));
    layer0_outputs(9660) <= not(inputs(218)) or (inputs(57));
    layer0_outputs(9661) <= not(inputs(24));
    layer0_outputs(9662) <= (inputs(98)) xor (inputs(73));
    layer0_outputs(9663) <= (inputs(133)) and not (inputs(139));
    layer0_outputs(9664) <= not(inputs(203)) or (inputs(99));
    layer0_outputs(9665) <= not(inputs(11)) or (inputs(146));
    layer0_outputs(9666) <= not(inputs(224));
    layer0_outputs(9667) <= not((inputs(11)) xor (inputs(43)));
    layer0_outputs(9668) <= (inputs(88)) and not (inputs(87));
    layer0_outputs(9669) <= not((inputs(92)) and (inputs(22)));
    layer0_outputs(9670) <= not(inputs(209));
    layer0_outputs(9671) <= (inputs(58)) and not (inputs(78));
    layer0_outputs(9672) <= inputs(241);
    layer0_outputs(9673) <= (inputs(205)) or (inputs(222));
    layer0_outputs(9674) <= not(inputs(9));
    layer0_outputs(9675) <= not(inputs(144)) or (inputs(54));
    layer0_outputs(9676) <= (inputs(1)) or (inputs(245));
    layer0_outputs(9677) <= (inputs(239)) or (inputs(180));
    layer0_outputs(9678) <= not(inputs(85));
    layer0_outputs(9679) <= inputs(237);
    layer0_outputs(9680) <= inputs(34);
    layer0_outputs(9681) <= '1';
    layer0_outputs(9682) <= (inputs(2)) or (inputs(43));
    layer0_outputs(9683) <= (inputs(165)) and not (inputs(20));
    layer0_outputs(9684) <= (inputs(192)) and not (inputs(118));
    layer0_outputs(9685) <= (inputs(85)) or (inputs(240));
    layer0_outputs(9686) <= not(inputs(182)) or (inputs(60));
    layer0_outputs(9687) <= inputs(60);
    layer0_outputs(9688) <= (inputs(71)) and not (inputs(179));
    layer0_outputs(9689) <= (inputs(108)) and (inputs(1));
    layer0_outputs(9690) <= not(inputs(20));
    layer0_outputs(9691) <= not((inputs(183)) xor (inputs(171)));
    layer0_outputs(9692) <= (inputs(233)) xor (inputs(208));
    layer0_outputs(9693) <= not((inputs(34)) xor (inputs(126)));
    layer0_outputs(9694) <= not((inputs(204)) xor (inputs(29)));
    layer0_outputs(9695) <= inputs(178);
    layer0_outputs(9696) <= (inputs(25)) or (inputs(238));
    layer0_outputs(9697) <= not(inputs(17)) or (inputs(201));
    layer0_outputs(9698) <= not((inputs(49)) or (inputs(148)));
    layer0_outputs(9699) <= (inputs(245)) and not (inputs(119));
    layer0_outputs(9700) <= not((inputs(115)) or (inputs(84)));
    layer0_outputs(9701) <= not(inputs(152));
    layer0_outputs(9702) <= inputs(149);
    layer0_outputs(9703) <= inputs(124);
    layer0_outputs(9704) <= not(inputs(167)) or (inputs(48));
    layer0_outputs(9705) <= (inputs(53)) and not (inputs(108));
    layer0_outputs(9706) <= not((inputs(188)) or (inputs(255)));
    layer0_outputs(9707) <= inputs(105);
    layer0_outputs(9708) <= not(inputs(95)) or (inputs(126));
    layer0_outputs(9709) <= not((inputs(241)) xor (inputs(58)));
    layer0_outputs(9710) <= not((inputs(177)) or (inputs(193)));
    layer0_outputs(9711) <= inputs(48);
    layer0_outputs(9712) <= (inputs(78)) or (inputs(192));
    layer0_outputs(9713) <= not((inputs(198)) xor (inputs(80)));
    layer0_outputs(9714) <= '1';
    layer0_outputs(9715) <= (inputs(233)) and not (inputs(58));
    layer0_outputs(9716) <= not(inputs(38));
    layer0_outputs(9717) <= '1';
    layer0_outputs(9718) <= (inputs(247)) or (inputs(77));
    layer0_outputs(9719) <= not(inputs(8));
    layer0_outputs(9720) <= not((inputs(65)) xor (inputs(98)));
    layer0_outputs(9721) <= inputs(46);
    layer0_outputs(9722) <= not(inputs(26));
    layer0_outputs(9723) <= not(inputs(47)) or (inputs(243));
    layer0_outputs(9724) <= (inputs(196)) xor (inputs(132));
    layer0_outputs(9725) <= not(inputs(188)) or (inputs(159));
    layer0_outputs(9726) <= not(inputs(213)) or (inputs(57));
    layer0_outputs(9727) <= inputs(114);
    layer0_outputs(9728) <= not(inputs(173));
    layer0_outputs(9729) <= (inputs(9)) and not (inputs(32));
    layer0_outputs(9730) <= not((inputs(97)) or (inputs(8)));
    layer0_outputs(9731) <= inputs(77);
    layer0_outputs(9732) <= not((inputs(172)) xor (inputs(210)));
    layer0_outputs(9733) <= inputs(230);
    layer0_outputs(9734) <= not(inputs(102));
    layer0_outputs(9735) <= not(inputs(231));
    layer0_outputs(9736) <= (inputs(226)) and not (inputs(139));
    layer0_outputs(9737) <= (inputs(7)) and (inputs(69));
    layer0_outputs(9738) <= inputs(69);
    layer0_outputs(9739) <= not((inputs(10)) or (inputs(5)));
    layer0_outputs(9740) <= inputs(175);
    layer0_outputs(9741) <= (inputs(110)) and (inputs(166));
    layer0_outputs(9742) <= '1';
    layer0_outputs(9743) <= (inputs(23)) or (inputs(151));
    layer0_outputs(9744) <= (inputs(100)) and not (inputs(163));
    layer0_outputs(9745) <= not(inputs(18)) or (inputs(169));
    layer0_outputs(9746) <= not(inputs(100)) or (inputs(233));
    layer0_outputs(9747) <= (inputs(172)) and not (inputs(64));
    layer0_outputs(9748) <= inputs(85);
    layer0_outputs(9749) <= not(inputs(140)) or (inputs(145));
    layer0_outputs(9750) <= not((inputs(208)) or (inputs(242)));
    layer0_outputs(9751) <= not(inputs(178));
    layer0_outputs(9752) <= not(inputs(242)) or (inputs(19));
    layer0_outputs(9753) <= not((inputs(216)) and (inputs(210)));
    layer0_outputs(9754) <= (inputs(122)) and not (inputs(165));
    layer0_outputs(9755) <= (inputs(114)) or (inputs(99));
    layer0_outputs(9756) <= (inputs(17)) and (inputs(106));
    layer0_outputs(9757) <= (inputs(47)) xor (inputs(18));
    layer0_outputs(9758) <= (inputs(103)) xor (inputs(164));
    layer0_outputs(9759) <= not(inputs(74));
    layer0_outputs(9760) <= inputs(117);
    layer0_outputs(9761) <= (inputs(27)) xor (inputs(78));
    layer0_outputs(9762) <= (inputs(63)) or (inputs(23));
    layer0_outputs(9763) <= (inputs(101)) and not (inputs(20));
    layer0_outputs(9764) <= (inputs(108)) and not (inputs(20));
    layer0_outputs(9765) <= (inputs(99)) xor (inputs(99));
    layer0_outputs(9766) <= not(inputs(245));
    layer0_outputs(9767) <= (inputs(106)) and not (inputs(220));
    layer0_outputs(9768) <= '0';
    layer0_outputs(9769) <= not((inputs(221)) or (inputs(149)));
    layer0_outputs(9770) <= not(inputs(72)) or (inputs(165));
    layer0_outputs(9771) <= not(inputs(217));
    layer0_outputs(9772) <= not(inputs(103));
    layer0_outputs(9773) <= (inputs(207)) and not (inputs(201));
    layer0_outputs(9774) <= not(inputs(91));
    layer0_outputs(9775) <= '0';
    layer0_outputs(9776) <= not(inputs(29)) or (inputs(90));
    layer0_outputs(9777) <= (inputs(193)) or (inputs(54));
    layer0_outputs(9778) <= not(inputs(156));
    layer0_outputs(9779) <= inputs(110);
    layer0_outputs(9780) <= not(inputs(97));
    layer0_outputs(9781) <= not((inputs(133)) xor (inputs(38)));
    layer0_outputs(9782) <= inputs(212);
    layer0_outputs(9783) <= (inputs(64)) xor (inputs(248));
    layer0_outputs(9784) <= (inputs(205)) and (inputs(122));
    layer0_outputs(9785) <= inputs(85);
    layer0_outputs(9786) <= (inputs(233)) or (inputs(113));
    layer0_outputs(9787) <= not((inputs(149)) xor (inputs(115)));
    layer0_outputs(9788) <= (inputs(47)) and not (inputs(213));
    layer0_outputs(9789) <= (inputs(208)) xor (inputs(37));
    layer0_outputs(9790) <= inputs(120);
    layer0_outputs(9791) <= (inputs(235)) and (inputs(200));
    layer0_outputs(9792) <= not(inputs(49)) or (inputs(6));
    layer0_outputs(9793) <= not(inputs(165));
    layer0_outputs(9794) <= (inputs(101)) and not (inputs(161));
    layer0_outputs(9795) <= (inputs(49)) or (inputs(182));
    layer0_outputs(9796) <= inputs(132);
    layer0_outputs(9797) <= (inputs(219)) or (inputs(225));
    layer0_outputs(9798) <= (inputs(248)) and (inputs(184));
    layer0_outputs(9799) <= inputs(62);
    layer0_outputs(9800) <= inputs(6);
    layer0_outputs(9801) <= inputs(123);
    layer0_outputs(9802) <= inputs(163);
    layer0_outputs(9803) <= inputs(96);
    layer0_outputs(9804) <= not((inputs(87)) or (inputs(225)));
    layer0_outputs(9805) <= (inputs(47)) and (inputs(227));
    layer0_outputs(9806) <= not((inputs(232)) and (inputs(26)));
    layer0_outputs(9807) <= not((inputs(117)) or (inputs(15)));
    layer0_outputs(9808) <= inputs(130);
    layer0_outputs(9809) <= '0';
    layer0_outputs(9810) <= not(inputs(53)) or (inputs(240));
    layer0_outputs(9811) <= inputs(83);
    layer0_outputs(9812) <= not(inputs(173));
    layer0_outputs(9813) <= (inputs(239)) xor (inputs(2));
    layer0_outputs(9814) <= not(inputs(237));
    layer0_outputs(9815) <= not(inputs(168));
    layer0_outputs(9816) <= not(inputs(7)) or (inputs(89));
    layer0_outputs(9817) <= '1';
    layer0_outputs(9818) <= not(inputs(169)) or (inputs(233));
    layer0_outputs(9819) <= not(inputs(156));
    layer0_outputs(9820) <= inputs(103);
    layer0_outputs(9821) <= (inputs(171)) or (inputs(179));
    layer0_outputs(9822) <= not((inputs(69)) xor (inputs(49)));
    layer0_outputs(9823) <= (inputs(10)) and (inputs(99));
    layer0_outputs(9824) <= not(inputs(9)) or (inputs(114));
    layer0_outputs(9825) <= not((inputs(212)) or (inputs(208)));
    layer0_outputs(9826) <= (inputs(94)) or (inputs(230));
    layer0_outputs(9827) <= not((inputs(48)) xor (inputs(224)));
    layer0_outputs(9828) <= (inputs(95)) xor (inputs(18));
    layer0_outputs(9829) <= (inputs(60)) xor (inputs(45));
    layer0_outputs(9830) <= not(inputs(31));
    layer0_outputs(9831) <= '0';
    layer0_outputs(9832) <= not(inputs(174));
    layer0_outputs(9833) <= (inputs(213)) and not (inputs(34));
    layer0_outputs(9834) <= not(inputs(195));
    layer0_outputs(9835) <= not(inputs(105));
    layer0_outputs(9836) <= not(inputs(132));
    layer0_outputs(9837) <= inputs(63);
    layer0_outputs(9838) <= (inputs(52)) xor (inputs(87));
    layer0_outputs(9839) <= (inputs(97)) xor (inputs(235));
    layer0_outputs(9840) <= not(inputs(185));
    layer0_outputs(9841) <= not(inputs(73)) or (inputs(81));
    layer0_outputs(9842) <= inputs(130);
    layer0_outputs(9843) <= (inputs(56)) or (inputs(200));
    layer0_outputs(9844) <= inputs(208);
    layer0_outputs(9845) <= not(inputs(140)) or (inputs(177));
    layer0_outputs(9846) <= '1';
    layer0_outputs(9847) <= (inputs(34)) or (inputs(76));
    layer0_outputs(9848) <= not(inputs(213)) or (inputs(45));
    layer0_outputs(9849) <= (inputs(13)) xor (inputs(212));
    layer0_outputs(9850) <= inputs(122);
    layer0_outputs(9851) <= not(inputs(117)) or (inputs(106));
    layer0_outputs(9852) <= not((inputs(56)) or (inputs(220)));
    layer0_outputs(9853) <= not((inputs(41)) or (inputs(57)));
    layer0_outputs(9854) <= not((inputs(193)) or (inputs(109)));
    layer0_outputs(9855) <= '0';
    layer0_outputs(9856) <= not(inputs(164));
    layer0_outputs(9857) <= not(inputs(114));
    layer0_outputs(9858) <= inputs(19);
    layer0_outputs(9859) <= not((inputs(222)) or (inputs(192)));
    layer0_outputs(9860) <= not((inputs(191)) or (inputs(212)));
    layer0_outputs(9861) <= not(inputs(92)) or (inputs(42));
    layer0_outputs(9862) <= not(inputs(10)) or (inputs(148));
    layer0_outputs(9863) <= (inputs(117)) and not (inputs(113));
    layer0_outputs(9864) <= (inputs(20)) xor (inputs(155));
    layer0_outputs(9865) <= not((inputs(148)) xor (inputs(160)));
    layer0_outputs(9866) <= (inputs(212)) and not (inputs(64));
    layer0_outputs(9867) <= inputs(89);
    layer0_outputs(9868) <= not(inputs(136)) or (inputs(59));
    layer0_outputs(9869) <= not(inputs(190));
    layer0_outputs(9870) <= (inputs(162)) xor (inputs(188));
    layer0_outputs(9871) <= not((inputs(174)) xor (inputs(226)));
    layer0_outputs(9872) <= '0';
    layer0_outputs(9873) <= not((inputs(233)) xor (inputs(62)));
    layer0_outputs(9874) <= '0';
    layer0_outputs(9875) <= not((inputs(254)) or (inputs(43)));
    layer0_outputs(9876) <= not(inputs(8)) or (inputs(103));
    layer0_outputs(9877) <= inputs(33);
    layer0_outputs(9878) <= not(inputs(129));
    layer0_outputs(9879) <= not((inputs(48)) or (inputs(89)));
    layer0_outputs(9880) <= inputs(59);
    layer0_outputs(9881) <= inputs(213);
    layer0_outputs(9882) <= not((inputs(203)) or (inputs(224)));
    layer0_outputs(9883) <= (inputs(17)) and not (inputs(95));
    layer0_outputs(9884) <= not(inputs(36)) or (inputs(184));
    layer0_outputs(9885) <= not(inputs(137)) or (inputs(24));
    layer0_outputs(9886) <= not(inputs(138));
    layer0_outputs(9887) <= not((inputs(94)) or (inputs(209)));
    layer0_outputs(9888) <= not(inputs(19)) or (inputs(234));
    layer0_outputs(9889) <= not(inputs(212));
    layer0_outputs(9890) <= (inputs(15)) or (inputs(125));
    layer0_outputs(9891) <= not((inputs(67)) xor (inputs(78)));
    layer0_outputs(9892) <= (inputs(146)) or (inputs(177));
    layer0_outputs(9893) <= not((inputs(96)) and (inputs(206)));
    layer0_outputs(9894) <= not((inputs(162)) and (inputs(93)));
    layer0_outputs(9895) <= (inputs(253)) or (inputs(151));
    layer0_outputs(9896) <= '0';
    layer0_outputs(9897) <= not(inputs(223)) or (inputs(23));
    layer0_outputs(9898) <= not((inputs(247)) or (inputs(245)));
    layer0_outputs(9899) <= not(inputs(82));
    layer0_outputs(9900) <= (inputs(68)) and not (inputs(190));
    layer0_outputs(9901) <= inputs(109);
    layer0_outputs(9902) <= inputs(47);
    layer0_outputs(9903) <= not(inputs(123));
    layer0_outputs(9904) <= not((inputs(236)) or (inputs(207)));
    layer0_outputs(9905) <= inputs(231);
    layer0_outputs(9906) <= not(inputs(61)) or (inputs(92));
    layer0_outputs(9907) <= not(inputs(25)) or (inputs(209));
    layer0_outputs(9908) <= not((inputs(7)) or (inputs(202)));
    layer0_outputs(9909) <= not(inputs(230));
    layer0_outputs(9910) <= '1';
    layer0_outputs(9911) <= (inputs(11)) and not (inputs(1));
    layer0_outputs(9912) <= (inputs(75)) or (inputs(210));
    layer0_outputs(9913) <= inputs(170);
    layer0_outputs(9914) <= inputs(99);
    layer0_outputs(9915) <= inputs(193);
    layer0_outputs(9916) <= (inputs(177)) and (inputs(35));
    layer0_outputs(9917) <= not(inputs(178)) or (inputs(15));
    layer0_outputs(9918) <= (inputs(240)) or (inputs(151));
    layer0_outputs(9919) <= not((inputs(252)) xor (inputs(186)));
    layer0_outputs(9920) <= not(inputs(86));
    layer0_outputs(9921) <= (inputs(148)) and not (inputs(226));
    layer0_outputs(9922) <= not((inputs(2)) and (inputs(40)));
    layer0_outputs(9923) <= not(inputs(182));
    layer0_outputs(9924) <= (inputs(31)) and not (inputs(239));
    layer0_outputs(9925) <= not(inputs(149)) or (inputs(123));
    layer0_outputs(9926) <= inputs(40);
    layer0_outputs(9927) <= not(inputs(93));
    layer0_outputs(9928) <= not((inputs(114)) or (inputs(99)));
    layer0_outputs(9929) <= (inputs(161)) xor (inputs(48));
    layer0_outputs(9930) <= (inputs(105)) and not (inputs(249));
    layer0_outputs(9931) <= not(inputs(250)) or (inputs(99));
    layer0_outputs(9932) <= (inputs(120)) and not (inputs(50));
    layer0_outputs(9933) <= '0';
    layer0_outputs(9934) <= not(inputs(9));
    layer0_outputs(9935) <= not((inputs(146)) xor (inputs(104)));
    layer0_outputs(9936) <= (inputs(101)) or (inputs(246));
    layer0_outputs(9937) <= not(inputs(27));
    layer0_outputs(9938) <= not(inputs(153)) or (inputs(135));
    layer0_outputs(9939) <= inputs(47);
    layer0_outputs(9940) <= not(inputs(179));
    layer0_outputs(9941) <= (inputs(129)) or (inputs(138));
    layer0_outputs(9942) <= not((inputs(20)) and (inputs(215)));
    layer0_outputs(9943) <= not(inputs(187));
    layer0_outputs(9944) <= '1';
    layer0_outputs(9945) <= not(inputs(185));
    layer0_outputs(9946) <= not(inputs(161));
    layer0_outputs(9947) <= not((inputs(200)) xor (inputs(232)));
    layer0_outputs(9948) <= not((inputs(126)) or (inputs(254)));
    layer0_outputs(9949) <= inputs(130);
    layer0_outputs(9950) <= (inputs(127)) and not (inputs(112));
    layer0_outputs(9951) <= inputs(54);
    layer0_outputs(9952) <= not((inputs(80)) xor (inputs(248)));
    layer0_outputs(9953) <= inputs(150);
    layer0_outputs(9954) <= (inputs(202)) and not (inputs(95));
    layer0_outputs(9955) <= not(inputs(168)) or (inputs(193));
    layer0_outputs(9956) <= (inputs(122)) and not (inputs(218));
    layer0_outputs(9957) <= (inputs(141)) and (inputs(162));
    layer0_outputs(9958) <= not((inputs(218)) and (inputs(147)));
    layer0_outputs(9959) <= not(inputs(177));
    layer0_outputs(9960) <= inputs(56);
    layer0_outputs(9961) <= (inputs(196)) and not (inputs(20));
    layer0_outputs(9962) <= not((inputs(102)) and (inputs(53)));
    layer0_outputs(9963) <= not(inputs(65));
    layer0_outputs(9964) <= not(inputs(215));
    layer0_outputs(9965) <= inputs(9);
    layer0_outputs(9966) <= (inputs(123)) and (inputs(40));
    layer0_outputs(9967) <= not(inputs(214)) or (inputs(48));
    layer0_outputs(9968) <= not(inputs(214)) or (inputs(113));
    layer0_outputs(9969) <= (inputs(133)) or (inputs(68));
    layer0_outputs(9970) <= not(inputs(59));
    layer0_outputs(9971) <= not(inputs(26));
    layer0_outputs(9972) <= not((inputs(124)) and (inputs(93)));
    layer0_outputs(9973) <= inputs(74);
    layer0_outputs(9974) <= inputs(61);
    layer0_outputs(9975) <= (inputs(68)) and not (inputs(120));
    layer0_outputs(9976) <= not((inputs(5)) xor (inputs(70)));
    layer0_outputs(9977) <= (inputs(92)) or (inputs(31));
    layer0_outputs(9978) <= inputs(100);
    layer0_outputs(9979) <= (inputs(109)) xor (inputs(237));
    layer0_outputs(9980) <= not((inputs(130)) or (inputs(172)));
    layer0_outputs(9981) <= (inputs(86)) and not (inputs(32));
    layer0_outputs(9982) <= (inputs(194)) and not (inputs(6));
    layer0_outputs(9983) <= inputs(89);
    layer0_outputs(9984) <= inputs(88);
    layer0_outputs(9985) <= (inputs(180)) or (inputs(158));
    layer0_outputs(9986) <= inputs(142);
    layer0_outputs(9987) <= '0';
    layer0_outputs(9988) <= (inputs(223)) xor (inputs(9));
    layer0_outputs(9989) <= not(inputs(26)) or (inputs(222));
    layer0_outputs(9990) <= '0';
    layer0_outputs(9991) <= (inputs(54)) or (inputs(82));
    layer0_outputs(9992) <= not(inputs(214));
    layer0_outputs(9993) <= not(inputs(141)) or (inputs(13));
    layer0_outputs(9994) <= (inputs(34)) or (inputs(83));
    layer0_outputs(9995) <= (inputs(5)) xor (inputs(214));
    layer0_outputs(9996) <= inputs(204);
    layer0_outputs(9997) <= inputs(28);
    layer0_outputs(9998) <= inputs(68);
    layer0_outputs(9999) <= (inputs(94)) and not (inputs(51));
    layer0_outputs(10000) <= (inputs(62)) and not (inputs(187));
    layer0_outputs(10001) <= not((inputs(5)) or (inputs(224)));
    layer0_outputs(10002) <= not(inputs(82));
    layer0_outputs(10003) <= (inputs(176)) xor (inputs(222));
    layer0_outputs(10004) <= not(inputs(8)) or (inputs(13));
    layer0_outputs(10005) <= (inputs(29)) and not (inputs(141));
    layer0_outputs(10006) <= inputs(181);
    layer0_outputs(10007) <= not(inputs(249)) or (inputs(63));
    layer0_outputs(10008) <= not(inputs(202));
    layer0_outputs(10009) <= inputs(28);
    layer0_outputs(10010) <= (inputs(4)) or (inputs(187));
    layer0_outputs(10011) <= (inputs(250)) or (inputs(149));
    layer0_outputs(10012) <= not(inputs(69));
    layer0_outputs(10013) <= not(inputs(97));
    layer0_outputs(10014) <= not((inputs(123)) or (inputs(14)));
    layer0_outputs(10015) <= (inputs(68)) xor (inputs(81));
    layer0_outputs(10016) <= (inputs(198)) and not (inputs(27));
    layer0_outputs(10017) <= not((inputs(224)) xor (inputs(89)));
    layer0_outputs(10018) <= not(inputs(210));
    layer0_outputs(10019) <= not(inputs(31));
    layer0_outputs(10020) <= not(inputs(108));
    layer0_outputs(10021) <= (inputs(11)) and not (inputs(251));
    layer0_outputs(10022) <= (inputs(115)) xor (inputs(255));
    layer0_outputs(10023) <= (inputs(90)) and not (inputs(201));
    layer0_outputs(10024) <= inputs(103);
    layer0_outputs(10025) <= inputs(108);
    layer0_outputs(10026) <= (inputs(212)) and not (inputs(109));
    layer0_outputs(10027) <= (inputs(144)) or (inputs(211));
    layer0_outputs(10028) <= (inputs(103)) and not (inputs(116));
    layer0_outputs(10029) <= not(inputs(31)) or (inputs(11));
    layer0_outputs(10030) <= not(inputs(164));
    layer0_outputs(10031) <= inputs(130);
    layer0_outputs(10032) <= not(inputs(234));
    layer0_outputs(10033) <= not(inputs(252));
    layer0_outputs(10034) <= (inputs(137)) or (inputs(76));
    layer0_outputs(10035) <= not((inputs(41)) and (inputs(42)));
    layer0_outputs(10036) <= not(inputs(233));
    layer0_outputs(10037) <= not(inputs(29));
    layer0_outputs(10038) <= '1';
    layer0_outputs(10039) <= inputs(213);
    layer0_outputs(10040) <= not((inputs(48)) xor (inputs(84)));
    layer0_outputs(10041) <= inputs(132);
    layer0_outputs(10042) <= not((inputs(77)) xor (inputs(183)));
    layer0_outputs(10043) <= not(inputs(213));
    layer0_outputs(10044) <= not(inputs(37)) or (inputs(238));
    layer0_outputs(10045) <= not((inputs(88)) and (inputs(115)));
    layer0_outputs(10046) <= (inputs(120)) and not (inputs(74));
    layer0_outputs(10047) <= (inputs(134)) or (inputs(7));
    layer0_outputs(10048) <= inputs(99);
    layer0_outputs(10049) <= (inputs(23)) and not (inputs(31));
    layer0_outputs(10050) <= (inputs(190)) or (inputs(193));
    layer0_outputs(10051) <= inputs(84);
    layer0_outputs(10052) <= (inputs(41)) and not (inputs(102));
    layer0_outputs(10053) <= (inputs(175)) or (inputs(176));
    layer0_outputs(10054) <= (inputs(181)) xor (inputs(89));
    layer0_outputs(10055) <= not(inputs(124)) or (inputs(250));
    layer0_outputs(10056) <= not(inputs(236));
    layer0_outputs(10057) <= inputs(70);
    layer0_outputs(10058) <= (inputs(168)) and not (inputs(24));
    layer0_outputs(10059) <= (inputs(140)) and (inputs(43));
    layer0_outputs(10060) <= inputs(194);
    layer0_outputs(10061) <= not((inputs(62)) xor (inputs(107)));
    layer0_outputs(10062) <= not(inputs(140));
    layer0_outputs(10063) <= (inputs(122)) and not (inputs(19));
    layer0_outputs(10064) <= (inputs(167)) and not (inputs(93));
    layer0_outputs(10065) <= (inputs(160)) xor (inputs(122));
    layer0_outputs(10066) <= inputs(202);
    layer0_outputs(10067) <= (inputs(230)) or (inputs(210));
    layer0_outputs(10068) <= not(inputs(61));
    layer0_outputs(10069) <= not((inputs(231)) or (inputs(191)));
    layer0_outputs(10070) <= (inputs(184)) and not (inputs(215));
    layer0_outputs(10071) <= inputs(59);
    layer0_outputs(10072) <= not(inputs(140)) or (inputs(17));
    layer0_outputs(10073) <= not(inputs(226));
    layer0_outputs(10074) <= (inputs(237)) xor (inputs(141));
    layer0_outputs(10075) <= '1';
    layer0_outputs(10076) <= inputs(83);
    layer0_outputs(10077) <= '1';
    layer0_outputs(10078) <= not(inputs(63));
    layer0_outputs(10079) <= (inputs(51)) and not (inputs(16));
    layer0_outputs(10080) <= inputs(59);
    layer0_outputs(10081) <= '0';
    layer0_outputs(10082) <= not(inputs(160)) or (inputs(17));
    layer0_outputs(10083) <= (inputs(241)) or (inputs(180));
    layer0_outputs(10084) <= not(inputs(205));
    layer0_outputs(10085) <= not(inputs(133)) or (inputs(241));
    layer0_outputs(10086) <= not((inputs(183)) xor (inputs(1)));
    layer0_outputs(10087) <= (inputs(45)) or (inputs(160));
    layer0_outputs(10088) <= not(inputs(194)) or (inputs(118));
    layer0_outputs(10089) <= not(inputs(173));
    layer0_outputs(10090) <= '0';
    layer0_outputs(10091) <= not(inputs(248));
    layer0_outputs(10092) <= inputs(209);
    layer0_outputs(10093) <= not(inputs(158)) or (inputs(238));
    layer0_outputs(10094) <= '0';
    layer0_outputs(10095) <= not((inputs(48)) or (inputs(194)));
    layer0_outputs(10096) <= not(inputs(103));
    layer0_outputs(10097) <= inputs(35);
    layer0_outputs(10098) <= (inputs(211)) and not (inputs(13));
    layer0_outputs(10099) <= not(inputs(245)) or (inputs(255));
    layer0_outputs(10100) <= inputs(3);
    layer0_outputs(10101) <= inputs(110);
    layer0_outputs(10102) <= (inputs(192)) and not (inputs(165));
    layer0_outputs(10103) <= inputs(106);
    layer0_outputs(10104) <= (inputs(36)) or (inputs(81));
    layer0_outputs(10105) <= not(inputs(212));
    layer0_outputs(10106) <= not(inputs(88)) or (inputs(60));
    layer0_outputs(10107) <= inputs(20);
    layer0_outputs(10108) <= not((inputs(0)) or (inputs(210)));
    layer0_outputs(10109) <= not((inputs(254)) or (inputs(176)));
    layer0_outputs(10110) <= not(inputs(195)) or (inputs(98));
    layer0_outputs(10111) <= not((inputs(137)) or (inputs(107)));
    layer0_outputs(10112) <= inputs(238);
    layer0_outputs(10113) <= not(inputs(174));
    layer0_outputs(10114) <= not((inputs(176)) xor (inputs(80)));
    layer0_outputs(10115) <= (inputs(26)) or (inputs(111));
    layer0_outputs(10116) <= not((inputs(76)) and (inputs(132)));
    layer0_outputs(10117) <= (inputs(194)) and (inputs(162));
    layer0_outputs(10118) <= not((inputs(229)) or (inputs(205)));
    layer0_outputs(10119) <= (inputs(178)) and not (inputs(13));
    layer0_outputs(10120) <= inputs(102);
    layer0_outputs(10121) <= (inputs(180)) xor (inputs(145));
    layer0_outputs(10122) <= not(inputs(127));
    layer0_outputs(10123) <= (inputs(123)) and not (inputs(71));
    layer0_outputs(10124) <= inputs(194);
    layer0_outputs(10125) <= not(inputs(167));
    layer0_outputs(10126) <= (inputs(197)) or (inputs(110));
    layer0_outputs(10127) <= (inputs(104)) and not (inputs(193));
    layer0_outputs(10128) <= inputs(202);
    layer0_outputs(10129) <= not((inputs(122)) xor (inputs(61)));
    layer0_outputs(10130) <= inputs(189);
    layer0_outputs(10131) <= (inputs(54)) or (inputs(208));
    layer0_outputs(10132) <= not(inputs(169));
    layer0_outputs(10133) <= (inputs(7)) and not (inputs(134));
    layer0_outputs(10134) <= inputs(114);
    layer0_outputs(10135) <= (inputs(83)) and not (inputs(32));
    layer0_outputs(10136) <= not(inputs(20)) or (inputs(178));
    layer0_outputs(10137) <= (inputs(234)) and not (inputs(128));
    layer0_outputs(10138) <= not((inputs(35)) or (inputs(152)));
    layer0_outputs(10139) <= inputs(206);
    layer0_outputs(10140) <= (inputs(120)) and not (inputs(157));
    layer0_outputs(10141) <= (inputs(12)) and not (inputs(130));
    layer0_outputs(10142) <= (inputs(125)) and not (inputs(236));
    layer0_outputs(10143) <= not(inputs(41));
    layer0_outputs(10144) <= not(inputs(201)) or (inputs(98));
    layer0_outputs(10145) <= not(inputs(242)) or (inputs(66));
    layer0_outputs(10146) <= not(inputs(167));
    layer0_outputs(10147) <= not(inputs(227)) or (inputs(73));
    layer0_outputs(10148) <= not(inputs(40));
    layer0_outputs(10149) <= inputs(29);
    layer0_outputs(10150) <= (inputs(249)) and not (inputs(35));
    layer0_outputs(10151) <= (inputs(249)) or (inputs(94));
    layer0_outputs(10152) <= not(inputs(31));
    layer0_outputs(10153) <= (inputs(63)) and not (inputs(244));
    layer0_outputs(10154) <= not((inputs(112)) xor (inputs(63)));
    layer0_outputs(10155) <= '1';
    layer0_outputs(10156) <= '1';
    layer0_outputs(10157) <= not(inputs(30)) or (inputs(127));
    layer0_outputs(10158) <= (inputs(109)) and not (inputs(236));
    layer0_outputs(10159) <= (inputs(208)) or (inputs(88));
    layer0_outputs(10160) <= '1';
    layer0_outputs(10161) <= not((inputs(122)) or (inputs(186)));
    layer0_outputs(10162) <= inputs(83);
    layer0_outputs(10163) <= not((inputs(24)) xor (inputs(208)));
    layer0_outputs(10164) <= '0';
    layer0_outputs(10165) <= not(inputs(136)) or (inputs(220));
    layer0_outputs(10166) <= (inputs(10)) and (inputs(190));
    layer0_outputs(10167) <= not((inputs(27)) or (inputs(47)));
    layer0_outputs(10168) <= inputs(44);
    layer0_outputs(10169) <= inputs(41);
    layer0_outputs(10170) <= not(inputs(68));
    layer0_outputs(10171) <= inputs(209);
    layer0_outputs(10172) <= (inputs(25)) and not (inputs(44));
    layer0_outputs(10173) <= (inputs(99)) and not (inputs(62));
    layer0_outputs(10174) <= inputs(150);
    layer0_outputs(10175) <= (inputs(79)) xor (inputs(63));
    layer0_outputs(10176) <= not((inputs(154)) xor (inputs(22)));
    layer0_outputs(10177) <= (inputs(12)) or (inputs(50));
    layer0_outputs(10178) <= (inputs(224)) or (inputs(234));
    layer0_outputs(10179) <= (inputs(208)) or (inputs(169));
    layer0_outputs(10180) <= (inputs(219)) and (inputs(205));
    layer0_outputs(10181) <= (inputs(189)) xor (inputs(161));
    layer0_outputs(10182) <= (inputs(236)) or (inputs(237));
    layer0_outputs(10183) <= not(inputs(186)) or (inputs(42));
    layer0_outputs(10184) <= (inputs(183)) and not (inputs(69));
    layer0_outputs(10185) <= inputs(206);
    layer0_outputs(10186) <= not((inputs(12)) or (inputs(15)));
    layer0_outputs(10187) <= not(inputs(245)) or (inputs(221));
    layer0_outputs(10188) <= not(inputs(98));
    layer0_outputs(10189) <= not(inputs(142));
    layer0_outputs(10190) <= not((inputs(34)) or (inputs(61)));
    layer0_outputs(10191) <= inputs(193);
    layer0_outputs(10192) <= inputs(13);
    layer0_outputs(10193) <= not((inputs(247)) or (inputs(40)));
    layer0_outputs(10194) <= (inputs(29)) and not (inputs(170));
    layer0_outputs(10195) <= (inputs(116)) and not (inputs(207));
    layer0_outputs(10196) <= not((inputs(78)) or (inputs(67)));
    layer0_outputs(10197) <= (inputs(198)) and not (inputs(61));
    layer0_outputs(10198) <= '0';
    layer0_outputs(10199) <= (inputs(156)) and not (inputs(106));
    layer0_outputs(10200) <= inputs(8);
    layer0_outputs(10201) <= (inputs(215)) or (inputs(64));
    layer0_outputs(10202) <= inputs(51);
    layer0_outputs(10203) <= not((inputs(164)) or (inputs(179)));
    layer0_outputs(10204) <= (inputs(161)) and not (inputs(56));
    layer0_outputs(10205) <= not(inputs(182));
    layer0_outputs(10206) <= not((inputs(252)) and (inputs(51)));
    layer0_outputs(10207) <= '1';
    layer0_outputs(10208) <= not((inputs(16)) or (inputs(195)));
    layer0_outputs(10209) <= (inputs(190)) and not (inputs(13));
    layer0_outputs(10210) <= inputs(78);
    layer0_outputs(10211) <= not((inputs(234)) xor (inputs(218)));
    layer0_outputs(10212) <= inputs(42);
    layer0_outputs(10213) <= not(inputs(215));
    layer0_outputs(10214) <= not(inputs(32));
    layer0_outputs(10215) <= not((inputs(64)) or (inputs(224)));
    layer0_outputs(10216) <= not((inputs(160)) and (inputs(55)));
    layer0_outputs(10217) <= not((inputs(52)) or (inputs(155)));
    layer0_outputs(10218) <= not((inputs(110)) or (inputs(15)));
    layer0_outputs(10219) <= (inputs(22)) and not (inputs(252));
    layer0_outputs(10220) <= '1';
    layer0_outputs(10221) <= not((inputs(53)) xor (inputs(6)));
    layer0_outputs(10222) <= (inputs(176)) and not (inputs(91));
    layer0_outputs(10223) <= (inputs(208)) or (inputs(36));
    layer0_outputs(10224) <= inputs(23);
    layer0_outputs(10225) <= (inputs(115)) or (inputs(131));
    layer0_outputs(10226) <= (inputs(12)) and not (inputs(86));
    layer0_outputs(10227) <= inputs(209);
    layer0_outputs(10228) <= (inputs(188)) or (inputs(242));
    layer0_outputs(10229) <= not((inputs(92)) or (inputs(112)));
    layer0_outputs(10230) <= (inputs(80)) xor (inputs(242));
    layer0_outputs(10231) <= not(inputs(101)) or (inputs(102));
    layer0_outputs(10232) <= (inputs(202)) and not (inputs(59));
    layer0_outputs(10233) <= not(inputs(57)) or (inputs(129));
    layer0_outputs(10234) <= not(inputs(116)) or (inputs(251));
    layer0_outputs(10235) <= not(inputs(150));
    layer0_outputs(10236) <= not((inputs(87)) or (inputs(121)));
    layer0_outputs(10237) <= not(inputs(177)) or (inputs(49));
    layer0_outputs(10238) <= not((inputs(29)) or (inputs(208)));
    layer0_outputs(10239) <= not((inputs(174)) or (inputs(157)));
    layer1_outputs(0) <= not(layer0_outputs(8768)) or (layer0_outputs(7794));
    layer1_outputs(1) <= not(layer0_outputs(6401)) or (layer0_outputs(5457));
    layer1_outputs(2) <= (layer0_outputs(1339)) and (layer0_outputs(1729));
    layer1_outputs(3) <= (layer0_outputs(7313)) and not (layer0_outputs(2839));
    layer1_outputs(4) <= not(layer0_outputs(4582)) or (layer0_outputs(8833));
    layer1_outputs(5) <= (layer0_outputs(4735)) or (layer0_outputs(9262));
    layer1_outputs(6) <= (layer0_outputs(8831)) and not (layer0_outputs(789));
    layer1_outputs(7) <= (layer0_outputs(9504)) or (layer0_outputs(8137));
    layer1_outputs(8) <= not((layer0_outputs(6605)) and (layer0_outputs(3435)));
    layer1_outputs(9) <= (layer0_outputs(6438)) xor (layer0_outputs(5004));
    layer1_outputs(10) <= not((layer0_outputs(7413)) xor (layer0_outputs(4149)));
    layer1_outputs(11) <= layer0_outputs(1027);
    layer1_outputs(12) <= not((layer0_outputs(4877)) and (layer0_outputs(1907)));
    layer1_outputs(13) <= not(layer0_outputs(2956));
    layer1_outputs(14) <= not((layer0_outputs(2765)) and (layer0_outputs(8475)));
    layer1_outputs(15) <= layer0_outputs(6910);
    layer1_outputs(16) <= not((layer0_outputs(8779)) or (layer0_outputs(9751)));
    layer1_outputs(17) <= not((layer0_outputs(5967)) and (layer0_outputs(8644)));
    layer1_outputs(18) <= layer0_outputs(9044);
    layer1_outputs(19) <= (layer0_outputs(7579)) and not (layer0_outputs(3953));
    layer1_outputs(20) <= not(layer0_outputs(4792));
    layer1_outputs(21) <= not((layer0_outputs(7458)) and (layer0_outputs(187)));
    layer1_outputs(22) <= (layer0_outputs(5621)) and (layer0_outputs(5643));
    layer1_outputs(23) <= (layer0_outputs(8847)) or (layer0_outputs(8870));
    layer1_outputs(24) <= not((layer0_outputs(2974)) or (layer0_outputs(9567)));
    layer1_outputs(25) <= not(layer0_outputs(1546));
    layer1_outputs(26) <= (layer0_outputs(1269)) and (layer0_outputs(1449));
    layer1_outputs(27) <= layer0_outputs(1550);
    layer1_outputs(28) <= not((layer0_outputs(3839)) or (layer0_outputs(4995)));
    layer1_outputs(29) <= not(layer0_outputs(6057));
    layer1_outputs(30) <= not(layer0_outputs(3950));
    layer1_outputs(31) <= (layer0_outputs(5460)) or (layer0_outputs(8103));
    layer1_outputs(32) <= not((layer0_outputs(5217)) xor (layer0_outputs(2404)));
    layer1_outputs(33) <= not(layer0_outputs(2776)) or (layer0_outputs(2607));
    layer1_outputs(34) <= layer0_outputs(5835);
    layer1_outputs(35) <= not(layer0_outputs(3944));
    layer1_outputs(36) <= not(layer0_outputs(10215));
    layer1_outputs(37) <= not(layer0_outputs(9469));
    layer1_outputs(38) <= not(layer0_outputs(7204));
    layer1_outputs(39) <= layer0_outputs(8830);
    layer1_outputs(40) <= (layer0_outputs(3927)) and not (layer0_outputs(226));
    layer1_outputs(41) <= (layer0_outputs(868)) or (layer0_outputs(8808));
    layer1_outputs(42) <= '1';
    layer1_outputs(43) <= (layer0_outputs(8856)) or (layer0_outputs(1833));
    layer1_outputs(44) <= not(layer0_outputs(6424));
    layer1_outputs(45) <= (layer0_outputs(2047)) and not (layer0_outputs(10050));
    layer1_outputs(46) <= not(layer0_outputs(9438));
    layer1_outputs(47) <= not((layer0_outputs(1327)) and (layer0_outputs(3413)));
    layer1_outputs(48) <= not(layer0_outputs(5150));
    layer1_outputs(49) <= layer0_outputs(6291);
    layer1_outputs(50) <= '1';
    layer1_outputs(51) <= (layer0_outputs(9806)) and (layer0_outputs(7551));
    layer1_outputs(52) <= (layer0_outputs(3761)) and (layer0_outputs(8377));
    layer1_outputs(53) <= (layer0_outputs(8864)) or (layer0_outputs(2987));
    layer1_outputs(54) <= layer0_outputs(6307);
    layer1_outputs(55) <= layer0_outputs(111);
    layer1_outputs(56) <= not(layer0_outputs(2222));
    layer1_outputs(57) <= not(layer0_outputs(8092)) or (layer0_outputs(6243));
    layer1_outputs(58) <= not(layer0_outputs(263));
    layer1_outputs(59) <= (layer0_outputs(9331)) or (layer0_outputs(5466));
    layer1_outputs(60) <= layer0_outputs(6474);
    layer1_outputs(61) <= (layer0_outputs(4459)) xor (layer0_outputs(1375));
    layer1_outputs(62) <= not((layer0_outputs(6423)) and (layer0_outputs(3904)));
    layer1_outputs(63) <= (layer0_outputs(6278)) xor (layer0_outputs(4041));
    layer1_outputs(64) <= not(layer0_outputs(6776));
    layer1_outputs(65) <= not(layer0_outputs(6823));
    layer1_outputs(66) <= not((layer0_outputs(3813)) xor (layer0_outputs(2535)));
    layer1_outputs(67) <= not(layer0_outputs(6306)) or (layer0_outputs(7578));
    layer1_outputs(68) <= not(layer0_outputs(2474)) or (layer0_outputs(8489));
    layer1_outputs(69) <= layer0_outputs(9870);
    layer1_outputs(70) <= layer0_outputs(6451);
    layer1_outputs(71) <= layer0_outputs(9351);
    layer1_outputs(72) <= (layer0_outputs(8011)) and (layer0_outputs(6014));
    layer1_outputs(73) <= not((layer0_outputs(3147)) or (layer0_outputs(7307)));
    layer1_outputs(74) <= (layer0_outputs(4907)) and not (layer0_outputs(739));
    layer1_outputs(75) <= (layer0_outputs(7308)) and not (layer0_outputs(7259));
    layer1_outputs(76) <= not(layer0_outputs(6994)) or (layer0_outputs(4831));
    layer1_outputs(77) <= layer0_outputs(7612);
    layer1_outputs(78) <= not((layer0_outputs(1045)) and (layer0_outputs(6713)));
    layer1_outputs(79) <= not(layer0_outputs(4842));
    layer1_outputs(80) <= layer0_outputs(2969);
    layer1_outputs(81) <= not(layer0_outputs(8551)) or (layer0_outputs(7186));
    layer1_outputs(82) <= '0';
    layer1_outputs(83) <= not((layer0_outputs(2336)) or (layer0_outputs(9345)));
    layer1_outputs(84) <= not((layer0_outputs(306)) or (layer0_outputs(8950)));
    layer1_outputs(85) <= not(layer0_outputs(4982));
    layer1_outputs(86) <= layer0_outputs(3835);
    layer1_outputs(87) <= layer0_outputs(8678);
    layer1_outputs(88) <= not((layer0_outputs(8843)) or (layer0_outputs(1402)));
    layer1_outputs(89) <= not(layer0_outputs(802)) or (layer0_outputs(2466));
    layer1_outputs(90) <= (layer0_outputs(1719)) or (layer0_outputs(7192));
    layer1_outputs(91) <= layer0_outputs(833);
    layer1_outputs(92) <= (layer0_outputs(2791)) and (layer0_outputs(3950));
    layer1_outputs(93) <= not(layer0_outputs(6428));
    layer1_outputs(94) <= (layer0_outputs(9199)) and not (layer0_outputs(5791));
    layer1_outputs(95) <= (layer0_outputs(226)) xor (layer0_outputs(313));
    layer1_outputs(96) <= (layer0_outputs(1677)) and not (layer0_outputs(3538));
    layer1_outputs(97) <= (layer0_outputs(9453)) and not (layer0_outputs(6986));
    layer1_outputs(98) <= layer0_outputs(5210);
    layer1_outputs(99) <= (layer0_outputs(4709)) or (layer0_outputs(2986));
    layer1_outputs(100) <= (layer0_outputs(7653)) and (layer0_outputs(1587));
    layer1_outputs(101) <= not(layer0_outputs(1880)) or (layer0_outputs(3693));
    layer1_outputs(102) <= (layer0_outputs(2501)) and not (layer0_outputs(1427));
    layer1_outputs(103) <= not(layer0_outputs(7105));
    layer1_outputs(104) <= layer0_outputs(5483);
    layer1_outputs(105) <= '0';
    layer1_outputs(106) <= (layer0_outputs(8671)) and not (layer0_outputs(9638));
    layer1_outputs(107) <= not(layer0_outputs(3856)) or (layer0_outputs(3493));
    layer1_outputs(108) <= not(layer0_outputs(3183));
    layer1_outputs(109) <= (layer0_outputs(7523)) or (layer0_outputs(3474));
    layer1_outputs(110) <= not((layer0_outputs(5088)) and (layer0_outputs(1327)));
    layer1_outputs(111) <= (layer0_outputs(238)) and (layer0_outputs(1887));
    layer1_outputs(112) <= layer0_outputs(1233);
    layer1_outputs(113) <= layer0_outputs(4118);
    layer1_outputs(114) <= not((layer0_outputs(7761)) or (layer0_outputs(8963)));
    layer1_outputs(115) <= layer0_outputs(2689);
    layer1_outputs(116) <= not((layer0_outputs(1826)) xor (layer0_outputs(5996)));
    layer1_outputs(117) <= not((layer0_outputs(2761)) and (layer0_outputs(7001)));
    layer1_outputs(118) <= (layer0_outputs(2232)) xor (layer0_outputs(2677));
    layer1_outputs(119) <= not(layer0_outputs(6988));
    layer1_outputs(120) <= (layer0_outputs(6831)) and not (layer0_outputs(6646));
    layer1_outputs(121) <= (layer0_outputs(8456)) and not (layer0_outputs(6379));
    layer1_outputs(122) <= not((layer0_outputs(9289)) and (layer0_outputs(6601)));
    layer1_outputs(123) <= (layer0_outputs(8748)) and (layer0_outputs(1024));
    layer1_outputs(124) <= not(layer0_outputs(6426)) or (layer0_outputs(4833));
    layer1_outputs(125) <= not((layer0_outputs(4614)) and (layer0_outputs(8328)));
    layer1_outputs(126) <= layer0_outputs(5494);
    layer1_outputs(127) <= not((layer0_outputs(2669)) xor (layer0_outputs(6259)));
    layer1_outputs(128) <= not(layer0_outputs(4203));
    layer1_outputs(129) <= not(layer0_outputs(1929)) or (layer0_outputs(669));
    layer1_outputs(130) <= '0';
    layer1_outputs(131) <= layer0_outputs(116);
    layer1_outputs(132) <= not((layer0_outputs(3459)) xor (layer0_outputs(8625)));
    layer1_outputs(133) <= layer0_outputs(6760);
    layer1_outputs(134) <= (layer0_outputs(3681)) and (layer0_outputs(9785));
    layer1_outputs(135) <= not(layer0_outputs(7209));
    layer1_outputs(136) <= not((layer0_outputs(6645)) xor (layer0_outputs(9078)));
    layer1_outputs(137) <= layer0_outputs(8503);
    layer1_outputs(138) <= '0';
    layer1_outputs(139) <= not(layer0_outputs(2692));
    layer1_outputs(140) <= layer0_outputs(7436);
    layer1_outputs(141) <= (layer0_outputs(2710)) and (layer0_outputs(7561));
    layer1_outputs(142) <= not(layer0_outputs(8896));
    layer1_outputs(143) <= layer0_outputs(227);
    layer1_outputs(144) <= (layer0_outputs(851)) or (layer0_outputs(9916));
    layer1_outputs(145) <= '1';
    layer1_outputs(146) <= not((layer0_outputs(7852)) or (layer0_outputs(6871)));
    layer1_outputs(147) <= layer0_outputs(6358);
    layer1_outputs(148) <= layer0_outputs(4801);
    layer1_outputs(149) <= (layer0_outputs(7023)) and (layer0_outputs(3826));
    layer1_outputs(150) <= not(layer0_outputs(613));
    layer1_outputs(151) <= layer0_outputs(1682);
    layer1_outputs(152) <= not(layer0_outputs(4760));
    layer1_outputs(153) <= layer0_outputs(584);
    layer1_outputs(154) <= not(layer0_outputs(4563)) or (layer0_outputs(3234));
    layer1_outputs(155) <= layer0_outputs(1979);
    layer1_outputs(156) <= not(layer0_outputs(2420)) or (layer0_outputs(899));
    layer1_outputs(157) <= not(layer0_outputs(5718));
    layer1_outputs(158) <= not((layer0_outputs(1038)) xor (layer0_outputs(7356)));
    layer1_outputs(159) <= not((layer0_outputs(6617)) or (layer0_outputs(4824)));
    layer1_outputs(160) <= layer0_outputs(8450);
    layer1_outputs(161) <= not(layer0_outputs(7118));
    layer1_outputs(162) <= not(layer0_outputs(5606));
    layer1_outputs(163) <= '0';
    layer1_outputs(164) <= not((layer0_outputs(192)) xor (layer0_outputs(9614)));
    layer1_outputs(165) <= (layer0_outputs(10234)) or (layer0_outputs(3136));
    layer1_outputs(166) <= (layer0_outputs(6092)) and not (layer0_outputs(7180));
    layer1_outputs(167) <= layer0_outputs(4253);
    layer1_outputs(168) <= not(layer0_outputs(6913)) or (layer0_outputs(3734));
    layer1_outputs(169) <= not(layer0_outputs(1345));
    layer1_outputs(170) <= not((layer0_outputs(4698)) and (layer0_outputs(9670)));
    layer1_outputs(171) <= layer0_outputs(1994);
    layer1_outputs(172) <= layer0_outputs(6676);
    layer1_outputs(173) <= not(layer0_outputs(6436)) or (layer0_outputs(6101));
    layer1_outputs(174) <= not(layer0_outputs(40)) or (layer0_outputs(4488));
    layer1_outputs(175) <= layer0_outputs(2919);
    layer1_outputs(176) <= not((layer0_outputs(9708)) xor (layer0_outputs(4533)));
    layer1_outputs(177) <= layer0_outputs(4056);
    layer1_outputs(178) <= (layer0_outputs(8106)) or (layer0_outputs(8581));
    layer1_outputs(179) <= (layer0_outputs(1229)) xor (layer0_outputs(2026));
    layer1_outputs(180) <= (layer0_outputs(7029)) or (layer0_outputs(8230));
    layer1_outputs(181) <= '0';
    layer1_outputs(182) <= not((layer0_outputs(9297)) or (layer0_outputs(4856)));
    layer1_outputs(183) <= layer0_outputs(1710);
    layer1_outputs(184) <= layer0_outputs(8606);
    layer1_outputs(185) <= '1';
    layer1_outputs(186) <= not(layer0_outputs(9008)) or (layer0_outputs(9659));
    layer1_outputs(187) <= not((layer0_outputs(5654)) xor (layer0_outputs(377)));
    layer1_outputs(188) <= (layer0_outputs(10080)) and not (layer0_outputs(6063));
    layer1_outputs(189) <= layer0_outputs(1465);
    layer1_outputs(190) <= not(layer0_outputs(7026)) or (layer0_outputs(2790));
    layer1_outputs(191) <= (layer0_outputs(8933)) and not (layer0_outputs(8008));
    layer1_outputs(192) <= (layer0_outputs(5119)) and not (layer0_outputs(7385));
    layer1_outputs(193) <= (layer0_outputs(7430)) and (layer0_outputs(1310));
    layer1_outputs(194) <= not((layer0_outputs(2276)) and (layer0_outputs(6770)));
    layer1_outputs(195) <= not(layer0_outputs(9890));
    layer1_outputs(196) <= (layer0_outputs(4479)) or (layer0_outputs(4234));
    layer1_outputs(197) <= (layer0_outputs(3703)) or (layer0_outputs(439));
    layer1_outputs(198) <= (layer0_outputs(9152)) or (layer0_outputs(5316));
    layer1_outputs(199) <= layer0_outputs(2174);
    layer1_outputs(200) <= '1';
    layer1_outputs(201) <= (layer0_outputs(8096)) or (layer0_outputs(6726));
    layer1_outputs(202) <= layer0_outputs(4567);
    layer1_outputs(203) <= layer0_outputs(3701);
    layer1_outputs(204) <= not(layer0_outputs(6709));
    layer1_outputs(205) <= not(layer0_outputs(7916));
    layer1_outputs(206) <= layer0_outputs(5006);
    layer1_outputs(207) <= (layer0_outputs(1154)) or (layer0_outputs(6239));
    layer1_outputs(208) <= not((layer0_outputs(5349)) and (layer0_outputs(7715)));
    layer1_outputs(209) <= (layer0_outputs(1832)) or (layer0_outputs(1180));
    layer1_outputs(210) <= not(layer0_outputs(4603)) or (layer0_outputs(3162));
    layer1_outputs(211) <= (layer0_outputs(404)) and not (layer0_outputs(6458));
    layer1_outputs(212) <= layer0_outputs(9917);
    layer1_outputs(213) <= '1';
    layer1_outputs(214) <= layer0_outputs(843);
    layer1_outputs(215) <= not((layer0_outputs(7236)) or (layer0_outputs(9169)));
    layer1_outputs(216) <= not(layer0_outputs(3256)) or (layer0_outputs(6716));
    layer1_outputs(217) <= not(layer0_outputs(3734));
    layer1_outputs(218) <= not((layer0_outputs(437)) and (layer0_outputs(3898)));
    layer1_outputs(219) <= (layer0_outputs(4176)) and not (layer0_outputs(1226));
    layer1_outputs(220) <= not((layer0_outputs(3451)) or (layer0_outputs(1869)));
    layer1_outputs(221) <= layer0_outputs(1942);
    layer1_outputs(222) <= (layer0_outputs(1604)) xor (layer0_outputs(4903));
    layer1_outputs(223) <= layer0_outputs(6081);
    layer1_outputs(224) <= (layer0_outputs(3135)) and (layer0_outputs(8286));
    layer1_outputs(225) <= layer0_outputs(8682);
    layer1_outputs(226) <= not(layer0_outputs(9611));
    layer1_outputs(227) <= not((layer0_outputs(6450)) or (layer0_outputs(2420)));
    layer1_outputs(228) <= (layer0_outputs(6687)) and not (layer0_outputs(1373));
    layer1_outputs(229) <= not((layer0_outputs(3411)) and (layer0_outputs(9861)));
    layer1_outputs(230) <= not((layer0_outputs(9196)) or (layer0_outputs(9449)));
    layer1_outputs(231) <= layer0_outputs(2427);
    layer1_outputs(232) <= (layer0_outputs(5681)) or (layer0_outputs(9727));
    layer1_outputs(233) <= layer0_outputs(5134);
    layer1_outputs(234) <= not(layer0_outputs(9566));
    layer1_outputs(235) <= not(layer0_outputs(2713)) or (layer0_outputs(482));
    layer1_outputs(236) <= (layer0_outputs(7899)) and (layer0_outputs(6229));
    layer1_outputs(237) <= not(layer0_outputs(7910));
    layer1_outputs(238) <= not(layer0_outputs(8174));
    layer1_outputs(239) <= not(layer0_outputs(6304)) or (layer0_outputs(9282));
    layer1_outputs(240) <= not(layer0_outputs(3177));
    layer1_outputs(241) <= not(layer0_outputs(6179)) or (layer0_outputs(2031));
    layer1_outputs(242) <= not(layer0_outputs(5328)) or (layer0_outputs(9697));
    layer1_outputs(243) <= layer0_outputs(5381);
    layer1_outputs(244) <= not(layer0_outputs(7204));
    layer1_outputs(245) <= layer0_outputs(5836);
    layer1_outputs(246) <= (layer0_outputs(8167)) and not (layer0_outputs(6213));
    layer1_outputs(247) <= not((layer0_outputs(5828)) or (layer0_outputs(3707)));
    layer1_outputs(248) <= (layer0_outputs(1727)) or (layer0_outputs(10091));
    layer1_outputs(249) <= (layer0_outputs(7140)) and not (layer0_outputs(6951));
    layer1_outputs(250) <= layer0_outputs(5038);
    layer1_outputs(251) <= (layer0_outputs(2777)) and not (layer0_outputs(9475));
    layer1_outputs(252) <= (layer0_outputs(130)) and (layer0_outputs(8211));
    layer1_outputs(253) <= layer0_outputs(1693);
    layer1_outputs(254) <= (layer0_outputs(1866)) and not (layer0_outputs(9232));
    layer1_outputs(255) <= not((layer0_outputs(875)) or (layer0_outputs(2910)));
    layer1_outputs(256) <= not((layer0_outputs(4583)) xor (layer0_outputs(7719)));
    layer1_outputs(257) <= layer0_outputs(6727);
    layer1_outputs(258) <= not((layer0_outputs(863)) and (layer0_outputs(5032)));
    layer1_outputs(259) <= not(layer0_outputs(5310));
    layer1_outputs(260) <= not(layer0_outputs(8165));
    layer1_outputs(261) <= not(layer0_outputs(231));
    layer1_outputs(262) <= layer0_outputs(4855);
    layer1_outputs(263) <= (layer0_outputs(1258)) or (layer0_outputs(6867));
    layer1_outputs(264) <= (layer0_outputs(444)) or (layer0_outputs(4800));
    layer1_outputs(265) <= not((layer0_outputs(4416)) or (layer0_outputs(10196)));
    layer1_outputs(266) <= '1';
    layer1_outputs(267) <= not(layer0_outputs(83));
    layer1_outputs(268) <= '1';
    layer1_outputs(269) <= (layer0_outputs(3917)) xor (layer0_outputs(9220));
    layer1_outputs(270) <= layer0_outputs(72);
    layer1_outputs(271) <= not((layer0_outputs(4827)) and (layer0_outputs(2859)));
    layer1_outputs(272) <= (layer0_outputs(1079)) or (layer0_outputs(1698));
    layer1_outputs(273) <= not((layer0_outputs(5717)) and (layer0_outputs(4884)));
    layer1_outputs(274) <= not((layer0_outputs(2073)) and (layer0_outputs(3162)));
    layer1_outputs(275) <= (layer0_outputs(4859)) xor (layer0_outputs(9274));
    layer1_outputs(276) <= (layer0_outputs(1454)) and not (layer0_outputs(3582));
    layer1_outputs(277) <= (layer0_outputs(6174)) xor (layer0_outputs(1770));
    layer1_outputs(278) <= layer0_outputs(9265);
    layer1_outputs(279) <= not(layer0_outputs(4746)) or (layer0_outputs(5773));
    layer1_outputs(280) <= '1';
    layer1_outputs(281) <= (layer0_outputs(549)) or (layer0_outputs(4836));
    layer1_outputs(282) <= (layer0_outputs(7372)) and not (layer0_outputs(7915));
    layer1_outputs(283) <= layer0_outputs(7334);
    layer1_outputs(284) <= '1';
    layer1_outputs(285) <= layer0_outputs(832);
    layer1_outputs(286) <= (layer0_outputs(1358)) and not (layer0_outputs(10045));
    layer1_outputs(287) <= not(layer0_outputs(8832)) or (layer0_outputs(811));
    layer1_outputs(288) <= not(layer0_outputs(211));
    layer1_outputs(289) <= not(layer0_outputs(8990));
    layer1_outputs(290) <= not(layer0_outputs(2061));
    layer1_outputs(291) <= not((layer0_outputs(5171)) or (layer0_outputs(8869)));
    layer1_outputs(292) <= '1';
    layer1_outputs(293) <= layer0_outputs(8209);
    layer1_outputs(294) <= not(layer0_outputs(7919)) or (layer0_outputs(176));
    layer1_outputs(295) <= not((layer0_outputs(5172)) xor (layer0_outputs(716)));
    layer1_outputs(296) <= (layer0_outputs(4064)) and not (layer0_outputs(3831));
    layer1_outputs(297) <= not((layer0_outputs(640)) and (layer0_outputs(7553)));
    layer1_outputs(298) <= layer0_outputs(6524);
    layer1_outputs(299) <= (layer0_outputs(7157)) and not (layer0_outputs(1482));
    layer1_outputs(300) <= (layer0_outputs(8060)) and (layer0_outputs(8033));
    layer1_outputs(301) <= not(layer0_outputs(5620));
    layer1_outputs(302) <= (layer0_outputs(4885)) xor (layer0_outputs(4088));
    layer1_outputs(303) <= (layer0_outputs(7754)) and not (layer0_outputs(1021));
    layer1_outputs(304) <= (layer0_outputs(10187)) and not (layer0_outputs(5401));
    layer1_outputs(305) <= not(layer0_outputs(2052)) or (layer0_outputs(8070));
    layer1_outputs(306) <= (layer0_outputs(380)) and not (layer0_outputs(2273));
    layer1_outputs(307) <= layer0_outputs(1585);
    layer1_outputs(308) <= '1';
    layer1_outputs(309) <= not(layer0_outputs(5027)) or (layer0_outputs(7961));
    layer1_outputs(310) <= not(layer0_outputs(3212));
    layer1_outputs(311) <= not(layer0_outputs(6250)) or (layer0_outputs(3466));
    layer1_outputs(312) <= not((layer0_outputs(1937)) xor (layer0_outputs(8337)));
    layer1_outputs(313) <= (layer0_outputs(7580)) or (layer0_outputs(8720));
    layer1_outputs(314) <= not(layer0_outputs(1715));
    layer1_outputs(315) <= layer0_outputs(7134);
    layer1_outputs(316) <= (layer0_outputs(5147)) and not (layer0_outputs(8351));
    layer1_outputs(317) <= not(layer0_outputs(1032)) or (layer0_outputs(1732));
    layer1_outputs(318) <= (layer0_outputs(1850)) xor (layer0_outputs(4537));
    layer1_outputs(319) <= (layer0_outputs(881)) or (layer0_outputs(1149));
    layer1_outputs(320) <= not((layer0_outputs(5733)) xor (layer0_outputs(1612)));
    layer1_outputs(321) <= not(layer0_outputs(6126)) or (layer0_outputs(7572));
    layer1_outputs(322) <= layer0_outputs(9526);
    layer1_outputs(323) <= (layer0_outputs(157)) and (layer0_outputs(7256));
    layer1_outputs(324) <= not(layer0_outputs(7974)) or (layer0_outputs(4440));
    layer1_outputs(325) <= layer0_outputs(3673);
    layer1_outputs(326) <= '1';
    layer1_outputs(327) <= not((layer0_outputs(3148)) and (layer0_outputs(2727)));
    layer1_outputs(328) <= not(layer0_outputs(6228)) or (layer0_outputs(7157));
    layer1_outputs(329) <= (layer0_outputs(9739)) and (layer0_outputs(4976));
    layer1_outputs(330) <= layer0_outputs(7313);
    layer1_outputs(331) <= not(layer0_outputs(9599)) or (layer0_outputs(1775));
    layer1_outputs(332) <= layer0_outputs(9733);
    layer1_outputs(333) <= not((layer0_outputs(9333)) xor (layer0_outputs(8137)));
    layer1_outputs(334) <= not((layer0_outputs(4947)) or (layer0_outputs(7742)));
    layer1_outputs(335) <= (layer0_outputs(7607)) xor (layer0_outputs(1527));
    layer1_outputs(336) <= (layer0_outputs(14)) xor (layer0_outputs(4442));
    layer1_outputs(337) <= (layer0_outputs(8102)) xor (layer0_outputs(5226));
    layer1_outputs(338) <= (layer0_outputs(3038)) and (layer0_outputs(1623));
    layer1_outputs(339) <= not(layer0_outputs(254));
    layer1_outputs(340) <= (layer0_outputs(5260)) xor (layer0_outputs(3663));
    layer1_outputs(341) <= (layer0_outputs(1964)) and not (layer0_outputs(2926));
    layer1_outputs(342) <= layer0_outputs(3113);
    layer1_outputs(343) <= not(layer0_outputs(3848));
    layer1_outputs(344) <= not((layer0_outputs(3593)) xor (layer0_outputs(9699)));
    layer1_outputs(345) <= not((layer0_outputs(3405)) or (layer0_outputs(9821)));
    layer1_outputs(346) <= (layer0_outputs(10090)) or (layer0_outputs(1043));
    layer1_outputs(347) <= not(layer0_outputs(5895));
    layer1_outputs(348) <= not(layer0_outputs(7154)) or (layer0_outputs(9515));
    layer1_outputs(349) <= (layer0_outputs(4904)) and (layer0_outputs(336));
    layer1_outputs(350) <= not(layer0_outputs(3757)) or (layer0_outputs(8757));
    layer1_outputs(351) <= (layer0_outputs(1586)) or (layer0_outputs(1373));
    layer1_outputs(352) <= (layer0_outputs(3047)) and (layer0_outputs(2654));
    layer1_outputs(353) <= not(layer0_outputs(8360)) or (layer0_outputs(9855));
    layer1_outputs(354) <= not((layer0_outputs(3395)) or (layer0_outputs(3657)));
    layer1_outputs(355) <= not((layer0_outputs(87)) or (layer0_outputs(8609)));
    layer1_outputs(356) <= layer0_outputs(4994);
    layer1_outputs(357) <= (layer0_outputs(1958)) and not (layer0_outputs(3687));
    layer1_outputs(358) <= not((layer0_outputs(8780)) and (layer0_outputs(6007)));
    layer1_outputs(359) <= (layer0_outputs(8929)) or (layer0_outputs(9568));
    layer1_outputs(360) <= not(layer0_outputs(5685));
    layer1_outputs(361) <= '0';
    layer1_outputs(362) <= (layer0_outputs(317)) and not (layer0_outputs(7363));
    layer1_outputs(363) <= not(layer0_outputs(991));
    layer1_outputs(364) <= not(layer0_outputs(621)) or (layer0_outputs(5561));
    layer1_outputs(365) <= not((layer0_outputs(9927)) and (layer0_outputs(6692)));
    layer1_outputs(366) <= (layer0_outputs(4853)) and not (layer0_outputs(1758));
    layer1_outputs(367) <= not(layer0_outputs(2215)) or (layer0_outputs(7889));
    layer1_outputs(368) <= layer0_outputs(7041);
    layer1_outputs(369) <= not(layer0_outputs(6782));
    layer1_outputs(370) <= layer0_outputs(2592);
    layer1_outputs(371) <= (layer0_outputs(3130)) and (layer0_outputs(2498));
    layer1_outputs(372) <= not(layer0_outputs(8676));
    layer1_outputs(373) <= not((layer0_outputs(2041)) and (layer0_outputs(2631)));
    layer1_outputs(374) <= layer0_outputs(8739);
    layer1_outputs(375) <= (layer0_outputs(9669)) and (layer0_outputs(5920));
    layer1_outputs(376) <= not(layer0_outputs(4031));
    layer1_outputs(377) <= not(layer0_outputs(1235));
    layer1_outputs(378) <= (layer0_outputs(9581)) or (layer0_outputs(64));
    layer1_outputs(379) <= not(layer0_outputs(9716));
    layer1_outputs(380) <= not(layer0_outputs(4047));
    layer1_outputs(381) <= not(layer0_outputs(7799));
    layer1_outputs(382) <= (layer0_outputs(4661)) and not (layer0_outputs(1412));
    layer1_outputs(383) <= not((layer0_outputs(9798)) xor (layer0_outputs(9564)));
    layer1_outputs(384) <= not(layer0_outputs(6801));
    layer1_outputs(385) <= '1';
    layer1_outputs(386) <= not((layer0_outputs(6677)) and (layer0_outputs(1913)));
    layer1_outputs(387) <= (layer0_outputs(1767)) and not (layer0_outputs(9600));
    layer1_outputs(388) <= not((layer0_outputs(6128)) xor (layer0_outputs(5145)));
    layer1_outputs(389) <= not(layer0_outputs(494));
    layer1_outputs(390) <= layer0_outputs(549);
    layer1_outputs(391) <= not(layer0_outputs(4538)) or (layer0_outputs(2860));
    layer1_outputs(392) <= (layer0_outputs(5100)) and not (layer0_outputs(304));
    layer1_outputs(393) <= not((layer0_outputs(4021)) or (layer0_outputs(739)));
    layer1_outputs(394) <= '0';
    layer1_outputs(395) <= layer0_outputs(1810);
    layer1_outputs(396) <= (layer0_outputs(5325)) and not (layer0_outputs(1409));
    layer1_outputs(397) <= not(layer0_outputs(9067)) or (layer0_outputs(2422));
    layer1_outputs(398) <= layer0_outputs(4017);
    layer1_outputs(399) <= not((layer0_outputs(8910)) or (layer0_outputs(4839)));
    layer1_outputs(400) <= not(layer0_outputs(2896));
    layer1_outputs(401) <= (layer0_outputs(2104)) or (layer0_outputs(2377));
    layer1_outputs(402) <= layer0_outputs(5498);
    layer1_outputs(403) <= not(layer0_outputs(1542));
    layer1_outputs(404) <= not(layer0_outputs(4555));
    layer1_outputs(405) <= not(layer0_outputs(557)) or (layer0_outputs(8950));
    layer1_outputs(406) <= not((layer0_outputs(6528)) xor (layer0_outputs(6311)));
    layer1_outputs(407) <= (layer0_outputs(4536)) or (layer0_outputs(4856));
    layer1_outputs(408) <= not(layer0_outputs(3060)) or (layer0_outputs(10225));
    layer1_outputs(409) <= not(layer0_outputs(7847));
    layer1_outputs(410) <= layer0_outputs(7146);
    layer1_outputs(411) <= layer0_outputs(5796);
    layer1_outputs(412) <= not(layer0_outputs(6600));
    layer1_outputs(413) <= not(layer0_outputs(3573)) or (layer0_outputs(3541));
    layer1_outputs(414) <= layer0_outputs(3148);
    layer1_outputs(415) <= (layer0_outputs(1236)) and (layer0_outputs(8902));
    layer1_outputs(416) <= layer0_outputs(9434);
    layer1_outputs(417) <= not(layer0_outputs(8590)) or (layer0_outputs(5115));
    layer1_outputs(418) <= (layer0_outputs(4538)) and (layer0_outputs(8071));
    layer1_outputs(419) <= not(layer0_outputs(1431));
    layer1_outputs(420) <= layer0_outputs(9500);
    layer1_outputs(421) <= not(layer0_outputs(7643));
    layer1_outputs(422) <= (layer0_outputs(10056)) and not (layer0_outputs(4360));
    layer1_outputs(423) <= layer0_outputs(6364);
    layer1_outputs(424) <= layer0_outputs(6887);
    layer1_outputs(425) <= (layer0_outputs(7288)) or (layer0_outputs(6114));
    layer1_outputs(426) <= layer0_outputs(2481);
    layer1_outputs(427) <= not(layer0_outputs(3264));
    layer1_outputs(428) <= layer0_outputs(3050);
    layer1_outputs(429) <= (layer0_outputs(3760)) or (layer0_outputs(8603));
    layer1_outputs(430) <= (layer0_outputs(8108)) and not (layer0_outputs(5624));
    layer1_outputs(431) <= not(layer0_outputs(5636));
    layer1_outputs(432) <= (layer0_outputs(7725)) and not (layer0_outputs(8874));
    layer1_outputs(433) <= (layer0_outputs(5623)) or (layer0_outputs(8497));
    layer1_outputs(434) <= layer0_outputs(9464);
    layer1_outputs(435) <= layer0_outputs(6135);
    layer1_outputs(436) <= not(layer0_outputs(4471));
    layer1_outputs(437) <= not((layer0_outputs(5745)) xor (layer0_outputs(1453)));
    layer1_outputs(438) <= (layer0_outputs(3025)) and not (layer0_outputs(9042));
    layer1_outputs(439) <= not(layer0_outputs(2465)) or (layer0_outputs(7339));
    layer1_outputs(440) <= not((layer0_outputs(5884)) xor (layer0_outputs(3210)));
    layer1_outputs(441) <= not((layer0_outputs(3249)) xor (layer0_outputs(6109)));
    layer1_outputs(442) <= not((layer0_outputs(1782)) xor (layer0_outputs(5842)));
    layer1_outputs(443) <= '0';
    layer1_outputs(444) <= not(layer0_outputs(6284)) or (layer0_outputs(1460));
    layer1_outputs(445) <= not(layer0_outputs(2571)) or (layer0_outputs(2773));
    layer1_outputs(446) <= '1';
    layer1_outputs(447) <= not(layer0_outputs(1609)) or (layer0_outputs(7064));
    layer1_outputs(448) <= not(layer0_outputs(7057));
    layer1_outputs(449) <= (layer0_outputs(6850)) or (layer0_outputs(58));
    layer1_outputs(450) <= not((layer0_outputs(9701)) and (layer0_outputs(9991)));
    layer1_outputs(451) <= (layer0_outputs(6164)) or (layer0_outputs(7656));
    layer1_outputs(452) <= not(layer0_outputs(5413)) or (layer0_outputs(9007));
    layer1_outputs(453) <= (layer0_outputs(5376)) and (layer0_outputs(4659));
    layer1_outputs(454) <= not((layer0_outputs(3228)) and (layer0_outputs(5785)));
    layer1_outputs(455) <= not(layer0_outputs(1527)) or (layer0_outputs(8501));
    layer1_outputs(456) <= not(layer0_outputs(4975)) or (layer0_outputs(3768));
    layer1_outputs(457) <= (layer0_outputs(3224)) or (layer0_outputs(1814));
    layer1_outputs(458) <= not(layer0_outputs(8687));
    layer1_outputs(459) <= not(layer0_outputs(8759));
    layer1_outputs(460) <= '0';
    layer1_outputs(461) <= not(layer0_outputs(8670));
    layer1_outputs(462) <= not((layer0_outputs(8106)) and (layer0_outputs(5444)));
    layer1_outputs(463) <= not(layer0_outputs(3549));
    layer1_outputs(464) <= (layer0_outputs(1543)) and not (layer0_outputs(1624));
    layer1_outputs(465) <= (layer0_outputs(4738)) xor (layer0_outputs(4015));
    layer1_outputs(466) <= not((layer0_outputs(6815)) or (layer0_outputs(9984)));
    layer1_outputs(467) <= not(layer0_outputs(10233)) or (layer0_outputs(5546));
    layer1_outputs(468) <= (layer0_outputs(10059)) and (layer0_outputs(10152));
    layer1_outputs(469) <= not(layer0_outputs(1986));
    layer1_outputs(470) <= not((layer0_outputs(146)) xor (layer0_outputs(5986)));
    layer1_outputs(471) <= (layer0_outputs(3173)) and (layer0_outputs(7603));
    layer1_outputs(472) <= (layer0_outputs(9999)) xor (layer0_outputs(5685));
    layer1_outputs(473) <= (layer0_outputs(9731)) and (layer0_outputs(4415));
    layer1_outputs(474) <= not((layer0_outputs(2253)) xor (layer0_outputs(3774)));
    layer1_outputs(475) <= layer0_outputs(7530);
    layer1_outputs(476) <= not(layer0_outputs(7291));
    layer1_outputs(477) <= not((layer0_outputs(2991)) xor (layer0_outputs(3144)));
    layer1_outputs(478) <= (layer0_outputs(7677)) and not (layer0_outputs(8037));
    layer1_outputs(479) <= not(layer0_outputs(520)) or (layer0_outputs(8368));
    layer1_outputs(480) <= layer0_outputs(1753);
    layer1_outputs(481) <= not(layer0_outputs(6761));
    layer1_outputs(482) <= not(layer0_outputs(1947)) or (layer0_outputs(1501));
    layer1_outputs(483) <= (layer0_outputs(4017)) and not (layer0_outputs(1885));
    layer1_outputs(484) <= (layer0_outputs(3624)) and (layer0_outputs(2778));
    layer1_outputs(485) <= not(layer0_outputs(9981));
    layer1_outputs(486) <= layer0_outputs(2155);
    layer1_outputs(487) <= not(layer0_outputs(9373)) or (layer0_outputs(8352));
    layer1_outputs(488) <= not(layer0_outputs(7268));
    layer1_outputs(489) <= (layer0_outputs(2113)) and not (layer0_outputs(6201));
    layer1_outputs(490) <= (layer0_outputs(3494)) and not (layer0_outputs(5878));
    layer1_outputs(491) <= layer0_outputs(4016);
    layer1_outputs(492) <= layer0_outputs(5373);
    layer1_outputs(493) <= layer0_outputs(1623);
    layer1_outputs(494) <= not(layer0_outputs(3043));
    layer1_outputs(495) <= not((layer0_outputs(5126)) or (layer0_outputs(2272)));
    layer1_outputs(496) <= layer0_outputs(733);
    layer1_outputs(497) <= layer0_outputs(3699);
    layer1_outputs(498) <= layer0_outputs(1839);
    layer1_outputs(499) <= (layer0_outputs(4287)) and not (layer0_outputs(5865));
    layer1_outputs(500) <= layer0_outputs(9099);
    layer1_outputs(501) <= (layer0_outputs(4666)) and not (layer0_outputs(1382));
    layer1_outputs(502) <= not(layer0_outputs(4154)) or (layer0_outputs(9184));
    layer1_outputs(503) <= not(layer0_outputs(2409));
    layer1_outputs(504) <= (layer0_outputs(7678)) or (layer0_outputs(1588));
    layer1_outputs(505) <= (layer0_outputs(9962)) and (layer0_outputs(4540));
    layer1_outputs(506) <= not(layer0_outputs(8517));
    layer1_outputs(507) <= layer0_outputs(4737);
    layer1_outputs(508) <= layer0_outputs(1917);
    layer1_outputs(509) <= layer0_outputs(300);
    layer1_outputs(510) <= (layer0_outputs(5540)) xor (layer0_outputs(5465));
    layer1_outputs(511) <= (layer0_outputs(7943)) xor (layer0_outputs(7636));
    layer1_outputs(512) <= (layer0_outputs(7844)) and (layer0_outputs(1861));
    layer1_outputs(513) <= layer0_outputs(8821);
    layer1_outputs(514) <= not((layer0_outputs(4292)) xor (layer0_outputs(8260)));
    layer1_outputs(515) <= not(layer0_outputs(2098));
    layer1_outputs(516) <= not(layer0_outputs(5888)) or (layer0_outputs(2360));
    layer1_outputs(517) <= (layer0_outputs(2833)) and not (layer0_outputs(4657));
    layer1_outputs(518) <= not(layer0_outputs(8205));
    layer1_outputs(519) <= (layer0_outputs(9722)) and not (layer0_outputs(6902));
    layer1_outputs(520) <= '0';
    layer1_outputs(521) <= not(layer0_outputs(9315)) or (layer0_outputs(2485));
    layer1_outputs(522) <= not(layer0_outputs(633));
    layer1_outputs(523) <= (layer0_outputs(6993)) and not (layer0_outputs(6955));
    layer1_outputs(524) <= not(layer0_outputs(1744)) or (layer0_outputs(7751));
    layer1_outputs(525) <= not((layer0_outputs(186)) and (layer0_outputs(7458)));
    layer1_outputs(526) <= layer0_outputs(4140);
    layer1_outputs(527) <= not((layer0_outputs(2268)) and (layer0_outputs(2108)));
    layer1_outputs(528) <= not(layer0_outputs(6237));
    layer1_outputs(529) <= not((layer0_outputs(3525)) xor (layer0_outputs(3596)));
    layer1_outputs(530) <= not((layer0_outputs(7709)) xor (layer0_outputs(7023)));
    layer1_outputs(531) <= layer0_outputs(3905);
    layer1_outputs(532) <= (layer0_outputs(2647)) and not (layer0_outputs(8549));
    layer1_outputs(533) <= '1';
    layer1_outputs(534) <= layer0_outputs(3154);
    layer1_outputs(535) <= not(layer0_outputs(8483));
    layer1_outputs(536) <= '1';
    layer1_outputs(537) <= layer0_outputs(5082);
    layer1_outputs(538) <= layer0_outputs(9905);
    layer1_outputs(539) <= layer0_outputs(6412);
    layer1_outputs(540) <= layer0_outputs(288);
    layer1_outputs(541) <= not(layer0_outputs(3155));
    layer1_outputs(542) <= not(layer0_outputs(8413));
    layer1_outputs(543) <= (layer0_outputs(8)) and (layer0_outputs(8493));
    layer1_outputs(544) <= layer0_outputs(6398);
    layer1_outputs(545) <= not(layer0_outputs(3563));
    layer1_outputs(546) <= not(layer0_outputs(5398));
    layer1_outputs(547) <= not((layer0_outputs(5417)) xor (layer0_outputs(6515)));
    layer1_outputs(548) <= not(layer0_outputs(8422));
    layer1_outputs(549) <= not((layer0_outputs(6808)) or (layer0_outputs(7852)));
    layer1_outputs(550) <= not(layer0_outputs(5469));
    layer1_outputs(551) <= (layer0_outputs(9802)) or (layer0_outputs(4300));
    layer1_outputs(552) <= not(layer0_outputs(7134)) or (layer0_outputs(8424));
    layer1_outputs(553) <= (layer0_outputs(1897)) xor (layer0_outputs(10121));
    layer1_outputs(554) <= layer0_outputs(1872);
    layer1_outputs(555) <= layer0_outputs(9956);
    layer1_outputs(556) <= layer0_outputs(9887);
    layer1_outputs(557) <= layer0_outputs(8279);
    layer1_outputs(558) <= (layer0_outputs(8823)) and not (layer0_outputs(2237));
    layer1_outputs(559) <= layer0_outputs(3940);
    layer1_outputs(560) <= layer0_outputs(5073);
    layer1_outputs(561) <= (layer0_outputs(7851)) and not (layer0_outputs(3490));
    layer1_outputs(562) <= layer0_outputs(9856);
    layer1_outputs(563) <= (layer0_outputs(2618)) and (layer0_outputs(8198));
    layer1_outputs(564) <= not(layer0_outputs(5018));
    layer1_outputs(565) <= not(layer0_outputs(7728));
    layer1_outputs(566) <= layer0_outputs(2039);
    layer1_outputs(567) <= layer0_outputs(2223);
    layer1_outputs(568) <= (layer0_outputs(6094)) or (layer0_outputs(6088));
    layer1_outputs(569) <= layer0_outputs(3569);
    layer1_outputs(570) <= (layer0_outputs(5246)) and (layer0_outputs(1935));
    layer1_outputs(571) <= not(layer0_outputs(1761));
    layer1_outputs(572) <= not(layer0_outputs(6099));
    layer1_outputs(573) <= layer0_outputs(5431);
    layer1_outputs(574) <= not((layer0_outputs(7391)) or (layer0_outputs(9988)));
    layer1_outputs(575) <= not(layer0_outputs(2037));
    layer1_outputs(576) <= (layer0_outputs(9013)) xor (layer0_outputs(7857));
    layer1_outputs(577) <= layer0_outputs(4766);
    layer1_outputs(578) <= (layer0_outputs(7682)) and (layer0_outputs(8170));
    layer1_outputs(579) <= (layer0_outputs(4793)) xor (layer0_outputs(2327));
    layer1_outputs(580) <= not(layer0_outputs(604)) or (layer0_outputs(4898));
    layer1_outputs(581) <= not(layer0_outputs(8254));
    layer1_outputs(582) <= layer0_outputs(9426);
    layer1_outputs(583) <= layer0_outputs(6315);
    layer1_outputs(584) <= layer0_outputs(6242);
    layer1_outputs(585) <= not(layer0_outputs(214));
    layer1_outputs(586) <= not(layer0_outputs(1601));
    layer1_outputs(587) <= (layer0_outputs(8248)) and not (layer0_outputs(6479));
    layer1_outputs(588) <= (layer0_outputs(4301)) xor (layer0_outputs(6637));
    layer1_outputs(589) <= not(layer0_outputs(348));
    layer1_outputs(590) <= layer0_outputs(7343);
    layer1_outputs(591) <= (layer0_outputs(5512)) and not (layer0_outputs(8425));
    layer1_outputs(592) <= layer0_outputs(9492);
    layer1_outputs(593) <= (layer0_outputs(7407)) and not (layer0_outputs(834));
    layer1_outputs(594) <= not(layer0_outputs(9180));
    layer1_outputs(595) <= (layer0_outputs(3027)) or (layer0_outputs(3032));
    layer1_outputs(596) <= (layer0_outputs(8823)) and not (layer0_outputs(778));
    layer1_outputs(597) <= (layer0_outputs(6478)) or (layer0_outputs(3968));
    layer1_outputs(598) <= layer0_outputs(764);
    layer1_outputs(599) <= not(layer0_outputs(3610)) or (layer0_outputs(2711));
    layer1_outputs(600) <= (layer0_outputs(8989)) and not (layer0_outputs(5280));
    layer1_outputs(601) <= not(layer0_outputs(3463));
    layer1_outputs(602) <= not(layer0_outputs(152));
    layer1_outputs(603) <= (layer0_outputs(1090)) and not (layer0_outputs(4697));
    layer1_outputs(604) <= not(layer0_outputs(8688));
    layer1_outputs(605) <= (layer0_outputs(4452)) or (layer0_outputs(9732));
    layer1_outputs(606) <= not(layer0_outputs(6164));
    layer1_outputs(607) <= not(layer0_outputs(815));
    layer1_outputs(608) <= not((layer0_outputs(4435)) and (layer0_outputs(8286)));
    layer1_outputs(609) <= (layer0_outputs(5626)) and (layer0_outputs(394));
    layer1_outputs(610) <= not(layer0_outputs(8013)) or (layer0_outputs(1036));
    layer1_outputs(611) <= (layer0_outputs(8225)) and not (layer0_outputs(2478));
    layer1_outputs(612) <= layer0_outputs(167);
    layer1_outputs(613) <= not((layer0_outputs(2606)) and (layer0_outputs(7461)));
    layer1_outputs(614) <= not((layer0_outputs(164)) or (layer0_outputs(2438)));
    layer1_outputs(615) <= not(layer0_outputs(7879));
    layer1_outputs(616) <= not(layer0_outputs(243));
    layer1_outputs(617) <= (layer0_outputs(1253)) and (layer0_outputs(9279));
    layer1_outputs(618) <= not((layer0_outputs(5497)) xor (layer0_outputs(1243)));
    layer1_outputs(619) <= not(layer0_outputs(8813)) or (layer0_outputs(5284));
    layer1_outputs(620) <= not(layer0_outputs(8515));
    layer1_outputs(621) <= (layer0_outputs(2544)) and not (layer0_outputs(3135));
    layer1_outputs(622) <= not(layer0_outputs(3503));
    layer1_outputs(623) <= layer0_outputs(9261);
    layer1_outputs(624) <= (layer0_outputs(3161)) or (layer0_outputs(9221));
    layer1_outputs(625) <= (layer0_outputs(1073)) and not (layer0_outputs(9264));
    layer1_outputs(626) <= not((layer0_outputs(923)) and (layer0_outputs(9182)));
    layer1_outputs(627) <= (layer0_outputs(9804)) and not (layer0_outputs(238));
    layer1_outputs(628) <= not(layer0_outputs(1563)) or (layer0_outputs(9821));
    layer1_outputs(629) <= layer0_outputs(8541);
    layer1_outputs(630) <= (layer0_outputs(9731)) xor (layer0_outputs(3737));
    layer1_outputs(631) <= layer0_outputs(8521);
    layer1_outputs(632) <= layer0_outputs(5663);
    layer1_outputs(633) <= layer0_outputs(6452);
    layer1_outputs(634) <= not(layer0_outputs(8899)) or (layer0_outputs(2264));
    layer1_outputs(635) <= layer0_outputs(6578);
    layer1_outputs(636) <= not(layer0_outputs(38)) or (layer0_outputs(2892));
    layer1_outputs(637) <= (layer0_outputs(5505)) and (layer0_outputs(4644));
    layer1_outputs(638) <= (layer0_outputs(4473)) and not (layer0_outputs(7911));
    layer1_outputs(639) <= '1';
    layer1_outputs(640) <= not(layer0_outputs(8676)) or (layer0_outputs(9452));
    layer1_outputs(641) <= not(layer0_outputs(2849));
    layer1_outputs(642) <= (layer0_outputs(9607)) and (layer0_outputs(917));
    layer1_outputs(643) <= not(layer0_outputs(782));
    layer1_outputs(644) <= (layer0_outputs(1032)) and (layer0_outputs(8561));
    layer1_outputs(645) <= layer0_outputs(2745);
    layer1_outputs(646) <= layer0_outputs(10028);
    layer1_outputs(647) <= layer0_outputs(6212);
    layer1_outputs(648) <= layer0_outputs(9198);
    layer1_outputs(649) <= not(layer0_outputs(6694));
    layer1_outputs(650) <= '0';
    layer1_outputs(651) <= (layer0_outputs(7579)) and not (layer0_outputs(2309));
    layer1_outputs(652) <= not(layer0_outputs(797));
    layer1_outputs(653) <= not(layer0_outputs(6059));
    layer1_outputs(654) <= not((layer0_outputs(8640)) or (layer0_outputs(9075)));
    layer1_outputs(655) <= layer0_outputs(4027);
    layer1_outputs(656) <= layer0_outputs(9903);
    layer1_outputs(657) <= (layer0_outputs(9931)) and not (layer0_outputs(3384));
    layer1_outputs(658) <= layer0_outputs(7507);
    layer1_outputs(659) <= not((layer0_outputs(8467)) or (layer0_outputs(4272)));
    layer1_outputs(660) <= not(layer0_outputs(6051)) or (layer0_outputs(7980));
    layer1_outputs(661) <= not(layer0_outputs(7160));
    layer1_outputs(662) <= layer0_outputs(751);
    layer1_outputs(663) <= not((layer0_outputs(26)) xor (layer0_outputs(8878)));
    layer1_outputs(664) <= layer0_outputs(6649);
    layer1_outputs(665) <= '0';
    layer1_outputs(666) <= not(layer0_outputs(1644));
    layer1_outputs(667) <= not((layer0_outputs(524)) or (layer0_outputs(5626)));
    layer1_outputs(668) <= (layer0_outputs(8064)) and not (layer0_outputs(8227));
    layer1_outputs(669) <= (layer0_outputs(3583)) and not (layer0_outputs(4081));
    layer1_outputs(670) <= not(layer0_outputs(6127));
    layer1_outputs(671) <= layer0_outputs(31);
    layer1_outputs(672) <= not(layer0_outputs(7662));
    layer1_outputs(673) <= not(layer0_outputs(9107)) or (layer0_outputs(9480));
    layer1_outputs(674) <= not(layer0_outputs(9679)) or (layer0_outputs(9187));
    layer1_outputs(675) <= not(layer0_outputs(7240)) or (layer0_outputs(1738));
    layer1_outputs(676) <= not((layer0_outputs(8981)) xor (layer0_outputs(8242)));
    layer1_outputs(677) <= layer0_outputs(3959);
    layer1_outputs(678) <= (layer0_outputs(4133)) xor (layer0_outputs(9414));
    layer1_outputs(679) <= not(layer0_outputs(2521)) or (layer0_outputs(4913));
    layer1_outputs(680) <= '1';
    layer1_outputs(681) <= (layer0_outputs(6076)) and (layer0_outputs(7823));
    layer1_outputs(682) <= layer0_outputs(5241);
    layer1_outputs(683) <= not(layer0_outputs(7887));
    layer1_outputs(684) <= not(layer0_outputs(7650));
    layer1_outputs(685) <= (layer0_outputs(1503)) and not (layer0_outputs(6222));
    layer1_outputs(686) <= layer0_outputs(10124);
    layer1_outputs(687) <= not(layer0_outputs(4082));
    layer1_outputs(688) <= not(layer0_outputs(4844)) or (layer0_outputs(4966));
    layer1_outputs(689) <= not(layer0_outputs(1059));
    layer1_outputs(690) <= (layer0_outputs(5730)) and not (layer0_outputs(5595));
    layer1_outputs(691) <= (layer0_outputs(1553)) and not (layer0_outputs(8799));
    layer1_outputs(692) <= not(layer0_outputs(1975));
    layer1_outputs(693) <= (layer0_outputs(6870)) xor (layer0_outputs(2432));
    layer1_outputs(694) <= layer0_outputs(4209);
    layer1_outputs(695) <= not(layer0_outputs(9615)) or (layer0_outputs(3297));
    layer1_outputs(696) <= layer0_outputs(2338);
    layer1_outputs(697) <= not((layer0_outputs(6488)) or (layer0_outputs(8343)));
    layer1_outputs(698) <= not(layer0_outputs(6506));
    layer1_outputs(699) <= (layer0_outputs(8862)) xor (layer0_outputs(3191));
    layer1_outputs(700) <= not(layer0_outputs(1169)) or (layer0_outputs(7478));
    layer1_outputs(701) <= layer0_outputs(3404);
    layer1_outputs(702) <= not(layer0_outputs(5482));
    layer1_outputs(703) <= (layer0_outputs(6204)) and not (layer0_outputs(492));
    layer1_outputs(704) <= not(layer0_outputs(7228));
    layer1_outputs(705) <= not((layer0_outputs(4815)) and (layer0_outputs(1312)));
    layer1_outputs(706) <= not((layer0_outputs(4957)) and (layer0_outputs(7429)));
    layer1_outputs(707) <= not(layer0_outputs(6722));
    layer1_outputs(708) <= not((layer0_outputs(5504)) and (layer0_outputs(4235)));
    layer1_outputs(709) <= layer0_outputs(4988);
    layer1_outputs(710) <= (layer0_outputs(10181)) and not (layer0_outputs(4984));
    layer1_outputs(711) <= (layer0_outputs(6674)) or (layer0_outputs(7279));
    layer1_outputs(712) <= not(layer0_outputs(3433)) or (layer0_outputs(9357));
    layer1_outputs(713) <= (layer0_outputs(5029)) and not (layer0_outputs(7755));
    layer1_outputs(714) <= (layer0_outputs(3584)) and (layer0_outputs(3763));
    layer1_outputs(715) <= not(layer0_outputs(3705));
    layer1_outputs(716) <= not(layer0_outputs(1507));
    layer1_outputs(717) <= (layer0_outputs(776)) xor (layer0_outputs(4104));
    layer1_outputs(718) <= layer0_outputs(4579);
    layer1_outputs(719) <= layer0_outputs(6226);
    layer1_outputs(720) <= (layer0_outputs(7251)) and (layer0_outputs(8405));
    layer1_outputs(721) <= '1';
    layer1_outputs(722) <= layer0_outputs(4933);
    layer1_outputs(723) <= layer0_outputs(4785);
    layer1_outputs(724) <= not(layer0_outputs(1816)) or (layer0_outputs(8114));
    layer1_outputs(725) <= not(layer0_outputs(7181));
    layer1_outputs(726) <= (layer0_outputs(5267)) xor (layer0_outputs(5676));
    layer1_outputs(727) <= not(layer0_outputs(4366));
    layer1_outputs(728) <= not(layer0_outputs(6188)) or (layer0_outputs(2289));
    layer1_outputs(729) <= not(layer0_outputs(1342));
    layer1_outputs(730) <= (layer0_outputs(6562)) and not (layer0_outputs(8340));
    layer1_outputs(731) <= not(layer0_outputs(5169));
    layer1_outputs(732) <= (layer0_outputs(7484)) xor (layer0_outputs(4539));
    layer1_outputs(733) <= not(layer0_outputs(3408));
    layer1_outputs(734) <= not(layer0_outputs(883));
    layer1_outputs(735) <= layer0_outputs(7740);
    layer1_outputs(736) <= not(layer0_outputs(3506));
    layer1_outputs(737) <= layer0_outputs(109);
    layer1_outputs(738) <= not(layer0_outputs(10193)) or (layer0_outputs(10102));
    layer1_outputs(739) <= not((layer0_outputs(1213)) or (layer0_outputs(5757)));
    layer1_outputs(740) <= (layer0_outputs(460)) and not (layer0_outputs(699));
    layer1_outputs(741) <= (layer0_outputs(5980)) xor (layer0_outputs(2546));
    layer1_outputs(742) <= not(layer0_outputs(1832));
    layer1_outputs(743) <= (layer0_outputs(6108)) and not (layer0_outputs(4350));
    layer1_outputs(744) <= (layer0_outputs(4423)) and not (layer0_outputs(5550));
    layer1_outputs(745) <= layer0_outputs(2172);
    layer1_outputs(746) <= (layer0_outputs(4260)) and (layer0_outputs(511));
    layer1_outputs(747) <= layer0_outputs(4022);
    layer1_outputs(748) <= not((layer0_outputs(4915)) and (layer0_outputs(6798)));
    layer1_outputs(749) <= not(layer0_outputs(9024));
    layer1_outputs(750) <= not(layer0_outputs(4797));
    layer1_outputs(751) <= layer0_outputs(2903);
    layer1_outputs(752) <= not(layer0_outputs(10118));
    layer1_outputs(753) <= not((layer0_outputs(6612)) xor (layer0_outputs(9603)));
    layer1_outputs(754) <= layer0_outputs(5087);
    layer1_outputs(755) <= not(layer0_outputs(8876));
    layer1_outputs(756) <= '0';
    layer1_outputs(757) <= (layer0_outputs(2279)) xor (layer0_outputs(2271));
    layer1_outputs(758) <= layer0_outputs(7116);
    layer1_outputs(759) <= (layer0_outputs(5552)) and not (layer0_outputs(1431));
    layer1_outputs(760) <= not(layer0_outputs(726));
    layer1_outputs(761) <= not(layer0_outputs(5391));
    layer1_outputs(762) <= (layer0_outputs(7407)) or (layer0_outputs(9653));
    layer1_outputs(763) <= not((layer0_outputs(6833)) and (layer0_outputs(2448)));
    layer1_outputs(764) <= '0';
    layer1_outputs(765) <= not((layer0_outputs(9368)) and (layer0_outputs(2678)));
    layer1_outputs(766) <= not(layer0_outputs(8506));
    layer1_outputs(767) <= (layer0_outputs(3454)) and (layer0_outputs(2153));
    layer1_outputs(768) <= not((layer0_outputs(297)) xor (layer0_outputs(7224)));
    layer1_outputs(769) <= layer0_outputs(4408);
    layer1_outputs(770) <= layer0_outputs(4292);
    layer1_outputs(771) <= '1';
    layer1_outputs(772) <= not((layer0_outputs(988)) and (layer0_outputs(7768)));
    layer1_outputs(773) <= not(layer0_outputs(2381));
    layer1_outputs(774) <= not((layer0_outputs(938)) or (layer0_outputs(7200)));
    layer1_outputs(775) <= not(layer0_outputs(5158));
    layer1_outputs(776) <= layer0_outputs(8152);
    layer1_outputs(777) <= not(layer0_outputs(2744));
    layer1_outputs(778) <= (layer0_outputs(9627)) and (layer0_outputs(8749));
    layer1_outputs(779) <= not((layer0_outputs(6014)) xor (layer0_outputs(2766)));
    layer1_outputs(780) <= layer0_outputs(4753);
    layer1_outputs(781) <= (layer0_outputs(6423)) xor (layer0_outputs(4086));
    layer1_outputs(782) <= not(layer0_outputs(2218));
    layer1_outputs(783) <= (layer0_outputs(1916)) and not (layer0_outputs(9778));
    layer1_outputs(784) <= layer0_outputs(8249);
    layer1_outputs(785) <= (layer0_outputs(2597)) xor (layer0_outputs(6490));
    layer1_outputs(786) <= not(layer0_outputs(4882));
    layer1_outputs(787) <= not((layer0_outputs(2873)) or (layer0_outputs(4228)));
    layer1_outputs(788) <= not(layer0_outputs(4317));
    layer1_outputs(789) <= layer0_outputs(9490);
    layer1_outputs(790) <= layer0_outputs(66);
    layer1_outputs(791) <= (layer0_outputs(3000)) xor (layer0_outputs(5131));
    layer1_outputs(792) <= not(layer0_outputs(5395)) or (layer0_outputs(2259));
    layer1_outputs(793) <= not(layer0_outputs(1930));
    layer1_outputs(794) <= not((layer0_outputs(8962)) and (layer0_outputs(9184)));
    layer1_outputs(795) <= layer0_outputs(4870);
    layer1_outputs(796) <= layer0_outputs(8353);
    layer1_outputs(797) <= (layer0_outputs(1703)) or (layer0_outputs(6443));
    layer1_outputs(798) <= not((layer0_outputs(8495)) or (layer0_outputs(3739)));
    layer1_outputs(799) <= not(layer0_outputs(6185));
    layer1_outputs(800) <= not(layer0_outputs(2062));
    layer1_outputs(801) <= (layer0_outputs(5772)) and (layer0_outputs(6200));
    layer1_outputs(802) <= layer0_outputs(5999);
    layer1_outputs(803) <= not(layer0_outputs(4747));
    layer1_outputs(804) <= layer0_outputs(6420);
    layer1_outputs(805) <= (layer0_outputs(4071)) and not (layer0_outputs(5538));
    layer1_outputs(806) <= not(layer0_outputs(1401));
    layer1_outputs(807) <= layer0_outputs(9703);
    layer1_outputs(808) <= not(layer0_outputs(1439));
    layer1_outputs(809) <= not(layer0_outputs(6924));
    layer1_outputs(810) <= (layer0_outputs(6685)) and not (layer0_outputs(8593));
    layer1_outputs(811) <= not(layer0_outputs(7855)) or (layer0_outputs(5067));
    layer1_outputs(812) <= layer0_outputs(6296);
    layer1_outputs(813) <= not(layer0_outputs(2545));
    layer1_outputs(814) <= (layer0_outputs(6349)) and (layer0_outputs(4888));
    layer1_outputs(815) <= not(layer0_outputs(1209));
    layer1_outputs(816) <= not(layer0_outputs(681)) or (layer0_outputs(3616));
    layer1_outputs(817) <= (layer0_outputs(273)) and (layer0_outputs(6926));
    layer1_outputs(818) <= layer0_outputs(7962);
    layer1_outputs(819) <= '1';
    layer1_outputs(820) <= layer0_outputs(2688);
    layer1_outputs(821) <= not((layer0_outputs(4569)) and (layer0_outputs(5896)));
    layer1_outputs(822) <= layer0_outputs(8680);
    layer1_outputs(823) <= not(layer0_outputs(2459));
    layer1_outputs(824) <= not(layer0_outputs(8310)) or (layer0_outputs(1575));
    layer1_outputs(825) <= '0';
    layer1_outputs(826) <= not(layer0_outputs(3217));
    layer1_outputs(827) <= layer0_outputs(5996);
    layer1_outputs(828) <= not(layer0_outputs(9877));
    layer1_outputs(829) <= layer0_outputs(4631);
    layer1_outputs(830) <= not((layer0_outputs(8390)) and (layer0_outputs(8840)));
    layer1_outputs(831) <= layer0_outputs(6417);
    layer1_outputs(832) <= not((layer0_outputs(8032)) xor (layer0_outputs(8529)));
    layer1_outputs(833) <= (layer0_outputs(7141)) and not (layer0_outputs(8113));
    layer1_outputs(834) <= not(layer0_outputs(6460));
    layer1_outputs(835) <= (layer0_outputs(10163)) and not (layer0_outputs(10092));
    layer1_outputs(836) <= (layer0_outputs(8281)) and not (layer0_outputs(7565));
    layer1_outputs(837) <= layer0_outputs(9159);
    layer1_outputs(838) <= layer0_outputs(6396);
    layer1_outputs(839) <= not(layer0_outputs(268));
    layer1_outputs(840) <= '1';
    layer1_outputs(841) <= not(layer0_outputs(2294));
    layer1_outputs(842) <= not(layer0_outputs(3774)) or (layer0_outputs(570));
    layer1_outputs(843) <= (layer0_outputs(7598)) and not (layer0_outputs(7557));
    layer1_outputs(844) <= not(layer0_outputs(3488)) or (layer0_outputs(725));
    layer1_outputs(845) <= layer0_outputs(8616);
    layer1_outputs(846) <= not(layer0_outputs(5468));
    layer1_outputs(847) <= layer0_outputs(7609);
    layer1_outputs(848) <= not(layer0_outputs(3009));
    layer1_outputs(849) <= layer0_outputs(4548);
    layer1_outputs(850) <= (layer0_outputs(10152)) and not (layer0_outputs(733));
    layer1_outputs(851) <= (layer0_outputs(7706)) xor (layer0_outputs(9757));
    layer1_outputs(852) <= (layer0_outputs(7477)) and not (layer0_outputs(2230));
    layer1_outputs(853) <= not(layer0_outputs(4159)) or (layer0_outputs(2249));
    layer1_outputs(854) <= (layer0_outputs(6018)) xor (layer0_outputs(607));
    layer1_outputs(855) <= (layer0_outputs(10101)) or (layer0_outputs(7355));
    layer1_outputs(856) <= (layer0_outputs(9879)) and not (layer0_outputs(6232));
    layer1_outputs(857) <= (layer0_outputs(10239)) xor (layer0_outputs(5613));
    layer1_outputs(858) <= (layer0_outputs(1529)) or (layer0_outputs(7287));
    layer1_outputs(859) <= not(layer0_outputs(4268)) or (layer0_outputs(2633));
    layer1_outputs(860) <= (layer0_outputs(3)) or (layer0_outputs(6525));
    layer1_outputs(861) <= not(layer0_outputs(6513));
    layer1_outputs(862) <= (layer0_outputs(9112)) and (layer0_outputs(7373));
    layer1_outputs(863) <= not((layer0_outputs(6431)) xor (layer0_outputs(4481)));
    layer1_outputs(864) <= not(layer0_outputs(9942));
    layer1_outputs(865) <= layer0_outputs(6400);
    layer1_outputs(866) <= (layer0_outputs(2111)) and not (layer0_outputs(8594));
    layer1_outputs(867) <= not(layer0_outputs(9137));
    layer1_outputs(868) <= (layer0_outputs(980)) or (layer0_outputs(1735));
    layer1_outputs(869) <= (layer0_outputs(4212)) and not (layer0_outputs(8372));
    layer1_outputs(870) <= not((layer0_outputs(2293)) xor (layer0_outputs(2183)));
    layer1_outputs(871) <= not(layer0_outputs(2825));
    layer1_outputs(872) <= layer0_outputs(9118);
    layer1_outputs(873) <= layer0_outputs(7901);
    layer1_outputs(874) <= '0';
    layer1_outputs(875) <= (layer0_outputs(363)) and not (layer0_outputs(87));
    layer1_outputs(876) <= (layer0_outputs(7147)) and (layer0_outputs(2856));
    layer1_outputs(877) <= layer0_outputs(6832);
    layer1_outputs(878) <= layer0_outputs(6058);
    layer1_outputs(879) <= not(layer0_outputs(4565));
    layer1_outputs(880) <= layer0_outputs(5933);
    layer1_outputs(881) <= not(layer0_outputs(7013));
    layer1_outputs(882) <= (layer0_outputs(6980)) xor (layer0_outputs(8558));
    layer1_outputs(883) <= '0';
    layer1_outputs(884) <= not(layer0_outputs(5439)) or (layer0_outputs(8188));
    layer1_outputs(885) <= layer0_outputs(4941);
    layer1_outputs(886) <= not(layer0_outputs(9395));
    layer1_outputs(887) <= (layer0_outputs(3122)) xor (layer0_outputs(6976));
    layer1_outputs(888) <= (layer0_outputs(9168)) or (layer0_outputs(8725));
    layer1_outputs(889) <= not(layer0_outputs(4237)) or (layer0_outputs(9283));
    layer1_outputs(890) <= not(layer0_outputs(7430));
    layer1_outputs(891) <= layer0_outputs(5298);
    layer1_outputs(892) <= (layer0_outputs(4745)) and not (layer0_outputs(5075));
    layer1_outputs(893) <= not(layer0_outputs(7235));
    layer1_outputs(894) <= not(layer0_outputs(7219));
    layer1_outputs(895) <= not(layer0_outputs(8976));
    layer1_outputs(896) <= not(layer0_outputs(53)) or (layer0_outputs(1260));
    layer1_outputs(897) <= not(layer0_outputs(4851));
    layer1_outputs(898) <= layer0_outputs(9242);
    layer1_outputs(899) <= layer0_outputs(7471);
    layer1_outputs(900) <= not((layer0_outputs(1081)) xor (layer0_outputs(3505)));
    layer1_outputs(901) <= layer0_outputs(4065);
    layer1_outputs(902) <= layer0_outputs(8311);
    layer1_outputs(903) <= (layer0_outputs(463)) or (layer0_outputs(839));
    layer1_outputs(904) <= not(layer0_outputs(8190));
    layer1_outputs(905) <= not((layer0_outputs(979)) xor (layer0_outputs(7476)));
    layer1_outputs(906) <= not((layer0_outputs(3843)) and (layer0_outputs(2027)));
    layer1_outputs(907) <= not((layer0_outputs(7296)) or (layer0_outputs(1285)));
    layer1_outputs(908) <= not(layer0_outputs(1441));
    layer1_outputs(909) <= (layer0_outputs(3088)) and not (layer0_outputs(8089));
    layer1_outputs(910) <= (layer0_outputs(9233)) and not (layer0_outputs(969));
    layer1_outputs(911) <= not(layer0_outputs(8821));
    layer1_outputs(912) <= (layer0_outputs(8740)) and (layer0_outputs(1711));
    layer1_outputs(913) <= not(layer0_outputs(5456)) or (layer0_outputs(7942));
    layer1_outputs(914) <= not(layer0_outputs(4390)) or (layer0_outputs(2580));
    layer1_outputs(915) <= not(layer0_outputs(4528));
    layer1_outputs(916) <= not((layer0_outputs(1675)) or (layer0_outputs(2704)));
    layer1_outputs(917) <= (layer0_outputs(3519)) xor (layer0_outputs(8022));
    layer1_outputs(918) <= not(layer0_outputs(9306));
    layer1_outputs(919) <= not(layer0_outputs(4884)) or (layer0_outputs(4324));
    layer1_outputs(920) <= layer0_outputs(177);
    layer1_outputs(921) <= not((layer0_outputs(3559)) and (layer0_outputs(5083)));
    layer1_outputs(922) <= not((layer0_outputs(966)) and (layer0_outputs(281)));
    layer1_outputs(923) <= not(layer0_outputs(5809)) or (layer0_outputs(9696));
    layer1_outputs(924) <= not(layer0_outputs(2054)) or (layer0_outputs(9040));
    layer1_outputs(925) <= not(layer0_outputs(5078)) or (layer0_outputs(2359));
    layer1_outputs(926) <= layer0_outputs(3421);
    layer1_outputs(927) <= layer0_outputs(10170);
    layer1_outputs(928) <= layer0_outputs(9760);
    layer1_outputs(929) <= not((layer0_outputs(10089)) and (layer0_outputs(10113)));
    layer1_outputs(930) <= not((layer0_outputs(4524)) xor (layer0_outputs(1979)));
    layer1_outputs(931) <= not(layer0_outputs(8804)) or (layer0_outputs(3270));
    layer1_outputs(932) <= (layer0_outputs(6780)) and not (layer0_outputs(7398));
    layer1_outputs(933) <= (layer0_outputs(1760)) or (layer0_outputs(10101));
    layer1_outputs(934) <= not(layer0_outputs(7969)) or (layer0_outputs(7498));
    layer1_outputs(935) <= not(layer0_outputs(5299)) or (layer0_outputs(6514));
    layer1_outputs(936) <= layer0_outputs(3419);
    layer1_outputs(937) <= not(layer0_outputs(3146));
    layer1_outputs(938) <= (layer0_outputs(3961)) and not (layer0_outputs(2784));
    layer1_outputs(939) <= not(layer0_outputs(333));
    layer1_outputs(940) <= layer0_outputs(5303);
    layer1_outputs(941) <= not((layer0_outputs(1130)) and (layer0_outputs(5644)));
    layer1_outputs(942) <= not((layer0_outputs(1769)) or (layer0_outputs(9762)));
    layer1_outputs(943) <= layer0_outputs(5591);
    layer1_outputs(944) <= not(layer0_outputs(5598));
    layer1_outputs(945) <= (layer0_outputs(9678)) and (layer0_outputs(9835));
    layer1_outputs(946) <= not(layer0_outputs(4525));
    layer1_outputs(947) <= layer0_outputs(6667);
    layer1_outputs(948) <= layer0_outputs(4310);
    layer1_outputs(949) <= not(layer0_outputs(4192));
    layer1_outputs(950) <= layer0_outputs(1461);
    layer1_outputs(951) <= not(layer0_outputs(4599));
    layer1_outputs(952) <= (layer0_outputs(781)) and not (layer0_outputs(6814));
    layer1_outputs(953) <= not(layer0_outputs(133));
    layer1_outputs(954) <= not(layer0_outputs(7330));
    layer1_outputs(955) <= not((layer0_outputs(9569)) or (layer0_outputs(179)));
    layer1_outputs(956) <= not(layer0_outputs(9730));
    layer1_outputs(957) <= not(layer0_outputs(1988));
    layer1_outputs(958) <= (layer0_outputs(2861)) and not (layer0_outputs(897));
    layer1_outputs(959) <= (layer0_outputs(5048)) or (layer0_outputs(496));
    layer1_outputs(960) <= (layer0_outputs(3548)) or (layer0_outputs(1754));
    layer1_outputs(961) <= not((layer0_outputs(8844)) xor (layer0_outputs(1555)));
    layer1_outputs(962) <= (layer0_outputs(5044)) and (layer0_outputs(4380));
    layer1_outputs(963) <= not(layer0_outputs(3706)) or (layer0_outputs(8940));
    layer1_outputs(964) <= not(layer0_outputs(4242)) or (layer0_outputs(3038));
    layer1_outputs(965) <= layer0_outputs(9957);
    layer1_outputs(966) <= (layer0_outputs(48)) or (layer0_outputs(5727));
    layer1_outputs(967) <= not((layer0_outputs(8975)) and (layer0_outputs(6157)));
    layer1_outputs(968) <= not(layer0_outputs(10208));
    layer1_outputs(969) <= (layer0_outputs(5339)) and not (layer0_outputs(3722));
    layer1_outputs(970) <= layer0_outputs(9313);
    layer1_outputs(971) <= (layer0_outputs(222)) or (layer0_outputs(7642));
    layer1_outputs(972) <= layer0_outputs(5392);
    layer1_outputs(973) <= layer0_outputs(2540);
    layer1_outputs(974) <= not(layer0_outputs(1419));
    layer1_outputs(975) <= not(layer0_outputs(1539)) or (layer0_outputs(4081));
    layer1_outputs(976) <= layer0_outputs(6523);
    layer1_outputs(977) <= not(layer0_outputs(5036));
    layer1_outputs(978) <= (layer0_outputs(9646)) or (layer0_outputs(8497));
    layer1_outputs(979) <= not((layer0_outputs(88)) xor (layer0_outputs(460)));
    layer1_outputs(980) <= not(layer0_outputs(7902));
    layer1_outputs(981) <= not(layer0_outputs(8848));
    layer1_outputs(982) <= not(layer0_outputs(960));
    layer1_outputs(983) <= (layer0_outputs(5491)) and not (layer0_outputs(5421));
    layer1_outputs(984) <= not((layer0_outputs(5001)) or (layer0_outputs(3707)));
    layer1_outputs(985) <= not(layer0_outputs(9314));
    layer1_outputs(986) <= (layer0_outputs(9696)) or (layer0_outputs(9488));
    layer1_outputs(987) <= not(layer0_outputs(8655));
    layer1_outputs(988) <= not(layer0_outputs(10027));
    layer1_outputs(989) <= not((layer0_outputs(1610)) or (layer0_outputs(2781)));
    layer1_outputs(990) <= (layer0_outputs(1997)) and not (layer0_outputs(9791));
    layer1_outputs(991) <= (layer0_outputs(1355)) xor (layer0_outputs(3486));
    layer1_outputs(992) <= layer0_outputs(7228);
    layer1_outputs(993) <= not(layer0_outputs(4449)) or (layer0_outputs(9349));
    layer1_outputs(994) <= not(layer0_outputs(8534));
    layer1_outputs(995) <= layer0_outputs(7375);
    layer1_outputs(996) <= layer0_outputs(7018);
    layer1_outputs(997) <= not(layer0_outputs(3286));
    layer1_outputs(998) <= not(layer0_outputs(5324));
    layer1_outputs(999) <= layer0_outputs(1619);
    layer1_outputs(1000) <= not(layer0_outputs(5127));
    layer1_outputs(1001) <= not(layer0_outputs(8877));
    layer1_outputs(1002) <= not(layer0_outputs(8496));
    layer1_outputs(1003) <= (layer0_outputs(2485)) and not (layer0_outputs(7801));
    layer1_outputs(1004) <= (layer0_outputs(1689)) and not (layer0_outputs(3283));
    layer1_outputs(1005) <= layer0_outputs(7871);
    layer1_outputs(1006) <= not(layer0_outputs(1972)) or (layer0_outputs(3828));
    layer1_outputs(1007) <= (layer0_outputs(1268)) and not (layer0_outputs(4849));
    layer1_outputs(1008) <= not(layer0_outputs(8128));
    layer1_outputs(1009) <= (layer0_outputs(1371)) and (layer0_outputs(7466));
    layer1_outputs(1010) <= (layer0_outputs(848)) or (layer0_outputs(1061));
    layer1_outputs(1011) <= not((layer0_outputs(5695)) or (layer0_outputs(9458)));
    layer1_outputs(1012) <= not(layer0_outputs(8865)) or (layer0_outputs(4699));
    layer1_outputs(1013) <= not(layer0_outputs(5177));
    layer1_outputs(1014) <= (layer0_outputs(1041)) or (layer0_outputs(10220));
    layer1_outputs(1015) <= (layer0_outputs(2856)) and not (layer0_outputs(3014));
    layer1_outputs(1016) <= not((layer0_outputs(7859)) and (layer0_outputs(3615)));
    layer1_outputs(1017) <= (layer0_outputs(7690)) and (layer0_outputs(7893));
    layer1_outputs(1018) <= not((layer0_outputs(9342)) and (layer0_outputs(1046)));
    layer1_outputs(1019) <= '0';
    layer1_outputs(1020) <= (layer0_outputs(6385)) xor (layer0_outputs(5640));
    layer1_outputs(1021) <= not((layer0_outputs(3040)) and (layer0_outputs(5471)));
    layer1_outputs(1022) <= not((layer0_outputs(1835)) xor (layer0_outputs(3012)));
    layer1_outputs(1023) <= (layer0_outputs(8025)) or (layer0_outputs(638));
    layer1_outputs(1024) <= not(layer0_outputs(9067)) or (layer0_outputs(4797));
    layer1_outputs(1025) <= (layer0_outputs(6805)) and (layer0_outputs(7606));
    layer1_outputs(1026) <= (layer0_outputs(8280)) or (layer0_outputs(8972));
    layer1_outputs(1027) <= (layer0_outputs(7858)) and not (layer0_outputs(4254));
    layer1_outputs(1028) <= (layer0_outputs(2470)) and not (layer0_outputs(5851));
    layer1_outputs(1029) <= (layer0_outputs(2421)) or (layer0_outputs(6609));
    layer1_outputs(1030) <= layer0_outputs(3188);
    layer1_outputs(1031) <= not(layer0_outputs(8517));
    layer1_outputs(1032) <= not((layer0_outputs(6402)) or (layer0_outputs(5811)));
    layer1_outputs(1033) <= (layer0_outputs(8765)) or (layer0_outputs(7880));
    layer1_outputs(1034) <= not(layer0_outputs(1518));
    layer1_outputs(1035) <= (layer0_outputs(8391)) and not (layer0_outputs(5570));
    layer1_outputs(1036) <= not((layer0_outputs(2486)) and (layer0_outputs(2426)));
    layer1_outputs(1037) <= (layer0_outputs(9867)) and (layer0_outputs(5304));
    layer1_outputs(1038) <= not(layer0_outputs(3648)) or (layer0_outputs(8204));
    layer1_outputs(1039) <= (layer0_outputs(6610)) and not (layer0_outputs(2452));
    layer1_outputs(1040) <= not(layer0_outputs(10228));
    layer1_outputs(1041) <= not(layer0_outputs(5912));
    layer1_outputs(1042) <= not((layer0_outputs(1189)) and (layer0_outputs(4819)));
    layer1_outputs(1043) <= not((layer0_outputs(5146)) xor (layer0_outputs(4028)));
    layer1_outputs(1044) <= '0';
    layer1_outputs(1045) <= not(layer0_outputs(2226));
    layer1_outputs(1046) <= not(layer0_outputs(2288)) or (layer0_outputs(6869));
    layer1_outputs(1047) <= not(layer0_outputs(7504));
    layer1_outputs(1048) <= (layer0_outputs(644)) and (layer0_outputs(4972));
    layer1_outputs(1049) <= not(layer0_outputs(4818)) or (layer0_outputs(9203));
    layer1_outputs(1050) <= (layer0_outputs(2591)) and (layer0_outputs(5205));
    layer1_outputs(1051) <= not((layer0_outputs(9081)) xor (layer0_outputs(8952)));
    layer1_outputs(1052) <= not((layer0_outputs(6147)) or (layer0_outputs(1355)));
    layer1_outputs(1053) <= '1';
    layer1_outputs(1054) <= '0';
    layer1_outputs(1055) <= not((layer0_outputs(7431)) and (layer0_outputs(46)));
    layer1_outputs(1056) <= not((layer0_outputs(5222)) and (layer0_outputs(4315)));
    layer1_outputs(1057) <= '0';
    layer1_outputs(1058) <= (layer0_outputs(8526)) and not (layer0_outputs(7640));
    layer1_outputs(1059) <= not(layer0_outputs(4938)) or (layer0_outputs(2561));
    layer1_outputs(1060) <= not((layer0_outputs(3580)) xor (layer0_outputs(7491)));
    layer1_outputs(1061) <= not(layer0_outputs(353));
    layer1_outputs(1062) <= not(layer0_outputs(3857)) or (layer0_outputs(1375));
    layer1_outputs(1063) <= not(layer0_outputs(9699));
    layer1_outputs(1064) <= not(layer0_outputs(9712));
    layer1_outputs(1065) <= not(layer0_outputs(2072)) or (layer0_outputs(5133));
    layer1_outputs(1066) <= layer0_outputs(10083);
    layer1_outputs(1067) <= not(layer0_outputs(1661)) or (layer0_outputs(1712));
    layer1_outputs(1068) <= (layer0_outputs(7283)) or (layer0_outputs(5737));
    layer1_outputs(1069) <= (layer0_outputs(6363)) and (layer0_outputs(9827));
    layer1_outputs(1070) <= layer0_outputs(1238);
    layer1_outputs(1071) <= not(layer0_outputs(3847)) or (layer0_outputs(804));
    layer1_outputs(1072) <= not(layer0_outputs(8741));
    layer1_outputs(1073) <= layer0_outputs(5449);
    layer1_outputs(1074) <= (layer0_outputs(8951)) and not (layer0_outputs(3588));
    layer1_outputs(1075) <= not(layer0_outputs(9085));
    layer1_outputs(1076) <= (layer0_outputs(7886)) xor (layer0_outputs(7536));
    layer1_outputs(1077) <= layer0_outputs(3290);
    layer1_outputs(1078) <= not(layer0_outputs(6216));
    layer1_outputs(1079) <= not(layer0_outputs(9366));
    layer1_outputs(1080) <= not((layer0_outputs(5769)) and (layer0_outputs(6774)));
    layer1_outputs(1081) <= not(layer0_outputs(8819));
    layer1_outputs(1082) <= layer0_outputs(286);
    layer1_outputs(1083) <= not(layer0_outputs(4516)) or (layer0_outputs(7789));
    layer1_outputs(1084) <= (layer0_outputs(7876)) or (layer0_outputs(3149));
    layer1_outputs(1085) <= not(layer0_outputs(9393));
    layer1_outputs(1086) <= (layer0_outputs(2063)) and (layer0_outputs(3814));
    layer1_outputs(1087) <= not(layer0_outputs(4756));
    layer1_outputs(1088) <= not(layer0_outputs(8069));
    layer1_outputs(1089) <= (layer0_outputs(7590)) or (layer0_outputs(10076));
    layer1_outputs(1090) <= not(layer0_outputs(149));
    layer1_outputs(1091) <= not((layer0_outputs(1862)) or (layer0_outputs(6350)));
    layer1_outputs(1092) <= not(layer0_outputs(8078));
    layer1_outputs(1093) <= not(layer0_outputs(7377));
    layer1_outputs(1094) <= not((layer0_outputs(6627)) xor (layer0_outputs(9329)));
    layer1_outputs(1095) <= not(layer0_outputs(9365));
    layer1_outputs(1096) <= not(layer0_outputs(1250)) or (layer0_outputs(4488));
    layer1_outputs(1097) <= not(layer0_outputs(2387)) or (layer0_outputs(10092));
    layer1_outputs(1098) <= not(layer0_outputs(2212)) or (layer0_outputs(7185));
    layer1_outputs(1099) <= (layer0_outputs(5341)) and (layer0_outputs(8218));
    layer1_outputs(1100) <= not(layer0_outputs(6383));
    layer1_outputs(1101) <= layer0_outputs(2139);
    layer1_outputs(1102) <= (layer0_outputs(8611)) and (layer0_outputs(6348));
    layer1_outputs(1103) <= layer0_outputs(9055);
    layer1_outputs(1104) <= layer0_outputs(7999);
    layer1_outputs(1105) <= (layer0_outputs(2961)) or (layer0_outputs(7263));
    layer1_outputs(1106) <= not(layer0_outputs(4554)) or (layer0_outputs(10171));
    layer1_outputs(1107) <= (layer0_outputs(3678)) and not (layer0_outputs(616));
    layer1_outputs(1108) <= not(layer0_outputs(5609)) or (layer0_outputs(2600));
    layer1_outputs(1109) <= (layer0_outputs(9219)) and (layer0_outputs(2560));
    layer1_outputs(1110) <= (layer0_outputs(7586)) and not (layer0_outputs(4446));
    layer1_outputs(1111) <= (layer0_outputs(6415)) xor (layer0_outputs(7964));
    layer1_outputs(1112) <= not((layer0_outputs(4891)) xor (layer0_outputs(9268)));
    layer1_outputs(1113) <= not((layer0_outputs(1659)) and (layer0_outputs(1751)));
    layer1_outputs(1114) <= not((layer0_outputs(3291)) xor (layer0_outputs(6085)));
    layer1_outputs(1115) <= layer0_outputs(334);
    layer1_outputs(1116) <= (layer0_outputs(9988)) or (layer0_outputs(1144));
    layer1_outputs(1117) <= (layer0_outputs(5462)) or (layer0_outputs(8294));
    layer1_outputs(1118) <= layer0_outputs(6654);
    layer1_outputs(1119) <= (layer0_outputs(10011)) or (layer0_outputs(7021));
    layer1_outputs(1120) <= (layer0_outputs(3649)) and not (layer0_outputs(1244));
    layer1_outputs(1121) <= (layer0_outputs(1360)) and (layer0_outputs(4125));
    layer1_outputs(1122) <= (layer0_outputs(10055)) or (layer0_outputs(3266));
    layer1_outputs(1123) <= not((layer0_outputs(2497)) or (layer0_outputs(5188)));
    layer1_outputs(1124) <= layer0_outputs(6058);
    layer1_outputs(1125) <= not((layer0_outputs(6579)) and (layer0_outputs(1228)));
    layer1_outputs(1126) <= (layer0_outputs(5575)) or (layer0_outputs(9303));
    layer1_outputs(1127) <= (layer0_outputs(6130)) or (layer0_outputs(2639));
    layer1_outputs(1128) <= (layer0_outputs(4758)) and not (layer0_outputs(10119));
    layer1_outputs(1129) <= (layer0_outputs(5551)) and not (layer0_outputs(5123));
    layer1_outputs(1130) <= not(layer0_outputs(1882)) or (layer0_outputs(3516));
    layer1_outputs(1131) <= layer0_outputs(1621);
    layer1_outputs(1132) <= layer0_outputs(7137);
    layer1_outputs(1133) <= not((layer0_outputs(5820)) or (layer0_outputs(1799)));
    layer1_outputs(1134) <= not(layer0_outputs(608));
    layer1_outputs(1135) <= (layer0_outputs(6615)) and not (layer0_outputs(7264));
    layer1_outputs(1136) <= layer0_outputs(2764);
    layer1_outputs(1137) <= not(layer0_outputs(703)) or (layer0_outputs(425));
    layer1_outputs(1138) <= not(layer0_outputs(2528));
    layer1_outputs(1139) <= not(layer0_outputs(9943));
    layer1_outputs(1140) <= (layer0_outputs(10072)) or (layer0_outputs(1331));
    layer1_outputs(1141) <= (layer0_outputs(8693)) or (layer0_outputs(3414));
    layer1_outputs(1142) <= not((layer0_outputs(4935)) or (layer0_outputs(4588)));
    layer1_outputs(1143) <= (layer0_outputs(2496)) and (layer0_outputs(459));
    layer1_outputs(1144) <= not((layer0_outputs(4753)) and (layer0_outputs(1733)));
    layer1_outputs(1145) <= not((layer0_outputs(3308)) xor (layer0_outputs(9050)));
    layer1_outputs(1146) <= (layer0_outputs(4560)) and (layer0_outputs(2493));
    layer1_outputs(1147) <= (layer0_outputs(4805)) and not (layer0_outputs(9610));
    layer1_outputs(1148) <= (layer0_outputs(6992)) and not (layer0_outputs(7701));
    layer1_outputs(1149) <= not((layer0_outputs(6121)) and (layer0_outputs(659)));
    layer1_outputs(1150) <= not(layer0_outputs(8256)) or (layer0_outputs(1687));
    layer1_outputs(1151) <= layer0_outputs(10072);
    layer1_outputs(1152) <= (layer0_outputs(3967)) and not (layer0_outputs(8432));
    layer1_outputs(1153) <= not(layer0_outputs(2412));
    layer1_outputs(1154) <= '0';
    layer1_outputs(1155) <= '0';
    layer1_outputs(1156) <= (layer0_outputs(2995)) and not (layer0_outputs(8189));
    layer1_outputs(1157) <= not(layer0_outputs(8097)) or (layer0_outputs(656));
    layer1_outputs(1158) <= not(layer0_outputs(2592));
    layer1_outputs(1159) <= (layer0_outputs(8356)) xor (layer0_outputs(4614));
    layer1_outputs(1160) <= not(layer0_outputs(3269));
    layer1_outputs(1161) <= layer0_outputs(3232);
    layer1_outputs(1162) <= not(layer0_outputs(4102)) or (layer0_outputs(598));
    layer1_outputs(1163) <= not((layer0_outputs(5101)) or (layer0_outputs(6172)));
    layer1_outputs(1164) <= layer0_outputs(3140);
    layer1_outputs(1165) <= not(layer0_outputs(3598));
    layer1_outputs(1166) <= layer0_outputs(337);
    layer1_outputs(1167) <= layer0_outputs(9976);
    layer1_outputs(1168) <= (layer0_outputs(5586)) and not (layer0_outputs(8444));
    layer1_outputs(1169) <= not(layer0_outputs(7925));
    layer1_outputs(1170) <= (layer0_outputs(4364)) and (layer0_outputs(3873));
    layer1_outputs(1171) <= not((layer0_outputs(6407)) or (layer0_outputs(1058)));
    layer1_outputs(1172) <= not((layer0_outputs(8615)) or (layer0_outputs(8292)));
    layer1_outputs(1173) <= '1';
    layer1_outputs(1174) <= not(layer0_outputs(5478));
    layer1_outputs(1175) <= not(layer0_outputs(4126)) or (layer0_outputs(580));
    layer1_outputs(1176) <= not(layer0_outputs(5719));
    layer1_outputs(1177) <= (layer0_outputs(7200)) and not (layer0_outputs(9227));
    layer1_outputs(1178) <= not(layer0_outputs(9804));
    layer1_outputs(1179) <= not(layer0_outputs(7234));
    layer1_outputs(1180) <= layer0_outputs(610);
    layer1_outputs(1181) <= (layer0_outputs(107)) and not (layer0_outputs(3149));
    layer1_outputs(1182) <= layer0_outputs(8618);
    layer1_outputs(1183) <= (layer0_outputs(7503)) and not (layer0_outputs(5454));
    layer1_outputs(1184) <= (layer0_outputs(6158)) xor (layer0_outputs(6696));
    layer1_outputs(1185) <= (layer0_outputs(6739)) xor (layer0_outputs(294));
    layer1_outputs(1186) <= not(layer0_outputs(629)) or (layer0_outputs(9600));
    layer1_outputs(1187) <= not(layer0_outputs(5287));
    layer1_outputs(1188) <= not(layer0_outputs(3556));
    layer1_outputs(1189) <= not((layer0_outputs(1206)) or (layer0_outputs(10012)));
    layer1_outputs(1190) <= not(layer0_outputs(9563)) or (layer0_outputs(1329));
    layer1_outputs(1191) <= (layer0_outputs(1633)) xor (layer0_outputs(6700));
    layer1_outputs(1192) <= not((layer0_outputs(1427)) xor (layer0_outputs(6296)));
    layer1_outputs(1193) <= not((layer0_outputs(4740)) and (layer0_outputs(1672)));
    layer1_outputs(1194) <= not(layer0_outputs(7043));
    layer1_outputs(1195) <= '1';
    layer1_outputs(1196) <= (layer0_outputs(1316)) and not (layer0_outputs(8616));
    layer1_outputs(1197) <= not(layer0_outputs(4346)) or (layer0_outputs(5616));
    layer1_outputs(1198) <= (layer0_outputs(907)) and (layer0_outputs(5700));
    layer1_outputs(1199) <= (layer0_outputs(4723)) and (layer0_outputs(3994));
    layer1_outputs(1200) <= layer0_outputs(7934);
    layer1_outputs(1201) <= not(layer0_outputs(8979)) or (layer0_outputs(5163));
    layer1_outputs(1202) <= not(layer0_outputs(1777)) or (layer0_outputs(8539));
    layer1_outputs(1203) <= layer0_outputs(5699);
    layer1_outputs(1204) <= not(layer0_outputs(8451)) or (layer0_outputs(5361));
    layer1_outputs(1205) <= not((layer0_outputs(7121)) xor (layer0_outputs(2160)));
    layer1_outputs(1206) <= layer0_outputs(5511);
    layer1_outputs(1207) <= (layer0_outputs(3361)) and not (layer0_outputs(6784));
    layer1_outputs(1208) <= not(layer0_outputs(4211));
    layer1_outputs(1209) <= not(layer0_outputs(3497));
    layer1_outputs(1210) <= (layer0_outputs(5780)) and not (layer0_outputs(8913));
    layer1_outputs(1211) <= layer0_outputs(4778);
    layer1_outputs(1212) <= not(layer0_outputs(3963)) or (layer0_outputs(5213));
    layer1_outputs(1213) <= not(layer0_outputs(1804));
    layer1_outputs(1214) <= (layer0_outputs(2789)) and not (layer0_outputs(5569));
    layer1_outputs(1215) <= not(layer0_outputs(3406)) or (layer0_outputs(10141));
    layer1_outputs(1216) <= (layer0_outputs(2575)) and (layer0_outputs(773));
    layer1_outputs(1217) <= (layer0_outputs(6472)) xor (layer0_outputs(10133));
    layer1_outputs(1218) <= not(layer0_outputs(2973));
    layer1_outputs(1219) <= not((layer0_outputs(6256)) or (layer0_outputs(1602)));
    layer1_outputs(1220) <= layer0_outputs(7935);
    layer1_outputs(1221) <= layer0_outputs(1407);
    layer1_outputs(1222) <= not((layer0_outputs(9588)) and (layer0_outputs(2708)));
    layer1_outputs(1223) <= not(layer0_outputs(3163));
    layer1_outputs(1224) <= not((layer0_outputs(3424)) and (layer0_outputs(8637)));
    layer1_outputs(1225) <= not((layer0_outputs(5343)) and (layer0_outputs(4902)));
    layer1_outputs(1226) <= layer0_outputs(2097);
    layer1_outputs(1227) <= (layer0_outputs(9884)) xor (layer0_outputs(5118));
    layer1_outputs(1228) <= layer0_outputs(1557);
    layer1_outputs(1229) <= layer0_outputs(943);
    layer1_outputs(1230) <= layer0_outputs(10232);
    layer1_outputs(1231) <= not(layer0_outputs(3326));
    layer1_outputs(1232) <= not(layer0_outputs(1302)) or (layer0_outputs(9683));
    layer1_outputs(1233) <= layer0_outputs(6273);
    layer1_outputs(1234) <= (layer0_outputs(1014)) and (layer0_outputs(8771));
    layer1_outputs(1235) <= (layer0_outputs(5350)) and not (layer0_outputs(1523));
    layer1_outputs(1236) <= not((layer0_outputs(4105)) and (layer0_outputs(3250)));
    layer1_outputs(1237) <= layer0_outputs(8978);
    layer1_outputs(1238) <= layer0_outputs(5641);
    layer1_outputs(1239) <= (layer0_outputs(9012)) xor (layer0_outputs(1971));
    layer1_outputs(1240) <= (layer0_outputs(3737)) or (layer0_outputs(6105));
    layer1_outputs(1241) <= '0';
    layer1_outputs(1242) <= (layer0_outputs(5213)) or (layer0_outputs(9593));
    layer1_outputs(1243) <= (layer0_outputs(4976)) or (layer0_outputs(3174));
    layer1_outputs(1244) <= (layer0_outputs(7838)) and (layer0_outputs(4497));
    layer1_outputs(1245) <= not((layer0_outputs(3976)) xor (layer0_outputs(9222)));
    layer1_outputs(1246) <= not(layer0_outputs(2123));
    layer1_outputs(1247) <= not(layer0_outputs(3377));
    layer1_outputs(1248) <= layer0_outputs(2573);
    layer1_outputs(1249) <= '1';
    layer1_outputs(1250) <= (layer0_outputs(6196)) and not (layer0_outputs(9741));
    layer1_outputs(1251) <= (layer0_outputs(5162)) or (layer0_outputs(713));
    layer1_outputs(1252) <= not(layer0_outputs(7305)) or (layer0_outputs(5676));
    layer1_outputs(1253) <= not((layer0_outputs(9643)) and (layer0_outputs(976)));
    layer1_outputs(1254) <= (layer0_outputs(763)) and not (layer0_outputs(4223));
    layer1_outputs(1255) <= not((layer0_outputs(1912)) and (layer0_outputs(4937)));
    layer1_outputs(1256) <= not(layer0_outputs(8810));
    layer1_outputs(1257) <= not((layer0_outputs(2775)) or (layer0_outputs(828)));
    layer1_outputs(1258) <= (layer0_outputs(4265)) and not (layer0_outputs(4729));
    layer1_outputs(1259) <= (layer0_outputs(5205)) and (layer0_outputs(8960));
    layer1_outputs(1260) <= layer0_outputs(5592);
    layer1_outputs(1261) <= not((layer0_outputs(9077)) or (layer0_outputs(1990)));
    layer1_outputs(1262) <= not((layer0_outputs(2061)) xor (layer0_outputs(464)));
    layer1_outputs(1263) <= layer0_outputs(7202);
    layer1_outputs(1264) <= not(layer0_outputs(2238));
    layer1_outputs(1265) <= not(layer0_outputs(7712)) or (layer0_outputs(2906));
    layer1_outputs(1266) <= layer0_outputs(788);
    layer1_outputs(1267) <= not(layer0_outputs(5312)) or (layer0_outputs(348));
    layer1_outputs(1268) <= not((layer0_outputs(2439)) and (layer0_outputs(5699)));
    layer1_outputs(1269) <= not((layer0_outputs(4609)) or (layer0_outputs(6180)));
    layer1_outputs(1270) <= (layer0_outputs(2022)) or (layer0_outputs(8229));
    layer1_outputs(1271) <= (layer0_outputs(6934)) xor (layer0_outputs(5291));
    layer1_outputs(1272) <= layer0_outputs(922);
    layer1_outputs(1273) <= not(layer0_outputs(2580));
    layer1_outputs(1274) <= not(layer0_outputs(3068)) or (layer0_outputs(903));
    layer1_outputs(1275) <= layer0_outputs(2015);
    layer1_outputs(1276) <= (layer0_outputs(6156)) or (layer0_outputs(8912));
    layer1_outputs(1277) <= layer0_outputs(5987);
    layer1_outputs(1278) <= layer0_outputs(9240);
    layer1_outputs(1279) <= not(layer0_outputs(415));
    layer1_outputs(1280) <= not(layer0_outputs(8512));
    layer1_outputs(1281) <= (layer0_outputs(10001)) and not (layer0_outputs(6933));
    layer1_outputs(1282) <= not((layer0_outputs(1281)) xor (layer0_outputs(3844)));
    layer1_outputs(1283) <= not(layer0_outputs(2476)) or (layer0_outputs(6914));
    layer1_outputs(1284) <= (layer0_outputs(2270)) or (layer0_outputs(3014));
    layer1_outputs(1285) <= layer0_outputs(1160);
    layer1_outputs(1286) <= not((layer0_outputs(10112)) and (layer0_outputs(7788)));
    layer1_outputs(1287) <= (layer0_outputs(1852)) or (layer0_outputs(9102));
    layer1_outputs(1288) <= layer0_outputs(3614);
    layer1_outputs(1289) <= not((layer0_outputs(1242)) xor (layer0_outputs(7322)));
    layer1_outputs(1290) <= layer0_outputs(2889);
    layer1_outputs(1291) <= (layer0_outputs(7084)) xor (layer0_outputs(4014));
    layer1_outputs(1292) <= (layer0_outputs(9439)) and not (layer0_outputs(8488));
    layer1_outputs(1293) <= '0';
    layer1_outputs(1294) <= not(layer0_outputs(2588));
    layer1_outputs(1295) <= layer0_outputs(2257);
    layer1_outputs(1296) <= layer0_outputs(7711);
    layer1_outputs(1297) <= '1';
    layer1_outputs(1298) <= not(layer0_outputs(9791));
    layer1_outputs(1299) <= not(layer0_outputs(989));
    layer1_outputs(1300) <= not(layer0_outputs(2167));
    layer1_outputs(1301) <= layer0_outputs(1805);
    layer1_outputs(1302) <= not(layer0_outputs(1784)) or (layer0_outputs(8192));
    layer1_outputs(1303) <= layer0_outputs(6706);
    layer1_outputs(1304) <= not(layer0_outputs(609));
    layer1_outputs(1305) <= '0';
    layer1_outputs(1306) <= not(layer0_outputs(5855));
    layer1_outputs(1307) <= (layer0_outputs(4165)) and not (layer0_outputs(4979));
    layer1_outputs(1308) <= (layer0_outputs(9391)) and not (layer0_outputs(4727));
    layer1_outputs(1309) <= not(layer0_outputs(6766)) or (layer0_outputs(8396));
    layer1_outputs(1310) <= (layer0_outputs(9116)) xor (layer0_outputs(6391));
    layer1_outputs(1311) <= not((layer0_outputs(8636)) or (layer0_outputs(8479)));
    layer1_outputs(1312) <= (layer0_outputs(2860)) or (layer0_outputs(5872));
    layer1_outputs(1313) <= not(layer0_outputs(89)) or (layer0_outputs(8316));
    layer1_outputs(1314) <= layer0_outputs(7681);
    layer1_outputs(1315) <= layer0_outputs(5097);
    layer1_outputs(1316) <= layer0_outputs(10212);
    layer1_outputs(1317) <= (layer0_outputs(4141)) xor (layer0_outputs(8566));
    layer1_outputs(1318) <= (layer0_outputs(3768)) and (layer0_outputs(6862));
    layer1_outputs(1319) <= layer0_outputs(3439);
    layer1_outputs(1320) <= not((layer0_outputs(2808)) or (layer0_outputs(6770)));
    layer1_outputs(1321) <= (layer0_outputs(9423)) xor (layer0_outputs(10087));
    layer1_outputs(1322) <= not(layer0_outputs(702));
    layer1_outputs(1323) <= not(layer0_outputs(9820));
    layer1_outputs(1324) <= not((layer0_outputs(6405)) and (layer0_outputs(2674)));
    layer1_outputs(1325) <= (layer0_outputs(8419)) or (layer0_outputs(7906));
    layer1_outputs(1326) <= not(layer0_outputs(7361)) or (layer0_outputs(6477));
    layer1_outputs(1327) <= '0';
    layer1_outputs(1328) <= not(layer0_outputs(8515));
    layer1_outputs(1329) <= not(layer0_outputs(4141));
    layer1_outputs(1330) <= (layer0_outputs(1947)) and (layer0_outputs(9976));
    layer1_outputs(1331) <= layer0_outputs(3476);
    layer1_outputs(1332) <= '1';
    layer1_outputs(1333) <= layer0_outputs(7604);
    layer1_outputs(1334) <= layer0_outputs(8759);
    layer1_outputs(1335) <= not((layer0_outputs(196)) xor (layer0_outputs(4255)));
    layer1_outputs(1336) <= not(layer0_outputs(3769));
    layer1_outputs(1337) <= layer0_outputs(7188);
    layer1_outputs(1338) <= layer0_outputs(5347);
    layer1_outputs(1339) <= not((layer0_outputs(1900)) and (layer0_outputs(9497)));
    layer1_outputs(1340) <= layer0_outputs(2209);
    layer1_outputs(1341) <= layer0_outputs(440);
    layer1_outputs(1342) <= not(layer0_outputs(6546));
    layer1_outputs(1343) <= (layer0_outputs(1251)) and (layer0_outputs(4637));
    layer1_outputs(1344) <= not((layer0_outputs(618)) and (layer0_outputs(4115)));
    layer1_outputs(1345) <= not(layer0_outputs(1968));
    layer1_outputs(1346) <= not(layer0_outputs(9134)) or (layer0_outputs(9914));
    layer1_outputs(1347) <= (layer0_outputs(1762)) and (layer0_outputs(2467));
    layer1_outputs(1348) <= not(layer0_outputs(1817));
    layer1_outputs(1349) <= '0';
    layer1_outputs(1350) <= (layer0_outputs(6966)) or (layer0_outputs(443));
    layer1_outputs(1351) <= not(layer0_outputs(3825));
    layer1_outputs(1352) <= not(layer0_outputs(7442)) or (layer0_outputs(7613));
    layer1_outputs(1353) <= (layer0_outputs(6654)) or (layer0_outputs(1996));
    layer1_outputs(1354) <= not(layer0_outputs(60)) or (layer0_outputs(5301));
    layer1_outputs(1355) <= (layer0_outputs(4477)) and (layer0_outputs(8105));
    layer1_outputs(1356) <= not((layer0_outputs(4519)) or (layer0_outputs(2907)));
    layer1_outputs(1357) <= not(layer0_outputs(6963)) or (layer0_outputs(1974));
    layer1_outputs(1358) <= not((layer0_outputs(3883)) or (layer0_outputs(6353)));
    layer1_outputs(1359) <= not((layer0_outputs(9175)) or (layer0_outputs(5012)));
    layer1_outputs(1360) <= not(layer0_outputs(2999));
    layer1_outputs(1361) <= layer0_outputs(7501);
    layer1_outputs(1362) <= not(layer0_outputs(3001)) or (layer0_outputs(2427));
    layer1_outputs(1363) <= (layer0_outputs(7565)) and (layer0_outputs(6764));
    layer1_outputs(1364) <= not(layer0_outputs(3675));
    layer1_outputs(1365) <= not(layer0_outputs(1955));
    layer1_outputs(1366) <= not(layer0_outputs(9755));
    layer1_outputs(1367) <= (layer0_outputs(9194)) xor (layer0_outputs(7555));
    layer1_outputs(1368) <= not(layer0_outputs(44));
    layer1_outputs(1369) <= layer0_outputs(8919);
    layer1_outputs(1370) <= (layer0_outputs(9556)) and not (layer0_outputs(1064));
    layer1_outputs(1371) <= not(layer0_outputs(2679));
    layer1_outputs(1372) <= not(layer0_outputs(10125));
    layer1_outputs(1373) <= '1';
    layer1_outputs(1374) <= layer0_outputs(102);
    layer1_outputs(1375) <= (layer0_outputs(3336)) and not (layer0_outputs(353));
    layer1_outputs(1376) <= not(layer0_outputs(6186));
    layer1_outputs(1377) <= not(layer0_outputs(7610));
    layer1_outputs(1378) <= (layer0_outputs(2969)) and not (layer0_outputs(261));
    layer1_outputs(1379) <= (layer0_outputs(7560)) and (layer0_outputs(4679));
    layer1_outputs(1380) <= not((layer0_outputs(4199)) or (layer0_outputs(2613)));
    layer1_outputs(1381) <= layer0_outputs(749);
    layer1_outputs(1382) <= not(layer0_outputs(705));
    layer1_outputs(1383) <= not(layer0_outputs(5625)) or (layer0_outputs(3386));
    layer1_outputs(1384) <= layer0_outputs(2044);
    layer1_outputs(1385) <= not(layer0_outputs(5741));
    layer1_outputs(1386) <= not((layer0_outputs(2616)) or (layer0_outputs(4218)));
    layer1_outputs(1387) <= (layer0_outputs(835)) and not (layer0_outputs(4168));
    layer1_outputs(1388) <= (layer0_outputs(6430)) or (layer0_outputs(1955));
    layer1_outputs(1389) <= not((layer0_outputs(3674)) xor (layer0_outputs(10090)));
    layer1_outputs(1390) <= (layer0_outputs(2151)) and (layer0_outputs(6347));
    layer1_outputs(1391) <= (layer0_outputs(4330)) and (layer0_outputs(810));
    layer1_outputs(1392) <= not(layer0_outputs(5706)) or (layer0_outputs(5910));
    layer1_outputs(1393) <= not((layer0_outputs(1663)) and (layer0_outputs(6797)));
    layer1_outputs(1394) <= layer0_outputs(8076);
    layer1_outputs(1395) <= not(layer0_outputs(10026)) or (layer0_outputs(6142));
    layer1_outputs(1396) <= (layer0_outputs(6053)) or (layer0_outputs(9829));
    layer1_outputs(1397) <= layer0_outputs(1128);
    layer1_outputs(1398) <= layer0_outputs(7761);
    layer1_outputs(1399) <= (layer0_outputs(5112)) or (layer0_outputs(3302));
    layer1_outputs(1400) <= (layer0_outputs(91)) and not (layer0_outputs(1003));
    layer1_outputs(1401) <= not(layer0_outputs(10239));
    layer1_outputs(1402) <= not(layer0_outputs(10074)) or (layer0_outputs(5222));
    layer1_outputs(1403) <= not((layer0_outputs(7747)) xor (layer0_outputs(10210)));
    layer1_outputs(1404) <= not(layer0_outputs(6727));
    layer1_outputs(1405) <= layer0_outputs(2114);
    layer1_outputs(1406) <= not(layer0_outputs(5285)) or (layer0_outputs(3897));
    layer1_outputs(1407) <= (layer0_outputs(7234)) or (layer0_outputs(295));
    layer1_outputs(1408) <= not(layer0_outputs(9326));
    layer1_outputs(1409) <= not(layer0_outputs(7073));
    layer1_outputs(1410) <= (layer0_outputs(3487)) and (layer0_outputs(5850));
    layer1_outputs(1411) <= (layer0_outputs(7745)) or (layer0_outputs(5854));
    layer1_outputs(1412) <= not((layer0_outputs(8006)) or (layer0_outputs(6407)));
    layer1_outputs(1413) <= layer0_outputs(1138);
    layer1_outputs(1414) <= layer0_outputs(1585);
    layer1_outputs(1415) <= not((layer0_outputs(1343)) xor (layer0_outputs(4347)));
    layer1_outputs(1416) <= not(layer0_outputs(1975));
    layer1_outputs(1417) <= '1';
    layer1_outputs(1418) <= not((layer0_outputs(5493)) and (layer0_outputs(3867)));
    layer1_outputs(1419) <= not(layer0_outputs(3979));
    layer1_outputs(1420) <= layer0_outputs(4006);
    layer1_outputs(1421) <= not(layer0_outputs(4710)) or (layer0_outputs(116));
    layer1_outputs(1422) <= (layer0_outputs(6888)) and not (layer0_outputs(8288));
    layer1_outputs(1423) <= not(layer0_outputs(3322)) or (layer0_outputs(7769));
    layer1_outputs(1424) <= not(layer0_outputs(8853));
    layer1_outputs(1425) <= not(layer0_outputs(9884));
    layer1_outputs(1426) <= '1';
    layer1_outputs(1427) <= not(layer0_outputs(225));
    layer1_outputs(1428) <= '1';
    layer1_outputs(1429) <= not(layer0_outputs(1526)) or (layer0_outputs(1824));
    layer1_outputs(1430) <= (layer0_outputs(2719)) and (layer0_outputs(3000));
    layer1_outputs(1431) <= not(layer0_outputs(6616)) or (layer0_outputs(774));
    layer1_outputs(1432) <= layer0_outputs(32);
    layer1_outputs(1433) <= not(layer0_outputs(2570));
    layer1_outputs(1434) <= (layer0_outputs(3782)) xor (layer0_outputs(268));
    layer1_outputs(1435) <= (layer0_outputs(3884)) and not (layer0_outputs(2270));
    layer1_outputs(1436) <= (layer0_outputs(2219)) and (layer0_outputs(8603));
    layer1_outputs(1437) <= not(layer0_outputs(8401));
    layer1_outputs(1438) <= '0';
    layer1_outputs(1439) <= not(layer0_outputs(8577));
    layer1_outputs(1440) <= not(layer0_outputs(8730));
    layer1_outputs(1441) <= (layer0_outputs(3966)) and not (layer0_outputs(9522));
    layer1_outputs(1442) <= layer0_outputs(5704);
    layer1_outputs(1443) <= not((layer0_outputs(2203)) xor (layer0_outputs(5192)));
    layer1_outputs(1444) <= (layer0_outputs(3249)) and (layer0_outputs(6105));
    layer1_outputs(1445) <= not(layer0_outputs(7597));
    layer1_outputs(1446) <= not(layer0_outputs(1690)) or (layer0_outputs(5691));
    layer1_outputs(1447) <= (layer0_outputs(4461)) xor (layer0_outputs(741));
    layer1_outputs(1448) <= not(layer0_outputs(6716));
    layer1_outputs(1449) <= (layer0_outputs(4215)) and not (layer0_outputs(5740));
    layer1_outputs(1450) <= (layer0_outputs(7214)) xor (layer0_outputs(1407));
    layer1_outputs(1451) <= not((layer0_outputs(890)) and (layer0_outputs(8485)));
    layer1_outputs(1452) <= not(layer0_outputs(6780));
    layer1_outputs(1453) <= not(layer0_outputs(3725)) or (layer0_outputs(4508));
    layer1_outputs(1454) <= not(layer0_outputs(3431));
    layer1_outputs(1455) <= (layer0_outputs(7796)) or (layer0_outputs(5502));
    layer1_outputs(1456) <= not(layer0_outputs(342)) or (layer0_outputs(6314));
    layer1_outputs(1457) <= (layer0_outputs(1258)) and (layer0_outputs(1033));
    layer1_outputs(1458) <= (layer0_outputs(9549)) xor (layer0_outputs(1483));
    layer1_outputs(1459) <= (layer0_outputs(5961)) and (layer0_outputs(9003));
    layer1_outputs(1460) <= (layer0_outputs(3881)) xor (layer0_outputs(8242));
    layer1_outputs(1461) <= (layer0_outputs(6246)) and not (layer0_outputs(7016));
    layer1_outputs(1462) <= (layer0_outputs(9854)) or (layer0_outputs(8696));
    layer1_outputs(1463) <= (layer0_outputs(5921)) or (layer0_outputs(1704));
    layer1_outputs(1464) <= layer0_outputs(7784);
    layer1_outputs(1465) <= (layer0_outputs(7894)) xor (layer0_outputs(3619));
    layer1_outputs(1466) <= not(layer0_outputs(255));
    layer1_outputs(1467) <= (layer0_outputs(2650)) and not (layer0_outputs(5772));
    layer1_outputs(1468) <= not(layer0_outputs(10117)) or (layer0_outputs(5216));
    layer1_outputs(1469) <= not(layer0_outputs(9863));
    layer1_outputs(1470) <= not((layer0_outputs(2046)) and (layer0_outputs(1216)));
    layer1_outputs(1471) <= not(layer0_outputs(2330)) or (layer0_outputs(2090));
    layer1_outputs(1472) <= (layer0_outputs(1845)) xor (layer0_outputs(27));
    layer1_outputs(1473) <= not(layer0_outputs(2035)) or (layer0_outputs(6254));
    layer1_outputs(1474) <= not(layer0_outputs(4887)) or (layer0_outputs(3865));
    layer1_outputs(1475) <= not(layer0_outputs(6015)) or (layer0_outputs(5096));
    layer1_outputs(1476) <= not(layer0_outputs(1491));
    layer1_outputs(1477) <= not(layer0_outputs(4241));
    layer1_outputs(1478) <= layer0_outputs(6836);
    layer1_outputs(1479) <= '1';
    layer1_outputs(1480) <= not(layer0_outputs(9069));
    layer1_outputs(1481) <= not(layer0_outputs(23));
    layer1_outputs(1482) <= not((layer0_outputs(6505)) or (layer0_outputs(6537)));
    layer1_outputs(1483) <= not(layer0_outputs(5477)) or (layer0_outputs(6119));
    layer1_outputs(1484) <= not((layer0_outputs(3138)) or (layer0_outputs(2583)));
    layer1_outputs(1485) <= layer0_outputs(9502);
    layer1_outputs(1486) <= (layer0_outputs(6050)) xor (layer0_outputs(9429));
    layer1_outputs(1487) <= not(layer0_outputs(2344));
    layer1_outputs(1488) <= (layer0_outputs(7924)) xor (layer0_outputs(6290));
    layer1_outputs(1489) <= layer0_outputs(10045);
    layer1_outputs(1490) <= not((layer0_outputs(8478)) and (layer0_outputs(7432)));
    layer1_outputs(1491) <= layer0_outputs(2663);
    layer1_outputs(1492) <= not(layer0_outputs(9758));
    layer1_outputs(1493) <= not(layer0_outputs(2924)) or (layer0_outputs(2405));
    layer1_outputs(1494) <= layer0_outputs(8845);
    layer1_outputs(1495) <= not(layer0_outputs(36)) or (layer0_outputs(9671));
    layer1_outputs(1496) <= (layer0_outputs(9018)) or (layer0_outputs(9335));
    layer1_outputs(1497) <= not(layer0_outputs(5976));
    layer1_outputs(1498) <= layer0_outputs(8284);
    layer1_outputs(1499) <= not(layer0_outputs(3756)) or (layer0_outputs(4252));
    layer1_outputs(1500) <= not((layer0_outputs(2954)) and (layer0_outputs(4772)));
    layer1_outputs(1501) <= (layer0_outputs(3928)) and (layer0_outputs(1168));
    layer1_outputs(1502) <= not(layer0_outputs(6604));
    layer1_outputs(1503) <= not(layer0_outputs(9496));
    layer1_outputs(1504) <= not(layer0_outputs(6377)) or (layer0_outputs(401));
    layer1_outputs(1505) <= not(layer0_outputs(6138));
    layer1_outputs(1506) <= layer0_outputs(2863);
    layer1_outputs(1507) <= layer0_outputs(2407);
    layer1_outputs(1508) <= not(layer0_outputs(2226)) or (layer0_outputs(8406));
    layer1_outputs(1509) <= not(layer0_outputs(7317)) or (layer0_outputs(2188));
    layer1_outputs(1510) <= (layer0_outputs(6182)) and not (layer0_outputs(3383));
    layer1_outputs(1511) <= (layer0_outputs(6778)) and not (layer0_outputs(8034));
    layer1_outputs(1512) <= layer0_outputs(9960);
    layer1_outputs(1513) <= (layer0_outputs(1251)) or (layer0_outputs(1886));
    layer1_outputs(1514) <= not(layer0_outputs(9741)) or (layer0_outputs(642));
    layer1_outputs(1515) <= (layer0_outputs(3332)) xor (layer0_outputs(1377));
    layer1_outputs(1516) <= not((layer0_outputs(6552)) and (layer0_outputs(1646)));
    layer1_outputs(1517) <= '1';
    layer1_outputs(1518) <= not(layer0_outputs(7938)) or (layer0_outputs(9796));
    layer1_outputs(1519) <= not((layer0_outputs(2324)) or (layer0_outputs(8303)));
    layer1_outputs(1520) <= not((layer0_outputs(6683)) or (layer0_outputs(174)));
    layer1_outputs(1521) <= not(layer0_outputs(3321)) or (layer0_outputs(7008));
    layer1_outputs(1522) <= layer0_outputs(421);
    layer1_outputs(1523) <= (layer0_outputs(6133)) and (layer0_outputs(2422));
    layer1_outputs(1524) <= '1';
    layer1_outputs(1525) <= not(layer0_outputs(2077)) or (layer0_outputs(3356));
    layer1_outputs(1526) <= (layer0_outputs(6534)) xor (layer0_outputs(4388));
    layer1_outputs(1527) <= layer0_outputs(7182);
    layer1_outputs(1528) <= not((layer0_outputs(7967)) xor (layer0_outputs(8601)));
    layer1_outputs(1529) <= not(layer0_outputs(3870));
    layer1_outputs(1530) <= not((layer0_outputs(2522)) or (layer0_outputs(8755)));
    layer1_outputs(1531) <= layer0_outputs(3796);
    layer1_outputs(1532) <= (layer0_outputs(1869)) or (layer0_outputs(6134));
    layer1_outputs(1533) <= not((layer0_outputs(6173)) or (layer0_outputs(1435)));
    layer1_outputs(1534) <= layer0_outputs(6842);
    layer1_outputs(1535) <= (layer0_outputs(8446)) and not (layer0_outputs(534));
    layer1_outputs(1536) <= layer0_outputs(1387);
    layer1_outputs(1537) <= not(layer0_outputs(5734));
    layer1_outputs(1538) <= not(layer0_outputs(8695));
    layer1_outputs(1539) <= (layer0_outputs(9133)) xor (layer0_outputs(1452));
    layer1_outputs(1540) <= (layer0_outputs(1015)) xor (layer0_outputs(5542));
    layer1_outputs(1541) <= not(layer0_outputs(8024)) or (layer0_outputs(3215));
    layer1_outputs(1542) <= not((layer0_outputs(3714)) or (layer0_outputs(2670)));
    layer1_outputs(1543) <= not(layer0_outputs(6135)) or (layer0_outputs(4466));
    layer1_outputs(1544) <= not(layer0_outputs(657));
    layer1_outputs(1545) <= not(layer0_outputs(2952));
    layer1_outputs(1546) <= layer0_outputs(6805);
    layer1_outputs(1547) <= layer0_outputs(4959);
    layer1_outputs(1548) <= (layer0_outputs(8148)) and (layer0_outputs(5361));
    layer1_outputs(1549) <= layer0_outputs(8612);
    layer1_outputs(1550) <= layer0_outputs(8713);
    layer1_outputs(1551) <= not(layer0_outputs(5843));
    layer1_outputs(1552) <= (layer0_outputs(9367)) and not (layer0_outputs(1667));
    layer1_outputs(1553) <= not(layer0_outputs(7735)) or (layer0_outputs(8620));
    layer1_outputs(1554) <= not(layer0_outputs(6580)) or (layer0_outputs(8709));
    layer1_outputs(1555) <= (layer0_outputs(9753)) and not (layer0_outputs(5737));
    layer1_outputs(1556) <= not(layer0_outputs(7546)) or (layer0_outputs(6440));
    layer1_outputs(1557) <= (layer0_outputs(7006)) and not (layer0_outputs(10024));
    layer1_outputs(1558) <= layer0_outputs(1502);
    layer1_outputs(1559) <= (layer0_outputs(8211)) xor (layer0_outputs(961));
    layer1_outputs(1560) <= (layer0_outputs(10226)) and (layer0_outputs(7172));
    layer1_outputs(1561) <= not(layer0_outputs(7508));
    layer1_outputs(1562) <= layer0_outputs(1976);
    layer1_outputs(1563) <= not(layer0_outputs(4811)) or (layer0_outputs(9764));
    layer1_outputs(1564) <= (layer0_outputs(339)) or (layer0_outputs(3006));
    layer1_outputs(1565) <= not(layer0_outputs(1107)) or (layer0_outputs(6144));
    layer1_outputs(1566) <= layer0_outputs(8536);
    layer1_outputs(1567) <= (layer0_outputs(4461)) and not (layer0_outputs(4428));
    layer1_outputs(1568) <= not((layer0_outputs(1472)) and (layer0_outputs(7921)));
    layer1_outputs(1569) <= layer0_outputs(7525);
    layer1_outputs(1570) <= not(layer0_outputs(2945)) or (layer0_outputs(3416));
    layer1_outputs(1571) <= not(layer0_outputs(7166));
    layer1_outputs(1572) <= not(layer0_outputs(7171));
    layer1_outputs(1573) <= '1';
    layer1_outputs(1574) <= not((layer0_outputs(5710)) or (layer0_outputs(10165)));
    layer1_outputs(1575) <= (layer0_outputs(7752)) and not (layer0_outputs(8102));
    layer1_outputs(1576) <= layer0_outputs(2977);
    layer1_outputs(1577) <= not(layer0_outputs(895)) or (layer0_outputs(9230));
    layer1_outputs(1578) <= (layer0_outputs(10140)) and not (layer0_outputs(2291));
    layer1_outputs(1579) <= layer0_outputs(4129);
    layer1_outputs(1580) <= layer0_outputs(1583);
    layer1_outputs(1581) <= not(layer0_outputs(1843)) or (layer0_outputs(570));
    layer1_outputs(1582) <= (layer0_outputs(3449)) or (layer0_outputs(3797));
    layer1_outputs(1583) <= not(layer0_outputs(4165));
    layer1_outputs(1584) <= (layer0_outputs(2954)) and not (layer0_outputs(1737));
    layer1_outputs(1585) <= not(layer0_outputs(8455));
    layer1_outputs(1586) <= not(layer0_outputs(9017));
    layer1_outputs(1587) <= layer0_outputs(3992);
    layer1_outputs(1588) <= (layer0_outputs(8689)) or (layer0_outputs(9052));
    layer1_outputs(1589) <= not((layer0_outputs(694)) and (layer0_outputs(3565)));
    layer1_outputs(1590) <= layer0_outputs(2004);
    layer1_outputs(1591) <= not(layer0_outputs(3392));
    layer1_outputs(1592) <= not(layer0_outputs(5473)) or (layer0_outputs(9698));
    layer1_outputs(1593) <= (layer0_outputs(5062)) or (layer0_outputs(4014));
    layer1_outputs(1594) <= layer0_outputs(10154);
    layer1_outputs(1595) <= (layer0_outputs(5735)) and not (layer0_outputs(4037));
    layer1_outputs(1596) <= not(layer0_outputs(8170));
    layer1_outputs(1597) <= (layer0_outputs(8718)) or (layer0_outputs(4767));
    layer1_outputs(1598) <= not(layer0_outputs(5584)) or (layer0_outputs(7781));
    layer1_outputs(1599) <= layer0_outputs(4852);
    layer1_outputs(1600) <= (layer0_outputs(6652)) and not (layer0_outputs(1728));
    layer1_outputs(1601) <= not((layer0_outputs(2000)) and (layer0_outputs(4667)));
    layer1_outputs(1602) <= layer0_outputs(3017);
    layer1_outputs(1603) <= not((layer0_outputs(2194)) and (layer0_outputs(9740)));
    layer1_outputs(1604) <= not(layer0_outputs(233));
    layer1_outputs(1605) <= layer0_outputs(5647);
    layer1_outputs(1606) <= layer0_outputs(3255);
    layer1_outputs(1607) <= not((layer0_outputs(3319)) or (layer0_outputs(9212)));
    layer1_outputs(1608) <= layer0_outputs(7811);
    layer1_outputs(1609) <= (layer0_outputs(8661)) and not (layer0_outputs(8730));
    layer1_outputs(1610) <= not(layer0_outputs(6106)) or (layer0_outputs(3468));
    layer1_outputs(1611) <= layer0_outputs(3178);
    layer1_outputs(1612) <= (layer0_outputs(2005)) and (layer0_outputs(7626));
    layer1_outputs(1613) <= layer0_outputs(1871);
    layer1_outputs(1614) <= layer0_outputs(146);
    layer1_outputs(1615) <= '1';
    layer1_outputs(1616) <= (layer0_outputs(1025)) and (layer0_outputs(3134));
    layer1_outputs(1617) <= (layer0_outputs(9583)) or (layer0_outputs(8841));
    layer1_outputs(1618) <= (layer0_outputs(6253)) or (layer0_outputs(9059));
    layer1_outputs(1619) <= layer0_outputs(3925);
    layer1_outputs(1620) <= (layer0_outputs(7711)) and (layer0_outputs(1275));
    layer1_outputs(1621) <= not((layer0_outputs(9723)) xor (layer0_outputs(5770)));
    layer1_outputs(1622) <= (layer0_outputs(8024)) and not (layer0_outputs(3110));
    layer1_outputs(1623) <= (layer0_outputs(2445)) xor (layer0_outputs(10131));
    layer1_outputs(1624) <= not(layer0_outputs(182));
    layer1_outputs(1625) <= (layer0_outputs(6444)) and (layer0_outputs(9308));
    layer1_outputs(1626) <= '0';
    layer1_outputs(1627) <= not((layer0_outputs(4054)) or (layer0_outputs(3447)));
    layer1_outputs(1628) <= layer0_outputs(825);
    layer1_outputs(1629) <= (layer0_outputs(7432)) or (layer0_outputs(3279));
    layer1_outputs(1630) <= not(layer0_outputs(8900)) or (layer0_outputs(2460));
    layer1_outputs(1631) <= layer0_outputs(8970);
    layer1_outputs(1632) <= not(layer0_outputs(6959)) or (layer0_outputs(6996));
    layer1_outputs(1633) <= (layer0_outputs(8014)) or (layer0_outputs(2040));
    layer1_outputs(1634) <= not(layer0_outputs(5621)) or (layer0_outputs(5077));
    layer1_outputs(1635) <= not(layer0_outputs(9127));
    layer1_outputs(1636) <= not(layer0_outputs(6328));
    layer1_outputs(1637) <= (layer0_outputs(4372)) xor (layer0_outputs(2077));
    layer1_outputs(1638) <= not(layer0_outputs(2933)) or (layer0_outputs(9409));
    layer1_outputs(1639) <= (layer0_outputs(6480)) and (layer0_outputs(8679));
    layer1_outputs(1640) <= layer0_outputs(232);
    layer1_outputs(1641) <= not(layer0_outputs(2069));
    layer1_outputs(1642) <= '0';
    layer1_outputs(1643) <= (layer0_outputs(6606)) and not (layer0_outputs(4058));
    layer1_outputs(1644) <= '0';
    layer1_outputs(1645) <= (layer0_outputs(4528)) and not (layer0_outputs(7105));
    layer1_outputs(1646) <= (layer0_outputs(4086)) xor (layer0_outputs(9182));
    layer1_outputs(1647) <= not((layer0_outputs(5524)) xor (layer0_outputs(577)));
    layer1_outputs(1648) <= not(layer0_outputs(6662)) or (layer0_outputs(486));
    layer1_outputs(1649) <= not(layer0_outputs(290));
    layer1_outputs(1650) <= layer0_outputs(9983);
    layer1_outputs(1651) <= not(layer0_outputs(2193));
    layer1_outputs(1652) <= not(layer0_outputs(2468)) or (layer0_outputs(1998));
    layer1_outputs(1653) <= layer0_outputs(4453);
    layer1_outputs(1654) <= not((layer0_outputs(8457)) xor (layer0_outputs(483)));
    layer1_outputs(1655) <= (layer0_outputs(3036)) and (layer0_outputs(10086));
    layer1_outputs(1656) <= not((layer0_outputs(9637)) and (layer0_outputs(1543)));
    layer1_outputs(1657) <= not(layer0_outputs(1865)) or (layer0_outputs(9881));
    layer1_outputs(1658) <= not(layer0_outputs(5616));
    layer1_outputs(1659) <= not(layer0_outputs(970));
    layer1_outputs(1660) <= '1';
    layer1_outputs(1661) <= not((layer0_outputs(9058)) or (layer0_outputs(5839)));
    layer1_outputs(1662) <= (layer0_outputs(914)) and not (layer0_outputs(4172));
    layer1_outputs(1663) <= not((layer0_outputs(9657)) and (layer0_outputs(9022)));
    layer1_outputs(1664) <= '1';
    layer1_outputs(1665) <= not(layer0_outputs(7057));
    layer1_outputs(1666) <= not(layer0_outputs(8083)) or (layer0_outputs(7529));
    layer1_outputs(1667) <= (layer0_outputs(9862)) and (layer0_outputs(1659));
    layer1_outputs(1668) <= not((layer0_outputs(4137)) and (layer0_outputs(412)));
    layer1_outputs(1669) <= (layer0_outputs(2978)) or (layer0_outputs(2971));
    layer1_outputs(1670) <= not(layer0_outputs(8734));
    layer1_outputs(1671) <= not(layer0_outputs(2555)) or (layer0_outputs(6155));
    layer1_outputs(1672) <= (layer0_outputs(722)) and (layer0_outputs(5500));
    layer1_outputs(1673) <= not((layer0_outputs(7443)) or (layer0_outputs(8492)));
    layer1_outputs(1674) <= not(layer0_outputs(5913));
    layer1_outputs(1675) <= not((layer0_outputs(5934)) and (layer0_outputs(3141)));
    layer1_outputs(1676) <= layer0_outputs(2547);
    layer1_outputs(1677) <= not(layer0_outputs(977)) or (layer0_outputs(8481));
    layer1_outputs(1678) <= layer0_outputs(2315);
    layer1_outputs(1679) <= layer0_outputs(5582);
    layer1_outputs(1680) <= not(layer0_outputs(4395)) or (layer0_outputs(4942));
    layer1_outputs(1681) <= not((layer0_outputs(183)) or (layer0_outputs(6345)));
    layer1_outputs(1682) <= not(layer0_outputs(649));
    layer1_outputs(1683) <= (layer0_outputs(349)) and not (layer0_outputs(10086));
    layer1_outputs(1684) <= not(layer0_outputs(3937));
    layer1_outputs(1685) <= not(layer0_outputs(1631));
    layer1_outputs(1686) <= not((layer0_outputs(252)) and (layer0_outputs(2299)));
    layer1_outputs(1687) <= (layer0_outputs(6735)) and not (layer0_outputs(9572));
    layer1_outputs(1688) <= not(layer0_outputs(4672));
    layer1_outputs(1689) <= not((layer0_outputs(8149)) or (layer0_outputs(4934)));
    layer1_outputs(1690) <= not(layer0_outputs(3119));
    layer1_outputs(1691) <= layer0_outputs(3477);
    layer1_outputs(1692) <= (layer0_outputs(2242)) and (layer0_outputs(7068));
    layer1_outputs(1693) <= not((layer0_outputs(9538)) xor (layer0_outputs(3897)));
    layer1_outputs(1694) <= not(layer0_outputs(970));
    layer1_outputs(1695) <= not((layer0_outputs(7817)) xor (layer0_outputs(10081)));
    layer1_outputs(1696) <= layer0_outputs(3687);
    layer1_outputs(1697) <= not((layer0_outputs(10158)) xor (layer0_outputs(7737)));
    layer1_outputs(1698) <= layer0_outputs(869);
    layer1_outputs(1699) <= not(layer0_outputs(10039)) or (layer0_outputs(4237));
    layer1_outputs(1700) <= (layer0_outputs(2060)) and not (layer0_outputs(9378));
    layer1_outputs(1701) <= layer0_outputs(6268);
    layer1_outputs(1702) <= layer0_outputs(4622);
    layer1_outputs(1703) <= not((layer0_outputs(5694)) and (layer0_outputs(4492)));
    layer1_outputs(1704) <= layer0_outputs(1960);
    layer1_outputs(1705) <= layer0_outputs(7390);
    layer1_outputs(1706) <= not(layer0_outputs(219));
    layer1_outputs(1707) <= not((layer0_outputs(6112)) xor (layer0_outputs(5366)));
    layer1_outputs(1708) <= layer0_outputs(6161);
    layer1_outputs(1709) <= (layer0_outputs(3806)) and (layer0_outputs(246));
    layer1_outputs(1710) <= (layer0_outputs(5984)) or (layer0_outputs(2504));
    layer1_outputs(1711) <= layer0_outputs(4007);
    layer1_outputs(1712) <= not(layer0_outputs(4755));
    layer1_outputs(1713) <= (layer0_outputs(2587)) xor (layer0_outputs(5281));
    layer1_outputs(1714) <= not(layer0_outputs(1162));
    layer1_outputs(1715) <= not(layer0_outputs(5303));
    layer1_outputs(1716) <= not(layer0_outputs(4762));
    layer1_outputs(1717) <= layer0_outputs(3373);
    layer1_outputs(1718) <= not(layer0_outputs(4029)) or (layer0_outputs(2820));
    layer1_outputs(1719) <= not((layer0_outputs(1165)) and (layer0_outputs(658)));
    layer1_outputs(1720) <= not(layer0_outputs(5308)) or (layer0_outputs(3142));
    layer1_outputs(1721) <= not(layer0_outputs(4676));
    layer1_outputs(1722) <= not(layer0_outputs(9483));
    layer1_outputs(1723) <= (layer0_outputs(1834)) and not (layer0_outputs(4498));
    layer1_outputs(1724) <= (layer0_outputs(3180)) xor (layer0_outputs(6995));
    layer1_outputs(1725) <= (layer0_outputs(6497)) and not (layer0_outputs(4310));
    layer1_outputs(1726) <= (layer0_outputs(4986)) and not (layer0_outputs(2920));
    layer1_outputs(1727) <= not(layer0_outputs(7274));
    layer1_outputs(1728) <= '0';
    layer1_outputs(1729) <= not(layer0_outputs(354));
    layer1_outputs(1730) <= (layer0_outputs(1115)) or (layer0_outputs(5645));
    layer1_outputs(1731) <= (layer0_outputs(3858)) and not (layer0_outputs(6669));
    layer1_outputs(1732) <= not((layer0_outputs(6075)) or (layer0_outputs(9403)));
    layer1_outputs(1733) <= layer0_outputs(5014);
    layer1_outputs(1734) <= layer0_outputs(8058);
    layer1_outputs(1735) <= not(layer0_outputs(6594));
    layer1_outputs(1736) <= (layer0_outputs(1928)) or (layer0_outputs(4256));
    layer1_outputs(1737) <= '1';
    layer1_outputs(1738) <= not((layer0_outputs(158)) xor (layer0_outputs(990)));
    layer1_outputs(1739) <= layer0_outputs(4502);
    layer1_outputs(1740) <= layer0_outputs(9171);
    layer1_outputs(1741) <= not((layer0_outputs(5845)) or (layer0_outputs(2663)));
    layer1_outputs(1742) <= not(layer0_outputs(2890)) or (layer0_outputs(8305));
    layer1_outputs(1743) <= not((layer0_outputs(9019)) or (layer0_outputs(8232)));
    layer1_outputs(1744) <= not(layer0_outputs(1533));
    layer1_outputs(1745) <= not(layer0_outputs(4674));
    layer1_outputs(1746) <= not((layer0_outputs(153)) xor (layer0_outputs(3986)));
    layer1_outputs(1747) <= not(layer0_outputs(316));
    layer1_outputs(1748) <= layer0_outputs(8052);
    layer1_outputs(1749) <= (layer0_outputs(8546)) and (layer0_outputs(2836));
    layer1_outputs(1750) <= (layer0_outputs(5315)) xor (layer0_outputs(1191));
    layer1_outputs(1751) <= not((layer0_outputs(3414)) or (layer0_outputs(2694)));
    layer1_outputs(1752) <= (layer0_outputs(5238)) and not (layer0_outputs(2544));
    layer1_outputs(1753) <= (layer0_outputs(138)) and not (layer0_outputs(2406));
    layer1_outputs(1754) <= (layer0_outputs(8356)) or (layer0_outputs(9682));
    layer1_outputs(1755) <= not((layer0_outputs(7497)) and (layer0_outputs(269)));
    layer1_outputs(1756) <= (layer0_outputs(488)) and (layer0_outputs(2833));
    layer1_outputs(1757) <= layer0_outputs(3021);
    layer1_outputs(1758) <= not(layer0_outputs(3678));
    layer1_outputs(1759) <= (layer0_outputs(7722)) or (layer0_outputs(6306));
    layer1_outputs(1760) <= (layer0_outputs(7210)) and not (layer0_outputs(5635));
    layer1_outputs(1761) <= (layer0_outputs(6025)) and not (layer0_outputs(9254));
    layer1_outputs(1762) <= not(layer0_outputs(7957)) or (layer0_outputs(2282));
    layer1_outputs(1763) <= layer0_outputs(747);
    layer1_outputs(1764) <= not((layer0_outputs(9608)) xor (layer0_outputs(4938)));
    layer1_outputs(1765) <= not(layer0_outputs(8997)) or (layer0_outputs(2086));
    layer1_outputs(1766) <= (layer0_outputs(8875)) and not (layer0_outputs(2462));
    layer1_outputs(1767) <= not(layer0_outputs(2227)) or (layer0_outputs(7189));
    layer1_outputs(1768) <= layer0_outputs(2506);
    layer1_outputs(1769) <= (layer0_outputs(5201)) and (layer0_outputs(7044));
    layer1_outputs(1770) <= not(layer0_outputs(122));
    layer1_outputs(1771) <= layer0_outputs(3247);
    layer1_outputs(1772) <= (layer0_outputs(1763)) or (layer0_outputs(9702));
    layer1_outputs(1773) <= not(layer0_outputs(3928));
    layer1_outputs(1774) <= not((layer0_outputs(3276)) or (layer0_outputs(7527)));
    layer1_outputs(1775) <= not((layer0_outputs(9677)) or (layer0_outputs(1619)));
    layer1_outputs(1776) <= not(layer0_outputs(10030));
    layer1_outputs(1777) <= not(layer0_outputs(1084));
    layer1_outputs(1778) <= not((layer0_outputs(4667)) xor (layer0_outputs(7386)));
    layer1_outputs(1779) <= layer0_outputs(8061);
    layer1_outputs(1780) <= not(layer0_outputs(6804));
    layer1_outputs(1781) <= not(layer0_outputs(1655)) or (layer0_outputs(7391));
    layer1_outputs(1782) <= not(layer0_outputs(2126));
    layer1_outputs(1783) <= (layer0_outputs(245)) or (layer0_outputs(6405));
    layer1_outputs(1784) <= not(layer0_outputs(7412));
    layer1_outputs(1785) <= not(layer0_outputs(274)) or (layer0_outputs(4754));
    layer1_outputs(1786) <= (layer0_outputs(2247)) or (layer0_outputs(2283));
    layer1_outputs(1787) <= layer0_outputs(1379);
    layer1_outputs(1788) <= not(layer0_outputs(1653));
    layer1_outputs(1789) <= '1';
    layer1_outputs(1790) <= (layer0_outputs(402)) and not (layer0_outputs(2127));
    layer1_outputs(1791) <= not((layer0_outputs(9826)) and (layer0_outputs(7526)));
    layer1_outputs(1792) <= not((layer0_outputs(2789)) or (layer0_outputs(1891)));
    layer1_outputs(1793) <= layer0_outputs(1749);
    layer1_outputs(1794) <= not(layer0_outputs(3439)) or (layer0_outputs(10027));
    layer1_outputs(1795) <= layer0_outputs(1740);
    layer1_outputs(1796) <= (layer0_outputs(407)) and not (layer0_outputs(2248));
    layer1_outputs(1797) <= layer0_outputs(4304);
    layer1_outputs(1798) <= not(layer0_outputs(5781)) or (layer0_outputs(1252));
    layer1_outputs(1799) <= not((layer0_outputs(9352)) xor (layer0_outputs(9852)));
    layer1_outputs(1800) <= not(layer0_outputs(5884));
    layer1_outputs(1801) <= (layer0_outputs(5534)) and (layer0_outputs(8054));
    layer1_outputs(1802) <= (layer0_outputs(7914)) or (layer0_outputs(3550));
    layer1_outputs(1803) <= not(layer0_outputs(3760));
    layer1_outputs(1804) <= (layer0_outputs(7726)) or (layer0_outputs(5296));
    layer1_outputs(1805) <= (layer0_outputs(5372)) xor (layer0_outputs(10172));
    layer1_outputs(1806) <= (layer0_outputs(6948)) and not (layer0_outputs(4399));
    layer1_outputs(1807) <= not(layer0_outputs(8879));
    layer1_outputs(1808) <= (layer0_outputs(4840)) and not (layer0_outputs(6019));
    layer1_outputs(1809) <= '0';
    layer1_outputs(1810) <= layer0_outputs(4560);
    layer1_outputs(1811) <= not(layer0_outputs(1133));
    layer1_outputs(1812) <= '1';
    layer1_outputs(1813) <= layer0_outputs(4914);
    layer1_outputs(1814) <= (layer0_outputs(9859)) and not (layer0_outputs(2985));
    layer1_outputs(1815) <= not((layer0_outputs(7896)) or (layer0_outputs(3387)));
    layer1_outputs(1816) <= layer0_outputs(1804);
    layer1_outputs(1817) <= (layer0_outputs(114)) and (layer0_outputs(7771));
    layer1_outputs(1818) <= layer0_outputs(4294);
    layer1_outputs(1819) <= not(layer0_outputs(8706));
    layer1_outputs(1820) <= (layer0_outputs(4653)) and (layer0_outputs(4965));
    layer1_outputs(1821) <= not(layer0_outputs(9106));
    layer1_outputs(1822) <= not(layer0_outputs(1665));
    layer1_outputs(1823) <= not(layer0_outputs(780));
    layer1_outputs(1824) <= not(layer0_outputs(581));
    layer1_outputs(1825) <= (layer0_outputs(5328)) and not (layer0_outputs(3343));
    layer1_outputs(1826) <= not((layer0_outputs(1828)) xor (layer0_outputs(7618)));
    layer1_outputs(1827) <= not((layer0_outputs(2387)) or (layer0_outputs(5916)));
    layer1_outputs(1828) <= layer0_outputs(2356);
    layer1_outputs(1829) <= not(layer0_outputs(507));
    layer1_outputs(1830) <= (layer0_outputs(3900)) and not (layer0_outputs(9767));
    layer1_outputs(1831) <= not(layer0_outputs(4272));
    layer1_outputs(1832) <= (layer0_outputs(6686)) or (layer0_outputs(7983));
    layer1_outputs(1833) <= (layer0_outputs(8373)) and not (layer0_outputs(2115));
    layer1_outputs(1834) <= not(layer0_outputs(4315));
    layer1_outputs(1835) <= not((layer0_outputs(3401)) xor (layer0_outputs(2603)));
    layer1_outputs(1836) <= '0';
    layer1_outputs(1837) <= (layer0_outputs(4418)) and (layer0_outputs(7708));
    layer1_outputs(1838) <= (layer0_outputs(8183)) and (layer0_outputs(2138));
    layer1_outputs(1839) <= layer0_outputs(8895);
    layer1_outputs(1840) <= layer0_outputs(2028);
    layer1_outputs(1841) <= layer0_outputs(4049);
    layer1_outputs(1842) <= (layer0_outputs(902)) and (layer0_outputs(9072));
    layer1_outputs(1843) <= not(layer0_outputs(4175));
    layer1_outputs(1844) <= (layer0_outputs(8443)) xor (layer0_outputs(1434));
    layer1_outputs(1845) <= layer0_outputs(5326);
    layer1_outputs(1846) <= not((layer0_outputs(6181)) and (layer0_outputs(6360)));
    layer1_outputs(1847) <= not(layer0_outputs(1130));
    layer1_outputs(1848) <= not((layer0_outputs(4080)) or (layer0_outputs(3525)));
    layer1_outputs(1849) <= not(layer0_outputs(5318));
    layer1_outputs(1850) <= not(layer0_outputs(3356));
    layer1_outputs(1851) <= not(layer0_outputs(6207));
    layer1_outputs(1852) <= not(layer0_outputs(5468)) or (layer0_outputs(3396));
    layer1_outputs(1853) <= not(layer0_outputs(10051));
    layer1_outputs(1854) <= not(layer0_outputs(5865));
    layer1_outputs(1855) <= '1';
    layer1_outputs(1856) <= not((layer0_outputs(1562)) or (layer0_outputs(9166)));
    layer1_outputs(1857) <= (layer0_outputs(7666)) and (layer0_outputs(8500));
    layer1_outputs(1858) <= not(layer0_outputs(3359));
    layer1_outputs(1859) <= layer0_outputs(6476);
    layer1_outputs(1860) <= not(layer0_outputs(3719)) or (layer0_outputs(642));
    layer1_outputs(1861) <= (layer0_outputs(9382)) and (layer0_outputs(6005));
    layer1_outputs(1862) <= (layer0_outputs(7733)) and (layer0_outputs(8623));
    layer1_outputs(1863) <= layer0_outputs(5435);
    layer1_outputs(1864) <= not(layer0_outputs(3822));
    layer1_outputs(1865) <= not(layer0_outputs(5340));
    layer1_outputs(1866) <= (layer0_outputs(2042)) xor (layer0_outputs(1972));
    layer1_outputs(1867) <= not(layer0_outputs(3617));
    layer1_outputs(1868) <= not(layer0_outputs(9408)) or (layer0_outputs(6813));
    layer1_outputs(1869) <= (layer0_outputs(4055)) or (layer0_outputs(2372));
    layer1_outputs(1870) <= layer0_outputs(4062);
    layer1_outputs(1871) <= layer0_outputs(6634);
    layer1_outputs(1872) <= layer0_outputs(6837);
    layer1_outputs(1873) <= not((layer0_outputs(5950)) and (layer0_outputs(3631)));
    layer1_outputs(1874) <= not((layer0_outputs(2786)) or (layer0_outputs(8393)));
    layer1_outputs(1875) <= layer0_outputs(1196);
    layer1_outputs(1876) <= not((layer0_outputs(3839)) xor (layer0_outputs(7276)));
    layer1_outputs(1877) <= not(layer0_outputs(4177)) or (layer0_outputs(8267));
    layer1_outputs(1878) <= (layer0_outputs(9705)) xor (layer0_outputs(1498));
    layer1_outputs(1879) <= not(layer0_outputs(8056)) or (layer0_outputs(10192));
    layer1_outputs(1880) <= not(layer0_outputs(7961));
    layer1_outputs(1881) <= not((layer0_outputs(4564)) and (layer0_outputs(8323)));
    layer1_outputs(1882) <= not((layer0_outputs(4147)) or (layer0_outputs(5310)));
    layer1_outputs(1883) <= layer0_outputs(9486);
    layer1_outputs(1884) <= not((layer0_outputs(8482)) or (layer0_outputs(1834)));
    layer1_outputs(1885) <= (layer0_outputs(6044)) xor (layer0_outputs(5450));
    layer1_outputs(1886) <= not((layer0_outputs(9531)) and (layer0_outputs(1757)));
    layer1_outputs(1887) <= not(layer0_outputs(1426)) or (layer0_outputs(6958));
    layer1_outputs(1888) <= '1';
    layer1_outputs(1889) <= not((layer0_outputs(3670)) xor (layer0_outputs(3623)));
    layer1_outputs(1890) <= not((layer0_outputs(4620)) and (layer0_outputs(9166)));
    layer1_outputs(1891) <= layer0_outputs(7879);
    layer1_outputs(1892) <= not(layer0_outputs(4327)) or (layer0_outputs(1559));
    layer1_outputs(1893) <= not((layer0_outputs(5594)) xor (layer0_outputs(5899)));
    layer1_outputs(1894) <= (layer0_outputs(4886)) and not (layer0_outputs(5972));
    layer1_outputs(1895) <= not(layer0_outputs(615));
    layer1_outputs(1896) <= layer0_outputs(4368);
    layer1_outputs(1897) <= not((layer0_outputs(7872)) or (layer0_outputs(2400)));
    layer1_outputs(1898) <= (layer0_outputs(1724)) and not (layer0_outputs(3607));
    layer1_outputs(1899) <= layer0_outputs(2169);
    layer1_outputs(1900) <= (layer0_outputs(8992)) and (layer0_outputs(4246));
    layer1_outputs(1901) <= layer0_outputs(1100);
    layer1_outputs(1902) <= not(layer0_outputs(9043));
    layer1_outputs(1903) <= not((layer0_outputs(829)) and (layer0_outputs(4773)));
    layer1_outputs(1904) <= not(layer0_outputs(669));
    layer1_outputs(1905) <= not(layer0_outputs(9120));
    layer1_outputs(1906) <= layer0_outputs(9786);
    layer1_outputs(1907) <= not(layer0_outputs(5420));
    layer1_outputs(1908) <= not((layer0_outputs(5323)) and (layer0_outputs(1495)));
    layer1_outputs(1909) <= '0';
    layer1_outputs(1910) <= layer0_outputs(6431);
    layer1_outputs(1911) <= not(layer0_outputs(2998));
    layer1_outputs(1912) <= layer0_outputs(8846);
    layer1_outputs(1913) <= not(layer0_outputs(9857)) or (layer0_outputs(7938));
    layer1_outputs(1914) <= '0';
    layer1_outputs(1915) <= not(layer0_outputs(1015));
    layer1_outputs(1916) <= not(layer0_outputs(6769));
    layer1_outputs(1917) <= not((layer0_outputs(2830)) and (layer0_outputs(9151)));
    layer1_outputs(1918) <= (layer0_outputs(8265)) and (layer0_outputs(8893));
    layer1_outputs(1919) <= not((layer0_outputs(8424)) or (layer0_outputs(17)));
    layer1_outputs(1920) <= not(layer0_outputs(10103)) or (layer0_outputs(1143));
    layer1_outputs(1921) <= (layer0_outputs(3803)) and not (layer0_outputs(2311));
    layer1_outputs(1922) <= not(layer0_outputs(309));
    layer1_outputs(1923) <= (layer0_outputs(4728)) and not (layer0_outputs(9867));
    layer1_outputs(1924) <= not(layer0_outputs(7980));
    layer1_outputs(1925) <= not(layer0_outputs(6319)) or (layer0_outputs(9492));
    layer1_outputs(1926) <= (layer0_outputs(6132)) and not (layer0_outputs(7958));
    layer1_outputs(1927) <= (layer0_outputs(3209)) and not (layer0_outputs(6087));
    layer1_outputs(1928) <= layer0_outputs(5230);
    layer1_outputs(1929) <= layer0_outputs(790);
    layer1_outputs(1930) <= not(layer0_outputs(9425)) or (layer0_outputs(7258));
    layer1_outputs(1931) <= (layer0_outputs(2707)) xor (layer0_outputs(2336));
    layer1_outputs(1932) <= not(layer0_outputs(8394));
    layer1_outputs(1933) <= not(layer0_outputs(2853)) or (layer0_outputs(2245));
    layer1_outputs(1934) <= not(layer0_outputs(6264));
    layer1_outputs(1935) <= '0';
    layer1_outputs(1936) <= (layer0_outputs(6311)) and (layer0_outputs(10044));
    layer1_outputs(1937) <= layer0_outputs(5424);
    layer1_outputs(1938) <= (layer0_outputs(856)) and not (layer0_outputs(3248));
    layer1_outputs(1939) <= not(layer0_outputs(8007)) or (layer0_outputs(4180));
    layer1_outputs(1940) <= not(layer0_outputs(10184));
    layer1_outputs(1941) <= not((layer0_outputs(3237)) xor (layer0_outputs(3889)));
    layer1_outputs(1942) <= (layer0_outputs(9365)) and not (layer0_outputs(9133));
    layer1_outputs(1943) <= (layer0_outputs(6142)) and not (layer0_outputs(533));
    layer1_outputs(1944) <= (layer0_outputs(9324)) and not (layer0_outputs(3795));
    layer1_outputs(1945) <= not(layer0_outputs(9434));
    layer1_outputs(1946) <= not((layer0_outputs(43)) and (layer0_outputs(8091)));
    layer1_outputs(1947) <= not(layer0_outputs(8272)) or (layer0_outputs(2020));
    layer1_outputs(1948) <= not(layer0_outputs(6908));
    layer1_outputs(1949) <= (layer0_outputs(4330)) and not (layer0_outputs(7220));
    layer1_outputs(1950) <= (layer0_outputs(7284)) or (layer0_outputs(2998));
    layer1_outputs(1951) <= not((layer0_outputs(9786)) and (layer0_outputs(4660)));
    layer1_outputs(1952) <= (layer0_outputs(8186)) or (layer0_outputs(8354));
    layer1_outputs(1953) <= layer0_outputs(5208);
    layer1_outputs(1954) <= not(layer0_outputs(4057));
    layer1_outputs(1955) <= (layer0_outputs(5653)) or (layer0_outputs(6881));
    layer1_outputs(1956) <= (layer0_outputs(707)) xor (layer0_outputs(9275));
    layer1_outputs(1957) <= not((layer0_outputs(9757)) xor (layer0_outputs(6922)));
    layer1_outputs(1958) <= layer0_outputs(2056);
    layer1_outputs(1959) <= not((layer0_outputs(401)) xor (layer0_outputs(5881)));
    layer1_outputs(1960) <= not(layer0_outputs(321));
    layer1_outputs(1961) <= not((layer0_outputs(3317)) or (layer0_outputs(9663)));
    layer1_outputs(1962) <= not(layer0_outputs(7819));
    layer1_outputs(1963) <= (layer0_outputs(67)) and not (layer0_outputs(5411));
    layer1_outputs(1964) <= layer0_outputs(1076);
    layer1_outputs(1965) <= layer0_outputs(1603);
    layer1_outputs(1966) <= not(layer0_outputs(6089));
    layer1_outputs(1967) <= not(layer0_outputs(2260));
    layer1_outputs(1968) <= not(layer0_outputs(10109));
    layer1_outputs(1969) <= (layer0_outputs(8490)) and (layer0_outputs(299));
    layer1_outputs(1970) <= not((layer0_outputs(5029)) xor (layer0_outputs(1647)));
    layer1_outputs(1971) <= (layer0_outputs(8787)) and (layer0_outputs(9114));
    layer1_outputs(1972) <= (layer0_outputs(9529)) and (layer0_outputs(9073));
    layer1_outputs(1973) <= layer0_outputs(4215);
    layer1_outputs(1974) <= layer0_outputs(1865);
    layer1_outputs(1975) <= layer0_outputs(378);
    layer1_outputs(1976) <= layer0_outputs(7238);
    layer1_outputs(1977) <= (layer0_outputs(6265)) and (layer0_outputs(5430));
    layer1_outputs(1978) <= not(layer0_outputs(4029));
    layer1_outputs(1979) <= (layer0_outputs(4061)) and (layer0_outputs(3464));
    layer1_outputs(1980) <= not((layer0_outputs(3814)) xor (layer0_outputs(521)));
    layer1_outputs(1981) <= '1';
    layer1_outputs(1982) <= layer0_outputs(10195);
    layer1_outputs(1983) <= layer0_outputs(9745);
    layer1_outputs(1984) <= layer0_outputs(1689);
    layer1_outputs(1985) <= (layer0_outputs(8203)) or (layer0_outputs(5893));
    layer1_outputs(1986) <= (layer0_outputs(22)) or (layer0_outputs(9981));
    layer1_outputs(1987) <= (layer0_outputs(1026)) or (layer0_outputs(9622));
    layer1_outputs(1988) <= layer0_outputs(7848);
    layer1_outputs(1989) <= not((layer0_outputs(8755)) or (layer0_outputs(1808)));
    layer1_outputs(1990) <= layer0_outputs(6102);
    layer1_outputs(1991) <= not(layer0_outputs(8144)) or (layer0_outputs(7960));
    layer1_outputs(1992) <= layer0_outputs(5062);
    layer1_outputs(1993) <= not(layer0_outputs(3374));
    layer1_outputs(1994) <= not(layer0_outputs(9336));
    layer1_outputs(1995) <= not(layer0_outputs(6938)) or (layer0_outputs(5455));
    layer1_outputs(1996) <= (layer0_outputs(6287)) or (layer0_outputs(6024));
    layer1_outputs(1997) <= not(layer0_outputs(4457)) or (layer0_outputs(634));
    layer1_outputs(1998) <= not(layer0_outputs(4939)) or (layer0_outputs(1945));
    layer1_outputs(1999) <= not(layer0_outputs(8525));
    layer1_outputs(2000) <= (layer0_outputs(709)) and not (layer0_outputs(8168));
    layer1_outputs(2001) <= not((layer0_outputs(6815)) and (layer0_outputs(9563)));
    layer1_outputs(2002) <= (layer0_outputs(4398)) and (layer0_outputs(3729));
    layer1_outputs(2003) <= layer0_outputs(1212);
    layer1_outputs(2004) <= layer0_outputs(2320);
    layer1_outputs(2005) <= (layer0_outputs(6255)) or (layer0_outputs(1940));
    layer1_outputs(2006) <= '0';
    layer1_outputs(2007) <= layer0_outputs(832);
    layer1_outputs(2008) <= layer0_outputs(9428);
    layer1_outputs(2009) <= not(layer0_outputs(8105)) or (layer0_outputs(7029));
    layer1_outputs(2010) <= not(layer0_outputs(8789)) or (layer0_outputs(3233));
    layer1_outputs(2011) <= layer0_outputs(6184);
    layer1_outputs(2012) <= not(layer0_outputs(4602));
    layer1_outputs(2013) <= (layer0_outputs(723)) and not (layer0_outputs(3260));
    layer1_outputs(2014) <= not((layer0_outputs(738)) xor (layer0_outputs(8050)));
    layer1_outputs(2015) <= (layer0_outputs(4352)) and not (layer0_outputs(3946));
    layer1_outputs(2016) <= not(layer0_outputs(4459));
    layer1_outputs(2017) <= not((layer0_outputs(9550)) xor (layer0_outputs(939)));
    layer1_outputs(2018) <= not(layer0_outputs(4485));
    layer1_outputs(2019) <= not((layer0_outputs(5762)) and (layer0_outputs(6768)));
    layer1_outputs(2020) <= (layer0_outputs(3691)) and (layer0_outputs(8123));
    layer1_outputs(2021) <= (layer0_outputs(882)) or (layer0_outputs(4651));
    layer1_outputs(2022) <= not(layer0_outputs(6521));
    layer1_outputs(2023) <= layer0_outputs(2938);
    layer1_outputs(2024) <= not((layer0_outputs(7929)) and (layer0_outputs(1429)));
    layer1_outputs(2025) <= layer0_outputs(2939);
    layer1_outputs(2026) <= (layer0_outputs(3994)) and not (layer0_outputs(3862));
    layer1_outputs(2027) <= layer0_outputs(8930);
    layer1_outputs(2028) <= not(layer0_outputs(7404)) or (layer0_outputs(7124));
    layer1_outputs(2029) <= not(layer0_outputs(7866));
    layer1_outputs(2030) <= layer0_outputs(9082);
    layer1_outputs(2031) <= layer0_outputs(3938);
    layer1_outputs(2032) <= (layer0_outputs(6719)) xor (layer0_outputs(418));
    layer1_outputs(2033) <= not(layer0_outputs(8155)) or (layer0_outputs(8240));
    layer1_outputs(2034) <= not((layer0_outputs(7509)) and (layer0_outputs(2705)));
    layer1_outputs(2035) <= (layer0_outputs(10219)) xor (layer0_outputs(8955));
    layer1_outputs(2036) <= (layer0_outputs(2770)) xor (layer0_outputs(3784));
    layer1_outputs(2037) <= not(layer0_outputs(3370));
    layer1_outputs(2038) <= (layer0_outputs(1630)) or (layer0_outputs(4894));
    layer1_outputs(2039) <= '0';
    layer1_outputs(2040) <= (layer0_outputs(165)) and not (layer0_outputs(569));
    layer1_outputs(2041) <= not(layer0_outputs(2828));
    layer1_outputs(2042) <= (layer0_outputs(10068)) and not (layer0_outputs(8469));
    layer1_outputs(2043) <= not(layer0_outputs(6099));
    layer1_outputs(2044) <= layer0_outputs(8885);
    layer1_outputs(2045) <= not(layer0_outputs(985)) or (layer0_outputs(4579));
    layer1_outputs(2046) <= not(layer0_outputs(4144)) or (layer0_outputs(5197));
    layer1_outputs(2047) <= (layer0_outputs(3435)) and not (layer0_outputs(6648));
    layer1_outputs(2048) <= (layer0_outputs(3547)) xor (layer0_outputs(445));
    layer1_outputs(2049) <= not(layer0_outputs(5993)) or (layer0_outputs(5450));
    layer1_outputs(2050) <= not((layer0_outputs(3022)) and (layer0_outputs(3910)));
    layer1_outputs(2051) <= not((layer0_outputs(3156)) or (layer0_outputs(6702)));
    layer1_outputs(2052) <= layer0_outputs(2852);
    layer1_outputs(2053) <= layer0_outputs(8808);
    layer1_outputs(2054) <= not(layer0_outputs(5000));
    layer1_outputs(2055) <= not((layer0_outputs(8387)) or (layer0_outputs(7655)));
    layer1_outputs(2056) <= layer0_outputs(2525);
    layer1_outputs(2057) <= layer0_outputs(9231);
    layer1_outputs(2058) <= not(layer0_outputs(9706));
    layer1_outputs(2059) <= not(layer0_outputs(4248));
    layer1_outputs(2060) <= '1';
    layer1_outputs(2061) <= not((layer0_outputs(7474)) and (layer0_outputs(5209)));
    layer1_outputs(2062) <= not((layer0_outputs(7691)) and (layer0_outputs(6749)));
    layer1_outputs(2063) <= layer0_outputs(9270);
    layer1_outputs(2064) <= not((layer0_outputs(5722)) and (layer0_outputs(9671)));
    layer1_outputs(2065) <= '0';
    layer1_outputs(2066) <= (layer0_outputs(4036)) and not (layer0_outputs(8597));
    layer1_outputs(2067) <= (layer0_outputs(2141)) and (layer0_outputs(9668));
    layer1_outputs(2068) <= not(layer0_outputs(10190));
    layer1_outputs(2069) <= '1';
    layer1_outputs(2070) <= layer0_outputs(4683);
    layer1_outputs(2071) <= not((layer0_outputs(9281)) xor (layer0_outputs(6955)));
    layer1_outputs(2072) <= (layer0_outputs(5692)) and (layer0_outputs(7092));
    layer1_outputs(2073) <= (layer0_outputs(5746)) and not (layer0_outputs(2455));
    layer1_outputs(2074) <= layer0_outputs(5423);
    layer1_outputs(2075) <= not(layer0_outputs(4344));
    layer1_outputs(2076) <= (layer0_outputs(7302)) and not (layer0_outputs(426));
    layer1_outputs(2077) <= layer0_outputs(8802);
    layer1_outputs(2078) <= not((layer0_outputs(3194)) and (layer0_outputs(6834)));
    layer1_outputs(2079) <= not(layer0_outputs(398)) or (layer0_outputs(971));
    layer1_outputs(2080) <= '1';
    layer1_outputs(2081) <= (layer0_outputs(615)) and (layer0_outputs(5244));
    layer1_outputs(2082) <= not(layer0_outputs(358)) or (layer0_outputs(6860));
    layer1_outputs(2083) <= (layer0_outputs(3218)) or (layer0_outputs(1304));
    layer1_outputs(2084) <= layer0_outputs(6113);
    layer1_outputs(2085) <= not(layer0_outputs(3870)) or (layer0_outputs(3066));
    layer1_outputs(2086) <= layer0_outputs(697);
    layer1_outputs(2087) <= not(layer0_outputs(6864)) or (layer0_outputs(9301));
    layer1_outputs(2088) <= not((layer0_outputs(4514)) and (layer0_outputs(6490)));
    layer1_outputs(2089) <= not(layer0_outputs(7299));
    layer1_outputs(2090) <= layer0_outputs(1753);
    layer1_outputs(2091) <= not((layer0_outputs(2687)) or (layer0_outputs(6901)));
    layer1_outputs(2092) <= (layer0_outputs(8297)) and not (layer0_outputs(6061));
    layer1_outputs(2093) <= (layer0_outputs(8557)) and not (layer0_outputs(2269));
    layer1_outputs(2094) <= (layer0_outputs(7396)) and (layer0_outputs(2196));
    layer1_outputs(2095) <= not((layer0_outputs(5783)) and (layer0_outputs(8658)));
    layer1_outputs(2096) <= (layer0_outputs(8633)) and not (layer0_outputs(4849));
    layer1_outputs(2097) <= not(layer0_outputs(2862)) or (layer0_outputs(9401));
    layer1_outputs(2098) <= not(layer0_outputs(2707)) or (layer0_outputs(1359));
    layer1_outputs(2099) <= '1';
    layer1_outputs(2100) <= layer0_outputs(764);
    layer1_outputs(2101) <= (layer0_outputs(6052)) or (layer0_outputs(1078));
    layer1_outputs(2102) <= '0';
    layer1_outputs(2103) <= layer0_outputs(4640);
    layer1_outputs(2104) <= (layer0_outputs(9228)) or (layer0_outputs(189));
    layer1_outputs(2105) <= layer0_outputs(6814);
    layer1_outputs(2106) <= not(layer0_outputs(7595));
    layer1_outputs(2107) <= not((layer0_outputs(1338)) or (layer0_outputs(7107)));
    layer1_outputs(2108) <= not((layer0_outputs(9015)) and (layer0_outputs(7456)));
    layer1_outputs(2109) <= not((layer0_outputs(6663)) or (layer0_outputs(7670)));
    layer1_outputs(2110) <= not(layer0_outputs(738));
    layer1_outputs(2111) <= '1';
    layer1_outputs(2112) <= (layer0_outputs(1028)) and not (layer0_outputs(9322));
    layer1_outputs(2113) <= layer0_outputs(389);
    layer1_outputs(2114) <= (layer0_outputs(9255)) and not (layer0_outputs(3070));
    layer1_outputs(2115) <= not((layer0_outputs(1016)) and (layer0_outputs(9927)));
    layer1_outputs(2116) <= (layer0_outputs(3301)) and not (layer0_outputs(8911));
    layer1_outputs(2117) <= not((layer0_outputs(266)) and (layer0_outputs(8006)));
    layer1_outputs(2118) <= layer0_outputs(7316);
    layer1_outputs(2119) <= not(layer0_outputs(7021));
    layer1_outputs(2120) <= (layer0_outputs(7035)) and (layer0_outputs(8081));
    layer1_outputs(2121) <= (layer0_outputs(6753)) xor (layer0_outputs(8535));
    layer1_outputs(2122) <= (layer0_outputs(3344)) xor (layer0_outputs(3744));
    layer1_outputs(2123) <= not(layer0_outputs(9394));
    layer1_outputs(2124) <= not(layer0_outputs(7273)) or (layer0_outputs(7870));
    layer1_outputs(2125) <= not(layer0_outputs(6700));
    layer1_outputs(2126) <= layer0_outputs(5933);
    layer1_outputs(2127) <= not((layer0_outputs(384)) and (layer0_outputs(428)));
    layer1_outputs(2128) <= not(layer0_outputs(7115)) or (layer0_outputs(6914));
    layer1_outputs(2129) <= not(layer0_outputs(4704)) or (layer0_outputs(305));
    layer1_outputs(2130) <= not(layer0_outputs(7149)) or (layer0_outputs(8388));
    layer1_outputs(2131) <= layer0_outputs(3627);
    layer1_outputs(2132) <= (layer0_outputs(3589)) and not (layer0_outputs(9591));
    layer1_outputs(2133) <= (layer0_outputs(8548)) and not (layer0_outputs(1615));
    layer1_outputs(2134) <= not(layer0_outputs(2252));
    layer1_outputs(2135) <= (layer0_outputs(2068)) or (layer0_outputs(5445));
    layer1_outputs(2136) <= not(layer0_outputs(1390));
    layer1_outputs(2137) <= layer0_outputs(7920);
    layer1_outputs(2138) <= (layer0_outputs(5762)) and not (layer0_outputs(1915));
    layer1_outputs(2139) <= not(layer0_outputs(6475)) or (layer0_outputs(4557));
    layer1_outputs(2140) <= not(layer0_outputs(8514)) or (layer0_outputs(9204));
    layer1_outputs(2141) <= (layer0_outputs(2538)) and not (layer0_outputs(559));
    layer1_outputs(2142) <= not((layer0_outputs(248)) or (layer0_outputs(9325)));
    layer1_outputs(2143) <= not(layer0_outputs(9241));
    layer1_outputs(2144) <= '1';
    layer1_outputs(2145) <= not(layer0_outputs(7734)) or (layer0_outputs(5490));
    layer1_outputs(2146) <= (layer0_outputs(9180)) xor (layer0_outputs(4683));
    layer1_outputs(2147) <= layer0_outputs(783);
    layer1_outputs(2148) <= (layer0_outputs(6167)) and (layer0_outputs(6788));
    layer1_outputs(2149) <= (layer0_outputs(5519)) or (layer0_outputs(7637));
    layer1_outputs(2150) <= (layer0_outputs(4458)) and not (layer0_outputs(8151));
    layer1_outputs(2151) <= (layer0_outputs(8766)) or (layer0_outputs(208));
    layer1_outputs(2152) <= not((layer0_outputs(6590)) and (layer0_outputs(4645)));
    layer1_outputs(2153) <= layer0_outputs(10171);
    layer1_outputs(2154) <= not((layer0_outputs(7777)) or (layer0_outputs(6916)));
    layer1_outputs(2155) <= not(layer0_outputs(5472)) or (layer0_outputs(551));
    layer1_outputs(2156) <= layer0_outputs(75);
    layer1_outputs(2157) <= '0';
    layer1_outputs(2158) <= layer0_outputs(10051);
    layer1_outputs(2159) <= not(layer0_outputs(6531)) or (layer0_outputs(4342));
    layer1_outputs(2160) <= layer0_outputs(1103);
    layer1_outputs(2161) <= not((layer0_outputs(10134)) xor (layer0_outputs(8019)));
    layer1_outputs(2162) <= layer0_outputs(6559);
    layer1_outputs(2163) <= not((layer0_outputs(5924)) and (layer0_outputs(5922)));
    layer1_outputs(2164) <= layer0_outputs(2044);
    layer1_outputs(2165) <= not(layer0_outputs(8615));
    layer1_outputs(2166) <= not(layer0_outputs(9296));
    layer1_outputs(2167) <= '0';
    layer1_outputs(2168) <= layer0_outputs(2931);
    layer1_outputs(2169) <= not(layer0_outputs(2318)) or (layer0_outputs(6872));
    layer1_outputs(2170) <= not((layer0_outputs(3343)) or (layer0_outputs(5903)));
    layer1_outputs(2171) <= '1';
    layer1_outputs(2172) <= not((layer0_outputs(8857)) or (layer0_outputs(2398)));
    layer1_outputs(2173) <= (layer0_outputs(6548)) and (layer0_outputs(108));
    layer1_outputs(2174) <= (layer0_outputs(1282)) xor (layer0_outputs(2093));
    layer1_outputs(2175) <= not(layer0_outputs(6252)) or (layer0_outputs(6521));
    layer1_outputs(2176) <= not((layer0_outputs(1866)) and (layer0_outputs(2596)));
    layer1_outputs(2177) <= (layer0_outputs(7093)) xor (layer0_outputs(7335));
    layer1_outputs(2178) <= not(layer0_outputs(4584));
    layer1_outputs(2179) <= not(layer0_outputs(2912)) or (layer0_outputs(10093));
    layer1_outputs(2180) <= not(layer0_outputs(6827));
    layer1_outputs(2181) <= not((layer0_outputs(5581)) and (layer0_outputs(2200)));
    layer1_outputs(2182) <= not(layer0_outputs(4515));
    layer1_outputs(2183) <= not(layer0_outputs(3586)) or (layer0_outputs(1246));
    layer1_outputs(2184) <= not(layer0_outputs(5664));
    layer1_outputs(2185) <= (layer0_outputs(3479)) and not (layer0_outputs(1532));
    layer1_outputs(2186) <= layer0_outputs(4529);
    layer1_outputs(2187) <= not((layer0_outputs(2304)) xor (layer0_outputs(6069)));
    layer1_outputs(2188) <= not(layer0_outputs(505));
    layer1_outputs(2189) <= not(layer0_outputs(7966));
    layer1_outputs(2190) <= not(layer0_outputs(1270)) or (layer0_outputs(8721));
    layer1_outputs(2191) <= not((layer0_outputs(4919)) and (layer0_outputs(1674)));
    layer1_outputs(2192) <= not(layer0_outputs(7203));
    layer1_outputs(2193) <= not(layer0_outputs(3459));
    layer1_outputs(2194) <= not(layer0_outputs(2642));
    layer1_outputs(2195) <= layer0_outputs(3510);
    layer1_outputs(2196) <= not((layer0_outputs(8423)) and (layer0_outputs(3833)));
    layer1_outputs(2197) <= not(layer0_outputs(6123));
    layer1_outputs(2198) <= not(layer0_outputs(2919));
    layer1_outputs(2199) <= not((layer0_outputs(3143)) xor (layer0_outputs(4535)));
    layer1_outputs(2200) <= (layer0_outputs(7164)) or (layer0_outputs(9738));
    layer1_outputs(2201) <= not((layer0_outputs(1729)) xor (layer0_outputs(8635)));
    layer1_outputs(2202) <= layer0_outputs(9511);
    layer1_outputs(2203) <= (layer0_outputs(8473)) and (layer0_outputs(1809));
    layer1_outputs(2204) <= not(layer0_outputs(1482));
    layer1_outputs(2205) <= (layer0_outputs(3306)) xor (layer0_outputs(2894));
    layer1_outputs(2206) <= not(layer0_outputs(8526));
    layer1_outputs(2207) <= '1';
    layer1_outputs(2208) <= (layer0_outputs(10075)) and not (layer0_outputs(2665));
    layer1_outputs(2209) <= layer0_outputs(9622);
    layer1_outputs(2210) <= not(layer0_outputs(5799)) or (layer0_outputs(2736));
    layer1_outputs(2211) <= not((layer0_outputs(4584)) and (layer0_outputs(2927)));
    layer1_outputs(2212) <= not(layer0_outputs(3145));
    layer1_outputs(2213) <= (layer0_outputs(3216)) and (layer0_outputs(9451));
    layer1_outputs(2214) <= (layer0_outputs(3951)) and (layer0_outputs(6666));
    layer1_outputs(2215) <= not((layer0_outputs(3231)) and (layer0_outputs(5476)));
    layer1_outputs(2216) <= not(layer0_outputs(874));
    layer1_outputs(2217) <= not(layer0_outputs(4904)) or (layer0_outputs(4343));
    layer1_outputs(2218) <= (layer0_outputs(8956)) xor (layer0_outputs(6165));
    layer1_outputs(2219) <= not((layer0_outputs(5441)) xor (layer0_outputs(5828)));
    layer1_outputs(2220) <= (layer0_outputs(2161)) or (layer0_outputs(4775));
    layer1_outputs(2221) <= not(layer0_outputs(169)) or (layer0_outputs(4048));
    layer1_outputs(2222) <= (layer0_outputs(1626)) or (layer0_outputs(2846));
    layer1_outputs(2223) <= layer0_outputs(5129);
    layer1_outputs(2224) <= not((layer0_outputs(5189)) or (layer0_outputs(6310)));
    layer1_outputs(2225) <= layer0_outputs(4267);
    layer1_outputs(2226) <= layer0_outputs(4993);
    layer1_outputs(2227) <= not((layer0_outputs(2370)) xor (layer0_outputs(2450)));
    layer1_outputs(2228) <= layer0_outputs(6969);
    layer1_outputs(2229) <= not(layer0_outputs(1484)) or (layer0_outputs(4541));
    layer1_outputs(2230) <= layer0_outputs(9865);
    layer1_outputs(2231) <= layer0_outputs(1601);
    layer1_outputs(2232) <= not((layer0_outputs(857)) or (layer0_outputs(343)));
    layer1_outputs(2233) <= layer0_outputs(6543);
    layer1_outputs(2234) <= not(layer0_outputs(7795)) or (layer0_outputs(9250));
    layer1_outputs(2235) <= not(layer0_outputs(2551));
    layer1_outputs(2236) <= (layer0_outputs(5230)) and (layer0_outputs(3194));
    layer1_outputs(2237) <= not(layer0_outputs(4905));
    layer1_outputs(2238) <= layer0_outputs(3924);
    layer1_outputs(2239) <= (layer0_outputs(1637)) and (layer0_outputs(2689));
    layer1_outputs(2240) <= (layer0_outputs(9290)) and not (layer0_outputs(4453));
    layer1_outputs(2241) <= not((layer0_outputs(6084)) and (layer0_outputs(3453)));
    layer1_outputs(2242) <= not(layer0_outputs(4393));
    layer1_outputs(2243) <= layer0_outputs(8277);
    layer1_outputs(2244) <= layer0_outputs(3501);
    layer1_outputs(2245) <= not((layer0_outputs(8628)) or (layer0_outputs(161)));
    layer1_outputs(2246) <= not(layer0_outputs(36));
    layer1_outputs(2247) <= layer0_outputs(2435);
    layer1_outputs(2248) <= not((layer0_outputs(1692)) or (layer0_outputs(623)));
    layer1_outputs(2249) <= not((layer0_outputs(7062)) xor (layer0_outputs(6079)));
    layer1_outputs(2250) <= (layer0_outputs(195)) and not (layer0_outputs(1688));
    layer1_outputs(2251) <= '0';
    layer1_outputs(2252) <= layer0_outputs(2885);
    layer1_outputs(2253) <= not(layer0_outputs(3451));
    layer1_outputs(2254) <= not(layer0_outputs(2513));
    layer1_outputs(2255) <= layer0_outputs(2529);
    layer1_outputs(2256) <= layer0_outputs(3880);
    layer1_outputs(2257) <= not((layer0_outputs(2686)) or (layer0_outputs(498)));
    layer1_outputs(2258) <= not(layer0_outputs(6661)) or (layer0_outputs(1769));
    layer1_outputs(2259) <= not(layer0_outputs(482));
    layer1_outputs(2260) <= '0';
    layer1_outputs(2261) <= not((layer0_outputs(3132)) and (layer0_outputs(7774)));
    layer1_outputs(2262) <= not(layer0_outputs(5078));
    layer1_outputs(2263) <= not((layer0_outputs(4184)) xor (layer0_outputs(7773)));
    layer1_outputs(2264) <= (layer0_outputs(5849)) and not (layer0_outputs(7713));
    layer1_outputs(2265) <= not(layer0_outputs(3117));
    layer1_outputs(2266) <= not(layer0_outputs(1286)) or (layer0_outputs(4203));
    layer1_outputs(2267) <= not((layer0_outputs(3969)) or (layer0_outputs(1207)));
    layer1_outputs(2268) <= (layer0_outputs(7619)) or (layer0_outputs(1631));
    layer1_outputs(2269) <= not((layer0_outputs(10094)) and (layer0_outputs(1314)));
    layer1_outputs(2270) <= (layer0_outputs(4789)) or (layer0_outputs(4513));
    layer1_outputs(2271) <= (layer0_outputs(8028)) and not (layer0_outputs(9926));
    layer1_outputs(2272) <= layer0_outputs(4865);
    layer1_outputs(2273) <= layer0_outputs(6634);
    layer1_outputs(2274) <= (layer0_outputs(15)) or (layer0_outputs(8199));
    layer1_outputs(2275) <= (layer0_outputs(5355)) or (layer0_outputs(9847));
    layer1_outputs(2276) <= not(layer0_outputs(9618));
    layer1_outputs(2277) <= layer0_outputs(4536);
    layer1_outputs(2278) <= not((layer0_outputs(7410)) xor (layer0_outputs(9148)));
    layer1_outputs(2279) <= layer0_outputs(6052);
    layer1_outputs(2280) <= not((layer0_outputs(2682)) or (layer0_outputs(3448)));
    layer1_outputs(2281) <= not((layer0_outputs(3097)) or (layer0_outputs(2215)));
    layer1_outputs(2282) <= (layer0_outputs(7634)) xor (layer0_outputs(5126));
    layer1_outputs(2283) <= layer0_outputs(5763);
    layer1_outputs(2284) <= not(layer0_outputs(554));
    layer1_outputs(2285) <= layer0_outputs(3743);
    layer1_outputs(2286) <= layer0_outputs(7315);
    layer1_outputs(2287) <= layer0_outputs(8020);
    layer1_outputs(2288) <= (layer0_outputs(2585)) and not (layer0_outputs(2802));
    layer1_outputs(2289) <= not(layer0_outputs(6266)) or (layer0_outputs(603));
    layer1_outputs(2290) <= (layer0_outputs(9636)) or (layer0_outputs(7915));
    layer1_outputs(2291) <= not((layer0_outputs(424)) or (layer0_outputs(8594)));
    layer1_outputs(2292) <= not(layer0_outputs(2671));
    layer1_outputs(2293) <= layer0_outputs(3087);
    layer1_outputs(2294) <= not(layer0_outputs(4906)) or (layer0_outputs(1150));
    layer1_outputs(2295) <= not((layer0_outputs(5849)) and (layer0_outputs(10088)));
    layer1_outputs(2296) <= not(layer0_outputs(4598)) or (layer0_outputs(8983));
    layer1_outputs(2297) <= not((layer0_outputs(2152)) or (layer0_outputs(4571)));
    layer1_outputs(2298) <= '0';
    layer1_outputs(2299) <= layer0_outputs(3495);
    layer1_outputs(2300) <= not(layer0_outputs(4749));
    layer1_outputs(2301) <= layer0_outputs(5913);
    layer1_outputs(2302) <= not(layer0_outputs(6359));
    layer1_outputs(2303) <= layer0_outputs(468);
    layer1_outputs(2304) <= (layer0_outputs(8111)) and not (layer0_outputs(3509));
    layer1_outputs(2305) <= not(layer0_outputs(8549)) or (layer0_outputs(9045));
    layer1_outputs(2306) <= not((layer0_outputs(1490)) and (layer0_outputs(4309)));
    layer1_outputs(2307) <= not((layer0_outputs(3114)) and (layer0_outputs(4689)));
    layer1_outputs(2308) <= not((layer0_outputs(5501)) or (layer0_outputs(5399)));
    layer1_outputs(2309) <= layer0_outputs(7720);
    layer1_outputs(2310) <= layer0_outputs(7352);
    layer1_outputs(2311) <= layer0_outputs(34);
    layer1_outputs(2312) <= not(layer0_outputs(4879));
    layer1_outputs(2313) <= not(layer0_outputs(273));
    layer1_outputs(2314) <= not((layer0_outputs(3154)) xor (layer0_outputs(6717)));
    layer1_outputs(2315) <= not((layer0_outputs(884)) or (layer0_outputs(867)));
    layer1_outputs(2316) <= not(layer0_outputs(1161));
    layer1_outputs(2317) <= not(layer0_outputs(4355));
    layer1_outputs(2318) <= not((layer0_outputs(7009)) or (layer0_outputs(4585)));
    layer1_outputs(2319) <= layer0_outputs(4358);
    layer1_outputs(2320) <= not(layer0_outputs(8673)) or (layer0_outputs(6408));
    layer1_outputs(2321) <= (layer0_outputs(2759)) and not (layer0_outputs(2680));
    layer1_outputs(2322) <= layer0_outputs(859);
    layer1_outputs(2323) <= not(layer0_outputs(8949)) or (layer0_outputs(4706));
    layer1_outputs(2324) <= (layer0_outputs(7176)) and (layer0_outputs(7732));
    layer1_outputs(2325) <= (layer0_outputs(2554)) or (layer0_outputs(9398));
    layer1_outputs(2326) <= layer0_outputs(1332);
    layer1_outputs(2327) <= not((layer0_outputs(4939)) and (layer0_outputs(2074)));
    layer1_outputs(2328) <= layer0_outputs(905);
    layer1_outputs(2329) <= layer0_outputs(3021);
    layer1_outputs(2330) <= not(layer0_outputs(484)) or (layer0_outputs(1758));
    layer1_outputs(2331) <= not(layer0_outputs(566)) or (layer0_outputs(4362));
    layer1_outputs(2332) <= not((layer0_outputs(6830)) or (layer0_outputs(8557)));
    layer1_outputs(2333) <= layer0_outputs(6541);
    layer1_outputs(2334) <= not((layer0_outputs(2662)) and (layer0_outputs(7888)));
    layer1_outputs(2335) <= not((layer0_outputs(1476)) and (layer0_outputs(1167)));
    layer1_outputs(2336) <= '1';
    layer1_outputs(2337) <= layer0_outputs(3114);
    layer1_outputs(2338) <= layer0_outputs(4530);
    layer1_outputs(2339) <= not(layer0_outputs(3741)) or (layer0_outputs(7860));
    layer1_outputs(2340) <= not((layer0_outputs(56)) and (layer0_outputs(2997)));
    layer1_outputs(2341) <= layer0_outputs(10179);
    layer1_outputs(2342) <= '0';
    layer1_outputs(2343) <= '0';
    layer1_outputs(2344) <= (layer0_outputs(5043)) and not (layer0_outputs(8344));
    layer1_outputs(2345) <= (layer0_outputs(981)) or (layer0_outputs(5110));
    layer1_outputs(2346) <= not((layer0_outputs(1459)) and (layer0_outputs(2881)));
    layer1_outputs(2347) <= not((layer0_outputs(9316)) xor (layer0_outputs(9029)));
    layer1_outputs(2348) <= (layer0_outputs(589)) and not (layer0_outputs(1307));
    layer1_outputs(2349) <= (layer0_outputs(1340)) and not (layer0_outputs(1524));
    layer1_outputs(2350) <= not(layer0_outputs(6642));
    layer1_outputs(2351) <= not(layer0_outputs(7177));
    layer1_outputs(2352) <= (layer0_outputs(9775)) and not (layer0_outputs(3496));
    layer1_outputs(2353) <= (layer0_outputs(7211)) or (layer0_outputs(4368));
    layer1_outputs(2354) <= (layer0_outputs(5026)) xor (layer0_outputs(9487));
    layer1_outputs(2355) <= not(layer0_outputs(4526)) or (layer0_outputs(5615));
    layer1_outputs(2356) <= not((layer0_outputs(8845)) xor (layer0_outputs(976)));
    layer1_outputs(2357) <= not(layer0_outputs(6543));
    layer1_outputs(2358) <= layer0_outputs(1686);
    layer1_outputs(2359) <= not(layer0_outputs(1083)) or (layer0_outputs(7692));
    layer1_outputs(2360) <= layer0_outputs(7763);
    layer1_outputs(2361) <= not(layer0_outputs(2784));
    layer1_outputs(2362) <= not(layer0_outputs(8300)) or (layer0_outputs(1799));
    layer1_outputs(2363) <= (layer0_outputs(1441)) xor (layer0_outputs(1371));
    layer1_outputs(2364) <= layer0_outputs(6882);
    layer1_outputs(2365) <= (layer0_outputs(4733)) and not (layer0_outputs(436));
    layer1_outputs(2366) <= '0';
    layer1_outputs(2367) <= (layer0_outputs(3926)) xor (layer0_outputs(7195));
    layer1_outputs(2368) <= layer0_outputs(3919);
    layer1_outputs(2369) <= layer0_outputs(6751);
    layer1_outputs(2370) <= (layer0_outputs(2149)) and not (layer0_outputs(1554));
    layer1_outputs(2371) <= layer0_outputs(5342);
    layer1_outputs(2372) <= layer0_outputs(9774);
    layer1_outputs(2373) <= (layer0_outputs(9344)) xor (layer0_outputs(3909));
    layer1_outputs(2374) <= not(layer0_outputs(7556));
    layer1_outputs(2375) <= not(layer0_outputs(8731));
    layer1_outputs(2376) <= (layer0_outputs(3867)) and (layer0_outputs(4941));
    layer1_outputs(2377) <= not(layer0_outputs(10041));
    layer1_outputs(2378) <= not((layer0_outputs(2066)) and (layer0_outputs(10222)));
    layer1_outputs(2379) <= (layer0_outputs(9899)) and (layer0_outputs(4024));
    layer1_outputs(2380) <= not((layer0_outputs(761)) xor (layer0_outputs(2560)));
    layer1_outputs(2381) <= layer0_outputs(5809);
    layer1_outputs(2382) <= not((layer0_outputs(201)) or (layer0_outputs(3641)));
    layer1_outputs(2383) <= not((layer0_outputs(7151)) xor (layer0_outputs(2337)));
    layer1_outputs(2384) <= (layer0_outputs(8737)) or (layer0_outputs(4348));
    layer1_outputs(2385) <= layer0_outputs(9360);
    layer1_outputs(2386) <= layer0_outputs(2788);
    layer1_outputs(2387) <= not(layer0_outputs(5566));
    layer1_outputs(2388) <= not((layer0_outputs(7082)) xor (layer0_outputs(6261)));
    layer1_outputs(2389) <= not((layer0_outputs(3568)) xor (layer0_outputs(6201)));
    layer1_outputs(2390) <= not((layer0_outputs(8830)) and (layer0_outputs(9832)));
    layer1_outputs(2391) <= layer0_outputs(10047);
    layer1_outputs(2392) <= layer0_outputs(5955);
    layer1_outputs(2393) <= layer0_outputs(4714);
    layer1_outputs(2394) <= layer0_outputs(4279);
    layer1_outputs(2395) <= not(layer0_outputs(3958));
    layer1_outputs(2396) <= not(layer0_outputs(5821)) or (layer0_outputs(9617));
    layer1_outputs(2397) <= (layer0_outputs(7380)) xor (layer0_outputs(5409));
    layer1_outputs(2398) <= not(layer0_outputs(5130));
    layer1_outputs(2399) <= not(layer0_outputs(8379)) or (layer0_outputs(9581));
    layer1_outputs(2400) <= (layer0_outputs(1899)) and not (layer0_outputs(3268));
    layer1_outputs(2401) <= (layer0_outputs(5156)) and (layer0_outputs(20));
    layer1_outputs(2402) <= not(layer0_outputs(8686)) or (layer0_outputs(6824));
    layer1_outputs(2403) <= layer0_outputs(5394);
    layer1_outputs(2404) <= (layer0_outputs(8784)) or (layer0_outputs(135));
    layer1_outputs(2405) <= (layer0_outputs(9073)) and not (layer0_outputs(4393));
    layer1_outputs(2406) <= not((layer0_outputs(6974)) or (layer0_outputs(2958)));
    layer1_outputs(2407) <= not(layer0_outputs(10004));
    layer1_outputs(2408) <= not(layer0_outputs(9477)) or (layer0_outputs(4042));
    layer1_outputs(2409) <= (layer0_outputs(2539)) xor (layer0_outputs(1993));
    layer1_outputs(2410) <= layer0_outputs(6476);
    layer1_outputs(2411) <= layer0_outputs(7219);
    layer1_outputs(2412) <= not(layer0_outputs(3764)) or (layer0_outputs(4496));
    layer1_outputs(2413) <= (layer0_outputs(2264)) and not (layer0_outputs(7539));
    layer1_outputs(2414) <= (layer0_outputs(9448)) and (layer0_outputs(3402));
    layer1_outputs(2415) <= not(layer0_outputs(9881));
    layer1_outputs(2416) <= not(layer0_outputs(2480)) or (layer0_outputs(2880));
    layer1_outputs(2417) <= not((layer0_outputs(8770)) or (layer0_outputs(5611)));
    layer1_outputs(2418) <= layer0_outputs(6845);
    layer1_outputs(2419) <= layer0_outputs(1338);
    layer1_outputs(2420) <= (layer0_outputs(7096)) and (layer0_outputs(5823));
    layer1_outputs(2421) <= not(layer0_outputs(10013));
    layer1_outputs(2422) <= not((layer0_outputs(4925)) xor (layer0_outputs(1466)));
    layer1_outputs(2423) <= not((layer0_outputs(6351)) or (layer0_outputs(871)));
    layer1_outputs(2424) <= layer0_outputs(3082);
    layer1_outputs(2425) <= layer0_outputs(5568);
    layer1_outputs(2426) <= (layer0_outputs(7790)) and (layer0_outputs(6126));
    layer1_outputs(2427) <= layer0_outputs(247);
    layer1_outputs(2428) <= not(layer0_outputs(607));
    layer1_outputs(2429) <= not(layer0_outputs(8798));
    layer1_outputs(2430) <= (layer0_outputs(9421)) and not (layer0_outputs(7532));
    layer1_outputs(2431) <= '0';
    layer1_outputs(2432) <= not(layer0_outputs(3698));
    layer1_outputs(2433) <= not((layer0_outputs(6072)) xor (layer0_outputs(1228)));
    layer1_outputs(2434) <= not(layer0_outputs(1708));
    layer1_outputs(2435) <= (layer0_outputs(3844)) or (layer0_outputs(8868));
    layer1_outputs(2436) <= not(layer0_outputs(1510));
    layer1_outputs(2437) <= not(layer0_outputs(7544)) or (layer0_outputs(7037));
    layer1_outputs(2438) <= (layer0_outputs(7046)) and (layer0_outputs(8301));
    layer1_outputs(2439) <= not(layer0_outputs(5240));
    layer1_outputs(2440) <= not(layer0_outputs(9855));
    layer1_outputs(2441) <= (layer0_outputs(6967)) and not (layer0_outputs(2502));
    layer1_outputs(2442) <= (layer0_outputs(6374)) and not (layer0_outputs(7773));
    layer1_outputs(2443) <= (layer0_outputs(6390)) xor (layer0_outputs(368));
    layer1_outputs(2444) <= not(layer0_outputs(5905));
    layer1_outputs(2445) <= not(layer0_outputs(8897)) or (layer0_outputs(7580));
    layer1_outputs(2446) <= not(layer0_outputs(258)) or (layer0_outputs(910));
    layer1_outputs(2447) <= layer0_outputs(1385);
    layer1_outputs(2448) <= not(layer0_outputs(8165));
    layer1_outputs(2449) <= (layer0_outputs(3034)) xor (layer0_outputs(151));
    layer1_outputs(2450) <= not(layer0_outputs(7372));
    layer1_outputs(2451) <= layer0_outputs(3989);
    layer1_outputs(2452) <= not(layer0_outputs(3017));
    layer1_outputs(2453) <= not(layer0_outputs(5829)) or (layer0_outputs(2802));
    layer1_outputs(2454) <= layer0_outputs(9049);
    layer1_outputs(2455) <= not((layer0_outputs(5338)) and (layer0_outputs(5232)));
    layer1_outputs(2456) <= (layer0_outputs(8599)) or (layer0_outputs(3846));
    layer1_outputs(2457) <= (layer0_outputs(8595)) and (layer0_outputs(2794));
    layer1_outputs(2458) <= not(layer0_outputs(8916));
    layer1_outputs(2459) <= layer0_outputs(5301);
    layer1_outputs(2460) <= not((layer0_outputs(6050)) and (layer0_outputs(8797)));
    layer1_outputs(2461) <= not((layer0_outputs(636)) and (layer0_outputs(5802)));
    layer1_outputs(2462) <= layer0_outputs(8877);
    layer1_outputs(2463) <= layer0_outputs(8796);
    layer1_outputs(2464) <= not((layer0_outputs(1313)) and (layer0_outputs(4172)));
    layer1_outputs(2465) <= layer0_outputs(988);
    layer1_outputs(2466) <= layer0_outputs(4952);
    layer1_outputs(2467) <= not((layer0_outputs(3217)) or (layer0_outputs(2772)));
    layer1_outputs(2468) <= (layer0_outputs(9251)) and (layer0_outputs(3623));
    layer1_outputs(2469) <= not((layer0_outputs(7545)) and (layer0_outputs(5268)));
    layer1_outputs(2470) <= not(layer0_outputs(157));
    layer1_outputs(2471) <= (layer0_outputs(2234)) and (layer0_outputs(5998));
    layer1_outputs(2472) <= (layer0_outputs(9261)) and not (layer0_outputs(4866));
    layer1_outputs(2473) <= (layer0_outputs(3260)) and (layer0_outputs(6453));
    layer1_outputs(2474) <= layer0_outputs(3068);
    layer1_outputs(2475) <= layer0_outputs(8791);
    layer1_outputs(2476) <= not(layer0_outputs(7188)) or (layer0_outputs(5755));
    layer1_outputs(2477) <= not(layer0_outputs(6912));
    layer1_outputs(2478) <= (layer0_outputs(3915)) and not (layer0_outputs(839));
    layer1_outputs(2479) <= (layer0_outputs(6970)) and not (layer0_outputs(3662));
    layer1_outputs(2480) <= (layer0_outputs(7848)) and (layer0_outputs(5590));
    layer1_outputs(2481) <= layer0_outputs(6607);
    layer1_outputs(2482) <= (layer0_outputs(4318)) and not (layer0_outputs(2599));
    layer1_outputs(2483) <= not((layer0_outputs(339)) xor (layer0_outputs(8610)));
    layer1_outputs(2484) <= (layer0_outputs(3187)) and not (layer0_outputs(8015));
    layer1_outputs(2485) <= not((layer0_outputs(6831)) or (layer0_outputs(6627)));
    layer1_outputs(2486) <= not(layer0_outputs(29)) or (layer0_outputs(5483));
    layer1_outputs(2487) <= layer0_outputs(6874);
    layer1_outputs(2488) <= not(layer0_outputs(6836)) or (layer0_outputs(8187));
    layer1_outputs(2489) <= not(layer0_outputs(5025));
    layer1_outputs(2490) <= not((layer0_outputs(8988)) and (layer0_outputs(4491)));
    layer1_outputs(2491) <= not((layer0_outputs(4660)) or (layer0_outputs(175)));
    layer1_outputs(2492) <= not(layer0_outputs(2866)) or (layer0_outputs(4493));
    layer1_outputs(2493) <= (layer0_outputs(974)) or (layer0_outputs(4779));
    layer1_outputs(2494) <= not(layer0_outputs(2177));
    layer1_outputs(2495) <= layer0_outputs(7142);
    layer1_outputs(2496) <= layer0_outputs(2066);
    layer1_outputs(2497) <= not((layer0_outputs(1020)) xor (layer0_outputs(8023)));
    layer1_outputs(2498) <= layer0_outputs(1230);
    layer1_outputs(2499) <= not(layer0_outputs(7845));
    layer1_outputs(2500) <= not((layer0_outputs(8124)) and (layer0_outputs(9017)));
    layer1_outputs(2501) <= layer0_outputs(2369);
    layer1_outputs(2502) <= (layer0_outputs(1841)) and not (layer0_outputs(6633));
    layer1_outputs(2503) <= not((layer0_outputs(5556)) or (layer0_outputs(3576)));
    layer1_outputs(2504) <= layer0_outputs(879);
    layer1_outputs(2505) <= not(layer0_outputs(9909));
    layer1_outputs(2506) <= not(layer0_outputs(1782)) or (layer0_outputs(9105));
    layer1_outputs(2507) <= layer0_outputs(1109);
    layer1_outputs(2508) <= not((layer0_outputs(8085)) xor (layer0_outputs(3528)));
    layer1_outputs(2509) <= not(layer0_outputs(3226));
    layer1_outputs(2510) <= not((layer0_outputs(1324)) or (layer0_outputs(2326)));
    layer1_outputs(2511) <= not((layer0_outputs(1117)) or (layer0_outputs(9538)));
    layer1_outputs(2512) <= not(layer0_outputs(7344));
    layer1_outputs(2513) <= not(layer0_outputs(8760));
    layer1_outputs(2514) <= layer0_outputs(9812);
    layer1_outputs(2515) <= layer0_outputs(6183);
    layer1_outputs(2516) <= not(layer0_outputs(3074));
    layer1_outputs(2517) <= not((layer0_outputs(3337)) and (layer0_outputs(9148)));
    layer1_outputs(2518) <= not(layer0_outputs(8711));
    layer1_outputs(2519) <= '0';
    layer1_outputs(2520) <= layer0_outputs(6712);
    layer1_outputs(2521) <= not((layer0_outputs(4642)) xor (layer0_outputs(4361)));
    layer1_outputs(2522) <= layer0_outputs(9035);
    layer1_outputs(2523) <= layer0_outputs(7373);
    layer1_outputs(2524) <= layer0_outputs(3201);
    layer1_outputs(2525) <= '0';
    layer1_outputs(2526) <= (layer0_outputs(6055)) or (layer0_outputs(3532));
    layer1_outputs(2527) <= (layer0_outputs(2994)) and not (layer0_outputs(8580));
    layer1_outputs(2528) <= not(layer0_outputs(836));
    layer1_outputs(2529) <= not(layer0_outputs(413));
    layer1_outputs(2530) <= not(layer0_outputs(7231));
    layer1_outputs(2531) <= not((layer0_outputs(3912)) and (layer0_outputs(7553)));
    layer1_outputs(2532) <= not((layer0_outputs(6987)) and (layer0_outputs(5863)));
    layer1_outputs(2533) <= not((layer0_outputs(9052)) or (layer0_outputs(3003)));
    layer1_outputs(2534) <= layer0_outputs(995);
    layer1_outputs(2535) <= (layer0_outputs(6358)) or (layer0_outputs(5617));
    layer1_outputs(2536) <= (layer0_outputs(9820)) and not (layer0_outputs(5102));
    layer1_outputs(2537) <= layer0_outputs(1889);
    layer1_outputs(2538) <= not(layer0_outputs(4916));
    layer1_outputs(2539) <= layer0_outputs(4289);
    layer1_outputs(2540) <= (layer0_outputs(4435)) and (layer0_outputs(1584));
    layer1_outputs(2541) <= (layer0_outputs(1289)) and (layer0_outputs(5229));
    layer1_outputs(2542) <= (layer0_outputs(9514)) and (layer0_outputs(9395));
    layer1_outputs(2543) <= not(layer0_outputs(7933));
    layer1_outputs(2544) <= '1';
    layer1_outputs(2545) <= layer0_outputs(6004);
    layer1_outputs(2546) <= not((layer0_outputs(9501)) or (layer0_outputs(6912)));
    layer1_outputs(2547) <= not(layer0_outputs(6366));
    layer1_outputs(2548) <= (layer0_outputs(5553)) and (layer0_outputs(6035));
    layer1_outputs(2549) <= (layer0_outputs(1771)) and not (layer0_outputs(10057));
    layer1_outputs(2550) <= not(layer0_outputs(3780)) or (layer0_outputs(8445));
    layer1_outputs(2551) <= layer0_outputs(7056);
    layer1_outputs(2552) <= (layer0_outputs(1381)) and not (layer0_outputs(3161));
    layer1_outputs(2553) <= not(layer0_outputs(1467));
    layer1_outputs(2554) <= (layer0_outputs(6455)) and (layer0_outputs(9185));
    layer1_outputs(2555) <= layer0_outputs(8851);
    layer1_outputs(2556) <= not(layer0_outputs(1127));
    layer1_outputs(2557) <= (layer0_outputs(3621)) and not (layer0_outputs(9332));
    layer1_outputs(2558) <= (layer0_outputs(2581)) and not (layer0_outputs(9405));
    layer1_outputs(2559) <= (layer0_outputs(3129)) xor (layer0_outputs(10095));
    layer1_outputs(2560) <= (layer0_outputs(9898)) and not (layer0_outputs(574));
    layer1_outputs(2561) <= layer0_outputs(10042);
    layer1_outputs(2562) <= not((layer0_outputs(5080)) or (layer0_outputs(4805)));
    layer1_outputs(2563) <= not((layer0_outputs(6899)) and (layer0_outputs(4892)));
    layer1_outputs(2564) <= not(layer0_outputs(5496));
    layer1_outputs(2565) <= layer0_outputs(787);
    layer1_outputs(2566) <= layer0_outputs(4043);
    layer1_outputs(2567) <= not((layer0_outputs(7394)) and (layer0_outputs(6174)));
    layer1_outputs(2568) <= not(layer0_outputs(1360));
    layer1_outputs(2569) <= not(layer0_outputs(3730));
    layer1_outputs(2570) <= not(layer0_outputs(7881));
    layer1_outputs(2571) <= (layer0_outputs(1896)) and not (layer0_outputs(2342));
    layer1_outputs(2572) <= (layer0_outputs(5380)) xor (layer0_outputs(7800));
    layer1_outputs(2573) <= not(layer0_outputs(2357));
    layer1_outputs(2574) <= '0';
    layer1_outputs(2575) <= layer0_outputs(1494);
    layer1_outputs(2576) <= not((layer0_outputs(6964)) and (layer0_outputs(2738)));
    layer1_outputs(2577) <= layer0_outputs(4068);
    layer1_outputs(2578) <= not(layer0_outputs(1891));
    layer1_outputs(2579) <= not(layer0_outputs(2309));
    layer1_outputs(2580) <= not((layer0_outputs(8329)) xor (layer0_outputs(6285)));
    layer1_outputs(2581) <= (layer0_outputs(4561)) xor (layer0_outputs(5964));
    layer1_outputs(2582) <= '1';
    layer1_outputs(2583) <= (layer0_outputs(249)) and (layer0_outputs(3866));
    layer1_outputs(2584) <= (layer0_outputs(7467)) or (layer0_outputs(5603));
    layer1_outputs(2585) <= (layer0_outputs(6074)) and not (layer0_outputs(9729));
    layer1_outputs(2586) <= not(layer0_outputs(4926));
    layer1_outputs(2587) <= layer0_outputs(6760);
    layer1_outputs(2588) <= layer0_outputs(1170);
    layer1_outputs(2589) <= not(layer0_outputs(4455));
    layer1_outputs(2590) <= not(layer0_outputs(1259)) or (layer0_outputs(1480));
    layer1_outputs(2591) <= not((layer0_outputs(7315)) or (layer0_outputs(8663)));
    layer1_outputs(2592) <= not(layer0_outputs(2448));
    layer1_outputs(2593) <= not((layer0_outputs(9495)) xor (layer0_outputs(3982)));
    layer1_outputs(2594) <= not(layer0_outputs(7864));
    layer1_outputs(2595) <= (layer0_outputs(2818)) and not (layer0_outputs(9454));
    layer1_outputs(2596) <= not((layer0_outputs(8639)) and (layer0_outputs(4929)));
    layer1_outputs(2597) <= layer0_outputs(8299);
    layer1_outputs(2598) <= '1';
    layer1_outputs(2599) <= (layer0_outputs(9886)) and not (layer0_outputs(3880));
    layer1_outputs(2600) <= not((layer0_outputs(3709)) or (layer0_outputs(1512)));
    layer1_outputs(2601) <= layer0_outputs(6100);
    layer1_outputs(2602) <= (layer0_outputs(2775)) and (layer0_outputs(5037));
    layer1_outputs(2603) <= (layer0_outputs(7288)) and not (layer0_outputs(1764));
    layer1_outputs(2604) <= layer0_outputs(6572);
    layer1_outputs(2605) <= not(layer0_outputs(7771)) or (layer0_outputs(6022));
    layer1_outputs(2606) <= (layer0_outputs(6384)) and (layer0_outputs(4810));
    layer1_outputs(2607) <= layer0_outputs(5851);
    layer1_outputs(2608) <= not((layer0_outputs(2908)) and (layer0_outputs(2673)));
    layer1_outputs(2609) <= not(layer0_outputs(4423));
    layer1_outputs(2610) <= not(layer0_outputs(7208)) or (layer0_outputs(5904));
    layer1_outputs(2611) <= (layer0_outputs(506)) or (layer0_outputs(2007));
    layer1_outputs(2612) <= (layer0_outputs(7733)) and (layer0_outputs(7793));
    layer1_outputs(2613) <= (layer0_outputs(3449)) and not (layer0_outputs(1224));
    layer1_outputs(2614) <= not(layer0_outputs(1681));
    layer1_outputs(2615) <= not((layer0_outputs(3457)) and (layer0_outputs(4336)));
    layer1_outputs(2616) <= layer0_outputs(4131);
    layer1_outputs(2617) <= not(layer0_outputs(3057));
    layer1_outputs(2618) <= (layer0_outputs(1212)) xor (layer0_outputs(2251));
    layer1_outputs(2619) <= not(layer0_outputs(3971)) or (layer0_outputs(1906));
    layer1_outputs(2620) <= (layer0_outputs(2959)) or (layer0_outputs(4085));
    layer1_outputs(2621) <= not(layer0_outputs(8842));
    layer1_outputs(2622) <= not(layer0_outputs(1458)) or (layer0_outputs(1380));
    layer1_outputs(2623) <= (layer0_outputs(320)) xor (layer0_outputs(9911));
    layer1_outputs(2624) <= not(layer0_outputs(497)) or (layer0_outputs(1785));
    layer1_outputs(2625) <= not((layer0_outputs(7536)) and (layer0_outputs(2156)));
    layer1_outputs(2626) <= not(layer0_outputs(3248));
    layer1_outputs(2627) <= not(layer0_outputs(4001)) or (layer0_outputs(9409));
    layer1_outputs(2628) <= (layer0_outputs(10009)) and not (layer0_outputs(8769));
    layer1_outputs(2629) <= (layer0_outputs(6067)) xor (layer0_outputs(1166));
    layer1_outputs(2630) <= (layer0_outputs(2737)) or (layer0_outputs(3364));
    layer1_outputs(2631) <= not((layer0_outputs(6427)) or (layer0_outputs(8888)));
    layer1_outputs(2632) <= (layer0_outputs(9283)) and not (layer0_outputs(9183));
    layer1_outputs(2633) <= not(layer0_outputs(3240)) or (layer0_outputs(4113));
    layer1_outputs(2634) <= not(layer0_outputs(2902));
    layer1_outputs(2635) <= layer0_outputs(9369);
    layer1_outputs(2636) <= (layer0_outputs(646)) and not (layer0_outputs(9381));
    layer1_outputs(2637) <= layer0_outputs(2945);
    layer1_outputs(2638) <= not(layer0_outputs(7601));
    layer1_outputs(2639) <= not((layer0_outputs(1406)) or (layer0_outputs(992)));
    layer1_outputs(2640) <= layer0_outputs(6064);
    layer1_outputs(2641) <= not(layer0_outputs(4422));
    layer1_outputs(2642) <= not(layer0_outputs(1013));
    layer1_outputs(2643) <= (layer0_outputs(6993)) and not (layer0_outputs(584));
    layer1_outputs(2644) <= (layer0_outputs(7198)) and (layer0_outputs(6260));
    layer1_outputs(2645) <= not(layer0_outputs(5375)) or (layer0_outputs(4383));
    layer1_outputs(2646) <= (layer0_outputs(6085)) and not (layer0_outputs(3303));
    layer1_outputs(2647) <= layer0_outputs(2486);
    layer1_outputs(2648) <= layer0_outputs(5930);
    layer1_outputs(2649) <= '0';
    layer1_outputs(2650) <= (layer0_outputs(494)) and (layer0_outputs(9104));
    layer1_outputs(2651) <= '1';
    layer1_outputs(2652) <= '0';
    layer1_outputs(2653) <= (layer0_outputs(1325)) and not (layer0_outputs(4974));
    layer1_outputs(2654) <= not((layer0_outputs(809)) or (layer0_outputs(686)));
    layer1_outputs(2655) <= (layer0_outputs(9772)) and not (layer0_outputs(5853));
    layer1_outputs(2656) <= not((layer0_outputs(9087)) or (layer0_outputs(6674)));
    layer1_outputs(2657) <= layer0_outputs(2639);
    layer1_outputs(2658) <= layer0_outputs(7362);
    layer1_outputs(2659) <= not(layer0_outputs(2631));
    layer1_outputs(2660) <= not((layer0_outputs(7543)) and (layer0_outputs(9350)));
    layer1_outputs(2661) <= (layer0_outputs(9887)) and (layer0_outputs(105));
    layer1_outputs(2662) <= (layer0_outputs(8848)) and not (layer0_outputs(8012));
    layer1_outputs(2663) <= (layer0_outputs(5630)) and not (layer0_outputs(3696));
    layer1_outputs(2664) <= not(layer0_outputs(8839));
    layer1_outputs(2665) <= not(layer0_outputs(4161));
    layer1_outputs(2666) <= '1';
    layer1_outputs(2667) <= not(layer0_outputs(3427)) or (layer0_outputs(1800));
    layer1_outputs(2668) <= (layer0_outputs(1422)) xor (layer0_outputs(7803));
    layer1_outputs(2669) <= not(layer0_outputs(6906));
    layer1_outputs(2670) <= layer0_outputs(7718);
    layer1_outputs(2671) <= (layer0_outputs(8349)) and (layer0_outputs(7159));
    layer1_outputs(2672) <= (layer0_outputs(4004)) and not (layer0_outputs(861));
    layer1_outputs(2673) <= not((layer0_outputs(2665)) and (layer0_outputs(6147)));
    layer1_outputs(2674) <= (layer0_outputs(2963)) and not (layer0_outputs(6929));
    layer1_outputs(2675) <= not(layer0_outputs(980));
    layer1_outputs(2676) <= not(layer0_outputs(5437));
    layer1_outputs(2677) <= layer0_outputs(5744);
    layer1_outputs(2678) <= not(layer0_outputs(1073));
    layer1_outputs(2679) <= (layer0_outputs(9288)) or (layer0_outputs(7821));
    layer1_outputs(2680) <= (layer0_outputs(2483)) or (layer0_outputs(1242));
    layer1_outputs(2681) <= layer0_outputs(616);
    layer1_outputs(2682) <= not(layer0_outputs(8736)) or (layer0_outputs(6047));
    layer1_outputs(2683) <= layer0_outputs(1232);
    layer1_outputs(2684) <= not(layer0_outputs(52));
    layer1_outputs(2685) <= not(layer0_outputs(9120));
    layer1_outputs(2686) <= not(layer0_outputs(6695));
    layer1_outputs(2687) <= not(layer0_outputs(5369));
    layer1_outputs(2688) <= (layer0_outputs(3490)) and not (layer0_outputs(7052));
    layer1_outputs(2689) <= not(layer0_outputs(9656));
    layer1_outputs(2690) <= not(layer0_outputs(7673)) or (layer0_outputs(1628));
    layer1_outputs(2691) <= not((layer0_outputs(359)) and (layer0_outputs(9034)));
    layer1_outputs(2692) <= layer0_outputs(6923);
    layer1_outputs(2693) <= (layer0_outputs(1794)) and not (layer0_outputs(9880));
    layer1_outputs(2694) <= not((layer0_outputs(8128)) or (layer0_outputs(8986)));
    layer1_outputs(2695) <= not(layer0_outputs(7464));
    layer1_outputs(2696) <= layer0_outputs(8792);
    layer1_outputs(2697) <= layer0_outputs(8613);
    layer1_outputs(2698) <= '0';
    layer1_outputs(2699) <= '0';
    layer1_outputs(2700) <= not((layer0_outputs(3833)) and (layer0_outputs(5111)));
    layer1_outputs(2701) <= (layer0_outputs(1153)) xor (layer0_outputs(6711));
    layer1_outputs(2702) <= (layer0_outputs(5962)) and (layer0_outputs(8762));
    layer1_outputs(2703) <= not(layer0_outputs(223));
    layer1_outputs(2704) <= not(layer0_outputs(7374));
    layer1_outputs(2705) <= not(layer0_outputs(8060));
    layer1_outputs(2706) <= (layer0_outputs(4263)) or (layer0_outputs(9458));
    layer1_outputs(2707) <= (layer0_outputs(5467)) and (layer0_outputs(1984));
    layer1_outputs(2708) <= (layer0_outputs(9512)) and not (layer0_outputs(9949));
    layer1_outputs(2709) <= (layer0_outputs(6234)) and not (layer0_outputs(6806));
    layer1_outputs(2710) <= (layer0_outputs(5920)) and not (layer0_outputs(7835));
    layer1_outputs(2711) <= layer0_outputs(5300);
    layer1_outputs(2712) <= (layer0_outputs(4256)) or (layer0_outputs(858));
    layer1_outputs(2713) <= layer0_outputs(9738);
    layer1_outputs(2714) <= not((layer0_outputs(5706)) and (layer0_outputs(8076)));
    layer1_outputs(2715) <= layer0_outputs(4283);
    layer1_outputs(2716) <= not(layer0_outputs(4673));
    layer1_outputs(2717) <= (layer0_outputs(2827)) xor (layer0_outputs(2980));
    layer1_outputs(2718) <= not(layer0_outputs(9264));
    layer1_outputs(2719) <= (layer0_outputs(197)) and not (layer0_outputs(2863));
    layer1_outputs(2720) <= '1';
    layer1_outputs(2721) <= not(layer0_outputs(4414));
    layer1_outputs(2722) <= layer0_outputs(5141);
    layer1_outputs(2723) <= layer0_outputs(441);
    layer1_outputs(2724) <= not((layer0_outputs(6197)) and (layer0_outputs(6828)));
    layer1_outputs(2725) <= (layer0_outputs(9258)) and not (layer0_outputs(6189));
    layer1_outputs(2726) <= not(layer0_outputs(4673));
    layer1_outputs(2727) <= layer0_outputs(4719);
    layer1_outputs(2728) <= (layer0_outputs(7872)) and not (layer0_outputs(2241));
    layer1_outputs(2729) <= (layer0_outputs(9851)) and not (layer0_outputs(5634));
    layer1_outputs(2730) <= not(layer0_outputs(7414));
    layer1_outputs(2731) <= not((layer0_outputs(1164)) and (layer0_outputs(3969)));
    layer1_outputs(2732) <= not((layer0_outputs(459)) and (layer0_outputs(5160)));
    layer1_outputs(2733) <= not(layer0_outputs(6075));
    layer1_outputs(2734) <= not(layer0_outputs(3085)) or (layer0_outputs(1225));
    layer1_outputs(2735) <= (layer0_outputs(2883)) and (layer0_outputs(703));
    layer1_outputs(2736) <= not((layer0_outputs(4760)) and (layer0_outputs(8052)));
    layer1_outputs(2737) <= not(layer0_outputs(855));
    layer1_outputs(2738) <= layer0_outputs(774);
    layer1_outputs(2739) <= not(layer0_outputs(9259));
    layer1_outputs(2740) <= (layer0_outputs(5156)) and not (layer0_outputs(9420));
    layer1_outputs(2741) <= not(layer0_outputs(1417));
    layer1_outputs(2742) <= not((layer0_outputs(8995)) and (layer0_outputs(9269)));
    layer1_outputs(2743) <= not((layer0_outputs(3013)) xor (layer0_outputs(3788)));
    layer1_outputs(2744) <= not(layer0_outputs(2353));
    layer1_outputs(2745) <= (layer0_outputs(5495)) and not (layer0_outputs(1712));
    layer1_outputs(2746) <= not((layer0_outputs(984)) and (layer0_outputs(4775)));
    layer1_outputs(2747) <= (layer0_outputs(5910)) and not (layer0_outputs(30));
    layer1_outputs(2748) <= (layer0_outputs(9780)) and not (layer0_outputs(3530));
    layer1_outputs(2749) <= (layer0_outputs(9531)) and (layer0_outputs(5159));
    layer1_outputs(2750) <= (layer0_outputs(9904)) and (layer0_outputs(9978));
    layer1_outputs(2751) <= not(layer0_outputs(5397)) or (layer0_outputs(9842));
    layer1_outputs(2752) <= (layer0_outputs(8750)) or (layer0_outputs(9407));
    layer1_outputs(2753) <= '0';
    layer1_outputs(2754) <= '1';
    layer1_outputs(2755) <= not(layer0_outputs(9894)) or (layer0_outputs(1825));
    layer1_outputs(2756) <= not(layer0_outputs(10148)) or (layer0_outputs(6447));
    layer1_outputs(2757) <= layer0_outputs(6595);
    layer1_outputs(2758) <= not(layer0_outputs(7094)) or (layer0_outputs(8681));
    layer1_outputs(2759) <= (layer0_outputs(2443)) or (layer0_outputs(1744));
    layer1_outputs(2760) <= (layer0_outputs(10053)) or (layer0_outputs(3628));
    layer1_outputs(2761) <= layer0_outputs(2605);
    layer1_outputs(2762) <= not((layer0_outputs(8402)) or (layer0_outputs(4222)));
    layer1_outputs(2763) <= not(layer0_outputs(1069));
    layer1_outputs(2764) <= not((layer0_outputs(400)) or (layer0_outputs(3142)));
    layer1_outputs(2765) <= (layer0_outputs(5373)) and (layer0_outputs(151));
    layer1_outputs(2766) <= layer0_outputs(10049);
    layer1_outputs(2767) <= layer0_outputs(5252);
    layer1_outputs(2768) <= not(layer0_outputs(7182));
    layer1_outputs(2769) <= layer0_outputs(6767);
    layer1_outputs(2770) <= '1';
    layer1_outputs(2771) <= not(layer0_outputs(9362));
    layer1_outputs(2772) <= (layer0_outputs(719)) and (layer0_outputs(2620));
    layer1_outputs(2773) <= layer0_outputs(452);
    layer1_outputs(2774) <= not((layer0_outputs(7409)) or (layer0_outputs(4128)));
    layer1_outputs(2775) <= not((layer0_outputs(8908)) xor (layer0_outputs(5099)));
    layer1_outputs(2776) <= (layer0_outputs(2529)) and (layer0_outputs(6798));
    layer1_outputs(2777) <= not((layer0_outputs(8380)) and (layer0_outputs(1520)));
    layer1_outputs(2778) <= not(layer0_outputs(5446)) or (layer0_outputs(2659));
    layer1_outputs(2779) <= not(layer0_outputs(6266)) or (layer0_outputs(2003));
    layer1_outputs(2780) <= not((layer0_outputs(9573)) or (layer0_outputs(8411)));
    layer1_outputs(2781) <= (layer0_outputs(6604)) and not (layer0_outputs(8046));
    layer1_outputs(2782) <= not((layer0_outputs(5026)) xor (layer0_outputs(7398)));
    layer1_outputs(2783) <= (layer0_outputs(5379)) and not (layer0_outputs(4627));
    layer1_outputs(2784) <= (layer0_outputs(106)) and (layer0_outputs(1978));
    layer1_outputs(2785) <= not((layer0_outputs(7359)) xor (layer0_outputs(7448)));
    layer1_outputs(2786) <= layer0_outputs(1568);
    layer1_outputs(2787) <= (layer0_outputs(2720)) and not (layer0_outputs(9541));
    layer1_outputs(2788) <= layer0_outputs(3550);
    layer1_outputs(2789) <= (layer0_outputs(2589)) and not (layer0_outputs(18));
    layer1_outputs(2790) <= not((layer0_outputs(5250)) and (layer0_outputs(747)));
    layer1_outputs(2791) <= (layer0_outputs(10224)) or (layer0_outputs(6048));
    layer1_outputs(2792) <= not(layer0_outputs(1949));
    layer1_outputs(2793) <= layer0_outputs(6257);
    layer1_outputs(2794) <= '1';
    layer1_outputs(2795) <= (layer0_outputs(1362)) and not (layer0_outputs(2411));
    layer1_outputs(2796) <= not(layer0_outputs(8451)) or (layer0_outputs(3361));
    layer1_outputs(2797) <= not(layer0_outputs(5860)) or (layer0_outputs(4432));
    layer1_outputs(2798) <= '1';
    layer1_outputs(2799) <= (layer0_outputs(5124)) and not (layer0_outputs(6648));
    layer1_outputs(2800) <= not((layer0_outputs(7117)) and (layer0_outputs(3854)));
    layer1_outputs(2801) <= (layer0_outputs(8627)) and not (layer0_outputs(8879));
    layer1_outputs(2802) <= layer0_outputs(5092);
    layer1_outputs(2803) <= (layer0_outputs(3726)) and not (layer0_outputs(4701));
    layer1_outputs(2804) <= (layer0_outputs(1732)) and (layer0_outputs(6425));
    layer1_outputs(2805) <= layer0_outputs(8986);
    layer1_outputs(2806) <= layer0_outputs(10048);
    layer1_outputs(2807) <= not(layer0_outputs(2897));
    layer1_outputs(2808) <= not(layer0_outputs(1941));
    layer1_outputs(2809) <= (layer0_outputs(7671)) and (layer0_outputs(8700));
    layer1_outputs(2810) <= not(layer0_outputs(9864));
    layer1_outputs(2811) <= not((layer0_outputs(4076)) xor (layer0_outputs(3878)));
    layer1_outputs(2812) <= (layer0_outputs(7260)) and not (layer0_outputs(5321));
    layer1_outputs(2813) <= not(layer0_outputs(8898));
    layer1_outputs(2814) <= not(layer0_outputs(7937)) or (layer0_outputs(5067));
    layer1_outputs(2815) <= (layer0_outputs(2340)) and not (layer0_outputs(324));
    layer1_outputs(2816) <= (layer0_outputs(1234)) or (layer0_outputs(9484));
    layer1_outputs(2817) <= (layer0_outputs(6983)) and not (layer0_outputs(284));
    layer1_outputs(2818) <= not((layer0_outputs(325)) and (layer0_outputs(9271)));
    layer1_outputs(2819) <= not(layer0_outputs(651));
    layer1_outputs(2820) <= (layer0_outputs(8441)) or (layer0_outputs(5166));
    layer1_outputs(2821) <= not(layer0_outputs(6820));
    layer1_outputs(2822) <= layer0_outputs(5484);
    layer1_outputs(2823) <= not((layer0_outputs(6060)) xor (layer0_outputs(5226)));
    layer1_outputs(2824) <= not(layer0_outputs(6803));
    layer1_outputs(2825) <= not(layer0_outputs(2723));
    layer1_outputs(2826) <= not(layer0_outputs(9452));
    layer1_outputs(2827) <= not((layer0_outputs(1563)) xor (layer0_outputs(6527)));
    layer1_outputs(2828) <= '1';
    layer1_outputs(2829) <= layer0_outputs(4960);
    layer1_outputs(2830) <= (layer0_outputs(5402)) and (layer0_outputs(2068));
    layer1_outputs(2831) <= layer0_outputs(2310);
    layer1_outputs(2832) <= not(layer0_outputs(57));
    layer1_outputs(2833) <= (layer0_outputs(5547)) or (layer0_outputs(7780));
    layer1_outputs(2834) <= not(layer0_outputs(1477));
    layer1_outputs(2835) <= not((layer0_outputs(6369)) and (layer0_outputs(5218)));
    layer1_outputs(2836) <= not((layer0_outputs(9004)) and (layer0_outputs(6773)));
    layer1_outputs(2837) <= not((layer0_outputs(6238)) or (layer0_outputs(1844)));
    layer1_outputs(2838) <= not(layer0_outputs(7555)) or (layer0_outputs(5137));
    layer1_outputs(2839) <= layer0_outputs(2400);
    layer1_outputs(2840) <= not(layer0_outputs(234)) or (layer0_outputs(1806));
    layer1_outputs(2841) <= not((layer0_outputs(6259)) or (layer0_outputs(9132)));
    layer1_outputs(2842) <= layer0_outputs(8250);
    layer1_outputs(2843) <= not((layer0_outputs(7435)) and (layer0_outputs(1017)));
    layer1_outputs(2844) <= '1';
    layer1_outputs(2845) <= (layer0_outputs(4578)) and not (layer0_outputs(4651));
    layer1_outputs(2846) <= layer0_outputs(4654);
    layer1_outputs(2847) <= not(layer0_outputs(10082)) or (layer0_outputs(3136));
    layer1_outputs(2848) <= not((layer0_outputs(5607)) or (layer0_outputs(3477)));
    layer1_outputs(2849) <= (layer0_outputs(6315)) and (layer0_outputs(344));
    layer1_outputs(2850) <= not((layer0_outputs(7618)) or (layer0_outputs(3727)));
    layer1_outputs(2851) <= (layer0_outputs(9410)) or (layer0_outputs(5136));
    layer1_outputs(2852) <= not(layer0_outputs(4209)) or (layer0_outputs(2535));
    layer1_outputs(2853) <= not(layer0_outputs(6479));
    layer1_outputs(2854) <= not((layer0_outputs(3155)) xor (layer0_outputs(6073)));
    layer1_outputs(2855) <= not(layer0_outputs(5045));
    layer1_outputs(2856) <= not((layer0_outputs(3437)) xor (layer0_outputs(3092)));
    layer1_outputs(2857) <= not(layer0_outputs(7191)) or (layer0_outputs(9237));
    layer1_outputs(2858) <= not(layer0_outputs(1706)) or (layer0_outputs(5293));
    layer1_outputs(2859) <= not(layer0_outputs(5065));
    layer1_outputs(2860) <= (layer0_outputs(862)) and not (layer0_outputs(3242));
    layer1_outputs(2861) <= layer0_outputs(2668);
    layer1_outputs(2862) <= (layer0_outputs(10151)) and not (layer0_outputs(8337));
    layer1_outputs(2863) <= (layer0_outputs(435)) or (layer0_outputs(8565));
    layer1_outputs(2864) <= (layer0_outputs(9921)) or (layer0_outputs(4950));
    layer1_outputs(2865) <= not(layer0_outputs(4554));
    layer1_outputs(2866) <= '1';
    layer1_outputs(2867) <= not(layer0_outputs(4694));
    layer1_outputs(2868) <= not(layer0_outputs(5211));
    layer1_outputs(2869) <= (layer0_outputs(8658)) and not (layer0_outputs(573));
    layer1_outputs(2870) <= (layer0_outputs(5956)) and not (layer0_outputs(3739));
    layer1_outputs(2871) <= layer0_outputs(6678);
    layer1_outputs(2872) <= layer0_outputs(7108);
    layer1_outputs(2873) <= not(layer0_outputs(1875));
    layer1_outputs(2874) <= not(layer0_outputs(10034)) or (layer0_outputs(2016));
    layer1_outputs(2875) <= (layer0_outputs(3624)) and not (layer0_outputs(2983));
    layer1_outputs(2876) <= (layer0_outputs(1669)) or (layer0_outputs(9470));
    layer1_outputs(2877) <= (layer0_outputs(2379)) and not (layer0_outputs(4050));
    layer1_outputs(2878) <= not(layer0_outputs(5873)) or (layer0_outputs(4610));
    layer1_outputs(2879) <= not((layer0_outputs(5007)) and (layer0_outputs(2686)));
    layer1_outputs(2880) <= not(layer0_outputs(218)) or (layer0_outputs(168));
    layer1_outputs(2881) <= layer0_outputs(8717);
    layer1_outputs(2882) <= not(layer0_outputs(9210));
    layer1_outputs(2883) <= not((layer0_outputs(3702)) and (layer0_outputs(9721)));
    layer1_outputs(2884) <= not(layer0_outputs(2307));
    layer1_outputs(2885) <= not(layer0_outputs(9310));
    layer1_outputs(2886) <= not(layer0_outputs(3936)) or (layer0_outputs(2611));
    layer1_outputs(2887) <= not((layer0_outputs(7998)) and (layer0_outputs(4386)));
    layer1_outputs(2888) <= not(layer0_outputs(2826)) or (layer0_outputs(308));
    layer1_outputs(2889) <= not(layer0_outputs(6491));
    layer1_outputs(2890) <= not(layer0_outputs(9667));
    layer1_outputs(2891) <= not(layer0_outputs(6403)) or (layer0_outputs(4931));
    layer1_outputs(2892) <= layer0_outputs(8839);
    layer1_outputs(2893) <= (layer0_outputs(7550)) and (layer0_outputs(3609));
    layer1_outputs(2894) <= layer0_outputs(5848);
    layer1_outputs(2895) <= not(layer0_outputs(8292));
    layer1_outputs(2896) <= not(layer0_outputs(6025)) or (layer0_outputs(8393));
    layer1_outputs(2897) <= (layer0_outputs(1944)) and not (layer0_outputs(2302));
    layer1_outputs(2898) <= layer0_outputs(4559);
    layer1_outputs(2899) <= (layer0_outputs(246)) and not (layer0_outputs(8969));
    layer1_outputs(2900) <= (layer0_outputs(185)) and not (layer0_outputs(418));
    layer1_outputs(2901) <= not(layer0_outputs(7306));
    layer1_outputs(2902) <= (layer0_outputs(9715)) or (layer0_outputs(2562));
    layer1_outputs(2903) <= not(layer0_outputs(2550)) or (layer0_outputs(8647));
    layer1_outputs(2904) <= (layer0_outputs(7518)) or (layer0_outputs(7570));
    layer1_outputs(2905) <= not((layer0_outputs(3508)) xor (layer0_outputs(4787)));
    layer1_outputs(2906) <= not((layer0_outputs(4983)) and (layer0_outputs(9689)));
    layer1_outputs(2907) <= not(layer0_outputs(9849)) or (layer0_outputs(5034));
    layer1_outputs(2908) <= not((layer0_outputs(7173)) or (layer0_outputs(4311)));
    layer1_outputs(2909) <= '0';
    layer1_outputs(2910) <= '1';
    layer1_outputs(2911) <= (layer0_outputs(191)) and not (layer0_outputs(2679));
    layer1_outputs(2912) <= layer0_outputs(4595);
    layer1_outputs(2913) <= not(layer0_outputs(9517));
    layer1_outputs(2914) <= layer0_outputs(6545);
    layer1_outputs(2915) <= (layer0_outputs(8639)) or (layer0_outputs(2246));
    layer1_outputs(2916) <= not((layer0_outputs(5182)) and (layer0_outputs(6316)));
    layer1_outputs(2917) <= layer0_outputs(4595);
    layer1_outputs(2918) <= layer0_outputs(5722);
    layer1_outputs(2919) <= (layer0_outputs(7289)) and (layer0_outputs(1888));
    layer1_outputs(2920) <= layer0_outputs(1873);
    layer1_outputs(2921) <= '1';
    layer1_outputs(2922) <= not(layer0_outputs(6287));
    layer1_outputs(2923) <= '1';
    layer1_outputs(2924) <= not(layer0_outputs(5109));
    layer1_outputs(2925) <= not(layer0_outputs(5437));
    layer1_outputs(2926) <= layer0_outputs(1019);
    layer1_outputs(2927) <= (layer0_outputs(2321)) and (layer0_outputs(9880));
    layer1_outputs(2928) <= not(layer0_outputs(2114)) or (layer0_outputs(3703));
    layer1_outputs(2929) <= not(layer0_outputs(6779));
    layer1_outputs(2930) <= not(layer0_outputs(237));
    layer1_outputs(2931) <= (layer0_outputs(6286)) or (layer0_outputs(209));
    layer1_outputs(2932) <= (layer0_outputs(1936)) and not (layer0_outputs(9553));
    layer1_outputs(2933) <= layer0_outputs(8588);
    layer1_outputs(2934) <= not(layer0_outputs(4441)) or (layer0_outputs(1500));
    layer1_outputs(2935) <= (layer0_outputs(3965)) and not (layer0_outputs(6586));
    layer1_outputs(2936) <= (layer0_outputs(1074)) and (layer0_outputs(6936));
    layer1_outputs(2937) <= not((layer0_outputs(1711)) xor (layer0_outputs(1160)));
    layer1_outputs(2938) <= layer0_outputs(4108);
    layer1_outputs(2939) <= not((layer0_outputs(149)) xor (layer0_outputs(9580)));
    layer1_outputs(2940) <= (layer0_outputs(1309)) xor (layer0_outputs(2975));
    layer1_outputs(2941) <= (layer0_outputs(1580)) and (layer0_outputs(6323));
    layer1_outputs(2942) <= not(layer0_outputs(6555));
    layer1_outputs(2943) <= (layer0_outputs(7684)) and not (layer0_outputs(4724));
    layer1_outputs(2944) <= (layer0_outputs(9084)) and (layer0_outputs(6409));
    layer1_outputs(2945) <= not((layer0_outputs(7512)) and (layer0_outputs(9160)));
    layer1_outputs(2946) <= not((layer0_outputs(4077)) or (layer0_outputs(3936)));
    layer1_outputs(2947) <= layer0_outputs(1336);
    layer1_outputs(2948) <= (layer0_outputs(8476)) and not (layer0_outputs(9645));
    layer1_outputs(2949) <= not(layer0_outputs(4186));
    layer1_outputs(2950) <= not(layer0_outputs(2456));
    layer1_outputs(2951) <= (layer0_outputs(10062)) or (layer0_outputs(3022));
    layer1_outputs(2952) <= not(layer0_outputs(4826)) or (layer0_outputs(4874));
    layer1_outputs(2953) <= not(layer0_outputs(3777));
    layer1_outputs(2954) <= layer0_outputs(10040);
    layer1_outputs(2955) <= layer0_outputs(9205);
    layer1_outputs(2956) <= not((layer0_outputs(9647)) xor (layer0_outputs(7487)));
    layer1_outputs(2957) <= layer0_outputs(7756);
    layer1_outputs(2958) <= layer0_outputs(3140);
    layer1_outputs(2959) <= layer0_outputs(5761);
    layer1_outputs(2960) <= layer0_outputs(10113);
    layer1_outputs(2961) <= not(layer0_outputs(6426));
    layer1_outputs(2962) <= (layer0_outputs(1033)) and not (layer0_outputs(7236));
    layer1_outputs(2963) <= not((layer0_outputs(7913)) or (layer0_outputs(478)));
    layer1_outputs(2964) <= (layer0_outputs(3736)) or (layer0_outputs(7238));
    layer1_outputs(2965) <= not(layer0_outputs(1400)) or (layer0_outputs(8586));
    layer1_outputs(2966) <= not(layer0_outputs(3608));
    layer1_outputs(2967) <= (layer0_outputs(3952)) and not (layer0_outputs(5051));
    layer1_outputs(2968) <= layer0_outputs(2514);
    layer1_outputs(2969) <= not(layer0_outputs(8347));
    layer1_outputs(2970) <= not(layer0_outputs(6992));
    layer1_outputs(2971) <= layer0_outputs(2830);
    layer1_outputs(2972) <= (layer0_outputs(4285)) or (layer0_outputs(9046));
    layer1_outputs(2973) <= (layer0_outputs(7459)) and not (layer0_outputs(3262));
    layer1_outputs(2974) <= (layer0_outputs(9440)) and (layer0_outputs(4371));
    layer1_outputs(2975) <= (layer0_outputs(114)) and not (layer0_outputs(9519));
    layer1_outputs(2976) <= not((layer0_outputs(6229)) xor (layer0_outputs(9948)));
    layer1_outputs(2977) <= not(layer0_outputs(1749));
    layer1_outputs(2978) <= layer0_outputs(8293);
    layer1_outputs(2979) <= not((layer0_outputs(10021)) or (layer0_outputs(9518)));
    layer1_outputs(2980) <= not((layer0_outputs(9383)) and (layer0_outputs(4948)));
    layer1_outputs(2981) <= not(layer0_outputs(2141));
    layer1_outputs(2982) <= layer0_outputs(4406);
    layer1_outputs(2983) <= layer0_outputs(6937);
    layer1_outputs(2984) <= not(layer0_outputs(5575)) or (layer0_outputs(3962));
    layer1_outputs(2985) <= (layer0_outputs(2649)) xor (layer0_outputs(6400));
    layer1_outputs(2986) <= not(layer0_outputs(7607)) or (layer0_outputs(2284));
    layer1_outputs(2987) <= (layer0_outputs(7088)) or (layer0_outputs(2951));
    layer1_outputs(2988) <= not(layer0_outputs(885)) or (layer0_outputs(7010));
    layer1_outputs(2989) <= (layer0_outputs(4501)) and not (layer0_outputs(8378));
    layer1_outputs(2990) <= not((layer0_outputs(4979)) or (layer0_outputs(1677)));
    layer1_outputs(2991) <= layer0_outputs(4862);
    layer1_outputs(2992) <= (layer0_outputs(8322)) and (layer0_outputs(1692));
    layer1_outputs(2993) <= not((layer0_outputs(9172)) and (layer0_outputs(1046)));
    layer1_outputs(2994) <= not(layer0_outputs(10061));
    layer1_outputs(2995) <= layer0_outputs(8935);
    layer1_outputs(2996) <= not((layer0_outputs(9014)) and (layer0_outputs(4920)));
    layer1_outputs(2997) <= not((layer0_outputs(8789)) and (layer0_outputs(6033)));
    layer1_outputs(2998) <= (layer0_outputs(6892)) and not (layer0_outputs(9763));
    layer1_outputs(2999) <= (layer0_outputs(1487)) and not (layer0_outputs(8011));
    layer1_outputs(3000) <= '0';
    layer1_outputs(3001) <= layer0_outputs(76);
    layer1_outputs(3002) <= (layer0_outputs(8796)) and not (layer0_outputs(6314));
    layer1_outputs(3003) <= not(layer0_outputs(2987));
    layer1_outputs(3004) <= not(layer0_outputs(5678));
    layer1_outputs(3005) <= (layer0_outputs(5320)) xor (layer0_outputs(2792));
    layer1_outputs(3006) <= not(layer0_outputs(362)) or (layer0_outputs(9381));
    layer1_outputs(3007) <= (layer0_outputs(5965)) and not (layer0_outputs(3565));
    layer1_outputs(3008) <= (layer0_outputs(6199)) and (layer0_outputs(8291));
    layer1_outputs(3009) <= not(layer0_outputs(4912));
    layer1_outputs(3010) <= not(layer0_outputs(10130));
    layer1_outputs(3011) <= layer0_outputs(4143);
    layer1_outputs(3012) <= not((layer0_outputs(2187)) or (layer0_outputs(509)));
    layer1_outputs(3013) <= not(layer0_outputs(9713));
    layer1_outputs(3014) <= layer0_outputs(1055);
    layer1_outputs(3015) <= not(layer0_outputs(2051)) or (layer0_outputs(8726));
    layer1_outputs(3016) <= not(layer0_outputs(6664));
    layer1_outputs(3017) <= (layer0_outputs(6251)) or (layer0_outputs(6941));
    layer1_outputs(3018) <= (layer0_outputs(672)) and not (layer0_outputs(7444));
    layer1_outputs(3019) <= not(layer0_outputs(4937));
    layer1_outputs(3020) <= layer0_outputs(2874);
    layer1_outputs(3021) <= (layer0_outputs(6699)) and (layer0_outputs(1455));
    layer1_outputs(3022) <= (layer0_outputs(4750)) and (layer0_outputs(4169));
    layer1_outputs(3023) <= not((layer0_outputs(3369)) or (layer0_outputs(565)));
    layer1_outputs(3024) <= not(layer0_outputs(9226));
    layer1_outputs(3025) <= (layer0_outputs(221)) or (layer0_outputs(2548));
    layer1_outputs(3026) <= layer0_outputs(9782);
    layer1_outputs(3027) <= (layer0_outputs(3334)) and not (layer0_outputs(5971));
    layer1_outputs(3028) <= layer0_outputs(5756);
    layer1_outputs(3029) <= not((layer0_outputs(3607)) or (layer0_outputs(2375)));
    layer1_outputs(3030) <= not(layer0_outputs(1933));
    layer1_outputs(3031) <= not(layer0_outputs(9111));
    layer1_outputs(3032) <= not((layer0_outputs(4963)) or (layer0_outputs(4246)));
    layer1_outputs(3033) <= not(layer0_outputs(3400));
    layer1_outputs(3034) <= not(layer0_outputs(9854)) or (layer0_outputs(711));
    layer1_outputs(3035) <= not((layer0_outputs(958)) xor (layer0_outputs(3283)));
    layer1_outputs(3036) <= not((layer0_outputs(7935)) xor (layer0_outputs(1924)));
    layer1_outputs(3037) <= layer0_outputs(9460);
    layer1_outputs(3038) <= (layer0_outputs(8698)) xor (layer0_outputs(2935));
    layer1_outputs(3039) <= not(layer0_outputs(9312));
    layer1_outputs(3040) <= not(layer0_outputs(7317));
    layer1_outputs(3041) <= (layer0_outputs(10146)) xor (layer0_outputs(9370));
    layer1_outputs(3042) <= not(layer0_outputs(4812));
    layer1_outputs(3043) <= not(layer0_outputs(8366)) or (layer0_outputs(5678));
    layer1_outputs(3044) <= not((layer0_outputs(5364)) or (layer0_outputs(1086)));
    layer1_outputs(3045) <= layer0_outputs(5138);
    layer1_outputs(3046) <= (layer0_outputs(9293)) xor (layer0_outputs(9764));
    layer1_outputs(3047) <= layer0_outputs(4812);
    layer1_outputs(3048) <= layer0_outputs(6860);
    layer1_outputs(3049) <= layer0_outputs(535);
    layer1_outputs(3050) <= layer0_outputs(9015);
    layer1_outputs(3051) <= not(layer0_outputs(9423));
    layer1_outputs(3052) <= (layer0_outputs(4901)) and not (layer0_outputs(429));
    layer1_outputs(3053) <= (layer0_outputs(2031)) xor (layer0_outputs(906));
    layer1_outputs(3054) <= not(layer0_outputs(5928));
    layer1_outputs(3055) <= not((layer0_outputs(958)) and (layer0_outputs(8534)));
    layer1_outputs(3056) <= (layer0_outputs(1423)) xor (layer0_outputs(6650));
    layer1_outputs(3057) <= layer0_outputs(4136);
    layer1_outputs(3058) <= layer0_outputs(8776);
    layer1_outputs(3059) <= layer0_outputs(4755);
    layer1_outputs(3060) <= not(layer0_outputs(4320));
    layer1_outputs(3061) <= (layer0_outputs(9684)) and not (layer0_outputs(1424));
    layer1_outputs(3062) <= (layer0_outputs(4496)) and not (layer0_outputs(5446));
    layer1_outputs(3063) <= layer0_outputs(2701);
    layer1_outputs(3064) <= layer0_outputs(117);
    layer1_outputs(3065) <= not((layer0_outputs(4890)) xor (layer0_outputs(3301)));
    layer1_outputs(3066) <= (layer0_outputs(6203)) xor (layer0_outputs(244));
    layer1_outputs(3067) <= layer0_outputs(3591);
    layer1_outputs(3068) <= (layer0_outputs(3368)) and (layer0_outputs(7244));
    layer1_outputs(3069) <= (layer0_outputs(3208)) and (layer0_outputs(718));
    layer1_outputs(3070) <= (layer0_outputs(2163)) xor (layer0_outputs(9528));
    layer1_outputs(3071) <= not(layer0_outputs(1646));
    layer1_outputs(3072) <= layer0_outputs(352);
    layer1_outputs(3073) <= not(layer0_outputs(9460)) or (layer0_outputs(7251));
    layer1_outputs(3074) <= not((layer0_outputs(68)) and (layer0_outputs(835)));
    layer1_outputs(3075) <= not((layer0_outputs(6313)) and (layer0_outputs(3241)));
    layer1_outputs(3076) <= not(layer0_outputs(1681));
    layer1_outputs(3077) <= not(layer0_outputs(8271));
    layer1_outputs(3078) <= layer0_outputs(7962);
    layer1_outputs(3079) <= layer0_outputs(3925);
    layer1_outputs(3080) <= not(layer0_outputs(3644)) or (layer0_outputs(695));
    layer1_outputs(3081) <= not(layer0_outputs(5617));
    layer1_outputs(3082) <= not((layer0_outputs(1314)) or (layer0_outputs(8618)));
    layer1_outputs(3083) <= not(layer0_outputs(8938));
    layer1_outputs(3084) <= not((layer0_outputs(9923)) or (layer0_outputs(5514)));
    layer1_outputs(3085) <= (layer0_outputs(1045)) and not (layer0_outputs(7723));
    layer1_outputs(3086) <= (layer0_outputs(7150)) and not (layer0_outputs(8280));
    layer1_outputs(3087) <= (layer0_outputs(2145)) or (layer0_outputs(2923));
    layer1_outputs(3088) <= layer0_outputs(6041);
    layer1_outputs(3089) <= layer0_outputs(4943);
    layer1_outputs(3090) <= not(layer0_outputs(6957));
    layer1_outputs(3091) <= not(layer0_outputs(317));
    layer1_outputs(3092) <= not(layer0_outputs(966)) or (layer0_outputs(2457));
    layer1_outputs(3093) <= (layer0_outputs(5986)) or (layer0_outputs(880));
    layer1_outputs(3094) <= (layer0_outputs(9897)) and not (layer0_outputs(525));
    layer1_outputs(3095) <= not(layer0_outputs(2135));
    layer1_outputs(3096) <= (layer0_outputs(4126)) and (layer0_outputs(2190));
    layer1_outputs(3097) <= not((layer0_outputs(9560)) xor (layer0_outputs(8649)));
    layer1_outputs(3098) <= (layer0_outputs(1147)) and not (layer0_outputs(2204));
    layer1_outputs(3099) <= not(layer0_outputs(1413));
    layer1_outputs(3100) <= not((layer0_outputs(3755)) or (layer0_outputs(5364)));
    layer1_outputs(3101) <= layer0_outputs(6995);
    layer1_outputs(3102) <= (layer0_outputs(4278)) and not (layer0_outputs(7254));
    layer1_outputs(3103) <= (layer0_outputs(233)) and not (layer0_outputs(9935));
    layer1_outputs(3104) <= (layer0_outputs(3229)) and not (layer0_outputs(8089));
    layer1_outputs(3105) <= not(layer0_outputs(1780));
    layer1_outputs(3106) <= (layer0_outputs(6090)) xor (layer0_outputs(4143));
    layer1_outputs(3107) <= layer0_outputs(3058);
    layer1_outputs(3108) <= (layer0_outputs(2568)) and (layer0_outputs(5484));
    layer1_outputs(3109) <= not((layer0_outputs(9307)) and (layer0_outputs(1065)));
    layer1_outputs(3110) <= not(layer0_outputs(8819)) or (layer0_outputs(5499));
    layer1_outputs(3111) <= not(layer0_outputs(1311));
    layer1_outputs(3112) <= not(layer0_outputs(9940)) or (layer0_outputs(919));
    layer1_outputs(3113) <= (layer0_outputs(3132)) and not (layer0_outputs(6857));
    layer1_outputs(3114) <= not(layer0_outputs(9083));
    layer1_outputs(3115) <= not(layer0_outputs(7460)) or (layer0_outputs(8115));
    layer1_outputs(3116) <= not(layer0_outputs(3865));
    layer1_outputs(3117) <= layer0_outputs(4178);
    layer1_outputs(3118) <= not(layer0_outputs(1996));
    layer1_outputs(3119) <= not((layer0_outputs(2171)) or (layer0_outputs(6376)));
    layer1_outputs(3120) <= not(layer0_outputs(9915));
    layer1_outputs(3121) <= (layer0_outputs(3526)) xor (layer0_outputs(9200));
    layer1_outputs(3122) <= (layer0_outputs(9075)) or (layer0_outputs(8202));
    layer1_outputs(3123) <= (layer0_outputs(5712)) or (layer0_outputs(6508));
    layer1_outputs(3124) <= not(layer0_outputs(3133));
    layer1_outputs(3125) <= not(layer0_outputs(390));
    layer1_outputs(3126) <= (layer0_outputs(2287)) or (layer0_outputs(6060));
    layer1_outputs(3127) <= not(layer0_outputs(4869)) or (layer0_outputs(8787));
    layer1_outputs(3128) <= layer0_outputs(9466);
    layer1_outputs(3129) <= (layer0_outputs(9831)) or (layer0_outputs(4155));
    layer1_outputs(3130) <= not(layer0_outputs(3581)) or (layer0_outputs(9412));
    layer1_outputs(3131) <= not(layer0_outputs(8466)) or (layer0_outputs(2973));
    layer1_outputs(3132) <= not(layer0_outputs(2811)) or (layer0_outputs(1982));
    layer1_outputs(3133) <= (layer0_outputs(7420)) and (layer0_outputs(123));
    layer1_outputs(3134) <= layer0_outputs(118);
    layer1_outputs(3135) <= not((layer0_outputs(2812)) xor (layer0_outputs(7816)));
    layer1_outputs(3136) <= not(layer0_outputs(3358)) or (layer0_outputs(9982));
    layer1_outputs(3137) <= not(layer0_outputs(9466));
    layer1_outputs(3138) <= layer0_outputs(1053);
    layer1_outputs(3139) <= not(layer0_outputs(7097));
    layer1_outputs(3140) <= not(layer0_outputs(9491)) or (layer0_outputs(8172));
    layer1_outputs(3141) <= not((layer0_outputs(8300)) or (layer0_outputs(8121)));
    layer1_outputs(3142) <= not(layer0_outputs(3930));
    layer1_outputs(3143) <= (layer0_outputs(5989)) and not (layer0_outputs(8788));
    layer1_outputs(3144) <= not(layer0_outputs(9914));
    layer1_outputs(3145) <= (layer0_outputs(2102)) xor (layer0_outputs(8178));
    layer1_outputs(3146) <= (layer0_outputs(3594)) and not (layer0_outputs(6820));
    layer1_outputs(3147) <= not(layer0_outputs(3007));
    layer1_outputs(3148) <= layer0_outputs(9703);
    layer1_outputs(3149) <= not(layer0_outputs(10142));
    layer1_outputs(3150) <= not((layer0_outputs(2354)) and (layer0_outputs(5807)));
    layer1_outputs(3151) <= layer0_outputs(2828);
    layer1_outputs(3152) <= (layer0_outputs(3787)) and (layer0_outputs(6858));
    layer1_outputs(3153) <= not((layer0_outputs(5173)) or (layer0_outputs(3512)));
    layer1_outputs(3154) <= layer0_outputs(9947);
    layer1_outputs(3155) <= layer0_outputs(3080);
    layer1_outputs(3156) <= (layer0_outputs(8295)) and (layer0_outputs(1334));
    layer1_outputs(3157) <= not((layer0_outputs(7053)) or (layer0_outputs(2011)));
    layer1_outputs(3158) <= '0';
    layer1_outputs(3159) <= layer0_outputs(4171);
    layer1_outputs(3160) <= (layer0_outputs(6387)) and not (layer0_outputs(6684));
    layer1_outputs(3161) <= not(layer0_outputs(8434)) or (layer0_outputs(6241));
    layer1_outputs(3162) <= layer0_outputs(8064);
    layer1_outputs(3163) <= layer0_outputs(6640);
    layer1_outputs(3164) <= not((layer0_outputs(878)) and (layer0_outputs(1599)));
    layer1_outputs(3165) <= (layer0_outputs(1547)) and not (layer0_outputs(5875));
    layer1_outputs(3166) <= '1';
    layer1_outputs(3167) <= (layer0_outputs(416)) and (layer0_outputs(4083));
    layer1_outputs(3168) <= not((layer0_outputs(4266)) or (layer0_outputs(1620)));
    layer1_outputs(3169) <= (layer0_outputs(5256)) xor (layer0_outputs(2070));
    layer1_outputs(3170) <= (layer0_outputs(6553)) and (layer0_outputs(1472));
    layer1_outputs(3171) <= layer0_outputs(5105);
    layer1_outputs(3172) <= (layer0_outputs(10096)) and not (layer0_outputs(3004));
    layer1_outputs(3173) <= not((layer0_outputs(2157)) and (layer0_outputs(4424)));
    layer1_outputs(3174) <= layer0_outputs(6984);
    layer1_outputs(3175) <= '0';
    layer1_outputs(3176) <= layer0_outputs(2646);
    layer1_outputs(3177) <= not((layer0_outputs(4567)) xor (layer0_outputs(3026)));
    layer1_outputs(3178) <= (layer0_outputs(9604)) and not (layer0_outputs(291));
    layer1_outputs(3179) <= (layer0_outputs(5563)) and not (layer0_outputs(10128));
    layer1_outputs(3180) <= not(layer0_outputs(7585)) or (layer0_outputs(4074));
    layer1_outputs(3181) <= '1';
    layer1_outputs(3182) <= not(layer0_outputs(3139));
    layer1_outputs(3183) <= (layer0_outputs(7016)) or (layer0_outputs(6140));
    layer1_outputs(3184) <= layer0_outputs(9300);
    layer1_outputs(3185) <= not(layer0_outputs(4390)) or (layer0_outputs(7104));
    layer1_outputs(3186) <= not(layer0_outputs(8281));
    layer1_outputs(3187) <= layer0_outputs(4535);
    layer1_outputs(3188) <= not((layer0_outputs(1649)) and (layer0_outputs(750)));
    layer1_outputs(3189) <= (layer0_outputs(7667)) or (layer0_outputs(9145));
    layer1_outputs(3190) <= not(layer0_outputs(5227));
    layer1_outputs(3191) <= not(layer0_outputs(7064)) or (layer0_outputs(9902));
    layer1_outputs(3192) <= (layer0_outputs(558)) xor (layer0_outputs(1498));
    layer1_outputs(3193) <= not((layer0_outputs(945)) xor (layer0_outputs(3665)));
    layer1_outputs(3194) <= not(layer0_outputs(7702)) or (layer0_outputs(2776));
    layer1_outputs(3195) <= (layer0_outputs(8447)) or (layer0_outputs(2125));
    layer1_outputs(3196) <= not((layer0_outputs(4151)) xor (layer0_outputs(8384)));
    layer1_outputs(3197) <= layer0_outputs(2796);
    layer1_outputs(3198) <= not(layer0_outputs(3082)) or (layer0_outputs(2328));
    layer1_outputs(3199) <= layer0_outputs(8513);
    layer1_outputs(3200) <= not((layer0_outputs(6002)) or (layer0_outputs(6775)));
    layer1_outputs(3201) <= not(layer0_outputs(913));
    layer1_outputs(3202) <= not((layer0_outputs(5658)) and (layer0_outputs(6973)));
    layer1_outputs(3203) <= layer0_outputs(6630);
    layer1_outputs(3204) <= '0';
    layer1_outputs(3205) <= (layer0_outputs(9398)) and not (layer0_outputs(7235));
    layer1_outputs(3206) <= not(layer0_outputs(8761)) or (layer0_outputs(5151));
    layer1_outputs(3207) <= not(layer0_outputs(3037));
    layer1_outputs(3208) <= (layer0_outputs(2343)) or (layer0_outputs(3307));
    layer1_outputs(3209) <= not(layer0_outputs(6625));
    layer1_outputs(3210) <= not(layer0_outputs(7304));
    layer1_outputs(3211) <= not(layer0_outputs(959));
    layer1_outputs(3212) <= not(layer0_outputs(1374));
    layer1_outputs(3213) <= not(layer0_outputs(8896)) or (layer0_outputs(2128));
    layer1_outputs(3214) <= layer0_outputs(583);
    layer1_outputs(3215) <= (layer0_outputs(933)) and not (layer0_outputs(4328));
    layer1_outputs(3216) <= (layer0_outputs(2434)) or (layer0_outputs(9478));
    layer1_outputs(3217) <= not(layer0_outputs(3853));
    layer1_outputs(3218) <= (layer0_outputs(6838)) and (layer0_outputs(4949));
    layer1_outputs(3219) <= not(layer0_outputs(1547));
    layer1_outputs(3220) <= (layer0_outputs(769)) and not (layer0_outputs(9598));
    layer1_outputs(3221) <= (layer0_outputs(9512)) and not (layer0_outputs(6202));
    layer1_outputs(3222) <= not(layer0_outputs(6812));
    layer1_outputs(3223) <= (layer0_outputs(5187)) or (layer0_outputs(6765));
    layer1_outputs(3224) <= not(layer0_outputs(1748));
    layer1_outputs(3225) <= (layer0_outputs(2118)) and not (layer0_outputs(6312));
    layer1_outputs(3226) <= not(layer0_outputs(4629));
    layer1_outputs(3227) <= (layer0_outputs(4046)) xor (layer0_outputs(729));
    layer1_outputs(3228) <= layer0_outputs(8082);
    layer1_outputs(3229) <= not((layer0_outputs(2796)) and (layer0_outputs(4456)));
    layer1_outputs(3230) <= (layer0_outputs(9414)) or (layer0_outputs(9149));
    layer1_outputs(3231) <= layer0_outputs(4961);
    layer1_outputs(3232) <= layer0_outputs(6920);
    layer1_outputs(3233) <= not(layer0_outputs(9971));
    layer1_outputs(3234) <= (layer0_outputs(8595)) and (layer0_outputs(4020));
    layer1_outputs(3235) <= not((layer0_outputs(686)) or (layer0_outputs(9443)));
    layer1_outputs(3236) <= not(layer0_outputs(8601)) or (layer0_outputs(9147));
    layer1_outputs(3237) <= not((layer0_outputs(9071)) or (layer0_outputs(8680)));
    layer1_outputs(3238) <= not((layer0_outputs(2278)) or (layer0_outputs(1088)));
    layer1_outputs(3239) <= layer0_outputs(6599);
    layer1_outputs(3240) <= layer0_outputs(3902);
    layer1_outputs(3241) <= '0';
    layer1_outputs(3242) <= '0';
    layer1_outputs(3243) <= '1';
    layer1_outputs(3244) <= not(layer0_outputs(8186));
    layer1_outputs(3245) <= layer0_outputs(7382);
    layer1_outputs(3246) <= (layer0_outputs(5050)) and (layer0_outputs(4716));
    layer1_outputs(3247) <= layer0_outputs(5973);
    layer1_outputs(3248) <= '0';
    layer1_outputs(3249) <= layer0_outputs(3374);
    layer1_outputs(3250) <= (layer0_outputs(7511)) and not (layer0_outputs(474));
    layer1_outputs(3251) <= not((layer0_outputs(8679)) and (layer0_outputs(9553)));
    layer1_outputs(3252) <= not(layer0_outputs(9833));
    layer1_outputs(3253) <= layer0_outputs(8925);
    layer1_outputs(3254) <= layer0_outputs(3078);
    layer1_outputs(3255) <= layer0_outputs(326);
    layer1_outputs(3256) <= layer0_outputs(3103);
    layer1_outputs(3257) <= layer0_outputs(3846);
    layer1_outputs(3258) <= not(layer0_outputs(4926));
    layer1_outputs(3259) <= not((layer0_outputs(5294)) or (layer0_outputs(2753)));
    layer1_outputs(3260) <= layer0_outputs(4369);
    layer1_outputs(3261) <= layer0_outputs(4479);
    layer1_outputs(3262) <= (layer0_outputs(1878)) and (layer0_outputs(5138));
    layer1_outputs(3263) <= not((layer0_outputs(7181)) or (layer0_outputs(5319)));
    layer1_outputs(3264) <= not((layer0_outputs(7293)) or (layer0_outputs(9872)));
    layer1_outputs(3265) <= layer0_outputs(2390);
    layer1_outputs(3266) <= layer0_outputs(5563);
    layer1_outputs(3267) <= (layer0_outputs(7083)) and not (layer0_outputs(9720));
    layer1_outputs(3268) <= (layer0_outputs(9869)) and not (layer0_outputs(3948));
    layer1_outputs(3269) <= not(layer0_outputs(10073));
    layer1_outputs(3270) <= (layer0_outputs(338)) or (layer0_outputs(2079));
    layer1_outputs(3271) <= not(layer0_outputs(389));
    layer1_outputs(3272) <= (layer0_outputs(9489)) or (layer0_outputs(8824));
    layer1_outputs(3273) <= (layer0_outputs(1608)) and not (layer0_outputs(3738));
    layer1_outputs(3274) <= (layer0_outputs(8318)) and (layer0_outputs(1849));
    layer1_outputs(3275) <= not((layer0_outputs(4193)) or (layer0_outputs(9192)));
    layer1_outputs(3276) <= (layer0_outputs(807)) and not (layer0_outputs(921));
    layer1_outputs(3277) <= not(layer0_outputs(6320));
    layer1_outputs(3278) <= not(layer0_outputs(7822)) or (layer0_outputs(8233));
    layer1_outputs(3279) <= not(layer0_outputs(8547)) or (layer0_outputs(2819));
    layer1_outputs(3280) <= not(layer0_outputs(5054)) or (layer0_outputs(3263));
    layer1_outputs(3281) <= not(layer0_outputs(4432));
    layer1_outputs(3282) <= not(layer0_outputs(2766));
    layer1_outputs(3283) <= not(layer0_outputs(2008));
    layer1_outputs(3284) <= layer0_outputs(1116);
    layer1_outputs(3285) <= layer0_outputs(216);
    layer1_outputs(3286) <= (layer0_outputs(9645)) and not (layer0_outputs(5789));
    layer1_outputs(3287) <= not(layer0_outputs(2335)) or (layer0_outputs(4627));
    layer1_outputs(3288) <= layer0_outputs(6552);
    layer1_outputs(3289) <= not((layer0_outputs(5347)) xor (layer0_outputs(2250)));
    layer1_outputs(3290) <= (layer0_outputs(265)) xor (layer0_outputs(4189));
    layer1_outputs(3291) <= (layer0_outputs(3465)) and not (layer0_outputs(4668));
    layer1_outputs(3292) <= not((layer0_outputs(9476)) or (layer0_outputs(2868)));
    layer1_outputs(3293) <= (layer0_outputs(1892)) and (layer0_outputs(4276));
    layer1_outputs(3294) <= not((layer0_outputs(6653)) and (layer0_outputs(10176)));
    layer1_outputs(3295) <= (layer0_outputs(528)) and not (layer0_outputs(8790));
    layer1_outputs(3296) <= not(layer0_outputs(7049));
    layer1_outputs(3297) <= layer0_outputs(6647);
    layer1_outputs(3298) <= not(layer0_outputs(6810)) or (layer0_outputs(6096));
    layer1_outputs(3299) <= layer0_outputs(9584);
    layer1_outputs(3300) <= (layer0_outputs(8860)) and not (layer0_outputs(9043));
    layer1_outputs(3301) <= not(layer0_outputs(9606));
    layer1_outputs(3302) <= not(layer0_outputs(7033));
    layer1_outputs(3303) <= not(layer0_outputs(9383));
    layer1_outputs(3304) <= (layer0_outputs(4786)) and not (layer0_outputs(4619));
    layer1_outputs(3305) <= not(layer0_outputs(1607)) or (layer0_outputs(5870));
    layer1_outputs(3306) <= layer0_outputs(8236);
    layer1_outputs(3307) <= (layer0_outputs(2630)) and not (layer0_outputs(3010));
    layer1_outputs(3308) <= not(layer0_outputs(2191)) or (layer0_outputs(7081));
    layer1_outputs(3309) <= not((layer0_outputs(2491)) and (layer0_outputs(8881)));
    layer1_outputs(3310) <= '0';
    layer1_outputs(3311) <= layer0_outputs(6854);
    layer1_outputs(3312) <= layer0_outputs(2829);
    layer1_outputs(3313) <= (layer0_outputs(7173)) and not (layer0_outputs(5847));
    layer1_outputs(3314) <= not(layer0_outputs(605));
    layer1_outputs(3315) <= not(layer0_outputs(7469));
    layer1_outputs(3316) <= not((layer0_outputs(7333)) or (layer0_outputs(7517)));
    layer1_outputs(3317) <= not(layer0_outputs(9688));
    layer1_outputs(3318) <= (layer0_outputs(3357)) and (layer0_outputs(5408));
    layer1_outputs(3319) <= not(layer0_outputs(4371));
    layer1_outputs(3320) <= (layer0_outputs(7196)) and not (layer0_outputs(1634));
    layer1_outputs(3321) <= (layer0_outputs(7031)) and (layer0_outputs(5359));
    layer1_outputs(3322) <= (layer0_outputs(8772)) or (layer0_outputs(6958));
    layer1_outputs(3323) <= layer0_outputs(4326);
    layer1_outputs(3324) <= (layer0_outputs(6249)) and not (layer0_outputs(1183));
    layer1_outputs(3325) <= layer0_outputs(7865);
    layer1_outputs(3326) <= (layer0_outputs(9321)) xor (layer0_outputs(7987));
    layer1_outputs(3327) <= (layer0_outputs(2968)) and not (layer0_outputs(493));
    layer1_outputs(3328) <= (layer0_outputs(3307)) xor (layer0_outputs(3221));
    layer1_outputs(3329) <= (layer0_outputs(9828)) and (layer0_outputs(98));
    layer1_outputs(3330) <= not((layer0_outputs(5729)) and (layer0_outputs(7608)));
    layer1_outputs(3331) <= layer0_outputs(465);
    layer1_outputs(3332) <= (layer0_outputs(805)) and not (layer0_outputs(751));
    layer1_outputs(3333) <= (layer0_outputs(7499)) and (layer0_outputs(4757));
    layer1_outputs(3334) <= not(layer0_outputs(9364));
    layer1_outputs(3335) <= not((layer0_outputs(4544)) or (layer0_outputs(6690)));
    layer1_outputs(3336) <= (layer0_outputs(6856)) and not (layer0_outputs(92));
    layer1_outputs(3337) <= layer0_outputs(7748);
    layer1_outputs(3338) <= not(layer0_outputs(7815)) or (layer0_outputs(7226));
    layer1_outputs(3339) <= (layer0_outputs(5456)) or (layer0_outputs(1357));
    layer1_outputs(3340) <= layer0_outputs(5526);
    layer1_outputs(3341) <= layer0_outputs(8055);
    layer1_outputs(3342) <= not(layer0_outputs(7750)) or (layer0_outputs(4655));
    layer1_outputs(3343) <= layer0_outputs(8820);
    layer1_outputs(3344) <= not(layer0_outputs(5869)) or (layer0_outputs(6114));
    layer1_outputs(3345) <= not(layer0_outputs(514));
    layer1_outputs(3346) <= layer0_outputs(7487);
    layer1_outputs(3347) <= not((layer0_outputs(1284)) xor (layer0_outputs(9142)));
    layer1_outputs(3348) <= layer0_outputs(4666);
    layer1_outputs(3349) <= layer0_outputs(6041);
    layer1_outputs(3350) <= not(layer0_outputs(7912)) or (layer0_outputs(4202));
    layer1_outputs(3351) <= not((layer0_outputs(9404)) and (layer0_outputs(2352)));
    layer1_outputs(3352) <= not(layer0_outputs(1519));
    layer1_outputs(3353) <= not(layer0_outputs(2275));
    layer1_outputs(3354) <= (layer0_outputs(8597)) and not (layer0_outputs(4363));
    layer1_outputs(3355) <= not(layer0_outputs(7876));
    layer1_outputs(3356) <= not(layer0_outputs(7760));
    layer1_outputs(3357) <= layer0_outputs(1773);
    layer1_outputs(3358) <= (layer0_outputs(8947)) and (layer0_outputs(2380));
    layer1_outputs(3359) <= not(layer0_outputs(6826));
    layer1_outputs(3360) <= layer0_outputs(5703);
    layer1_outputs(3361) <= (layer0_outputs(5711)) xor (layer0_outputs(3808));
    layer1_outputs(3362) <= not(layer0_outputs(8005));
    layer1_outputs(3363) <= layer0_outputs(2432);
    layer1_outputs(3364) <= layer0_outputs(6594);
    layer1_outputs(3365) <= (layer0_outputs(2278)) xor (layer0_outputs(8991));
    layer1_outputs(3366) <= not((layer0_outputs(7367)) xor (layer0_outputs(2099)));
    layer1_outputs(3367) <= not((layer0_outputs(1632)) and (layer0_outputs(9841)));
    layer1_outputs(3368) <= not((layer0_outputs(155)) xor (layer0_outputs(8798)));
    layer1_outputs(3369) <= not(layer0_outputs(8724)) or (layer0_outputs(8849));
    layer1_outputs(3370) <= not(layer0_outputs(5137)) or (layer0_outputs(2711));
    layer1_outputs(3371) <= not(layer0_outputs(1645));
    layer1_outputs(3372) <= (layer0_outputs(6645)) or (layer0_outputs(3411));
    layer1_outputs(3373) <= not(layer0_outputs(7099));
    layer1_outputs(3374) <= layer0_outputs(2135);
    layer1_outputs(3375) <= (layer0_outputs(1990)) xor (layer0_outputs(7533));
    layer1_outputs(3376) <= not(layer0_outputs(8533)) or (layer0_outputs(4467));
    layer1_outputs(3377) <= layer0_outputs(3824);
    layer1_outputs(3378) <= (layer0_outputs(1428)) and not (layer0_outputs(2020));
    layer1_outputs(3379) <= not((layer0_outputs(1123)) and (layer0_outputs(900)));
    layer1_outputs(3380) <= layer0_outputs(4035);
    layer1_outputs(3381) <= layer0_outputs(5975);
    layer1_outputs(3382) <= not((layer0_outputs(2722)) and (layer0_outputs(2333)));
    layer1_outputs(3383) <= not(layer0_outputs(6166)) or (layer0_outputs(5559));
    layer1_outputs(3384) <= not(layer0_outputs(121));
    layer1_outputs(3385) <= not(layer0_outputs(2131));
    layer1_outputs(3386) <= layer0_outputs(4102);
    layer1_outputs(3387) <= layer0_outputs(4316);
    layer1_outputs(3388) <= not(layer0_outputs(2368));
    layer1_outputs(3389) <= layer0_outputs(7146);
    layer1_outputs(3390) <= '1';
    layer1_outputs(3391) <= not(layer0_outputs(6560));
    layer1_outputs(3392) <= (layer0_outputs(7)) or (layer0_outputs(1633));
    layer1_outputs(3393) <= not((layer0_outputs(5019)) and (layer0_outputs(2089)));
    layer1_outputs(3394) <= '1';
    layer1_outputs(3395) <= layer0_outputs(7599);
    layer1_outputs(3396) <= layer0_outputs(7177);
    layer1_outputs(3397) <= not(layer0_outputs(8909));
    layer1_outputs(3398) <= layer0_outputs(951);
    layer1_outputs(3399) <= (layer0_outputs(2021)) or (layer0_outputs(3887));
    layer1_outputs(3400) <= not(layer0_outputs(7395));
    layer1_outputs(3401) <= not(layer0_outputs(7829)) or (layer0_outputs(5024));
    layer1_outputs(3402) <= (layer0_outputs(7022)) and (layer0_outputs(3044));
    layer1_outputs(3403) <= not(layer0_outputs(4266)) or (layer0_outputs(2972));
    layer1_outputs(3404) <= layer0_outputs(1665);
    layer1_outputs(3405) <= (layer0_outputs(2879)) and not (layer0_outputs(5530));
    layer1_outputs(3406) <= not(layer0_outputs(6367));
    layer1_outputs(3407) <= not((layer0_outputs(5004)) and (layer0_outputs(1875)));
    layer1_outputs(3408) <= (layer0_outputs(7609)) or (layer0_outputs(1436));
    layer1_outputs(3409) <= not((layer0_outputs(772)) xor (layer0_outputs(7066)));
    layer1_outputs(3410) <= not((layer0_outputs(3124)) xor (layer0_outputs(9533)));
    layer1_outputs(3411) <= not((layer0_outputs(6876)) or (layer0_outputs(688)));
    layer1_outputs(3412) <= layer0_outputs(8104);
    layer1_outputs(3413) <= not(layer0_outputs(4200)) or (layer0_outputs(2739));
    layer1_outputs(3414) <= not((layer0_outputs(8867)) xor (layer0_outputs(429)));
    layer1_outputs(3415) <= layer0_outputs(4527);
    layer1_outputs(3416) <= (layer0_outputs(6372)) and not (layer0_outputs(8350));
    layer1_outputs(3417) <= layer0_outputs(4610);
    layer1_outputs(3418) <= (layer0_outputs(5607)) and not (layer0_outputs(8349));
    layer1_outputs(3419) <= (layer0_outputs(5756)) xor (layer0_outputs(1189));
    layer1_outputs(3420) <= '1';
    layer1_outputs(3421) <= (layer0_outputs(3011)) and not (layer0_outputs(3534));
    layer1_outputs(3422) <= (layer0_outputs(7138)) xor (layer0_outputs(4948));
    layer1_outputs(3423) <= not(layer0_outputs(6165));
    layer1_outputs(3424) <= (layer0_outputs(5831)) and (layer0_outputs(4406));
    layer1_outputs(3425) <= not(layer0_outputs(9498)) or (layer0_outputs(8449));
    layer1_outputs(3426) <= layer0_outputs(894);
    layer1_outputs(3427) <= not((layer0_outputs(1959)) xor (layer0_outputs(3860)));
    layer1_outputs(3428) <= not((layer0_outputs(6209)) and (layer0_outputs(1500)));
    layer1_outputs(3429) <= not((layer0_outputs(9123)) or (layer0_outputs(4273)));
    layer1_outputs(3430) <= layer0_outputs(9150);
    layer1_outputs(3431) <= not((layer0_outputs(2696)) or (layer0_outputs(6786)));
    layer1_outputs(3432) <= (layer0_outputs(3659)) and not (layer0_outputs(2083));
    layer1_outputs(3433) <= (layer0_outputs(5622)) and (layer0_outputs(5981));
    layer1_outputs(3434) <= not((layer0_outputs(6536)) or (layer0_outputs(5190)));
    layer1_outputs(3435) <= layer0_outputs(2957);
    layer1_outputs(3436) <= not(layer0_outputs(3353));
    layer1_outputs(3437) <= not((layer0_outputs(6154)) xor (layer0_outputs(1254)));
    layer1_outputs(3438) <= layer0_outputs(4121);
    layer1_outputs(3439) <= layer0_outputs(3748);
    layer1_outputs(3440) <= (layer0_outputs(8949)) and (layer0_outputs(76));
    layer1_outputs(3441) <= (layer0_outputs(1920)) or (layer0_outputs(3849));
    layer1_outputs(3442) <= not(layer0_outputs(3667)) or (layer0_outputs(1952));
    layer1_outputs(3443) <= (layer0_outputs(434)) or (layer0_outputs(1159));
    layer1_outputs(3444) <= (layer0_outputs(590)) and not (layer0_outputs(7809));
    layer1_outputs(3445) <= (layer0_outputs(3091)) or (layer0_outputs(6637));
    layer1_outputs(3446) <= not((layer0_outputs(1367)) and (layer0_outputs(9962)));
    layer1_outputs(3447) <= not(layer0_outputs(7751));
    layer1_outputs(3448) <= layer0_outputs(6139);
    layer1_outputs(3449) <= layer0_outputs(6430);
    layer1_outputs(3450) <= layer0_outputs(2868);
    layer1_outputs(3451) <= (layer0_outputs(8240)) and not (layer0_outputs(2671));
    layer1_outputs(3452) <= not(layer0_outputs(2271));
    layer1_outputs(3453) <= not(layer0_outputs(7698)) or (layer0_outputs(5240));
    layer1_outputs(3454) <= (layer0_outputs(4278)) and not (layer0_outputs(9384));
    layer1_outputs(3455) <= not(layer0_outputs(2412)) or (layer0_outputs(9634));
    layer1_outputs(3456) <= not((layer0_outputs(9870)) or (layer0_outputs(1556)));
    layer1_outputs(3457) <= not(layer0_outputs(2682));
    layer1_outputs(3458) <= not(layer0_outputs(8157)) or (layer0_outputs(9621));
    layer1_outputs(3459) <= (layer0_outputs(7969)) and (layer0_outputs(1755));
    layer1_outputs(3460) <= (layer0_outputs(2444)) and not (layer0_outputs(6737));
    layer1_outputs(3461) <= not(layer0_outputs(5775));
    layer1_outputs(3462) <= not((layer0_outputs(5118)) or (layer0_outputs(3263)));
    layer1_outputs(3463) <= layer0_outputs(2059);
    layer1_outputs(3464) <= layer0_outputs(4450);
    layer1_outputs(3465) <= not(layer0_outputs(2732));
    layer1_outputs(3466) <= (layer0_outputs(1883)) and (layer0_outputs(69));
    layer1_outputs(3467) <= layer0_outputs(9576);
    layer1_outputs(3468) <= not(layer0_outputs(7839)) or (layer0_outputs(10175));
    layer1_outputs(3469) <= not(layer0_outputs(3286));
    layer1_outputs(3470) <= not(layer0_outputs(10139)) or (layer0_outputs(8634));
    layer1_outputs(3471) <= (layer0_outputs(4177)) and not (layer0_outputs(9422));
    layer1_outputs(3472) <= not((layer0_outputs(7222)) and (layer0_outputs(9396)));
    layer1_outputs(3473) <= not(layer0_outputs(5008));
    layer1_outputs(3474) <= not(layer0_outputs(6742));
    layer1_outputs(3475) <= not(layer0_outputs(1845)) or (layer0_outputs(1231));
    layer1_outputs(3476) <= not(layer0_outputs(6063));
    layer1_outputs(3477) <= not(layer0_outputs(10233)) or (layer0_outputs(6909));
    layer1_outputs(3478) <= (layer0_outputs(4424)) and not (layer0_outputs(4572));
    layer1_outputs(3479) <= not(layer0_outputs(10084)) or (layer0_outputs(3608));
    layer1_outputs(3480) <= not(layer0_outputs(8952)) or (layer0_outputs(6784));
    layer1_outputs(3481) <= '1';
    layer1_outputs(3482) <= (layer0_outputs(3722)) and not (layer0_outputs(5794));
    layer1_outputs(3483) <= not(layer0_outputs(1396));
    layer1_outputs(3484) <= not(layer0_outputs(3689)) or (layer0_outputs(9020));
    layer1_outputs(3485) <= not(layer0_outputs(8223));
    layer1_outputs(3486) <= '0';
    layer1_outputs(3487) <= (layer0_outputs(7168)) xor (layer0_outputs(3005));
    layer1_outputs(3488) <= not((layer0_outputs(9403)) xor (layer0_outputs(5672)));
    layer1_outputs(3489) <= (layer0_outputs(8030)) and (layer0_outputs(1094));
    layer1_outputs(3490) <= (layer0_outputs(5526)) and not (layer0_outputs(9256));
    layer1_outputs(3491) <= not((layer0_outputs(1506)) xor (layer0_outputs(8408)));
    layer1_outputs(3492) <= (layer0_outputs(7975)) or (layer0_outputs(5332));
    layer1_outputs(3493) <= (layer0_outputs(6080)) and (layer0_outputs(5476));
    layer1_outputs(3494) <= layer0_outputs(4287);
    layer1_outputs(3495) <= not(layer0_outputs(8458)) or (layer0_outputs(1133));
    layer1_outputs(3496) <= layer0_outputs(4556);
    layer1_outputs(3497) <= not((layer0_outputs(5388)) and (layer0_outputs(526)));
    layer1_outputs(3498) <= not((layer0_outputs(8415)) or (layer0_outputs(8352)));
    layer1_outputs(3499) <= not(layer0_outputs(9895));
    layer1_outputs(3500) <= not((layer0_outputs(7946)) or (layer0_outputs(4260)));
    layer1_outputs(3501) <= not(layer0_outputs(5266));
    layer1_outputs(3502) <= layer0_outputs(5351);
    layer1_outputs(3503) <= not(layer0_outputs(8210));
    layer1_outputs(3504) <= layer0_outputs(6439);
    layer1_outputs(3505) <= not(layer0_outputs(9279)) or (layer0_outputs(8994));
    layer1_outputs(3506) <= layer0_outputs(2107);
    layer1_outputs(3507) <= not(layer0_outputs(3939));
    layer1_outputs(3508) <= not(layer0_outputs(5939));
    layer1_outputs(3509) <= layer0_outputs(8001);
    layer1_outputs(3510) <= (layer0_outputs(3736)) xor (layer0_outputs(203));
    layer1_outputs(3511) <= not(layer0_outputs(5747));
    layer1_outputs(3512) <= (layer0_outputs(10164)) and not (layer0_outputs(2804));
    layer1_outputs(3513) <= (layer0_outputs(10200)) and (layer0_outputs(1816));
    layer1_outputs(3514) <= layer0_outputs(132);
    layer1_outputs(3515) <= not((layer0_outputs(9064)) and (layer0_outputs(4267)));
    layer1_outputs(3516) <= (layer0_outputs(9592)) and not (layer0_outputs(6435));
    layer1_outputs(3517) <= not((layer0_outputs(4871)) and (layer0_outputs(1699)));
    layer1_outputs(3518) <= layer0_outputs(10071);
    layer1_outputs(3519) <= not(layer0_outputs(2092)) or (layer0_outputs(6577));
    layer1_outputs(3520) <= not((layer0_outputs(4956)) or (layer0_outputs(8567)));
    layer1_outputs(3521) <= (layer0_outputs(3876)) and (layer0_outputs(3545));
    layer1_outputs(3522) <= not(layer0_outputs(9687));
    layer1_outputs(3523) <= not(layer0_outputs(3821));
    layer1_outputs(3524) <= layer0_outputs(8977);
    layer1_outputs(3525) <= layer0_outputs(8698);
    layer1_outputs(3526) <= (layer0_outputs(366)) and not (layer0_outputs(8409));
    layer1_outputs(3527) <= not(layer0_outputs(6957));
    layer1_outputs(3528) <= (layer0_outputs(2076)) and not (layer0_outputs(2454));
    layer1_outputs(3529) <= not(layer0_outputs(5567)) or (layer0_outputs(3537));
    layer1_outputs(3530) <= (layer0_outputs(2797)) and not (layer0_outputs(6633));
    layer1_outputs(3531) <= layer0_outputs(6558);
    layer1_outputs(3532) <= layer0_outputs(2577);
    layer1_outputs(3533) <= layer0_outputs(5832);
    layer1_outputs(3534) <= (layer0_outputs(5919)) or (layer0_outputs(2236));
    layer1_outputs(3535) <= (layer0_outputs(3199)) and not (layer0_outputs(548));
    layer1_outputs(3536) <= not((layer0_outputs(8208)) and (layer0_outputs(2936)));
    layer1_outputs(3537) <= not(layer0_outputs(3993));
    layer1_outputs(3538) <= layer0_outputs(5480);
    layer1_outputs(3539) <= not(layer0_outputs(2852));
    layer1_outputs(3540) <= not((layer0_outputs(6756)) or (layer0_outputs(9802)));
    layer1_outputs(3541) <= not(layer0_outputs(2669));
    layer1_outputs(3542) <= not(layer0_outputs(4337));
    layer1_outputs(3543) <= '1';
    layer1_outputs(3544) <= layer0_outputs(1318);
    layer1_outputs(3545) <= layer0_outputs(6599);
    layer1_outputs(3546) <= not((layer0_outputs(4854)) xor (layer0_outputs(9649)));
    layer1_outputs(3547) <= (layer0_outputs(544)) and not (layer0_outputs(681));
    layer1_outputs(3548) <= layer0_outputs(8838);
    layer1_outputs(3549) <= not((layer0_outputs(5969)) xor (layer0_outputs(365)));
    layer1_outputs(3550) <= layer0_outputs(4855);
    layer1_outputs(3551) <= not(layer0_outputs(6129));
    layer1_outputs(3552) <= (layer0_outputs(1044)) and (layer0_outputs(1255));
    layer1_outputs(3553) <= (layer0_outputs(9624)) xor (layer0_outputs(6717));
    layer1_outputs(3554) <= (layer0_outputs(9770)) and (layer0_outputs(6294));
    layer1_outputs(3555) <= not(layer0_outputs(8021));
    layer1_outputs(3556) <= not((layer0_outputs(7611)) and (layer0_outputs(4802)));
    layer1_outputs(3557) <= layer0_outputs(7101);
    layer1_outputs(3558) <= not(layer0_outputs(7144));
    layer1_outputs(3559) <= (layer0_outputs(9225)) or (layer0_outputs(3502));
    layer1_outputs(3560) <= not(layer0_outputs(5668));
    layer1_outputs(3561) <= not((layer0_outputs(9093)) or (layer0_outputs(6288)));
    layer1_outputs(3562) <= not(layer0_outputs(5122));
    layer1_outputs(3563) <= layer0_outputs(3738);
    layer1_outputs(3564) <= not(layer0_outputs(8761));
    layer1_outputs(3565) <= (layer0_outputs(7522)) and not (layer0_outputs(7808));
    layer1_outputs(3566) <= not((layer0_outputs(8135)) or (layer0_outputs(3378)));
    layer1_outputs(3567) <= (layer0_outputs(9356)) xor (layer0_outputs(1497));
    layer1_outputs(3568) <= (layer0_outputs(1078)) and not (layer0_outputs(5814));
    layer1_outputs(3569) <= not((layer0_outputs(4244)) or (layer0_outputs(3922)));
    layer1_outputs(3570) <= layer0_outputs(820);
    layer1_outputs(3571) <= not(layer0_outputs(4518)) or (layer0_outputs(9456));
    layer1_outputs(3572) <= layer0_outputs(9285);
    layer1_outputs(3573) <= layer0_outputs(6688);
    layer1_outputs(3574) <= not(layer0_outputs(5249)) or (layer0_outputs(4038));
    layer1_outputs(3575) <= '1';
    layer1_outputs(3576) <= (layer0_outputs(9758)) and (layer0_outputs(3935));
    layer1_outputs(3577) <= not(layer0_outputs(7440)) or (layer0_outputs(2533));
    layer1_outputs(3578) <= layer0_outputs(3403);
    layer1_outputs(3579) <= not(layer0_outputs(1168));
    layer1_outputs(3580) <= (layer0_outputs(713)) and (layer0_outputs(2385));
    layer1_outputs(3581) <= not(layer0_outputs(3316));
    layer1_outputs(3582) <= not(layer0_outputs(6854));
    layer1_outputs(3583) <= not((layer0_outputs(7433)) xor (layer0_outputs(9793)));
    layer1_outputs(3584) <= layer0_outputs(3095);
    layer1_outputs(3585) <= layer0_outputs(9980);
    layer1_outputs(3586) <= layer0_outputs(9658);
    layer1_outputs(3587) <= not((layer0_outputs(8025)) xor (layer0_outputs(45)));
    layer1_outputs(3588) <= not((layer0_outputs(1337)) or (layer0_outputs(819)));
    layer1_outputs(3589) <= layer0_outputs(242);
    layer1_outputs(3590) <= (layer0_outputs(474)) xor (layer0_outputs(3278));
    layer1_outputs(3591) <= layer0_outputs(4150);
    layer1_outputs(3592) <= layer0_outputs(8504);
    layer1_outputs(3593) <= not((layer0_outputs(8675)) xor (layer0_outputs(74)));
    layer1_outputs(3594) <= layer0_outputs(7652);
    layer1_outputs(3595) <= not(layer0_outputs(4631));
    layer1_outputs(3596) <= not(layer0_outputs(3585));
    layer1_outputs(3597) <= (layer0_outputs(1778)) and not (layer0_outputs(5513));
    layer1_outputs(3598) <= layer0_outputs(3820);
    layer1_outputs(3599) <= (layer0_outputs(3824)) and (layer0_outputs(1675));
    layer1_outputs(3600) <= not(layer0_outputs(7156));
    layer1_outputs(3601) <= not((layer0_outputs(5827)) or (layer0_outputs(7017)));
    layer1_outputs(3602) <= not(layer0_outputs(8295)) or (layer0_outputs(6408));
    layer1_outputs(3603) <= (layer0_outputs(8660)) and not (layer0_outputs(5824));
    layer1_outputs(3604) <= not((layer0_outputs(3911)) and (layer0_outputs(5391)));
    layer1_outputs(3605) <= (layer0_outputs(9827)) xor (layer0_outputs(9753));
    layer1_outputs(3606) <= layer0_outputs(1296);
    layer1_outputs(3607) <= not(layer0_outputs(8215));
    layer1_outputs(3608) <= not((layer0_outputs(467)) xor (layer0_outputs(7809)));
    layer1_outputs(3609) <= layer0_outputs(8898);
    layer1_outputs(3610) <= layer0_outputs(8273);
    layer1_outputs(3611) <= not((layer0_outputs(1504)) or (layer0_outputs(8438)));
    layer1_outputs(3612) <= not(layer0_outputs(6768));
    layer1_outputs(3613) <= (layer0_outputs(568)) or (layer0_outputs(2121));
    layer1_outputs(3614) <= not(layer0_outputs(3169)) or (layer0_outputs(4340));
    layer1_outputs(3615) <= (layer0_outputs(4675)) and (layer0_outputs(895));
    layer1_outputs(3616) <= not(layer0_outputs(81));
    layer1_outputs(3617) <= layer0_outputs(2385);
    layer1_outputs(3618) <= (layer0_outputs(2660)) and not (layer0_outputs(797));
    layer1_outputs(3619) <= '0';
    layer1_outputs(3620) <= not(layer0_outputs(9530));
    layer1_outputs(3621) <= not((layer0_outputs(489)) and (layer0_outputs(6494)));
    layer1_outputs(3622) <= not(layer0_outputs(5315));
    layer1_outputs(3623) <= (layer0_outputs(9625)) and not (layer0_outputs(7140));
    layer1_outputs(3624) <= (layer0_outputs(9765)) and not (layer0_outputs(2458));
    layer1_outputs(3625) <= not(layer0_outputs(3797));
    layer1_outputs(3626) <= '1';
    layer1_outputs(3627) <= not(layer0_outputs(6231));
    layer1_outputs(3628) <= not(layer0_outputs(1595));
    layer1_outputs(3629) <= not(layer0_outputs(3062));
    layer1_outputs(3630) <= not((layer0_outputs(3708)) and (layer0_outputs(9421)));
    layer1_outputs(3631) <= '1';
    layer1_outputs(3632) <= not(layer0_outputs(9485));
    layer1_outputs(3633) <= (layer0_outputs(8880)) or (layer0_outputs(3518));
    layer1_outputs(3634) <= (layer0_outputs(9310)) and (layer0_outputs(6107));
    layer1_outputs(3635) <= not(layer0_outputs(9613));
    layer1_outputs(3636) <= not(layer0_outputs(5025));
    layer1_outputs(3637) <= not((layer0_outputs(3563)) and (layer0_outputs(7649)));
    layer1_outputs(3638) <= layer0_outputs(5305);
    layer1_outputs(3639) <= layer0_outputs(605);
    layer1_outputs(3640) <= not((layer0_outputs(759)) and (layer0_outputs(4257)));
    layer1_outputs(3641) <= layer0_outputs(4109);
    layer1_outputs(3642) <= '0';
    layer1_outputs(3643) <= layer0_outputs(9010);
    layer1_outputs(3644) <= (layer0_outputs(1645)) and (layer0_outputs(1925));
    layer1_outputs(3645) <= (layer0_outputs(866)) xor (layer0_outputs(9917));
    layer1_outputs(3646) <= not(layer0_outputs(3175));
    layer1_outputs(3647) <= not(layer0_outputs(8886)) or (layer0_outputs(3305));
    layer1_outputs(3648) <= not(layer0_outputs(8095));
    layer1_outputs(3649) <= layer0_outputs(4935);
    layer1_outputs(3650) <= '1';
    layer1_outputs(3651) <= not(layer0_outputs(8336)) or (layer0_outputs(8414));
    layer1_outputs(3652) <= not((layer0_outputs(1357)) or (layer0_outputs(2531)));
    layer1_outputs(3653) <= layer0_outputs(4263);
    layer1_outputs(3654) <= (layer0_outputs(10122)) and not (layer0_outputs(6983));
    layer1_outputs(3655) <= (layer0_outputs(5817)) or (layer0_outputs(6329));
    layer1_outputs(3656) <= not(layer0_outputs(6538));
    layer1_outputs(3657) <= layer0_outputs(688);
    layer1_outputs(3658) <= not((layer0_outputs(127)) and (layer0_outputs(6950)));
    layer1_outputs(3659) <= not((layer0_outputs(7102)) and (layer0_outputs(1793)));
    layer1_outputs(3660) <= not((layer0_outputs(6884)) or (layer0_outputs(4430)));
    layer1_outputs(3661) <= layer0_outputs(6028);
    layer1_outputs(3662) <= (layer0_outputs(5661)) and not (layer0_outputs(6608));
    layer1_outputs(3663) <= not(layer0_outputs(4682));
    layer1_outputs(3664) <= not(layer0_outputs(4799)) or (layer0_outputs(4783));
    layer1_outputs(3665) <= not(layer0_outputs(5169));
    layer1_outputs(3666) <= (layer0_outputs(1520)) and not (layer0_outputs(8090));
    layer1_outputs(3667) <= not(layer0_outputs(2750)) or (layer0_outputs(4843));
    layer1_outputs(3668) <= (layer0_outputs(3035)) and not (layer0_outputs(1618));
    layer1_outputs(3669) <= (layer0_outputs(5728)) and not (layer0_outputs(7683));
    layer1_outputs(3670) <= not((layer0_outputs(5631)) and (layer0_outputs(4217)));
    layer1_outputs(3671) <= '0';
    layer1_outputs(3672) <= (layer0_outputs(7063)) and not (layer0_outputs(2067));
    layer1_outputs(3673) <= layer0_outputs(1830);
    layer1_outputs(3674) <= not((layer0_outputs(4419)) or (layer0_outputs(3572)));
    layer1_outputs(3675) <= layer0_outputs(4189);
    layer1_outputs(3676) <= layer0_outputs(1838);
    layer1_outputs(3677) <= layer0_outputs(6544);
    layer1_outputs(3678) <= (layer0_outputs(1352)) and not (layer0_outputs(6068));
    layer1_outputs(3679) <= layer0_outputs(8090);
    layer1_outputs(3680) <= not((layer0_outputs(4056)) or (layer0_outputs(2471)));
    layer1_outputs(3681) <= layer0_outputs(1781);
    layer1_outputs(3682) <= layer0_outputs(1143);
    layer1_outputs(3683) <= '1';
    layer1_outputs(3684) <= not((layer0_outputs(8824)) or (layer0_outputs(4743)));
    layer1_outputs(3685) <= (layer0_outputs(5071)) or (layer0_outputs(4207));
    layer1_outputs(3686) <= not((layer0_outputs(8822)) or (layer0_outputs(1352)));
    layer1_outputs(3687) <= not(layer0_outputs(7892));
    layer1_outputs(3688) <= (layer0_outputs(5329)) or (layer0_outputs(5280));
    layer1_outputs(3689) <= '0';
    layer1_outputs(3690) <= not(layer0_outputs(4718)) or (layer0_outputs(8803));
    layer1_outputs(3691) <= (layer0_outputs(5330)) and (layer0_outputs(7942));
    layer1_outputs(3692) <= not(layer0_outputs(5314));
    layer1_outputs(3693) <= not(layer0_outputs(44)) or (layer0_outputs(6398));
    layer1_outputs(3694) <= (layer0_outputs(5533)) and not (layer0_outputs(9973));
    layer1_outputs(3695) <= not(layer0_outputs(5076)) or (layer0_outputs(7592));
    layer1_outputs(3696) <= (layer0_outputs(8387)) or (layer0_outputs(2583));
    layer1_outputs(3697) <= layer0_outputs(6894);
    layer1_outputs(3698) <= '1';
    layer1_outputs(3699) <= not((layer0_outputs(5192)) and (layer0_outputs(7667)));
    layer1_outputs(3700) <= (layer0_outputs(6012)) or (layer0_outputs(6624));
    layer1_outputs(3701) <= not(layer0_outputs(2503));
    layer1_outputs(3702) <= layer0_outputs(5527);
    layer1_outputs(3703) <= not((layer0_outputs(2078)) or (layer0_outputs(1671)));
    layer1_outputs(3704) <= not((layer0_outputs(9798)) and (layer0_outputs(1593)));
    layer1_outputs(3705) <= not(layer0_outputs(4774));
    layer1_outputs(3706) <= not(layer0_outputs(6271));
    layer1_outputs(3707) <= layer0_outputs(8377);
    layer1_outputs(3708) <= layer0_outputs(7042);
    layer1_outputs(3709) <= (layer0_outputs(9690)) and not (layer0_outputs(6843));
    layer1_outputs(3710) <= (layer0_outputs(791)) and not (layer0_outputs(312));
    layer1_outputs(3711) <= layer0_outputs(952);
    layer1_outputs(3712) <= layer0_outputs(6205);
    layer1_outputs(3713) <= not((layer0_outputs(2683)) and (layer0_outputs(6221)));
    layer1_outputs(3714) <= layer0_outputs(3561);
    layer1_outputs(3715) <= not(layer0_outputs(3603));
    layer1_outputs(3716) <= (layer0_outputs(5494)) xor (layer0_outputs(5203));
    layer1_outputs(3717) <= layer0_outputs(6374);
    layer1_outputs(3718) <= layer0_outputs(4931);
    layer1_outputs(3719) <= '1';
    layer1_outputs(3720) <= not((layer0_outputs(7196)) or (layer0_outputs(9633)));
    layer1_outputs(3721) <= layer0_outputs(3075);
    layer1_outputs(3722) <= not((layer0_outputs(7227)) xor (layer0_outputs(1484)));
    layer1_outputs(3723) <= layer0_outputs(7331);
    layer1_outputs(3724) <= not(layer0_outputs(8799));
    layer1_outputs(3725) <= (layer0_outputs(5295)) or (layer0_outputs(3499));
    layer1_outputs(3726) <= '0';
    layer1_outputs(3727) <= not(layer0_outputs(2733));
    layer1_outputs(3728) <= not(layer0_outputs(1877));
    layer1_outputs(3729) <= not((layer0_outputs(8118)) or (layer0_outputs(2094)));
    layer1_outputs(3730) <= layer0_outputs(9140);
    layer1_outputs(3731) <= layer0_outputs(9664);
    layer1_outputs(3732) <= '1';
    layer1_outputs(3733) <= '1';
    layer1_outputs(3734) <= not(layer0_outputs(721));
    layer1_outputs(3735) <= not(layer0_outputs(77)) or (layer0_outputs(4412));
    layer1_outputs(3736) <= not(layer0_outputs(8692)) or (layer0_outputs(9064));
    layer1_outputs(3737) <= not(layer0_outputs(6752)) or (layer0_outputs(5585));
    layer1_outputs(3738) <= not(layer0_outputs(8939)) or (layer0_outputs(3394));
    layer1_outputs(3739) <= layer0_outputs(2850);
    layer1_outputs(3740) <= (layer0_outputs(3337)) and not (layer0_outputs(7744));
    layer1_outputs(3741) <= (layer0_outputs(9178)) and (layer0_outputs(6352));
    layer1_outputs(3742) <= layer0_outputs(167);
    layer1_outputs(3743) <= layer0_outputs(4112);
    layer1_outputs(3744) <= not(layer0_outputs(9901)) or (layer0_outputs(2805));
    layer1_outputs(3745) <= (layer0_outputs(3806)) xor (layer0_outputs(3164));
    layer1_outputs(3746) <= not(layer0_outputs(143));
    layer1_outputs(3747) <= (layer0_outputs(4405)) xor (layer0_outputs(722));
    layer1_outputs(3748) <= layer0_outputs(10043);
    layer1_outputs(3749) <= not(layer0_outputs(5018));
    layer1_outputs(3750) <= (layer0_outputs(9994)) xor (layer0_outputs(8030));
    layer1_outputs(3751) <= not(layer0_outputs(8712)) or (layer0_outputs(4337));
    layer1_outputs(3752) <= (layer0_outputs(9649)) and not (layer0_outputs(4840));
    layer1_outputs(3753) <= not(layer0_outputs(2308)) or (layer0_outputs(9574));
    layer1_outputs(3754) <= (layer0_outputs(9535)) and not (layer0_outputs(5443));
    layer1_outputs(3755) <= '1';
    layer1_outputs(3756) <= not(layer0_outputs(9597));
    layer1_outputs(3757) <= (layer0_outputs(5564)) xor (layer0_outputs(8900));
    layer1_outputs(3758) <= layer0_outputs(5932);
    layer1_outputs(3759) <= not(layer0_outputs(2306));
    layer1_outputs(3760) <= (layer0_outputs(1998)) and (layer0_outputs(350));
    layer1_outputs(3761) <= (layer0_outputs(431)) and not (layer0_outputs(8223));
    layer1_outputs(3762) <= layer0_outputs(7737);
    layer1_outputs(3763) <= not(layer0_outputs(8995));
    layer1_outputs(3764) <= not((layer0_outputs(8496)) xor (layer0_outputs(1486)));
    layer1_outputs(3765) <= layer0_outputs(3201);
    layer1_outputs(3766) <= not((layer0_outputs(4499)) xor (layer0_outputs(4996)));
    layer1_outputs(3767) <= not(layer0_outputs(7253));
    layer1_outputs(3768) <= (layer0_outputs(4553)) and not (layer0_outputs(9961));
    layer1_outputs(3769) <= (layer0_outputs(9084)) or (layer0_outputs(6469));
    layer1_outputs(3770) <= layer0_outputs(8150);
    layer1_outputs(3771) <= layer0_outputs(7308);
    layer1_outputs(3772) <= layer0_outputs(2231);
    layer1_outputs(3773) <= (layer0_outputs(6816)) and (layer0_outputs(7596));
    layer1_outputs(3774) <= not((layer0_outputs(6933)) xor (layer0_outputs(9644)));
    layer1_outputs(3775) <= (layer0_outputs(3371)) or (layer0_outputs(10129));
    layer1_outputs(3776) <= (layer0_outputs(1611)) and not (layer0_outputs(7304));
    layer1_outputs(3777) <= layer0_outputs(9291);
    layer1_outputs(3778) <= layer0_outputs(1931);
    layer1_outputs(3779) <= layer0_outputs(759);
    layer1_outputs(3780) <= not(layer0_outputs(6496));
    layer1_outputs(3781) <= not((layer0_outputs(446)) or (layer0_outputs(9503)));
    layer1_outputs(3782) <= layer0_outputs(4771);
    layer1_outputs(3783) <= not(layer0_outputs(4068));
    layer1_outputs(3784) <= not(layer0_outputs(712));
    layer1_outputs(3785) <= layer0_outputs(7893);
    layer1_outputs(3786) <= layer0_outputs(9201);
    layer1_outputs(3787) <= (layer0_outputs(9096)) or (layer0_outputs(9626));
    layer1_outputs(3788) <= layer0_outputs(5932);
    layer1_outputs(3789) <= not((layer0_outputs(2375)) xor (layer0_outputs(1217)));
    layer1_outputs(3790) <= '0';
    layer1_outputs(3791) <= not(layer0_outputs(3369));
    layer1_outputs(3792) <= not((layer0_outputs(7730)) or (layer0_outputs(5952)));
    layer1_outputs(3793) <= (layer0_outputs(8614)) and (layer0_outputs(3769));
    layer1_outputs(3794) <= (layer0_outputs(3787)) and (layer0_outputs(1137));
    layer1_outputs(3795) <= (layer0_outputs(3139)) xor (layer0_outputs(3452));
    layer1_outputs(3796) <= layer0_outputs(5294);
    layer1_outputs(3797) <= (layer0_outputs(9604)) xor (layer0_outputs(174));
    layer1_outputs(3798) <= not(layer0_outputs(479)) or (layer0_outputs(1199));
    layer1_outputs(3799) <= not(layer0_outputs(5432));
    layer1_outputs(3800) <= not(layer0_outputs(5016)) or (layer0_outputs(6585));
    layer1_outputs(3801) <= (layer0_outputs(7746)) and not (layer0_outputs(6362));
    layer1_outputs(3802) <= layer0_outputs(1644);
    layer1_outputs(3803) <= layer0_outputs(2666);
    layer1_outputs(3804) <= (layer0_outputs(2488)) and not (layer0_outputs(10202));
    layer1_outputs(3805) <= not(layer0_outputs(2088));
    layer1_outputs(3806) <= layer0_outputs(1509);
    layer1_outputs(3807) <= '0';
    layer1_outputs(3808) <= not(layer0_outputs(6240)) or (layer0_outputs(7445));
    layer1_outputs(3809) <= layer0_outputs(7465);
    layer1_outputs(3810) <= layer0_outputs(6301);
    layer1_outputs(3811) <= layer0_outputs(2481);
    layer1_outputs(3812) <= not(layer0_outputs(4678));
    layer1_outputs(3813) <= (layer0_outputs(9257)) and not (layer0_outputs(4187));
    layer1_outputs(3814) <= layer0_outputs(5047);
    layer1_outputs(3815) <= not(layer0_outputs(7776));
    layer1_outputs(3816) <= not(layer0_outputs(7269));
    layer1_outputs(3817) <= (layer0_outputs(8598)) and (layer0_outputs(9743));
    layer1_outputs(3818) <= not(layer0_outputs(10134));
    layer1_outputs(3819) <= layer0_outputs(5008);
    layer1_outputs(3820) <= not(layer0_outputs(9946));
    layer1_outputs(3821) <= not(layer0_outputs(1970));
    layer1_outputs(3822) <= not(layer0_outputs(1283)) or (layer0_outputs(6698));
    layer1_outputs(3823) <= (layer0_outputs(7683)) or (layer0_outputs(5415));
    layer1_outputs(3824) <= '0';
    layer1_outputs(3825) <= layer0_outputs(9023);
    layer1_outputs(3826) <= not(layer0_outputs(59));
    layer1_outputs(3827) <= not(layer0_outputs(2948)) or (layer0_outputs(9136));
    layer1_outputs(3828) <= not(layer0_outputs(6658));
    layer1_outputs(3829) <= (layer0_outputs(4893)) and not (layer0_outputs(1152));
    layer1_outputs(3830) <= layer0_outputs(3861);
    layer1_outputs(3831) <= (layer0_outputs(2101)) and not (layer0_outputs(643));
    layer1_outputs(3832) <= not(layer0_outputs(1156));
    layer1_outputs(3833) <= (layer0_outputs(8674)) and not (layer0_outputs(5549));
    layer1_outputs(3834) <= not(layer0_outputs(6456));
    layer1_outputs(3835) <= not(layer0_outputs(8199));
    layer1_outputs(3836) <= not(layer0_outputs(6509));
    layer1_outputs(3837) <= not(layer0_outputs(2718));
    layer1_outputs(3838) <= (layer0_outputs(9361)) and not (layer0_outputs(6307));
    layer1_outputs(3839) <= (layer0_outputs(9250)) xor (layer0_outputs(2818));
    layer1_outputs(3840) <= (layer0_outputs(7905)) xor (layer0_outputs(6146));
    layer1_outputs(3841) <= not(layer0_outputs(5708));
    layer1_outputs(3842) <= layer0_outputs(973);
    layer1_outputs(3843) <= not((layer0_outputs(6835)) xor (layer0_outputs(1450)));
    layer1_outputs(3844) <= not(layer0_outputs(4124));
    layer1_outputs(3845) <= layer0_outputs(1002);
    layer1_outputs(3846) <= not((layer0_outputs(4257)) and (layer0_outputs(5352)));
    layer1_outputs(3847) <= not((layer0_outputs(9813)) and (layer0_outputs(3237)));
    layer1_outputs(3848) <= (layer0_outputs(7638)) or (layer0_outputs(7978));
    layer1_outputs(3849) <= (layer0_outputs(4305)) and (layer0_outputs(6215));
    layer1_outputs(3850) <= '1';
    layer1_outputs(3851) <= not(layer0_outputs(2214)) or (layer0_outputs(7438));
    layer1_outputs(3852) <= layer0_outputs(2680);
    layer1_outputs(3853) <= (layer0_outputs(3261)) or (layer0_outputs(665));
    layer1_outputs(3854) <= layer0_outputs(340);
    layer1_outputs(3855) <= layer0_outputs(5832);
    layer1_outputs(3856) <= layer0_outputs(2658);
    layer1_outputs(3857) <= not(layer0_outputs(4909));
    layer1_outputs(3858) <= not(layer0_outputs(6303));
    layer1_outputs(3859) <= layer0_outputs(7705);
    layer1_outputs(3860) <= not(layer0_outputs(7325));
    layer1_outputs(3861) <= layer0_outputs(2888);
    layer1_outputs(3862) <= layer0_outputs(9677);
    layer1_outputs(3863) <= (layer0_outputs(5120)) xor (layer0_outputs(8971));
    layer1_outputs(3864) <= not((layer0_outputs(2569)) and (layer0_outputs(9097)));
    layer1_outputs(3865) <= not(layer0_outputs(8547)) or (layer0_outputs(1946));
    layer1_outputs(3866) <= layer0_outputs(6404);
    layer1_outputs(3867) <= layer0_outputs(7844);
    layer1_outputs(3868) <= not(layer0_outputs(5020)) or (layer0_outputs(2821));
    layer1_outputs(3869) <= (layer0_outputs(9455)) or (layer0_outputs(5408));
    layer1_outputs(3870) <= '1';
    layer1_outputs(3871) <= not(layer0_outputs(6033));
    layer1_outputs(3872) <= layer0_outputs(5042);
    layer1_outputs(3873) <= '0';
    layer1_outputs(3874) <= layer0_outputs(5735);
    layer1_outputs(3875) <= not((layer0_outputs(10155)) xor (layer0_outputs(4328)));
    layer1_outputs(3876) <= (layer0_outputs(7923)) or (layer0_outputs(1468));
    layer1_outputs(3877) <= not((layer0_outputs(4945)) and (layer0_outputs(5188)));
    layer1_outputs(3878) <= layer0_outputs(6622);
    layer1_outputs(3879) <= (layer0_outputs(8307)) and not (layer0_outputs(3663));
    layer1_outputs(3880) <= not((layer0_outputs(2930)) or (layer0_outputs(2870)));
    layer1_outputs(3881) <= not(layer0_outputs(2030)) or (layer0_outputs(7753));
    layer1_outputs(3882) <= not(layer0_outputs(4183));
    layer1_outputs(3883) <= (layer0_outputs(6632)) or (layer0_outputs(3409));
    layer1_outputs(3884) <= (layer0_outputs(2096)) or (layer0_outputs(7945));
    layer1_outputs(3885) <= (layer0_outputs(7645)) and (layer0_outputs(9736));
    layer1_outputs(3886) <= not((layer0_outputs(8957)) and (layer0_outputs(7716)));
    layer1_outputs(3887) <= layer0_outputs(8430);
    layer1_outputs(3888) <= not(layer0_outputs(7043));
    layer1_outputs(3889) <= not(layer0_outputs(5764)) or (layer0_outputs(7671));
    layer1_outputs(3890) <= (layer0_outputs(8508)) and not (layer0_outputs(121));
    layer1_outputs(3891) <= not(layer0_outputs(4395));
    layer1_outputs(3892) <= layer0_outputs(9982);
    layer1_outputs(3893) <= (layer0_outputs(10041)) and not (layer0_outputs(3207));
    layer1_outputs(3894) <= not((layer0_outputs(3690)) or (layer0_outputs(10021)));
    layer1_outputs(3895) <= (layer0_outputs(1923)) and not (layer0_outputs(6540));
    layer1_outputs(3896) <= (layer0_outputs(7387)) and (layer0_outputs(2785));
    layer1_outputs(3897) <= not(layer0_outputs(6395));
    layer1_outputs(3898) <= (layer0_outputs(7425)) and not (layer0_outputs(8920));
    layer1_outputs(3899) <= (layer0_outputs(165)) or (layer0_outputs(6223));
    layer1_outputs(3900) <= (layer0_outputs(6867)) and (layer0_outputs(8705));
    layer1_outputs(3901) <= '1';
    layer1_outputs(3902) <= not(layer0_outputs(1961));
    layer1_outputs(3903) <= not(layer0_outputs(9350)) or (layer0_outputs(8136));
    layer1_outputs(3904) <= (layer0_outputs(2497)) and not (layer0_outputs(1006));
    layer1_outputs(3905) <= (layer0_outputs(1153)) and (layer0_outputs(5313));
    layer1_outputs(3906) <= (layer0_outputs(2989)) and (layer0_outputs(7594));
    layer1_outputs(3907) <= (layer0_outputs(9641)) or (layer0_outputs(935));
    layer1_outputs(3908) <= layer0_outputs(450);
    layer1_outputs(3909) <= layer0_outputs(3426);
    layer1_outputs(3910) <= (layer0_outputs(9839)) or (layer0_outputs(2361));
    layer1_outputs(3911) <= not(layer0_outputs(1025));
    layer1_outputs(3912) <= layer0_outputs(4835);
    layer1_outputs(3913) <= (layer0_outputs(7248)) or (layer0_outputs(9115));
    layer1_outputs(3914) <= (layer0_outputs(2231)) or (layer0_outputs(8883));
    layer1_outputs(3915) <= (layer0_outputs(8158)) or (layer0_outputs(6936));
    layer1_outputs(3916) <= (layer0_outputs(7091)) or (layer0_outputs(9047));
    layer1_outputs(3917) <= (layer0_outputs(5886)) or (layer0_outputs(8191));
    layer1_outputs(3918) <= not(layer0_outputs(3037));
    layer1_outputs(3919) <= not(layer0_outputs(5236));
    layer1_outputs(3920) <= not(layer0_outputs(3757)) or (layer0_outputs(7945));
    layer1_outputs(3921) <= (layer0_outputs(9952)) xor (layer0_outputs(2685));
    layer1_outputs(3922) <= (layer0_outputs(5159)) and not (layer0_outputs(6273));
    layer1_outputs(3923) <= layer0_outputs(3546);
    layer1_outputs(3924) <= (layer0_outputs(5877)) or (layer0_outputs(5433));
    layer1_outputs(3925) <= not(layer0_outputs(808));
    layer1_outputs(3926) <= not((layer0_outputs(9335)) or (layer0_outputs(9331)));
    layer1_outputs(3927) <= (layer0_outputs(1715)) and not (layer0_outputs(5406));
    layer1_outputs(3928) <= (layer0_outputs(6744)) or (layer0_outputs(1910));
    layer1_outputs(3929) <= not(layer0_outputs(2876));
    layer1_outputs(3930) <= layer0_outputs(6081);
    layer1_outputs(3931) <= layer0_outputs(2701);
    layer1_outputs(3932) <= layer0_outputs(419);
    layer1_outputs(3933) <= '1';
    layer1_outputs(3934) <= not((layer0_outputs(6030)) or (layer0_outputs(934)));
    layer1_outputs(3935) <= not(layer0_outputs(2955)) or (layer0_outputs(9689));
    layer1_outputs(3936) <= '0';
    layer1_outputs(3937) <= not((layer0_outputs(3422)) or (layer0_outputs(5021)));
    layer1_outputs(3938) <= not(layer0_outputs(6671)) or (layer0_outputs(7936));
    layer1_outputs(3939) <= not(layer0_outputs(5835)) or (layer0_outputs(6220));
    layer1_outputs(3940) <= layer0_outputs(8027);
    layer1_outputs(3941) <= layer0_outputs(1163);
    layer1_outputs(3942) <= (layer0_outputs(4839)) or (layer0_outputs(2338));
    layer1_outputs(3943) <= '1';
    layer1_outputs(3944) <= not(layer0_outputs(10138));
    layer1_outputs(3945) <= not((layer0_outputs(5599)) and (layer0_outputs(8354)));
    layer1_outputs(3946) <= layer0_outputs(5665);
    layer1_outputs(3947) <= not(layer0_outputs(4744));
    layer1_outputs(3948) <= not(layer0_outputs(9969));
    layer1_outputs(3949) <= '0';
    layer1_outputs(3950) <= not(layer0_outputs(9952));
    layer1_outputs(3951) <= layer0_outputs(462);
    layer1_outputs(3952) <= not((layer0_outputs(2922)) or (layer0_outputs(2988)));
    layer1_outputs(3953) <= (layer0_outputs(8390)) and not (layer0_outputs(5644));
    layer1_outputs(3954) <= not(layer0_outputs(9771));
    layer1_outputs(3955) <= not((layer0_outputs(8130)) or (layer0_outputs(2488)));
    layer1_outputs(3956) <= (layer0_outputs(2442)) xor (layer0_outputs(3008));
    layer1_outputs(3957) <= not((layer0_outputs(727)) and (layer0_outputs(3216)));
    layer1_outputs(3958) <= not(layer0_outputs(5890));
    layer1_outputs(3959) <= layer0_outputs(10138);
    layer1_outputs(3960) <= (layer0_outputs(8407)) and (layer0_outputs(7261));
    layer1_outputs(3961) <= not(layer0_outputs(7040));
    layer1_outputs(3962) <= not(layer0_outputs(3512)) or (layer0_outputs(7687));
    layer1_outputs(3963) <= not((layer0_outputs(8053)) or (layer0_outputs(6598)));
    layer1_outputs(3964) <= not(layer0_outputs(1181));
    layer1_outputs(3965) <= layer0_outputs(8829);
    layer1_outputs(3966) <= layer0_outputs(8846);
    layer1_outputs(3967) <= not(layer0_outputs(3900));
    layer1_outputs(3968) <= layer0_outputs(7150);
    layer1_outputs(3969) <= layer0_outputs(4603);
    layer1_outputs(3970) <= layer0_outputs(8159);
    layer1_outputs(3971) <= (layer0_outputs(8441)) and not (layer0_outputs(1750));
    layer1_outputs(3972) <= not(layer0_outputs(6318)) or (layer0_outputs(5157));
    layer1_outputs(3973) <= not(layer0_outputs(4832)) or (layer0_outputs(3664));
    layer1_outputs(3974) <= not(layer0_outputs(8132));
    layer1_outputs(3975) <= not((layer0_outputs(2383)) xor (layer0_outputs(2418)));
    layer1_outputs(3976) <= not(layer0_outputs(9144)) or (layer0_outputs(9032));
    layer1_outputs(3977) <= (layer0_outputs(1612)) or (layer0_outputs(2773));
    layer1_outputs(3978) <= '0';
    layer1_outputs(3979) <= not(layer0_outputs(8996));
    layer1_outputs(3980) <= (layer0_outputs(8648)) and (layer0_outputs(3527));
    layer1_outputs(3981) <= (layer0_outputs(3334)) and not (layer0_outputs(3831));
    layer1_outputs(3982) <= (layer0_outputs(6034)) and not (layer0_outputs(3772));
    layer1_outputs(3983) <= layer0_outputs(8834);
    layer1_outputs(3984) <= not(layer0_outputs(8700)) or (layer0_outputs(6225));
    layer1_outputs(3985) <= not(layer0_outputs(6844));
    layer1_outputs(3986) <= not(layer0_outputs(9405)) or (layer0_outputs(4820));
    layer1_outputs(3987) <= (layer0_outputs(8684)) and not (layer0_outputs(4259));
    layer1_outputs(3988) <= (layer0_outputs(2002)) and not (layer0_outputs(8039));
    layer1_outputs(3989) <= (layer0_outputs(2878)) and not (layer0_outputs(1134));
    layer1_outputs(3990) <= (layer0_outputs(253)) xor (layer0_outputs(35));
    layer1_outputs(3991) <= (layer0_outputs(5781)) or (layer0_outputs(8581));
    layer1_outputs(3992) <= (layer0_outputs(4048)) or (layer0_outputs(6350));
    layer1_outputs(3993) <= not(layer0_outputs(1292));
    layer1_outputs(3994) <= not((layer0_outputs(6762)) and (layer0_outputs(3672)));
    layer1_outputs(3995) <= not(layer0_outputs(6520)) or (layer0_outputs(2984));
    layer1_outputs(3996) <= layer0_outputs(10158);
    layer1_outputs(3997) <= (layer0_outputs(3048)) and not (layer0_outputs(319));
    layer1_outputs(3998) <= not(layer0_outputs(8359));
    layer1_outputs(3999) <= not(layer0_outputs(9888));
    layer1_outputs(4000) <= (layer0_outputs(7970)) and not (layer0_outputs(3646));
    layer1_outputs(4001) <= not(layer0_outputs(7492)) or (layer0_outputs(7981));
    layer1_outputs(4002) <= not(layer0_outputs(7686));
    layer1_outputs(4003) <= (layer0_outputs(4736)) and not (layer0_outputs(925));
    layer1_outputs(4004) <= not((layer0_outputs(4981)) and (layer0_outputs(9995)));
    layer1_outputs(4005) <= (layer0_outputs(6519)) or (layer0_outputs(9928));
    layer1_outputs(4006) <= not(layer0_outputs(4380));
    layer1_outputs(4007) <= (layer0_outputs(8728)) xor (layer0_outputs(1641));
    layer1_outputs(4008) <= not(layer0_outputs(2234));
    layer1_outputs(4009) <= not(layer0_outputs(4478)) or (layer0_outputs(8706));
    layer1_outputs(4010) <= (layer0_outputs(3198)) or (layer0_outputs(1656));
    layer1_outputs(4011) <= layer0_outputs(5992);
    layer1_outputs(4012) <= not((layer0_outputs(3934)) or (layer0_outputs(9889)));
    layer1_outputs(4013) <= (layer0_outputs(1833)) xor (layer0_outputs(5358));
    layer1_outputs(4014) <= not(layer0_outputs(8955));
    layer1_outputs(4015) <= '1';
    layer1_outputs(4016) <= not(layer0_outputs(7378));
    layer1_outputs(4017) <= layer0_outputs(5947);
    layer1_outputs(4018) <= (layer0_outputs(2957)) and not (layer0_outputs(1184));
    layer1_outputs(4019) <= not(layer0_outputs(7933)) or (layer0_outputs(1155));
    layer1_outputs(4020) <= (layer0_outputs(2455)) xor (layer0_outputs(668));
    layer1_outputs(4021) <= not(layer0_outputs(3299));
    layer1_outputs(4022) <= not(layer0_outputs(5228));
    layer1_outputs(4023) <= (layer0_outputs(7991)) and not (layer0_outputs(6577));
    layer1_outputs(4024) <= (layer0_outputs(4151)) and not (layer0_outputs(5680));
    layer1_outputs(4025) <= layer0_outputs(7392);
    layer1_outputs(4026) <= not((layer0_outputs(1372)) and (layer0_outputs(5152)));
    layer1_outputs(4027) <= not((layer0_outputs(8431)) and (layer0_outputs(4601)));
    layer1_outputs(4028) <= not(layer0_outputs(700)) or (layer0_outputs(10078));
    layer1_outputs(4029) <= not(layer0_outputs(37));
    layer1_outputs(4030) <= (layer0_outputs(3385)) and (layer0_outputs(9953));
    layer1_outputs(4031) <= layer0_outputs(4501);
    layer1_outputs(4032) <= layer0_outputs(8470);
    layer1_outputs(4033) <= not(layer0_outputs(17));
    layer1_outputs(4034) <= layer0_outputs(361);
    layer1_outputs(4035) <= (layer0_outputs(1678)) and not (layer0_outputs(3553));
    layer1_outputs(4036) <= layer0_outputs(253);
    layer1_outputs(4037) <= not(layer0_outputs(5413)) or (layer0_outputs(5679));
    layer1_outputs(4038) <= not(layer0_outputs(1134)) or (layer0_outputs(5479));
    layer1_outputs(4039) <= not(layer0_outputs(3035));
    layer1_outputs(4040) <= layer0_outputs(2197);
    layer1_outputs(4041) <= '0';
    layer1_outputs(4042) <= not((layer0_outputs(4242)) and (layer0_outputs(4429)));
    layer1_outputs(4043) <= layer0_outputs(4992);
    layer1_outputs(4044) <= (layer0_outputs(9892)) or (layer0_outputs(2301));
    layer1_outputs(4045) <= not(layer0_outputs(4792));
    layer1_outputs(4046) <= not(layer0_outputs(9748));
    layer1_outputs(4047) <= layer0_outputs(3647);
    layer1_outputs(4048) <= (layer0_outputs(9431)) and not (layer0_outputs(9734));
    layer1_outputs(4049) <= layer0_outputs(4338);
    layer1_outputs(4050) <= layer0_outputs(7207);
    layer1_outputs(4051) <= '1';
    layer1_outputs(4052) <= layer0_outputs(257);
    layer1_outputs(4053) <= not((layer0_outputs(2889)) and (layer0_outputs(2084)));
    layer1_outputs(4054) <= not(layer0_outputs(6872));
    layer1_outputs(4055) <= (layer0_outputs(10078)) and (layer0_outputs(2071));
    layer1_outputs(4056) <= layer0_outputs(912);
    layer1_outputs(4057) <= not(layer0_outputs(7069));
    layer1_outputs(4058) <= not(layer0_outputs(10228));
    layer1_outputs(4059) <= not(layer0_outputs(3346));
    layer1_outputs(4060) <= layer0_outputs(5145);
    layer1_outputs(4061) <= (layer0_outputs(6718)) and (layer0_outputs(3267));
    layer1_outputs(4062) <= (layer0_outputs(7441)) or (layer0_outputs(1854));
    layer1_outputs(4063) <= layer0_outputs(5943);
    layer1_outputs(4064) <= not((layer0_outputs(2058)) or (layer0_outputs(5370)));
    layer1_outputs(4065) <= '0';
    layer1_outputs(4066) <= not(layer0_outputs(8111));
    layer1_outputs(4067) <= not(layer0_outputs(2373));
    layer1_outputs(4068) <= (layer0_outputs(4733)) and not (layer0_outputs(4186));
    layer1_outputs(4069) <= (layer0_outputs(5938)) and not (layer0_outputs(1296));
    layer1_outputs(4070) <= not(layer0_outputs(7050));
    layer1_outputs(4071) <= not(layer0_outputs(283)) or (layer0_outputs(8325));
    layer1_outputs(4072) <= not(layer0_outputs(3542));
    layer1_outputs(4073) <= (layer0_outputs(8746)) xor (layer0_outputs(1372));
    layer1_outputs(4074) <= not((layer0_outputs(9173)) and (layer0_outputs(5220)));
    layer1_outputs(4075) <= (layer0_outputs(5819)) xor (layer0_outputs(3102));
    layer1_outputs(4076) <= not(layer0_outputs(3569));
    layer1_outputs(4077) <= '0';
    layer1_outputs(4078) <= not(layer0_outputs(4104)) or (layer0_outputs(9560));
    layer1_outputs(4079) <= layer0_outputs(1341);
    layer1_outputs(4080) <= (layer0_outputs(8932)) or (layer0_outputs(9334));
    layer1_outputs(4081) <= not((layer0_outputs(3564)) or (layer0_outputs(7120)));
    layer1_outputs(4082) <= (layer0_outputs(2615)) and not (layer0_outputs(8374));
    layer1_outputs(4083) <= layer0_outputs(2466);
    layer1_outputs(4084) <= not((layer0_outputs(4834)) and (layer0_outputs(5666)));
    layer1_outputs(4085) <= not((layer0_outputs(8585)) and (layer0_outputs(898)));
    layer1_outputs(4086) <= layer0_outputs(2687);
    layer1_outputs(4087) <= layer0_outputs(5061);
    layer1_outputs(4088) <= (layer0_outputs(6663)) xor (layer0_outputs(4727));
    layer1_outputs(4089) <= not((layer0_outputs(9332)) or (layer0_outputs(5344)));
    layer1_outputs(4090) <= (layer0_outputs(3107)) and not (layer0_outputs(5807));
    layer1_outputs(4091) <= (layer0_outputs(6810)) and (layer0_outputs(4288));
    layer1_outputs(4092) <= (layer0_outputs(4359)) and not (layer0_outputs(3480));
    layer1_outputs(4093) <= not(layer0_outputs(6621)) or (layer0_outputs(4064));
    layer1_outputs(4094) <= not(layer0_outputs(4542));
    layer1_outputs(4095) <= not(layer0_outputs(9481)) or (layer0_outputs(8204));
    layer1_outputs(4096) <= not(layer0_outputs(9187));
    layer1_outputs(4097) <= not((layer0_outputs(7247)) and (layer0_outputs(8264)));
    layer1_outputs(4098) <= not((layer0_outputs(5195)) xor (layer0_outputs(2864)));
    layer1_outputs(4099) <= not((layer0_outputs(3420)) and (layer0_outputs(3724)));
    layer1_outputs(4100) <= (layer0_outputs(5125)) or (layer0_outputs(8416));
    layer1_outputs(4101) <= (layer0_outputs(470)) and (layer0_outputs(4210));
    layer1_outputs(4102) <= not(layer0_outputs(3841));
    layer1_outputs(4103) <= (layer0_outputs(4825)) and not (layer0_outputs(7368));
    layer1_outputs(4104) <= not((layer0_outputs(5246)) xor (layer0_outputs(9920)));
    layer1_outputs(4105) <= (layer0_outputs(366)) xor (layer0_outputs(5039));
    layer1_outputs(4106) <= not((layer0_outputs(1183)) and (layer0_outputs(1597)));
    layer1_outputs(4107) <= not((layer0_outputs(3349)) and (layer0_outputs(5064)));
    layer1_outputs(4108) <= (layer0_outputs(579)) or (layer0_outputs(5415));
    layer1_outputs(4109) <= not(layer0_outputs(4163));
    layer1_outputs(4110) <= not(layer0_outputs(6857));
    layer1_outputs(4111) <= not(layer0_outputs(2041)) or (layer0_outputs(1007));
    layer1_outputs(4112) <= (layer0_outputs(3125)) and (layer0_outputs(3499));
    layer1_outputs(4113) <= not(layer0_outputs(7189));
    layer1_outputs(4114) <= (layer0_outputs(3075)) and not (layer0_outputs(3540));
    layer1_outputs(4115) <= not((layer0_outputs(6602)) and (layer0_outputs(2366)));
    layer1_outputs(4116) <= not((layer0_outputs(277)) and (layer0_outputs(1302)));
    layer1_outputs(4117) <= (layer0_outputs(6997)) or (layer0_outputs(9816));
    layer1_outputs(4118) <= not(layer0_outputs(1881));
    layer1_outputs(4119) <= layer0_outputs(5566);
    layer1_outputs(4120) <= not((layer0_outputs(1993)) xor (layer0_outputs(9963)));
    layer1_outputs(4121) <= layer0_outputs(5320);
    layer1_outputs(4122) <= layer0_outputs(6734);
    layer1_outputs(4123) <= not(layer0_outputs(5279)) or (layer0_outputs(796));
    layer1_outputs(4124) <= not(layer0_outputs(2176));
    layer1_outputs(4125) <= (layer0_outputs(9397)) xor (layer0_outputs(9176));
    layer1_outputs(4126) <= not((layer0_outputs(9865)) xor (layer0_outputs(10221)));
    layer1_outputs(4127) <= not((layer0_outputs(9010)) and (layer0_outputs(698)));
    layer1_outputs(4128) <= not(layer0_outputs(9571));
    layer1_outputs(4129) <= layer0_outputs(10137);
    layer1_outputs(4130) <= not(layer0_outputs(3347));
    layer1_outputs(4131) <= not(layer0_outputs(833));
    layer1_outputs(4132) <= (layer0_outputs(1163)) and not (layer0_outputs(8505));
    layer1_outputs(4133) <= layer0_outputs(8901);
    layer1_outputs(4134) <= layer0_outputs(79);
    layer1_outputs(4135) <= layer0_outputs(2842);
    layer1_outputs(4136) <= '0';
    layer1_outputs(4137) <= (layer0_outputs(5486)) and (layer0_outputs(4008));
    layer1_outputs(4138) <= (layer0_outputs(3733)) and (layer0_outputs(4590));
    layer1_outputs(4139) <= not(layer0_outputs(5808));
    layer1_outputs(4140) <= layer0_outputs(1734);
    layer1_outputs(4141) <= layer0_outputs(5614);
    layer1_outputs(4142) <= layer0_outputs(6378);
    layer1_outputs(4143) <= layer0_outputs(6413);
    layer1_outputs(4144) <= not((layer0_outputs(2644)) xor (layer0_outputs(9127)));
    layer1_outputs(4145) <= layer0_outputs(7303);
    layer1_outputs(4146) <= not(layer0_outputs(7128)) or (layer0_outputs(2431));
    layer1_outputs(4147) <= not((layer0_outputs(6441)) and (layer0_outputs(6835)));
    layer1_outputs(4148) <= (layer0_outputs(6044)) and not (layer0_outputs(8410));
    layer1_outputs(4149) <= layer0_outputs(3513);
    layer1_outputs(4150) <= (layer0_outputs(5496)) and (layer0_outputs(5982));
    layer1_outputs(4151) <= layer0_outputs(3197);
    layer1_outputs(4152) <= (layer0_outputs(56)) or (layer0_outputs(7354));
    layer1_outputs(4153) <= layer0_outputs(8033);
    layer1_outputs(4154) <= not(layer0_outputs(2768));
    layer1_outputs(4155) <= (layer0_outputs(10177)) and not (layer0_outputs(2887));
    layer1_outputs(4156) <= (layer0_outputs(675)) and not (layer0_outputs(6951));
    layer1_outputs(4157) <= layer0_outputs(5267);
    layer1_outputs(4158) <= not((layer0_outputs(2763)) xor (layer0_outputs(3638)));
    layer1_outputs(4159) <= (layer0_outputs(8222)) and (layer0_outputs(6037));
    layer1_outputs(4160) <= (layer0_outputs(7725)) and not (layer0_outputs(8635));
    layer1_outputs(4161) <= not(layer0_outputs(1734));
    layer1_outputs(4162) <= layer0_outputs(5019);
    layer1_outputs(4163) <= (layer0_outputs(1900)) or (layer0_outputs(8331));
    layer1_outputs(4164) <= (layer0_outputs(7823)) and (layer0_outputs(1787));
    layer1_outputs(4165) <= not((layer0_outputs(1487)) and (layer0_outputs(5860)));
    layer1_outputs(4166) <= (layer0_outputs(9893)) and not (layer0_outputs(1309));
    layer1_outputs(4167) <= not(layer0_outputs(582)) or (layer0_outputs(5980));
    layer1_outputs(4168) <= not(layer0_outputs(6614));
    layer1_outputs(4169) <= layer0_outputs(3891);
    layer1_outputs(4170) <= layer0_outputs(7508);
    layer1_outputs(4171) <= not(layer0_outputs(360));
    layer1_outputs(4172) <= not((layer0_outputs(2652)) and (layer0_outputs(3819)));
    layer1_outputs(4173) <= not(layer0_outputs(9110)) or (layer0_outputs(9750));
    layer1_outputs(4174) <= (layer0_outputs(6388)) and not (layer0_outputs(8418));
    layer1_outputs(4175) <= not((layer0_outputs(6897)) or (layer0_outputs(64)));
    layer1_outputs(4176) <= not(layer0_outputs(9575));
    layer1_outputs(4177) <= layer0_outputs(9122);
    layer1_outputs(4178) <= not(layer0_outputs(294));
    layer1_outputs(4179) <= layer0_outputs(8814);
    layer1_outputs(4180) <= not(layer0_outputs(3579)) or (layer0_outputs(2402));
    layer1_outputs(4181) <= layer0_outputs(8931);
    layer1_outputs(4182) <= (layer0_outputs(5175)) xor (layer0_outputs(2838));
    layer1_outputs(4183) <= layer0_outputs(4462);
    layer1_outputs(4184) <= not((layer0_outputs(4504)) and (layer0_outputs(6809)));
    layer1_outputs(4185) <= not(layer0_outputs(6188));
    layer1_outputs(4186) <= not(layer0_outputs(765)) or (layer0_outputs(9544));
    layer1_outputs(4187) <= layer0_outputs(9362);
    layer1_outputs(4188) <= not(layer0_outputs(4454));
    layer1_outputs(4189) <= not(layer0_outputs(2617));
    layer1_outputs(4190) <= layer0_outputs(5109);
    layer1_outputs(4191) <= not((layer0_outputs(944)) and (layer0_outputs(369)));
    layer1_outputs(4192) <= (layer0_outputs(6639)) or (layer0_outputs(9610));
    layer1_outputs(4193) <= not((layer0_outputs(7471)) or (layer0_outputs(5765)));
    layer1_outputs(4194) <= (layer0_outputs(4011)) and (layer0_outputs(8822));
    layer1_outputs(4195) <= (layer0_outputs(3960)) and (layer0_outputs(117));
    layer1_outputs(4196) <= layer0_outputs(2011);
    layer1_outputs(4197) <= '1';
    layer1_outputs(4198) <= not(layer0_outputs(9161)) or (layer0_outputs(8704));
    layer1_outputs(4199) <= (layer0_outputs(1811)) and not (layer0_outputs(4720));
    layer1_outputs(4200) <= layer0_outputs(8026);
    layer1_outputs(4201) <= not((layer0_outputs(9385)) and (layer0_outputs(9733)));
    layer1_outputs(4202) <= not(layer0_outputs(7392)) or (layer0_outputs(3312));
    layer1_outputs(4203) <= not(layer0_outputs(4438));
    layer1_outputs(4204) <= layer0_outputs(7991);
    layer1_outputs(4205) <= not(layer0_outputs(928));
    layer1_outputs(4206) <= not(layer0_outputs(9816));
    layer1_outputs(4207) <= not(layer0_outputs(1312));
    layer1_outputs(4208) <= not((layer0_outputs(8338)) xor (layer0_outputs(5178)));
    layer1_outputs(4209) <= layer0_outputs(6858);
    layer1_outputs(4210) <= (layer0_outputs(4145)) and (layer0_outputs(3628));
    layer1_outputs(4211) <= (layer0_outputs(529)) and (layer0_outputs(670));
    layer1_outputs(4212) <= not(layer0_outputs(4587)) or (layer0_outputs(8694));
    layer1_outputs(4213) <= (layer0_outputs(4748)) and (layer0_outputs(4908));
    layer1_outputs(4214) <= (layer0_outputs(8200)) and not (layer0_outputs(122));
    layer1_outputs(4215) <= (layer0_outputs(9998)) or (layer0_outputs(4788));
    layer1_outputs(4216) <= (layer0_outputs(1574)) xor (layer0_outputs(8110));
    layer1_outputs(4217) <= not(layer0_outputs(5194));
    layer1_outputs(4218) <= not(layer0_outputs(1370)) or (layer0_outputs(650));
    layer1_outputs(4219) <= not(layer0_outputs(9390));
    layer1_outputs(4220) <= not(layer0_outputs(692));
    layer1_outputs(4221) <= not(layer0_outputs(9215));
    layer1_outputs(4222) <= layer0_outputs(5308);
    layer1_outputs(4223) <= not((layer0_outputs(5384)) and (layer0_outputs(911)));
    layer1_outputs(4224) <= not(layer0_outputs(4837));
    layer1_outputs(4225) <= not(layer0_outputs(8558));
    layer1_outputs(4226) <= layer0_outputs(7158);
    layer1_outputs(4227) <= not(layer0_outputs(5774)) or (layer0_outputs(849));
    layer1_outputs(4228) <= not((layer0_outputs(7463)) or (layer0_outputs(1697)));
    layer1_outputs(4229) <= not(layer0_outputs(1702));
    layer1_outputs(4230) <= layer0_outputs(3527);
    layer1_outputs(4231) <= layer0_outputs(8816);
    layer1_outputs(4232) <= (layer0_outputs(736)) and not (layer0_outputs(6703));
    layer1_outputs(4233) <= layer0_outputs(1770);
    layer1_outputs(4234) <= not((layer0_outputs(5257)) or (layer0_outputs(7604)));
    layer1_outputs(4235) <= (layer0_outputs(490)) and not (layer0_outputs(8196));
    layer1_outputs(4236) <= not(layer0_outputs(4985));
    layer1_outputs(4237) <= (layer0_outputs(7131)) and not (layer0_outputs(3802));
    layer1_outputs(4238) <= layer0_outputs(5844);
    layer1_outputs(4239) <= layer0_outputs(5072);
    layer1_outputs(4240) <= not(layer0_outputs(3935));
    layer1_outputs(4241) <= layer0_outputs(1516);
    layer1_outputs(4242) <= (layer0_outputs(940)) and not (layer0_outputs(9109));
    layer1_outputs(4243) <= layer0_outputs(8607);
    layer1_outputs(4244) <= (layer0_outputs(662)) and not (layer0_outputs(3637));
    layer1_outputs(4245) <= (layer0_outputs(9)) and (layer0_outputs(8235));
    layer1_outputs(4246) <= layer0_outputs(5052);
    layer1_outputs(4247) <= not((layer0_outputs(6199)) and (layer0_outputs(9985)));
    layer1_outputs(4248) <= not(layer0_outputs(5991));
    layer1_outputs(4249) <= layer0_outputs(6522);
    layer1_outputs(4250) <= '0';
    layer1_outputs(4251) <= layer0_outputs(7034);
    layer1_outputs(4252) <= not(layer0_outputs(9905));
    layer1_outputs(4253) <= not(layer0_outputs(6054)) or (layer0_outputs(5545));
    layer1_outputs(4254) <= '1';
    layer1_outputs(4255) <= layer0_outputs(5522);
    layer1_outputs(4256) <= layer0_outputs(1685);
    layer1_outputs(4257) <= not(layer0_outputs(7073)) or (layer0_outputs(6237));
    layer1_outputs(4258) <= not(layer0_outputs(1240));
    layer1_outputs(4259) <= not(layer0_outputs(6104));
    layer1_outputs(4260) <= not((layer0_outputs(9612)) or (layer0_outputs(3509)));
    layer1_outputs(4261) <= not(layer0_outputs(275));
    layer1_outputs(4262) <= layer0_outputs(9716);
    layer1_outputs(4263) <= not(layer0_outputs(5995)) or (layer0_outputs(1847));
    layer1_outputs(4264) <= (layer0_outputs(7379)) and (layer0_outputs(7241));
    layer1_outputs(4265) <= not(layer0_outputs(8660));
    layer1_outputs(4266) <= layer0_outputs(10132);
    layer1_outputs(4267) <= (layer0_outputs(1271)) xor (layer0_outputs(8857));
    layer1_outputs(4268) <= not(layer0_outputs(9223));
    layer1_outputs(4269) <= layer0_outputs(6944);
    layer1_outputs(4270) <= layer0_outputs(7270);
    layer1_outputs(4271) <= not((layer0_outputs(4899)) and (layer0_outputs(8262)));
    layer1_outputs(4272) <= layer0_outputs(7863);
    layer1_outputs(4273) <= not(layer0_outputs(6888));
    layer1_outputs(4274) <= (layer0_outputs(9551)) or (layer0_outputs(3430));
    layer1_outputs(4275) <= not(layer0_outputs(811));
    layer1_outputs(4276) <= not(layer0_outputs(9639));
    layer1_outputs(4277) <= (layer0_outputs(4446)) and not (layer0_outputs(9113));
    layer1_outputs(4278) <= (layer0_outputs(6679)) xor (layer0_outputs(7255));
    layer1_outputs(4279) <= not(layer0_outputs(9121));
    layer1_outputs(4280) <= layer0_outputs(6683);
    layer1_outputs(4281) <= layer0_outputs(2795);
    layer1_outputs(4282) <= '0';
    layer1_outputs(4283) <= not((layer0_outputs(5605)) xor (layer0_outputs(7909)));
    layer1_outputs(4284) <= layer0_outputs(5436);
    layer1_outputs(4285) <= not(layer0_outputs(7468));
    layer1_outputs(4286) <= not(layer0_outputs(4413));
    layer1_outputs(4287) <= (layer0_outputs(7403)) or (layer0_outputs(727));
    layer1_outputs(4288) <= (layer0_outputs(1378)) and (layer0_outputs(4669));
    layer1_outputs(4289) <= (layer0_outputs(3780)) and not (layer0_outputs(6865));
    layer1_outputs(4290) <= not(layer0_outputs(5471));
    layer1_outputs(4291) <= not(layer0_outputs(8225));
    layer1_outputs(4292) <= (layer0_outputs(2415)) or (layer0_outputs(6593));
    layer1_outputs(4293) <= layer0_outputs(6498);
    layer1_outputs(4294) <= not(layer0_outputs(112));
    layer1_outputs(4295) <= layer0_outputs(1995);
    layer1_outputs(4296) <= not((layer0_outputs(3397)) or (layer0_outputs(8236)));
    layer1_outputs(4297) <= (layer0_outputs(3479)) or (layer0_outputs(1238));
    layer1_outputs(4298) <= layer0_outputs(6123);
    layer1_outputs(4299) <= layer0_outputs(5915);
    layer1_outputs(4300) <= (layer0_outputs(3817)) xor (layer0_outputs(6801));
    layer1_outputs(4301) <= not((layer0_outputs(4024)) xor (layer0_outputs(8320)));
    layer1_outputs(4302) <= (layer0_outputs(7994)) or (layer0_outputs(8413));
    layer1_outputs(4303) <= layer0_outputs(4822);
    layer1_outputs(4304) <= not((layer0_outputs(6261)) and (layer0_outputs(8207)));
    layer1_outputs(4305) <= (layer0_outputs(4484)) xor (layer0_outputs(458));
    layer1_outputs(4306) <= (layer0_outputs(10198)) and not (layer0_outputs(7926));
    layer1_outputs(4307) <= not(layer0_outputs(8828));
    layer1_outputs(4308) <= (layer0_outputs(2425)) and (layer0_outputs(2343));
    layer1_outputs(4309) <= (layer0_outputs(632)) or (layer0_outputs(5265));
    layer1_outputs(4310) <= (layer0_outputs(7772)) and not (layer0_outputs(216));
    layer1_outputs(4311) <= '0';
    layer1_outputs(4312) <= not(layer0_outputs(3785));
    layer1_outputs(4313) <= (layer0_outputs(6789)) or (layer0_outputs(2173));
    layer1_outputs(4314) <= (layer0_outputs(6546)) and not (layer0_outputs(6289));
    layer1_outputs(4315) <= not(layer0_outputs(4464)) or (layer0_outputs(6131));
    layer1_outputs(4316) <= (layer0_outputs(7020)) and (layer0_outputs(3551));
    layer1_outputs(4317) <= not(layer0_outputs(287));
    layer1_outputs(4318) <= '0';
    layer1_outputs(4319) <= not(layer0_outputs(8083));
    layer1_outputs(4320) <= (layer0_outputs(1256)) and (layer0_outputs(2709));
    layer1_outputs(4321) <= not(layer0_outputs(5452));
    layer1_outputs(4322) <= layer0_outputs(5622);
    layer1_outputs(4323) <= (layer0_outputs(10218)) and not (layer0_outputs(3231));
    layer1_outputs(4324) <= not(layer0_outputs(6332));
    layer1_outputs(4325) <= not(layer0_outputs(7995)) or (layer0_outputs(779));
    layer1_outputs(4326) <= '0';
    layer1_outputs(4327) <= not(layer0_outputs(5417)) or (layer0_outputs(7153));
    layer1_outputs(4328) <= layer0_outputs(4686);
    layer1_outputs(4329) <= not(layer0_outputs(3597)) or (layer0_outputs(504));
    layer1_outputs(4330) <= (layer0_outputs(6448)) and not (layer0_outputs(1190));
    layer1_outputs(4331) <= not((layer0_outputs(7665)) xor (layer0_outputs(9003)));
    layer1_outputs(4332) <= layer0_outputs(645);
    layer1_outputs(4333) <= (layer0_outputs(6170)) and (layer0_outputs(4442));
    layer1_outputs(4334) <= not(layer0_outputs(9682));
    layer1_outputs(4335) <= (layer0_outputs(6669)) or (layer0_outputs(5263));
    layer1_outputs(4336) <= (layer0_outputs(8944)) or (layer0_outputs(8190));
    layer1_outputs(4337) <= not(layer0_outputs(1120));
    layer1_outputs(4338) <= not((layer0_outputs(5142)) and (layer0_outputs(7428)));
    layer1_outputs(4339) <= (layer0_outputs(1530)) and not (layer0_outputs(4305));
    layer1_outputs(4340) <= (layer0_outputs(9945)) xor (layer0_outputs(1295));
    layer1_outputs(4341) <= not(layer0_outputs(6207)) or (layer0_outputs(220));
    layer1_outputs(4342) <= layer0_outputs(3047);
    layer1_outputs(4343) <= (layer0_outputs(5388)) and (layer0_outputs(4570));
    layer1_outputs(4344) <= not(layer0_outputs(2103));
    layer1_outputs(4345) <= not((layer0_outputs(8402)) and (layer0_outputs(3854)));
    layer1_outputs(4346) <= layer0_outputs(10025);
    layer1_outputs(4347) <= not(layer0_outputs(1389));
    layer1_outputs(4348) <= (layer0_outputs(1842)) xor (layer0_outputs(9590));
    layer1_outputs(4349) <= not(layer0_outputs(2623));
    layer1_outputs(4350) <= (layer0_outputs(1512)) and (layer0_outputs(4439));
    layer1_outputs(4351) <= not((layer0_outputs(3003)) and (layer0_outputs(4813)));
    layer1_outputs(4352) <= (layer0_outputs(5725)) and (layer0_outputs(68));
    layer1_outputs(4353) <= not((layer0_outputs(3222)) and (layer0_outputs(5682)));
    layer1_outputs(4354) <= (layer0_outputs(611)) and (layer0_outputs(2881));
    layer1_outputs(4355) <= (layer0_outputs(6840)) and (layer0_outputs(7567));
    layer1_outputs(4356) <= not((layer0_outputs(9012)) or (layer0_outputs(6397)));
    layer1_outputs(4357) <= '0';
    layer1_outputs(4358) <= layer0_outputs(50);
    layer1_outputs(4359) <= not((layer0_outputs(5880)) and (layer0_outputs(6357)));
    layer1_outputs(4360) <= not(layer0_outputs(2322));
    layer1_outputs(4361) <= (layer0_outputs(1308)) or (layer0_outputs(10096));
    layer1_outputs(4362) <= not((layer0_outputs(901)) and (layer0_outputs(8753)));
    layer1_outputs(4363) <= not(layer0_outputs(485));
    layer1_outputs(4364) <= not(layer0_outputs(1656));
    layer1_outputs(4365) <= not(layer0_outputs(1552));
    layer1_outputs(4366) <= (layer0_outputs(9430)) and not (layer0_outputs(2178));
    layer1_outputs(4367) <= (layer0_outputs(8406)) and not (layer0_outputs(6626));
    layer1_outputs(4368) <= (layer0_outputs(2090)) and not (layer0_outputs(469));
    layer1_outputs(4369) <= layer0_outputs(2901);
    layer1_outputs(4370) <= (layer0_outputs(3354)) or (layer0_outputs(7949));
    layer1_outputs(4371) <= (layer0_outputs(7889)) and not (layer0_outputs(6640));
    layer1_outputs(4372) <= layer0_outputs(8251);
    layer1_outputs(4373) <= layer0_outputs(2783);
    layer1_outputs(4374) <= (layer0_outputs(10036)) or (layer0_outputs(5669));
    layer1_outputs(4375) <= layer0_outputs(9320);
    layer1_outputs(4376) <= (layer0_outputs(1879)) and (layer0_outputs(4617));
    layer1_outputs(4377) <= (layer0_outputs(7221)) and (layer0_outputs(3543));
    layer1_outputs(4378) <= layer0_outputs(5015);
    layer1_outputs(4379) <= not(layer0_outputs(3167)) or (layer0_outputs(8516));
    layer1_outputs(4380) <= not(layer0_outputs(8719)) or (layer0_outputs(4546));
    layer1_outputs(4381) <= layer0_outputs(5007);
    layer1_outputs(4382) <= layer0_outputs(9311);
    layer1_outputs(4383) <= (layer0_outputs(4190)) and (layer0_outputs(1809));
    layer1_outputs(4384) <= not(layer0_outputs(7990));
    layer1_outputs(4385) <= not(layer0_outputs(10127));
    layer1_outputs(4386) <= not((layer0_outputs(9318)) or (layer0_outputs(5562)));
    layer1_outputs(4387) <= (layer0_outputs(3371)) xor (layer0_outputs(6425));
    layer1_outputs(4388) <= layer0_outputs(2746);
    layer1_outputs(4389) <= layer0_outputs(1549);
    layer1_outputs(4390) <= layer0_outputs(3877);
    layer1_outputs(4391) <= not(layer0_outputs(770)) or (layer0_outputs(7573));
    layer1_outputs(4392) <= layer0_outputs(4798);
    layer1_outputs(4393) <= not(layer0_outputs(2217));
    layer1_outputs(4394) <= not((layer0_outputs(6573)) xor (layer0_outputs(7787)));
    layer1_outputs(4395) <= (layer0_outputs(7033)) and not (layer0_outputs(5822));
    layer1_outputs(4396) <= not(layer0_outputs(3694));
    layer1_outputs(4397) <= layer0_outputs(4808);
    layer1_outputs(4398) <= not(layer0_outputs(1299));
    layer1_outputs(4399) <= not(layer0_outputs(4980)) or (layer0_outputs(5858));
    layer1_outputs(4400) <= not(layer0_outputs(1508));
    layer1_outputs(4401) <= (layer0_outputs(7988)) and not (layer0_outputs(8874));
    layer1_outputs(4402) <= (layer0_outputs(9154)) and (layer0_outputs(6219));
    layer1_outputs(4403) <= not(layer0_outputs(6235));
    layer1_outputs(4404) <= layer0_outputs(141);
    layer1_outputs(4405) <= layer0_outputs(4566);
    layer1_outputs(4406) <= (layer0_outputs(5103)) and not (layer0_outputs(370));
    layer1_outputs(4407) <= not((layer0_outputs(3002)) or (layer0_outputs(3838)));
    layer1_outputs(4408) <= layer0_outputs(4298);
    layer1_outputs(4409) <= (layer0_outputs(7329)) and (layer0_outputs(5742));
    layer1_outputs(4410) <= not(layer0_outputs(302));
    layer1_outputs(4411) <= not(layer0_outputs(6985));
    layer1_outputs(4412) <= not(layer0_outputs(4897)) or (layer0_outputs(6651));
    layer1_outputs(4413) <= not((layer0_outputs(9932)) or (layer0_outputs(9059)));
    layer1_outputs(4414) <= not(layer0_outputs(8773));
    layer1_outputs(4415) <= not((layer0_outputs(6244)) xor (layer0_outputs(5390)));
    layer1_outputs(4416) <= (layer0_outputs(8508)) and not (layer0_outputs(1241));
    layer1_outputs(4417) <= not(layer0_outputs(3295));
    layer1_outputs(4418) <= layer0_outputs(7472);
    layer1_outputs(4419) <= '1';
    layer1_outputs(4420) <= (layer0_outputs(9387)) xor (layer0_outputs(439));
    layer1_outputs(4421) <= (layer0_outputs(5649)) and not (layer0_outputs(9545));
    layer1_outputs(4422) <= layer0_outputs(5162);
    layer1_outputs(4423) <= layer0_outputs(3113);
    layer1_outputs(4424) <= not(layer0_outputs(8343));
    layer1_outputs(4425) <= not(layer0_outputs(1017)) or (layer0_outputs(4451));
    layer1_outputs(4426) <= not((layer0_outputs(8316)) and (layer0_outputs(3108)));
    layer1_outputs(4427) <= not((layer0_outputs(6655)) and (layer0_outputs(2698)));
    layer1_outputs(4428) <= not((layer0_outputs(2899)) or (layer0_outputs(7087)));
    layer1_outputs(4429) <= not(layer0_outputs(3192));
    layer1_outputs(4430) <= (layer0_outputs(8709)) or (layer0_outputs(1949));
    layer1_outputs(4431) <= '0';
    layer1_outputs(4432) <= layer0_outputs(3328);
    layer1_outputs(4433) <= not(layer0_outputs(8075));
    layer1_outputs(4434) <= not(layer0_outputs(3007));
    layer1_outputs(4435) <= layer0_outputs(9349);
    layer1_outputs(4436) <= (layer0_outputs(1789)) and not (layer0_outputs(3222));
    layer1_outputs(4437) <= (layer0_outputs(7633)) or (layer0_outputs(3446));
    layer1_outputs(4438) <= (layer0_outputs(5297)) and not (layer0_outputs(5462));
    layer1_outputs(4439) <= not((layer0_outputs(9087)) and (layer0_outputs(5461)));
    layer1_outputs(4440) <= not((layer0_outputs(2164)) or (layer0_outputs(2809)));
    layer1_outputs(4441) <= (layer0_outputs(3422)) xor (layer0_outputs(2419));
    layer1_outputs(4442) <= not(layer0_outputs(9206));
    layer1_outputs(4443) <= (layer0_outputs(1489)) and (layer0_outputs(701));
    layer1_outputs(4444) <= '1';
    layer1_outputs(4445) <= (layer0_outputs(8487)) xor (layer0_outputs(2561));
    layer1_outputs(4446) <= (layer0_outputs(3170)) and not (layer0_outputs(5495));
    layer1_outputs(4447) <= (layer0_outputs(8945)) and not (layer0_outputs(6353));
    layer1_outputs(4448) <= not(layer0_outputs(7485));
    layer1_outputs(4449) <= not(layer0_outputs(7802));
    layer1_outputs(4450) <= not((layer0_outputs(7528)) and (layer0_outputs(7928)));
    layer1_outputs(4451) <= not(layer0_outputs(5511));
    layer1_outputs(4452) <= (layer0_outputs(7502)) and (layer0_outputs(8999));
    layer1_outputs(4453) <= not(layer0_outputs(8918));
    layer1_outputs(4454) <= (layer0_outputs(6154)) and (layer0_outputs(407));
    layer1_outputs(4455) <= not(layer0_outputs(2006));
    layer1_outputs(4456) <= not(layer0_outputs(4308)) or (layer0_outputs(8365));
    layer1_outputs(4457) <= (layer0_outputs(9769)) and not (layer0_outputs(546));
    layer1_outputs(4458) <= not(layer0_outputs(9450));
    layer1_outputs(4459) <= not(layer0_outputs(206));
    layer1_outputs(4460) <= layer0_outputs(8010);
    layer1_outputs(4461) <= layer0_outputs(5976);
    layer1_outputs(4462) <= not((layer0_outputs(176)) and (layer0_outputs(5243)));
    layer1_outputs(4463) <= not((layer0_outputs(2373)) or (layer0_outputs(8127)));
    layer1_outputs(4464) <= (layer0_outputs(653)) and not (layer0_outputs(5693));
    layer1_outputs(4465) <= not((layer0_outputs(3091)) and (layer0_outputs(2536)));
    layer1_outputs(4466) <= not(layer0_outputs(9837)) or (layer0_outputs(5363));
    layer1_outputs(4467) <= not(layer0_outputs(2779)) or (layer0_outputs(3311));
    layer1_outputs(4468) <= not((layer0_outputs(4303)) xor (layer0_outputs(9136)));
    layer1_outputs(4469) <= layer0_outputs(6224);
    layer1_outputs(4470) <= not(layer0_outputs(5836));
    layer1_outputs(4471) <= not(layer0_outputs(4469)) or (layer0_outputs(876));
    layer1_outputs(4472) <= not(layer0_outputs(600));
    layer1_outputs(4473) <= not((layer0_outputs(3168)) and (layer0_outputs(9463)));
    layer1_outputs(4474) <= (layer0_outputs(6226)) and not (layer0_outputs(8567));
    layer1_outputs(4475) <= layer0_outputs(1794);
    layer1_outputs(4476) <= not((layer0_outputs(3849)) or (layer0_outputs(2050)));
    layer1_outputs(4477) <= not(layer0_outputs(2735));
    layer1_outputs(4478) <= not(layer0_outputs(7464));
    layer1_outputs(4479) <= (layer0_outputs(6755)) or (layer0_outputs(4028));
    layer1_outputs(4480) <= not(layer0_outputs(6239));
    layer1_outputs(4481) <= not(layer0_outputs(6248));
    layer1_outputs(4482) <= not(layer0_outputs(5059)) or (layer0_outputs(2256));
    layer1_outputs(4483) <= not((layer0_outputs(987)) or (layer0_outputs(3036)));
    layer1_outputs(4484) <= (layer0_outputs(8657)) and not (layer0_outputs(120));
    layer1_outputs(4485) <= not((layer0_outputs(7169)) or (layer0_outputs(6503)));
    layer1_outputs(4486) <= not(layer0_outputs(8946)) or (layer0_outputs(9377));
    layer1_outputs(4487) <= layer0_outputs(9216);
    layer1_outputs(4488) <= layer0_outputs(3015);
    layer1_outputs(4489) <= not((layer0_outputs(109)) or (layer0_outputs(10050)));
    layer1_outputs(4490) <= not(layer0_outputs(6286));
    layer1_outputs(4491) <= not((layer0_outputs(4626)) or (layer0_outputs(6327)));
    layer1_outputs(4492) <= (layer0_outputs(32)) and not (layer0_outputs(7568));
    layer1_outputs(4493) <= layer0_outputs(7603);
    layer1_outputs(4494) <= (layer0_outputs(2418)) xor (layer0_outputs(5718));
    layer1_outputs(4495) <= not(layer0_outputs(8067)) or (layer0_outputs(10009));
    layer1_outputs(4496) <= layer0_outputs(8885);
    layer1_outputs(4497) <= (layer0_outputs(9537)) or (layer0_outputs(1505));
    layer1_outputs(4498) <= (layer0_outputs(1057)) xor (layer0_outputs(8391));
    layer1_outputs(4499) <= layer0_outputs(2262);
    layer1_outputs(4500) <= (layer0_outputs(1471)) and not (layer0_outputs(7783));
    layer1_outputs(4501) <= layer0_outputs(8226);
    layer1_outputs(4502) <= not((layer0_outputs(1821)) or (layer0_outputs(7194)));
    layer1_outputs(4503) <= not((layer0_outputs(2896)) xor (layer0_outputs(1974)));
    layer1_outputs(4504) <= (layer0_outputs(6740)) and not (layer0_outputs(4641));
    layer1_outputs(4505) <= (layer0_outputs(7139)) and not (layer0_outputs(6511));
    layer1_outputs(4506) <= not((layer0_outputs(3380)) or (layer0_outputs(4241)));
    layer1_outputs(4507) <= not(layer0_outputs(3366));
    layer1_outputs(4508) <= not((layer0_outputs(1877)) xor (layer0_outputs(8523)));
    layer1_outputs(4509) <= (layer0_outputs(7187)) or (layer0_outputs(1571));
    layer1_outputs(4510) <= (layer0_outputs(6466)) and not (layer0_outputs(4092));
    layer1_outputs(4511) <= (layer0_outputs(5663)) and (layer0_outputs(2990));
    layer1_outputs(4512) <= not(layer0_outputs(2564)) or (layer0_outputs(2643));
    layer1_outputs(4513) <= layer0_outputs(4407);
    layer1_outputs(4514) <= (layer0_outputs(406)) and not (layer0_outputs(5628));
    layer1_outputs(4515) <= layer0_outputs(9937);
    layer1_outputs(4516) <= not((layer0_outputs(1170)) and (layer0_outputs(10071)));
    layer1_outputs(4517) <= not(layer0_outputs(9915)) or (layer0_outputs(4875));
    layer1_outputs(4518) <= not(layer0_outputs(6589));
    layer1_outputs(4519) <= not((layer0_outputs(1089)) or (layer0_outputs(3272)));
    layer1_outputs(4520) <= not(layer0_outputs(1099));
    layer1_outputs(4521) <= (layer0_outputs(3327)) and not (layer0_outputs(6939));
    layer1_outputs(4522) <= '1';
    layer1_outputs(4523) <= not(layer0_outputs(2508));
    layer1_outputs(4524) <= not((layer0_outputs(5558)) or (layer0_outputs(9318)));
    layer1_outputs(4525) <= not(layer0_outputs(4181));
    layer1_outputs(4526) <= not((layer0_outputs(1425)) or (layer0_outputs(5056)));
    layer1_outputs(4527) <= not(layer0_outputs(10032));
    layer1_outputs(4528) <= not((layer0_outputs(9841)) or (layer0_outputs(104)));
    layer1_outputs(4529) <= (layer0_outputs(5934)) xor (layer0_outputs(3199));
    layer1_outputs(4530) <= not((layer0_outputs(1796)) xor (layer0_outputs(2959)));
    layer1_outputs(4531) <= not(layer0_outputs(6571)) or (layer0_outputs(8659));
    layer1_outputs(4532) <= layer0_outputs(1836);
    layer1_outputs(4533) <= layer0_outputs(7723);
    layer1_outputs(4534) <= not(layer0_outputs(3282)) or (layer0_outputs(9834));
    layer1_outputs(4535) <= not(layer0_outputs(1509));
    layer1_outputs(4536) <= (layer0_outputs(5690)) and (layer0_outputs(3460));
    layer1_outputs(4537) <= (layer0_outputs(5316)) and not (layer0_outputs(9068));
    layer1_outputs(4538) <= (layer0_outputs(831)) xor (layer0_outputs(5571));
    layer1_outputs(4539) <= not(layer0_outputs(1363));
    layer1_outputs(4540) <= not(layer0_outputs(8884)) or (layer0_outputs(7854));
    layer1_outputs(4541) <= not(layer0_outputs(3274));
    layer1_outputs(4542) <= not((layer0_outputs(8948)) xor (layer0_outputs(5154)));
    layer1_outputs(4543) <= '1';
    layer1_outputs(4544) <= not((layer0_outputs(2228)) or (layer0_outputs(9954)));
    layer1_outputs(4545) <= (layer0_outputs(6671)) and not (layer0_outputs(2105));
    layer1_outputs(4546) <= layer0_outputs(9159);
    layer1_outputs(4547) <= not(layer0_outputs(1350)) or (layer0_outputs(7358));
    layer1_outputs(4548) <= not(layer0_outputs(3157)) or (layer0_outputs(2724));
    layer1_outputs(4549) <= not(layer0_outputs(1447));
    layer1_outputs(4550) <= layer0_outputs(9737);
    layer1_outputs(4551) <= not(layer0_outputs(5902));
    layer1_outputs(4552) <= (layer0_outputs(6455)) and not (layer0_outputs(2109));
    layer1_outputs(4553) <= not(layer0_outputs(3372));
    layer1_outputs(4554) <= not(layer0_outputs(4991));
    layer1_outputs(4555) <= layer0_outputs(1743);
    layer1_outputs(4556) <= (layer0_outputs(4862)) and not (layer0_outputs(5334));
    layer1_outputs(4557) <= not(layer0_outputs(9379)) or (layer0_outputs(8429));
    layer1_outputs(4558) <= layer0_outputs(6016);
    layer1_outputs(4559) <= layer0_outputs(9302);
    layer1_outputs(4560) <= not(layer0_outputs(6326));
    layer1_outputs(4561) <= not((layer0_outputs(9129)) xor (layer0_outputs(2500)));
    layer1_outputs(4562) <= not((layer0_outputs(3424)) xor (layer0_outputs(3270)));
    layer1_outputs(4563) <= not(layer0_outputs(8029));
    layer1_outputs(4564) <= not(layer0_outputs(446));
    layer1_outputs(4565) <= layer0_outputs(6137);
    layer1_outputs(4566) <= (layer0_outputs(2402)) or (layer0_outputs(1454));
    layer1_outputs(4567) <= not((layer0_outputs(4713)) and (layer0_outputs(10203)));
    layer1_outputs(4568) <= (layer0_outputs(5602)) and not (layer0_outputs(1291));
    layer1_outputs(4569) <= not(layer0_outputs(6613));
    layer1_outputs(4570) <= not(layer0_outputs(5269));
    layer1_outputs(4571) <= layer0_outputs(3572);
    layer1_outputs(4572) <= layer0_outputs(7693);
    layer1_outputs(4573) <= not((layer0_outputs(5766)) xor (layer0_outputs(3138)));
    layer1_outputs(4574) <= (layer0_outputs(1916)) and not (layer0_outputs(84));
    layer1_outputs(4575) <= not(layer0_outputs(6088));
    layer1_outputs(4576) <= not(layer0_outputs(6269));
    layer1_outputs(4577) <= layer0_outputs(4077);
    layer1_outputs(4578) <= not((layer0_outputs(7701)) or (layer0_outputs(3728)));
    layer1_outputs(4579) <= layer0_outputs(8669);
    layer1_outputs(4580) <= layer0_outputs(1791);
    layer1_outputs(4581) <= not((layer0_outputs(4699)) or (layer0_outputs(4071)));
    layer1_outputs(4582) <= layer0_outputs(9550);
    layer1_outputs(4583) <= not(layer0_outputs(5350));
    layer1_outputs(4584) <= (layer0_outputs(3410)) and (layer0_outputs(9815));
    layer1_outputs(4585) <= not((layer0_outputs(9070)) xor (layer0_outputs(6492)));
    layer1_outputs(4586) <= not((layer0_outputs(2009)) xor (layer0_outputs(9200)));
    layer1_outputs(4587) <= (layer0_outputs(519)) xor (layer0_outputs(9901));
    layer1_outputs(4588) <= not(layer0_outputs(115));
    layer1_outputs(4589) <= not(layer0_outputs(6450)) or (layer0_outputs(8865));
    layer1_outputs(4590) <= (layer0_outputs(7704)) and not (layer0_outputs(9001));
    layer1_outputs(4591) <= layer0_outputs(5697);
    layer1_outputs(4592) <= layer0_outputs(2866);
    layer1_outputs(4593) <= not(layer0_outputs(1396));
    layer1_outputs(4594) <= not((layer0_outputs(8221)) and (layer0_outputs(8126)));
    layer1_outputs(4595) <= not(layer0_outputs(5625)) or (layer0_outputs(3122));
    layer1_outputs(4596) <= not(layer0_outputs(6930));
    layer1_outputs(4597) <= not(layer0_outputs(9735));
    layer1_outputs(4598) <= not(layer0_outputs(2754)) or (layer0_outputs(5866));
    layer1_outputs(4599) <= not((layer0_outputs(4344)) and (layer0_outputs(3898)));
    layer1_outputs(4600) <= (layer0_outputs(1886)) and not (layer0_outputs(5210));
    layer1_outputs(4601) <= not(layer0_outputs(926));
    layer1_outputs(4602) <= layer0_outputs(6734);
    layer1_outputs(4603) <= not(layer0_outputs(3556)) or (layer0_outputs(458));
    layer1_outputs(4604) <= not((layer0_outputs(735)) or (layer0_outputs(2328)));
    layer1_outputs(4605) <= not((layer0_outputs(1902)) xor (layer0_outputs(5290)));
    layer1_outputs(4606) <= not(layer0_outputs(9346)) or (layer0_outputs(3668));
    layer1_outputs(4607) <= not(layer0_outputs(996)) or (layer0_outputs(1277));
    layer1_outputs(4608) <= not(layer0_outputs(5579));
    layer1_outputs(4609) <= not(layer0_outputs(9374));
    layer1_outputs(4610) <= not(layer0_outputs(2514));
    layer1_outputs(4611) <= layer0_outputs(442);
    layer1_outputs(4612) <= (layer0_outputs(5946)) and (layer0_outputs(4150));
    layer1_outputs(4613) <= (layer0_outputs(643)) and (layer0_outputs(9983));
    layer1_outputs(4614) <= (layer0_outputs(5954)) xor (layer0_outputs(10010));
    layer1_outputs(4615) <= not((layer0_outputs(8156)) and (layer0_outputs(7632)));
    layer1_outputs(4616) <= not(layer0_outputs(7270));
    layer1_outputs(4617) <= layer0_outputs(5191);
    layer1_outputs(4618) <= not(layer0_outputs(586)) or (layer0_outputs(7963));
    layer1_outputs(4619) <= not((layer0_outputs(4548)) and (layer0_outputs(836)));
    layer1_outputs(4620) <= not(layer0_outputs(8622)) or (layer0_outputs(4283));
    layer1_outputs(4621) <= not(layer0_outputs(3995)) or (layer0_outputs(5041));
    layer1_outputs(4622) <= not((layer0_outputs(7641)) xor (layer0_outputs(6073)));
    layer1_outputs(4623) <= layer0_outputs(6697);
    layer1_outputs(4624) <= (layer0_outputs(10196)) xor (layer0_outputs(2616));
    layer1_outputs(4625) <= (layer0_outputs(1172)) or (layer0_outputs(1694));
    layer1_outputs(4626) <= not((layer0_outputs(8335)) or (layer0_outputs(9784)));
    layer1_outputs(4627) <= layer0_outputs(7648);
    layer1_outputs(4628) <= (layer0_outputs(1648)) and not (layer0_outputs(3461));
    layer1_outputs(4629) <= not(layer0_outputs(1400));
    layer1_outputs(4630) <= layer0_outputs(1518);
    layer1_outputs(4631) <= not(layer0_outputs(10214)) or (layer0_outputs(8531));
    layer1_outputs(4632) <= not(layer0_outputs(202));
    layer1_outputs(4633) <= layer0_outputs(6493);
    layer1_outputs(4634) <= layer0_outputs(7910);
    layer1_outputs(4635) <= not((layer0_outputs(3239)) and (layer0_outputs(5727)));
    layer1_outputs(4636) <= not(layer0_outputs(9216));
    layer1_outputs(4637) <= layer0_outputs(4867);
    layer1_outputs(4638) <= layer0_outputs(4599);
    layer1_outputs(4639) <= layer0_outputs(2699);
    layer1_outputs(4640) <= layer0_outputs(987);
    layer1_outputs(4641) <= layer0_outputs(9033);
    layer1_outputs(4642) <= layer0_outputs(956);
    layer1_outputs(4643) <= layer0_outputs(5895);
    layer1_outputs(4644) <= not(layer0_outputs(7868));
    layer1_outputs(4645) <= (layer0_outputs(9352)) and (layer0_outputs(3626));
    layer1_outputs(4646) <= (layer0_outputs(6724)) and (layer0_outputs(1882));
    layer1_outputs(4647) <= '0';
    layer1_outputs(4648) <= layer0_outputs(2315);
    layer1_outputs(4649) <= (layer0_outputs(10231)) and (layer0_outputs(2087));
    layer1_outputs(4650) <= not(layer0_outputs(1594));
    layer1_outputs(4651) <= not(layer0_outputs(1132));
    layer1_outputs(4652) <= not((layer0_outputs(4897)) and (layer0_outputs(7162)));
    layer1_outputs(4653) <= (layer0_outputs(1426)) or (layer0_outputs(1893));
    layer1_outputs(4654) <= (layer0_outputs(503)) xor (layer0_outputs(10186));
    layer1_outputs(4655) <= not(layer0_outputs(6004)) or (layer0_outputs(5782));
    layer1_outputs(4656) <= '1';
    layer1_outputs(4657) <= not(layer0_outputs(3118)) or (layer0_outputs(8417));
    layer1_outputs(4658) <= layer0_outputs(2655);
    layer1_outputs(4659) <= (layer0_outputs(5937)) and not (layer0_outputs(3630));
    layer1_outputs(4660) <= not((layer0_outputs(2038)) and (layer0_outputs(1579)));
    layer1_outputs(4661) <= not(layer0_outputs(1301));
    layer1_outputs(4662) <= (layer0_outputs(10216)) and not (layer0_outputs(4359));
    layer1_outputs(4663) <= not((layer0_outputs(7011)) and (layer0_outputs(5747)));
    layer1_outputs(4664) <= layer0_outputs(817);
    layer1_outputs(4665) <= not(layer0_outputs(1094));
    layer1_outputs(4666) <= not(layer0_outputs(9840));
    layer1_outputs(4667) <= not(layer0_outputs(1325));
    layer1_outputs(4668) <= layer0_outputs(4807);
    layer1_outputs(4669) <= not((layer0_outputs(3495)) or (layer0_outputs(2662)));
    layer1_outputs(4670) <= (layer0_outputs(3602)) and not (layer0_outputs(1801));
    layer1_outputs(4671) <= not((layer0_outputs(3396)) xor (layer0_outputs(6980)));
    layer1_outputs(4672) <= not(layer0_outputs(575));
    layer1_outputs(4673) <= not(layer0_outputs(5221));
    layer1_outputs(4674) <= not((layer0_outputs(6787)) and (layer0_outputs(3559)));
    layer1_outputs(4675) <= not((layer0_outputs(2750)) xor (layer0_outputs(5449)));
    layer1_outputs(4676) <= (layer0_outputs(9576)) and not (layer0_outputs(983));
    layer1_outputs(4677) <= not((layer0_outputs(4224)) or (layer0_outputs(4407)));
    layer1_outputs(4678) <= (layer0_outputs(7637)) and not (layer0_outputs(6288));
    layer1_outputs(4679) <= not(layer0_outputs(8138)) or (layer0_outputs(9630));
    layer1_outputs(4680) <= not(layer0_outputs(4682));
    layer1_outputs(4681) <= not(layer0_outputs(5084)) or (layer0_outputs(8579));
    layer1_outputs(4682) <= not(layer0_outputs(7877));
    layer1_outputs(4683) <= (layer0_outputs(9507)) or (layer0_outputs(8412));
    layer1_outputs(4684) <= (layer0_outputs(1138)) and not (layer0_outputs(9592));
    layer1_outputs(4685) <= not((layer0_outputs(2472)) and (layer0_outputs(4588)));
    layer1_outputs(4686) <= (layer0_outputs(7305)) and (layer0_outputs(3419));
    layer1_outputs(4687) <= (layer0_outputs(6928)) xor (layer0_outputs(3912));
    layer1_outputs(4688) <= layer0_outputs(978);
    layer1_outputs(4689) <= not(layer0_outputs(9389)) or (layer0_outputs(9528));
    layer1_outputs(4690) <= (layer0_outputs(5618)) and not (layer0_outputs(1774));
    layer1_outputs(4691) <= not(layer0_outputs(8021));
    layer1_outputs(4692) <= layer0_outputs(690);
    layer1_outputs(4693) <= layer0_outputs(2342);
    layer1_outputs(4694) <= not(layer0_outputs(8084));
    layer1_outputs(4695) <= not(layer0_outputs(5379));
    layer1_outputs(4696) <= (layer0_outputs(3570)) xor (layer0_outputs(1048));
    layer1_outputs(4697) <= layer0_outputs(3930);
    layer1_outputs(4698) <= (layer0_outputs(6210)) or (layer0_outputs(51));
    layer1_outputs(4699) <= not((layer0_outputs(4378)) xor (layer0_outputs(10135)));
    layer1_outputs(4700) <= not((layer0_outputs(3750)) xor (layer0_outputs(8590)));
    layer1_outputs(4701) <= not(layer0_outputs(5410));
    layer1_outputs(4702) <= not(layer0_outputs(5132));
    layer1_outputs(4703) <= layer0_outputs(5964);
    layer1_outputs(4704) <= (layer0_outputs(6730)) and (layer0_outputs(4121));
    layer1_outputs(4705) <= not(layer0_outputs(1605)) or (layer0_outputs(8524));
    layer1_outputs(4706) <= (layer0_outputs(8770)) or (layer0_outputs(91));
    layer1_outputs(4707) <= layer0_outputs(4520);
    layer1_outputs(4708) <= not(layer0_outputs(1546));
    layer1_outputs(4709) <= not((layer0_outputs(5705)) xor (layer0_outputs(7785)));
    layer1_outputs(4710) <= (layer0_outputs(8468)) and not (layer0_outputs(5461));
    layer1_outputs(4711) <= not(layer0_outputs(3681)) or (layer0_outputs(283));
    layer1_outputs(4712) <= not(layer0_outputs(2536)) or (layer0_outputs(3522));
    layer1_outputs(4713) <= not(layer0_outputs(1705));
    layer1_outputs(4714) <= (layer0_outputs(6913)) or (layer0_outputs(1649));
    layer1_outputs(4715) <= (layer0_outputs(4386)) and (layer0_outputs(5612));
    layer1_outputs(4716) <= layer0_outputs(732);
    layer1_outputs(4717) <= not(layer0_outputs(2434));
    layer1_outputs(4718) <= not((layer0_outputs(4026)) and (layer0_outputs(2469)));
    layer1_outputs(4719) <= not((layer0_outputs(965)) xor (layer0_outputs(674)));
    layer1_outputs(4720) <= '1';
    layer1_outputs(4721) <= not(layer0_outputs(3836));
    layer1_outputs(4722) <= layer0_outputs(1987);
    layer1_outputs(4723) <= layer0_outputs(4575);
    layer1_outputs(4724) <= not(layer0_outputs(1147));
    layer1_outputs(4725) <= (layer0_outputs(3852)) and (layer0_outputs(6619));
    layer1_outputs(4726) <= layer0_outputs(5128);
    layer1_outputs(4727) <= layer0_outputs(9128);
    layer1_outputs(4728) <= (layer0_outputs(5253)) and not (layer0_outputs(7326));
    layer1_outputs(4729) <= (layer0_outputs(1700)) and not (layer0_outputs(10006));
    layer1_outputs(4730) <= not(layer0_outputs(5382));
    layer1_outputs(4731) <= (layer0_outputs(7493)) or (layer0_outputs(3302));
    layer1_outputs(4732) <= (layer0_outputs(4541)) or (layer0_outputs(5451));
    layer1_outputs(4733) <= (layer0_outputs(10106)) and not (layer0_outputs(6984));
    layer1_outputs(4734) <= not(layer0_outputs(5157)) or (layer0_outputs(7024));
    layer1_outputs(4735) <= layer0_outputs(2992);
    layer1_outputs(4736) <= not((layer0_outputs(4675)) xor (layer0_outputs(8498)));
    layer1_outputs(4737) <= (layer0_outputs(1146)) and (layer0_outputs(3032));
    layer1_outputs(4738) <= (layer0_outputs(2575)) and (layer0_outputs(4408));
    layer1_outputs(4739) <= not(layer0_outputs(5968));
    layer1_outputs(4740) <= not(layer0_outputs(8782));
    layer1_outputs(4741) <= layer0_outputs(7756);
    layer1_outputs(4742) <= not(layer0_outputs(9446));
    layer1_outputs(4743) <= layer0_outputs(386);
    layer1_outputs(4744) <= layer0_outputs(1860);
    layer1_outputs(4745) <= '0';
    layer1_outputs(4746) <= layer0_outputs(7246);
    layer1_outputs(4747) <= (layer0_outputs(6921)) and (layer0_outputs(5089));
    layer1_outputs(4748) <= not((layer0_outputs(336)) and (layer0_outputs(10084)));
    layer1_outputs(4749) <= (layer0_outputs(9636)) or (layer0_outputs(4384));
    layer1_outputs(4750) <= not(layer0_outputs(8711));
    layer1_outputs(4751) <= (layer0_outputs(8376)) xor (layer0_outputs(1188));
    layer1_outputs(4752) <= not(layer0_outputs(1237)) or (layer0_outputs(9119));
    layer1_outputs(4753) <= not(layer0_outputs(8921));
    layer1_outputs(4754) <= (layer0_outputs(9309)) and (layer0_outputs(4063));
    layer1_outputs(4755) <= not((layer0_outputs(7130)) xor (layer0_outputs(2893)));
    layer1_outputs(4756) <= (layer0_outputs(1250)) or (layer0_outputs(2181));
    layer1_outputs(4757) <= layer0_outputs(6800);
    layer1_outputs(4758) <= not(layer0_outputs(3364)) or (layer0_outputs(9912));
    layer1_outputs(4759) <= not((layer0_outputs(3911)) and (layer0_outputs(8719)));
    layer1_outputs(4760) <= (layer0_outputs(3781)) and not (layer0_outputs(8835));
    layer1_outputs(4761) <= not(layer0_outputs(8335));
    layer1_outputs(4762) <= (layer0_outputs(8859)) and not (layer0_outputs(7496));
    layer1_outputs(4763) <= not(layer0_outputs(8268)) or (layer0_outputs(936));
    layer1_outputs(4764) <= not(layer0_outputs(4489));
    layer1_outputs(4765) <= layer0_outputs(1423);
    layer1_outputs(4766) <= layer0_outputs(2572);
    layer1_outputs(4767) <= (layer0_outputs(1943)) and (layer0_outputs(728));
    layer1_outputs(4768) <= not((layer0_outputs(7886)) xor (layer0_outputs(8268)));
    layer1_outputs(4769) <= (layer0_outputs(3397)) or (layer0_outputs(5656));
    layer1_outputs(4770) <= layer0_outputs(4962);
    layer1_outputs(4771) <= not(layer0_outputs(3918));
    layer1_outputs(4772) <= not(layer0_outputs(3987));
    layer1_outputs(4773) <= not(layer0_outputs(9453)) or (layer0_outputs(9856));
    layer1_outputs(4774) <= (layer0_outputs(49)) and not (layer0_outputs(5562));
    layer1_outputs(4775) <= not(layer0_outputs(5959)) or (layer0_outputs(8114));
    layer1_outputs(4776) <= '0';
    layer1_outputs(4777) <= (layer0_outputs(4244)) and not (layer0_outputs(66));
    layer1_outputs(4778) <= (layer0_outputs(4400)) and not (layer0_outputs(107));
    layer1_outputs(4779) <= (layer0_outputs(103)) xor (layer0_outputs(7544));
    layer1_outputs(4780) <= layer0_outputs(9214);
    layer1_outputs(4781) <= (layer0_outputs(8728)) and not (layer0_outputs(5973));
    layer1_outputs(4782) <= not(layer0_outputs(6438));
    layer1_outputs(4783) <= (layer0_outputs(4497)) or (layer0_outputs(565));
    layer1_outputs(4784) <= layer0_outputs(6968);
    layer1_outputs(4785) <= not((layer0_outputs(5759)) xor (layer0_outputs(3115)));
    layer1_outputs(4786) <= '0';
    layer1_outputs(4787) <= layer0_outputs(1040);
    layer1_outputs(4788) <= layer0_outputs(2064);
    layer1_outputs(4789) <= not(layer0_outputs(1009)) or (layer0_outputs(8858));
    layer1_outputs(4790) <= layer0_outputs(2649);
    layer1_outputs(4791) <= '1';
    layer1_outputs(4792) <= not(layer0_outputs(8502));
    layer1_outputs(4793) <= layer0_outputs(9885);
    layer1_outputs(4794) <= layer0_outputs(2801);
    layer1_outputs(4795) <= not(layer0_outputs(1667));
    layer1_outputs(4796) <= layer0_outputs(9769);
    layer1_outputs(4797) <= not(layer0_outputs(10190)) or (layer0_outputs(3894));
    layer1_outputs(4798) <= not(layer0_outputs(4366));
    layer1_outputs(4799) <= not((layer0_outputs(9411)) and (layer0_outputs(5179)));
    layer1_outputs(4800) <= layer0_outputs(7030);
    layer1_outputs(4801) <= layer0_outputs(6118);
    layer1_outputs(4802) <= layer0_outputs(4647);
    layer1_outputs(4803) <= (layer0_outputs(3292)) and not (layer0_outputs(9098));
    layer1_outputs(4804) <= not(layer0_outputs(6793));
    layer1_outputs(4805) <= (layer0_outputs(6225)) and not (layer0_outputs(2505));
    layer1_outputs(4806) <= not((layer0_outputs(275)) and (layer0_outputs(5140)));
    layer1_outputs(4807) <= not((layer0_outputs(804)) and (layer0_outputs(7769)));
    layer1_outputs(4808) <= not(layer0_outputs(8220));
    layer1_outputs(4809) <= layer0_outputs(8904);
    layer1_outputs(4810) <= '1';
    layer1_outputs(4811) <= (layer0_outputs(9206)) xor (layer0_outputs(5507));
    layer1_outputs(4812) <= not(layer0_outputs(10)) or (layer0_outputs(2332));
    layer1_outputs(4813) <= layer0_outputs(5777);
    layer1_outputs(4814) <= not((layer0_outputs(3974)) or (layer0_outputs(1191)));
    layer1_outputs(4815) <= not((layer0_outputs(3775)) or (layer0_outputs(5581)));
    layer1_outputs(4816) <= layer0_outputs(1560);
    layer1_outputs(4817) <= not((layer0_outputs(845)) and (layer0_outputs(9013)));
    layer1_outputs(4818) <= layer0_outputs(3305);
    layer1_outputs(4819) <= (layer0_outputs(1376)) and not (layer0_outputs(1730));
    layer1_outputs(4820) <= not((layer0_outputs(7450)) or (layer0_outputs(708)));
    layer1_outputs(4821) <= not(layer0_outputs(9239));
    layer1_outputs(4822) <= (layer0_outputs(5416)) xor (layer0_outputs(5684));
    layer1_outputs(4823) <= not(layer0_outputs(5862));
    layer1_outputs(4824) <= (layer0_outputs(394)) and (layer0_outputs(2456));
    layer1_outputs(4825) <= not(layer0_outputs(195));
    layer1_outputs(4826) <= (layer0_outputs(10209)) or (layer0_outputs(3650));
    layer1_outputs(4827) <= not((layer0_outputs(3524)) or (layer0_outputs(6299)));
    layer1_outputs(4828) <= not((layer0_outputs(9500)) and (layer0_outputs(3211)));
    layer1_outputs(4829) <= layer0_outputs(8194);
    layer1_outputs(4830) <= '0';
    layer1_outputs(4831) <= not((layer0_outputs(6471)) xor (layer0_outputs(6504)));
    layer1_outputs(4832) <= layer0_outputs(918);
    layer1_outputs(4833) <= not((layer0_outputs(5432)) or (layer0_outputs(4640)));
    layer1_outputs(4834) <= (layer0_outputs(1831)) and not (layer0_outputs(4270));
    layer1_outputs(4835) <= (layer0_outputs(942)) and not (layer0_outputs(5414));
    layer1_outputs(4836) <= not(layer0_outputs(861));
    layer1_outputs(4837) <= not((layer0_outputs(901)) or (layer0_outputs(4317)));
    layer1_outputs(4838) <= not((layer0_outputs(8648)) or (layer0_outputs(2582)));
    layer1_outputs(4839) <= not(layer0_outputs(5343));
    layer1_outputs(4840) <= not(layer0_outputs(6902)) or (layer0_outputs(6029));
    layer1_outputs(4841) <= layer0_outputs(6397);
    layer1_outputs(4842) <= (layer0_outputs(9057)) and (layer0_outputs(846));
    layer1_outputs(4843) <= not((layer0_outputs(5970)) xor (layer0_outputs(7426)));
    layer1_outputs(4844) <= not((layer0_outputs(5776)) xor (layer0_outputs(6672)));
    layer1_outputs(4845) <= not(layer0_outputs(10035)) or (layer0_outputs(4847));
    layer1_outputs(4846) <= not(layer0_outputs(7987)) or (layer0_outputs(3225));
    layer1_outputs(4847) <= not(layer0_outputs(3965)) or (layer0_outputs(5561));
    layer1_outputs(4848) <= layer0_outputs(9192);
    layer1_outputs(4849) <= layer0_outputs(5620);
    layer1_outputs(4850) <= (layer0_outputs(2050)) and not (layer0_outputs(9807));
    layer1_outputs(4851) <= layer0_outputs(579);
    layer1_outputs(4852) <= '1';
    layer1_outputs(4853) <= layer0_outputs(960);
    layer1_outputs(4854) <= not(layer0_outputs(5528));
    layer1_outputs(4855) <= layer0_outputs(7956);
    layer1_outputs(4856) <= not(layer0_outputs(7030));
    layer1_outputs(4857) <= not((layer0_outputs(9941)) or (layer0_outputs(1679)));
    layer1_outputs(4858) <= layer0_outputs(2196);
    layer1_outputs(4859) <= not(layer0_outputs(1672)) or (layer0_outputs(4955));
    layer1_outputs(4860) <= '0';
    layer1_outputs(4861) <= layer0_outputs(7661);
    layer1_outputs(4862) <= not(layer0_outputs(372)) or (layer0_outputs(100));
    layer1_outputs(4863) <= (layer0_outputs(8689)) and not (layer0_outputs(9558));
    layer1_outputs(4864) <= layer0_outputs(5528);
    layer1_outputs(4865) <= (layer0_outputs(25)) or (layer0_outputs(2368));
    layer1_outputs(4866) <= (layer0_outputs(7106)) and not (layer0_outputs(7122));
    layer1_outputs(4867) <= layer0_outputs(9168);
    layer1_outputs(4868) <= not(layer0_outputs(6685));
    layer1_outputs(4869) <= not(layer0_outputs(2148)) or (layer0_outputs(8214));
    layer1_outputs(4870) <= not((layer0_outputs(5393)) and (layer0_outputs(5340)));
    layer1_outputs(4871) <= (layer0_outputs(6597)) and (layer0_outputs(6781));
    layer1_outputs(4872) <= (layer0_outputs(9091)) and not (layer0_outputs(9860));
    layer1_outputs(4873) <= layer0_outputs(2819);
    layer1_outputs(4874) <= not((layer0_outputs(5010)) and (layer0_outputs(10022)));
    layer1_outputs(4875) <= not(layer0_outputs(5588));
    layer1_outputs(4876) <= (layer0_outputs(1502)) or (layer0_outputs(341));
    layer1_outputs(4877) <= (layer0_outputs(5805)) and not (layer0_outputs(3388));
    layer1_outputs(4878) <= layer0_outputs(7185);
    layer1_outputs(4879) <= (layer0_outputs(687)) and not (layer0_outputs(855));
    layer1_outputs(4880) <= '0';
    layer1_outputs(4881) <= not((layer0_outputs(7076)) and (layer0_outputs(8381)));
    layer1_outputs(4882) <= not(layer0_outputs(857));
    layer1_outputs(4883) <= layer0_outputs(6964);
    layer1_outputs(4884) <= layer0_outputs(6715);
    layer1_outputs(4885) <= layer0_outputs(4011);
    layer1_outputs(4886) <= layer0_outputs(1485);
    layer1_outputs(4887) <= not(layer0_outputs(4830));
    layer1_outputs(4888) <= not(layer0_outputs(6795)) or (layer0_outputs(9070));
    layer1_outputs(4889) <= (layer0_outputs(10221)) and not (layer0_outputs(7411));
    layer1_outputs(4890) <= not((layer0_outputs(9372)) or (layer0_outputs(3523)));
    layer1_outputs(4891) <= layer0_outputs(5810);
    layer1_outputs(4892) <= not(layer0_outputs(2180)) or (layer0_outputs(4224));
    layer1_outputs(4893) <= layer0_outputs(1432);
    layer1_outputs(4894) <= layer0_outputs(7321);
    layer1_outputs(4895) <= (layer0_outputs(1104)) xor (layer0_outputs(3523));
    layer1_outputs(4896) <= layer0_outputs(926);
    layer1_outputs(4897) <= (layer0_outputs(5586)) and (layer0_outputs(4196));
    layer1_outputs(4898) <= layer0_outputs(9665);
    layer1_outputs(4899) <= not((layer0_outputs(3213)) or (layer0_outputs(1703)));
    layer1_outputs(4900) <= (layer0_outputs(7124)) or (layer0_outputs(9631));
    layer1_outputs(4901) <= '1';
    layer1_outputs(4902) <= layer0_outputs(601);
    layer1_outputs(4903) <= '1';
    layer1_outputs(4904) <= layer0_outputs(475);
    layer1_outputs(4905) <= layer0_outputs(9246);
    layer1_outputs(4906) <= (layer0_outputs(433)) and not (layer0_outputs(3811));
    layer1_outputs(4907) <= layer0_outputs(8218);
    layer1_outputs(4908) <= layer0_outputs(672);
    layer1_outputs(4909) <= layer0_outputs(3615);
    layer1_outputs(4910) <= not(layer0_outputs(7888));
    layer1_outputs(4911) <= not((layer0_outputs(4357)) or (layer0_outputs(4147)));
    layer1_outputs(4912) <= layer0_outputs(7993);
    layer1_outputs(4913) <= not(layer0_outputs(3481)) or (layer0_outputs(4924));
    layer1_outputs(4914) <= '1';
    layer1_outputs(4915) <= '1';
    layer1_outputs(4916) <= layer0_outputs(9268);
    layer1_outputs(4917) <= (layer0_outputs(5419)) and (layer0_outputs(6136));
    layer1_outputs(4918) <= layer0_outputs(6702);
    layer1_outputs(4919) <= (layer0_outputs(2112)) and not (layer0_outputs(1855));
    layer1_outputs(4920) <= (layer0_outputs(8805)) or (layer0_outputs(5194));
    layer1_outputs(4921) <= layer0_outputs(826);
    layer1_outputs(4922) <= layer0_outputs(1745);
    layer1_outputs(4923) <= not((layer0_outputs(9668)) or (layer0_outputs(4869)));
    layer1_outputs(4924) <= (layer0_outputs(8271)) or (layer0_outputs(4425));
    layer1_outputs(4925) <= '0';
    layer1_outputs(4926) <= not((layer0_outputs(2401)) and (layer0_outputs(4815)));
    layer1_outputs(4927) <= not(layer0_outputs(9599));
    layer1_outputs(4928) <= not(layer0_outputs(7246)) or (layer0_outputs(1787));
    layer1_outputs(4929) <= not((layer0_outputs(2179)) or (layer0_outputs(9158)));
    layer1_outputs(4930) <= not((layer0_outputs(236)) or (layer0_outputs(8074)));
    layer1_outputs(4931) <= (layer0_outputs(9916)) and not (layer0_outputs(307));
    layer1_outputs(4932) <= not(layer0_outputs(8563));
    layer1_outputs(4933) <= (layer0_outputs(5750)) and not (layer0_outputs(5236));
    layer1_outputs(4934) <= (layer0_outputs(5212)) and not (layer0_outputs(2289));
    layer1_outputs(4935) <= layer0_outputs(1871);
    layer1_outputs(4936) <= layer0_outputs(5650);
    layer1_outputs(4937) <= not(layer0_outputs(4997));
    layer1_outputs(4938) <= not(layer0_outputs(7792));
    layer1_outputs(4939) <= not(layer0_outputs(3545));
    layer1_outputs(4940) <= not(layer0_outputs(7608));
    layer1_outputs(4941) <= (layer0_outputs(6707)) and not (layer0_outputs(6411));
    layer1_outputs(4942) <= not(layer0_outputs(2024));
    layer1_outputs(4943) <= not((layer0_outputs(7298)) and (layer0_outputs(8100)));
    layer1_outputs(4944) <= (layer0_outputs(3226)) and (layer0_outputs(3060));
    layer1_outputs(4945) <= layer0_outputs(8979);
    layer1_outputs(4946) <= (layer0_outputs(8454)) xor (layer0_outputs(9062));
    layer1_outputs(4947) <= layer0_outputs(7337);
    layer1_outputs(4948) <= layer0_outputs(9519);
    layer1_outputs(4949) <= not((layer0_outputs(2961)) or (layer0_outputs(1142)));
    layer1_outputs(4950) <= not(layer0_outputs(3050));
    layer1_outputs(4951) <= not(layer0_outputs(5215));
    layer1_outputs(4952) <= '1';
    layer1_outputs(4953) <= not(layer0_outputs(1201));
    layer1_outputs(4954) <= (layer0_outputs(6686)) xor (layer0_outputs(5431));
    layer1_outputs(4955) <= layer0_outputs(3432);
    layer1_outputs(4956) <= (layer0_outputs(6731)) and not (layer0_outputs(1609));
    layer1_outputs(4957) <= not(layer0_outputs(1477));
    layer1_outputs(4958) <= layer0_outputs(3016);
    layer1_outputs(4959) <= (layer0_outputs(662)) and not (layer0_outputs(9245));
    layer1_outputs(4960) <= layer0_outputs(2203);
    layer1_outputs(4961) <= '0';
    layer1_outputs(4962) <= not(layer0_outputs(5876));
    layer1_outputs(4963) <= not(layer0_outputs(4138)) or (layer0_outputs(8435));
    layer1_outputs(4964) <= not(layer0_outputs(2286));
    layer1_outputs(4965) <= layer0_outputs(8810);
    layer1_outputs(4966) <= (layer0_outputs(3168)) and (layer0_outputs(7730));
    layer1_outputs(4967) <= not(layer0_outputs(7820));
    layer1_outputs(4968) <= not(layer0_outputs(6442));
    layer1_outputs(4969) <= not(layer0_outputs(2189));
    layer1_outputs(4970) <= not(layer0_outputs(2847));
    layer1_outputs(4971) <= not(layer0_outputs(8889));
    layer1_outputs(4972) <= not((layer0_outputs(3869)) xor (layer0_outputs(2058)));
    layer1_outputs(4973) <= not((layer0_outputs(115)) and (layer0_outputs(5144)));
    layer1_outputs(4974) <= not((layer0_outputs(5915)) xor (layer0_outputs(8038)));
    layer1_outputs(4975) <= layer0_outputs(6416);
    layer1_outputs(4976) <= not(layer0_outputs(2960));
    layer1_outputs(4977) <= (layer0_outputs(3642)) xor (layer0_outputs(388));
    layer1_outputs(4978) <= layer0_outputs(9792);
    layer1_outputs(4979) <= (layer0_outputs(8495)) and not (layer0_outputs(5108));
    layer1_outputs(4980) <= not(layer0_outputs(5453)) or (layer0_outputs(430));
    layer1_outputs(4981) <= (layer0_outputs(7408)) and not (layer0_outputs(4149));
    layer1_outputs(4982) <= not(layer0_outputs(6422));
    layer1_outputs(4983) <= not(layer0_outputs(4007)) or (layer0_outputs(8853));
    layer1_outputs(4984) <= not((layer0_outputs(4026)) or (layer0_outputs(2634)));
    layer1_outputs(4985) <= not((layer0_outputs(6656)) xor (layer0_outputs(10210)));
    layer1_outputs(4986) <= not(layer0_outputs(2981)) or (layer0_outputs(784));
    layer1_outputs(4987) <= not((layer0_outputs(395)) xor (layer0_outputs(6297)));
    layer1_outputs(4988) <= layer0_outputs(9533);
    layer1_outputs(4989) <= not(layer0_outputs(198));
    layer1_outputs(4990) <= layer0_outputs(7132);
    layer1_outputs(4991) <= (layer0_outputs(3080)) and (layer0_outputs(2255));
    layer1_outputs(4992) <= not(layer0_outputs(5580));
    layer1_outputs(4993) <= not(layer0_outputs(3743));
    layer1_outputs(4994) <= '1';
    layer1_outputs(4995) <= '1';
    layer1_outputs(4996) <= (layer0_outputs(6364)) and (layer0_outputs(9058));
    layer1_outputs(4997) <= not((layer0_outputs(2640)) or (layer0_outputs(1037)));
    layer1_outputs(4998) <= not(layer0_outputs(1594)) or (layer0_outputs(330));
    layer1_outputs(4999) <= (layer0_outputs(7320)) and not (layer0_outputs(1351));
    layer1_outputs(5000) <= (layer0_outputs(1864)) and (layer0_outputs(7481));
    layer1_outputs(5001) <= not((layer0_outputs(7538)) and (layer0_outputs(7959)));
    layer1_outputs(5002) <= (layer0_outputs(3673)) or (layer0_outputs(7891));
    layer1_outputs(5003) <= (layer0_outputs(3939)) and (layer0_outputs(3539));
    layer1_outputs(5004) <= not(layer0_outputs(5998));
    layer1_outputs(5005) <= not(layer0_outputs(626)) or (layer0_outputs(9253));
    layer1_outputs(5006) <= layer0_outputs(5064);
    layer1_outputs(5007) <= layer0_outputs(4422);
    layer1_outputs(5008) <= (layer0_outputs(8598)) xor (layer0_outputs(7281));
    layer1_outputs(5009) <= not(layer0_outputs(7343));
    layer1_outputs(5010) <= (layer0_outputs(5352)) and not (layer0_outputs(6144));
    layer1_outputs(5011) <= not((layer0_outputs(983)) xor (layer0_outputs(1994)));
    layer1_outputs(5012) <= not(layer0_outputs(9309)) or (layer0_outputs(3973));
    layer1_outputs(5013) <= not((layer0_outputs(3187)) or (layer0_outputs(267)));
    layer1_outputs(5014) <= (layer0_outputs(5400)) or (layer0_outputs(6636));
    layer1_outputs(5015) <= not((layer0_outputs(678)) or (layer0_outputs(7357)));
    layer1_outputs(5016) <= not((layer0_outputs(9506)) or (layer0_outputs(2105)));
    layer1_outputs(5017) <= layer0_outputs(3578);
    layer1_outputs(5018) <= (layer0_outputs(6412)) and (layer0_outputs(4585));
    layer1_outputs(5019) <= (layer0_outputs(8410)) or (layer0_outputs(3618));
    layer1_outputs(5020) <= not(layer0_outputs(2313)) or (layer0_outputs(4958));
    layer1_outputs(5021) <= (layer0_outputs(8683)) and (layer0_outputs(134));
    layer1_outputs(5022) <= layer0_outputs(4546);
    layer1_outputs(5023) <= not(layer0_outputs(7505));
    layer1_outputs(5024) <= (layer0_outputs(6228)) and not (layer0_outputs(2273));
    layer1_outputs(5025) <= (layer0_outputs(2803)) or (layer0_outputs(746));
    layer1_outputs(5026) <= not(layer0_outputs(9818)) or (layer0_outputs(9789));
    layer1_outputs(5027) <= (layer0_outputs(6357)) and not (layer0_outputs(9427));
    layer1_outputs(5028) <= layer0_outputs(8442);
    layer1_outputs(5029) <= layer0_outputs(1491);
    layer1_outputs(5030) <= not(layer0_outputs(8723));
    layer1_outputs(5031) <= layer0_outputs(3097);
    layer1_outputs(5032) <= layer0_outputs(7123);
    layer1_outputs(5033) <= layer0_outputs(900);
    layer1_outputs(5034) <= layer0_outputs(8968);
    layer1_outputs(5035) <= not(layer0_outputs(9803));
    layer1_outputs(5036) <= not(layer0_outputs(10074)) or (layer0_outputs(4418));
    layer1_outputs(5037) <= not(layer0_outputs(1466));
    layer1_outputs(5038) <= not(layer0_outputs(8809)) or (layer0_outputs(3759));
    layer1_outputs(5039) <= (layer0_outputs(4846)) xor (layer0_outputs(10141));
    layer1_outputs(5040) <= layer0_outputs(4327);
    layer1_outputs(5041) <= not(layer0_outputs(9248));
    layer1_outputs(5042) <= (layer0_outputs(2355)) and not (layer0_outputs(691));
    layer1_outputs(5043) <= layer0_outputs(8383);
    layer1_outputs(5044) <= (layer0_outputs(3517)) and not (layer0_outputs(7920));
    layer1_outputs(5045) <= not((layer0_outputs(6141)) or (layer0_outputs(3431)));
    layer1_outputs(5046) <= (layer0_outputs(3127)) and not (layer0_outputs(1676));
    layer1_outputs(5047) <= layer0_outputs(6536);
    layer1_outputs(5048) <= not(layer0_outputs(8638)) or (layer0_outputs(4545));
    layer1_outputs(5049) <= layer0_outputs(5365);
    layer1_outputs(5050) <= layer0_outputs(7349);
    layer1_outputs(5051) <= '0';
    layer1_outputs(5052) <= not(layer0_outputs(7434));
    layer1_outputs(5053) <= '1';
    layer1_outputs(5054) <= layer0_outputs(4420);
    layer1_outputs(5055) <= '1';
    layer1_outputs(5056) <= '0';
    layer1_outputs(5057) <= layer0_outputs(8154);
    layer1_outputs(5058) <= (layer0_outputs(1684)) and not (layer0_outputs(9267));
    layer1_outputs(5059) <= (layer0_outputs(10203)) and (layer0_outputs(5555));
    layer1_outputs(5060) <= (layer0_outputs(809)) and not (layer0_outputs(4009));
    layer1_outputs(5061) <= not(layer0_outputs(977)) or (layer0_outputs(11));
    layer1_outputs(5062) <= not((layer0_outputs(1218)) or (layer0_outputs(856)));
    layer1_outputs(5063) <= not(layer0_outputs(490));
    layer1_outputs(5064) <= layer0_outputs(5374);
    layer1_outputs(5065) <= not((layer0_outputs(7807)) and (layer0_outputs(8016)));
    layer1_outputs(5066) <= (layer0_outputs(7055)) and not (layer0_outputs(6657));
    layer1_outputs(5067) <= not(layer0_outputs(3710)) or (layer0_outputs(1005));
    layer1_outputs(5068) <= (layer0_outputs(5011)) and not (layer0_outputs(2386));
    layer1_outputs(5069) <= '0';
    layer1_outputs(5070) <= layer0_outputs(7581);
    layer1_outputs(5071) <= not(layer0_outputs(7862));
    layer1_outputs(5072) <= not((layer0_outputs(9099)) or (layer0_outputs(4767)));
    layer1_outputs(5073) <= not(layer0_outputs(6421));
    layer1_outputs(5074) <= (layer0_outputs(2633)) or (layer0_outputs(2934));
    layer1_outputs(5075) <= (layer0_outputs(4854)) and (layer0_outputs(4859));
    layer1_outputs(5076) <= layer0_outputs(1830);
    layer1_outputs(5077) <= not(layer0_outputs(8871)) or (layer0_outputs(1925));
    layer1_outputs(5078) <= (layer0_outputs(8072)) and not (layer0_outputs(2950));
    layer1_outputs(5079) <= not((layer0_outputs(3008)) xor (layer0_outputs(9238)));
    layer1_outputs(5080) <= (layer0_outputs(7541)) and not (layer0_outputs(7480));
    layer1_outputs(5081) <= (layer0_outputs(1953)) and (layer0_outputs(9781));
    layer1_outputs(5082) <= not(layer0_outputs(10229));
    layer1_outputs(5083) <= not(layer0_outputs(1980)) or (layer0_outputs(2370));
    layer1_outputs(5084) <= not((layer0_outputs(7776)) or (layer0_outputs(9172)));
    layer1_outputs(5085) <= not((layer0_outputs(1294)) xor (layer0_outputs(6832)));
    layer1_outputs(5086) <= '1';
    layer1_outputs(5087) <= not(layer0_outputs(6763)) or (layer0_outputs(5012));
    layer1_outputs(5088) <= not((layer0_outputs(7085)) and (layer0_outputs(148)));
    layer1_outputs(5089) <= layer0_outputs(6811);
    layer1_outputs(5090) <= not((layer0_outputs(6211)) or (layer0_outputs(10130)));
    layer1_outputs(5091) <= not(layer0_outputs(10183));
    layer1_outputs(5092) <= layer0_outputs(1266);
    layer1_outputs(5093) <= not(layer0_outputs(3024));
    layer1_outputs(5094) <= '0';
    layer1_outputs(5095) <= (layer0_outputs(9539)) xor (layer0_outputs(2807));
    layer1_outputs(5096) <= not(layer0_outputs(5066));
    layer1_outputs(5097) <= (layer0_outputs(7513)) or (layer0_outputs(2899));
    layer1_outputs(5098) <= not(layer0_outputs(8708));
    layer1_outputs(5099) <= (layer0_outputs(1124)) and not (layer0_outputs(5198));
    layer1_outputs(5100) <= not(layer0_outputs(1590));
    layer1_outputs(5101) <= layer0_outputs(2364);
    layer1_outputs(5102) <= (layer0_outputs(9849)) and (layer0_outputs(10002));
    layer1_outputs(5103) <= layer0_outputs(4013);
    layer1_outputs(5104) <= layer0_outputs(7257);
    layer1_outputs(5105) <= layer0_outputs(3828);
    layer1_outputs(5106) <= (layer0_outputs(8886)) and (layer0_outputs(2198));
    layer1_outputs(5107) <= not((layer0_outputs(2487)) or (layer0_outputs(364)));
    layer1_outputs(5108) <= layer0_outputs(8914);
    layer1_outputs(5109) <= (layer0_outputs(3975)) xor (layer0_outputs(8478));
    layer1_outputs(5110) <= layer0_outputs(7296);
    layer1_outputs(5111) <= (layer0_outputs(9593)) and not (layer0_outputs(4312));
    layer1_outputs(5112) <= not(layer0_outputs(2904)) or (layer0_outputs(3732));
    layer1_outputs(5113) <= layer0_outputs(7454);
    layer1_outputs(5114) <= (layer0_outputs(4187)) or (layer0_outputs(3053));
    layer1_outputs(5115) <= not((layer0_outputs(3261)) or (layer0_outputs(10116)));
    layer1_outputs(5116) <= layer0_outputs(9002);
    layer1_outputs(5117) <= not((layer0_outputs(4521)) or (layer0_outputs(7503)));
    layer1_outputs(5118) <= not((layer0_outputs(2017)) and (layer0_outputs(3150)));
    layer1_outputs(5119) <= (layer0_outputs(2600)) xor (layer0_outputs(3558));
    layer1_outputs(5120) <= not((layer0_outputs(9930)) and (layer0_outputs(4090)));
    layer1_outputs(5121) <= not((layer0_outputs(9929)) xor (layer0_outputs(5180)));
    layer1_outputs(5122) <= not(layer0_outputs(1602)) or (layer0_outputs(877));
    layer1_outputs(5123) <= not((layer0_outputs(820)) or (layer0_outputs(1071)));
    layer1_outputs(5124) <= layer0_outputs(5538);
    layer1_outputs(5125) <= (layer0_outputs(271)) and not (layer0_outputs(1340));
    layer1_outputs(5126) <= layer0_outputs(4605);
    layer1_outputs(5127) <= not(layer0_outputs(3864));
    layer1_outputs(5128) <= (layer0_outputs(4136)) and (layer0_outputs(262));
    layer1_outputs(5129) <= not(layer0_outputs(7805)) or (layer0_outputs(4838));
    layer1_outputs(5130) <= not(layer0_outputs(7070)) or (layer0_outputs(631));
    layer1_outputs(5131) <= layer0_outputs(4441);
    layer1_outputs(5132) <= not(layer0_outputs(9074));
    layer1_outputs(5133) <= not(layer0_outputs(2878));
    layer1_outputs(5134) <= (layer0_outputs(3633)) or (layer0_outputs(6486));
    layer1_outputs(5135) <= (layer0_outputs(507)) and not (layer0_outputs(4726));
    layer1_outputs(5136) <= layer0_outputs(4016);
    layer1_outputs(5137) <= (layer0_outputs(593)) and not (layer0_outputs(5697));
    layer1_outputs(5138) <= layer0_outputs(2864);
    layer1_outputs(5139) <= not((layer0_outputs(6492)) xor (layer0_outputs(807)));
    layer1_outputs(5140) <= (layer0_outputs(9025)) and not (layer0_outputs(325));
    layer1_outputs(5141) <= not((layer0_outputs(6975)) or (layer0_outputs(1511)));
    layer1_outputs(5142) <= (layer0_outputs(1519)) and not (layer0_outputs(1346));
    layer1_outputs(5143) <= layer0_outputs(1185);
    layer1_outputs(5144) <= not((layer0_outputs(9042)) and (layer0_outputs(1548)));
    layer1_outputs(5145) <= (layer0_outputs(8491)) and not (layer0_outputs(5593));
    layer1_outputs(5146) <= not(layer0_outputs(8683));
    layer1_outputs(5147) <= (layer0_outputs(239)) or (layer0_outputs(2981));
    layer1_outputs(5148) <= not((layer0_outputs(7631)) xor (layer0_outputs(9971)));
    layer1_outputs(5149) <= (layer0_outputs(4850)) xor (layer0_outputs(10111));
    layer1_outputs(5150) <= (layer0_outputs(7972)) and not (layer0_outputs(7351));
    layer1_outputs(5151) <= not((layer0_outputs(7950)) or (layer0_outputs(6496)));
    layer1_outputs(5152) <= not(layer0_outputs(4098));
    layer1_outputs(5153) <= not(layer0_outputs(710)) or (layer0_outputs(6178));
    layer1_outputs(5154) <= not(layer0_outputs(9363));
    layer1_outputs(5155) <= not(layer0_outputs(10033)) or (layer0_outputs(591));
    layer1_outputs(5156) <= layer0_outputs(1395);
    layer1_outputs(5157) <= (layer0_outputs(3294)) and (layer0_outputs(4389));
    layer1_outputs(5158) <= (layer0_outputs(8)) and (layer0_outputs(5565));
    layer1_outputs(5159) <= not(layer0_outputs(3552)) or (layer0_outputs(6880));
    layer1_outputs(5160) <= (layer0_outputs(9795)) or (layer0_outputs(1713));
    layer1_outputs(5161) <= (layer0_outputs(3401)) xor (layer0_outputs(2874));
    layer1_outputs(5162) <= not((layer0_outputs(7174)) and (layer0_outputs(9934)));
    layer1_outputs(5163) <= layer0_outputs(2857);
    layer1_outputs(5164) <= (layer0_outputs(5124)) and not (layer0_outputs(7865));
    layer1_outputs(5165) <= layer0_outputs(1060);
    layer1_outputs(5166) <= not((layer0_outputs(4299)) and (layer0_outputs(2571)));
    layer1_outputs(5167) <= (layer0_outputs(10070)) xor (layer0_outputs(2761));
    layer1_outputs(5168) <= not(layer0_outputs(4403));
    layer1_outputs(5169) <= (layer0_outputs(6732)) and not (layer0_outputs(6653));
    layer1_outputs(5170) <= not(layer0_outputs(9658));
    layer1_outputs(5171) <= not((layer0_outputs(973)) and (layer0_outputs(4977)));
    layer1_outputs(5172) <= (layer0_outputs(8214)) xor (layer0_outputs(3236));
    layer1_outputs(5173) <= (layer0_outputs(7083)) and not (layer0_outputs(3938));
    layer1_outputs(5174) <= layer0_outputs(996);
    layer1_outputs(5175) <= not(layer0_outputs(7066));
    layer1_outputs(5176) <= (layer0_outputs(1827)) and not (layer0_outputs(7145));
    layer1_outputs(5177) <= layer0_outputs(3359);
    layer1_outputs(5178) <= layer0_outputs(5287);
    layer1_outputs(5179) <= not(layer0_outputs(1534)) or (layer0_outputs(2785));
    layer1_outputs(5180) <= layer0_outputs(9530);
    layer1_outputs(5181) <= (layer0_outputs(1562)) and not (layer0_outputs(6323));
    layer1_outputs(5182) <= (layer0_outputs(7680)) or (layer0_outputs(1870));
    layer1_outputs(5183) <= not(layer0_outputs(2629)) or (layer0_outputs(6625));
    layer1_outputs(5184) <= '1';
    layer1_outputs(5185) <= layer0_outputs(8605);
    layer1_outputs(5186) <= '0';
    layer1_outputs(5187) <= not(layer0_outputs(10235));
    layer1_outputs(5188) <= layer0_outputs(8944);
    layer1_outputs(5189) <= layer0_outputs(2542);
    layer1_outputs(5190) <= (layer0_outputs(413)) or (layer0_outputs(1951));
    layer1_outputs(5191) <= not((layer0_outputs(4842)) or (layer0_outputs(3389)));
    layer1_outputs(5192) <= not(layer0_outputs(5148)) or (layer0_outputs(5174));
    layer1_outputs(5193) <= not((layer0_outputs(1101)) xor (layer0_outputs(3219)));
    layer1_outputs(5194) <= (layer0_outputs(7704)) and (layer0_outputs(3456));
    layer1_outputs(5195) <= not(layer0_outputs(1636));
    layer1_outputs(5196) <= layer0_outputs(3184);
    layer1_outputs(5197) <= '1';
    layer1_outputs(5198) <= not(layer0_outputs(6420)) or (layer0_outputs(1345));
    layer1_outputs(5199) <= (layer0_outputs(6550)) and not (layer0_outputs(5936));
    layer1_outputs(5200) <= not(layer0_outputs(2841));
    layer1_outputs(5201) <= not(layer0_outputs(2181));
    layer1_outputs(5202) <= (layer0_outputs(10238)) xor (layer0_outputs(5072));
    layer1_outputs(5203) <= not(layer0_outputs(6336)) or (layer0_outputs(3314));
    layer1_outputs(5204) <= not(layer0_outputs(2414));
    layer1_outputs(5205) <= not((layer0_outputs(9965)) and (layer0_outputs(5768)));
    layer1_outputs(5206) <= not((layer0_outputs(3083)) xor (layer0_outputs(6852)));
    layer1_outputs(5207) <= not(layer0_outputs(4319));
    layer1_outputs(5208) <= not(layer0_outputs(5815));
    layer1_outputs(5209) <= (layer0_outputs(9292)) or (layer0_outputs(5655));
    layer1_outputs(5210) <= layer0_outputs(4417);
    layer1_outputs(5211) <= layer0_outputs(812);
    layer1_outputs(5212) <= not(layer0_outputs(7387));
    layer1_outputs(5213) <= not(layer0_outputs(8980));
    layer1_outputs(5214) <= not(layer0_outputs(4498));
    layer1_outputs(5215) <= layer0_outputs(4291);
    layer1_outputs(5216) <= layer0_outputs(7588);
    layer1_outputs(5217) <= (layer0_outputs(5517)) and not (layer0_outputs(1730));
    layer1_outputs(5218) <= layer0_outputs(10039);
    layer1_outputs(5219) <= (layer0_outputs(8600)) and not (layer0_outputs(9612));
    layer1_outputs(5220) <= not(layer0_outputs(1097));
    layer1_outputs(5221) <= not(layer0_outputs(9211));
    layer1_outputs(5222) <= not((layer0_outputs(7680)) or (layer0_outputs(6891)));
    layer1_outputs(5223) <= (layer0_outputs(9598)) and not (layer0_outputs(5653));
    layer1_outputs(5224) <= (layer0_outputs(3671)) or (layer0_outputs(1664));
    layer1_outputs(5225) <= not(layer0_outputs(885));
    layer1_outputs(5226) <= layer0_outputs(8569);
    layer1_outputs(5227) <= not(layer0_outputs(8840)) or (layer0_outputs(2229));
    layer1_outputs(5228) <= not(layer0_outputs(1047));
    layer1_outputs(5229) <= not((layer0_outputs(7775)) or (layer0_outputs(6979)));
    layer1_outputs(5230) <= (layer0_outputs(421)) or (layer0_outputs(6038));
    layer1_outputs(5231) <= not(layer0_outputs(3649));
    layer1_outputs(5232) <= not(layer0_outputs(3554)) or (layer0_outputs(6981));
    layer1_outputs(5233) <= not(layer0_outputs(9467));
    layer1_outputs(5234) <= not(layer0_outputs(2168)) or (layer0_outputs(8652));
    layer1_outputs(5235) <= not(layer0_outputs(7738)) or (layer0_outputs(699));
    layer1_outputs(5236) <= layer0_outputs(2351);
    layer1_outputs(5237) <= not(layer0_outputs(7190)) or (layer0_outputs(1444));
    layer1_outputs(5238) <= layer0_outputs(170);
    layer1_outputs(5239) <= not(layer0_outputs(7018)) or (layer0_outputs(9620));
    layer1_outputs(5240) <= (layer0_outputs(5369)) and (layer0_outputs(4491));
    layer1_outputs(5241) <= not(layer0_outputs(8920));
    layer1_outputs(5242) <= (layer0_outputs(6281)) and not (layer0_outputs(6234));
    layer1_outputs(5243) <= (layer0_outputs(405)) xor (layer0_outputs(3295));
    layer1_outputs(5244) <= '1';
    layer1_outputs(5245) <= layer0_outputs(4075);
    layer1_outputs(5246) <= not(layer0_outputs(4701)) or (layer0_outputs(1607));
    layer1_outputs(5247) <= not((layer0_outputs(1534)) or (layer0_outputs(902)));
    layer1_outputs(5248) <= layer0_outputs(8303);
    layer1_outputs(5249) <= (layer0_outputs(3300)) and not (layer0_outputs(3752));
    layer1_outputs(5250) <= layer0_outputs(3662);
    layer1_outputs(5251) <= layer0_outputs(7827);
    layer1_outputs(5252) <= (layer0_outputs(666)) xor (layer0_outputs(6297));
    layer1_outputs(5253) <= not(layer0_outputs(602));
    layer1_outputs(5254) <= '1';
    layer1_outputs(5255) <= not(layer0_outputs(8082));
    layer1_outputs(5256) <= not(layer0_outputs(5558));
    layer1_outputs(5257) <= not(layer0_outputs(6446));
    layer1_outputs(5258) <= not(layer0_outputs(6954));
    layer1_outputs(5259) <= layer0_outputs(5506);
    layer1_outputs(5260) <= not(layer0_outputs(3413));
    layer1_outputs(5261) <= not(layer0_outputs(3245));
    layer1_outputs(5262) <= not(layer0_outputs(2567));
    layer1_outputs(5263) <= '0';
    layer1_outputs(5264) <= not(layer0_outputs(6766)) or (layer0_outputs(8539));
    layer1_outputs(5265) <= (layer0_outputs(6138)) and not (layer0_outputs(9026));
    layer1_outputs(5266) <= not(layer0_outputs(9789)) or (layer0_outputs(9054));
    layer1_outputs(5267) <= not((layer0_outputs(799)) and (layer0_outputs(6878)));
    layer1_outputs(5268) <= not(layer0_outputs(8289));
    layer1_outputs(5269) <= layer0_outputs(2797);
    layer1_outputs(5270) <= not(layer0_outputs(5896));
    layer1_outputs(5271) <= not(layer0_outputs(1765));
    layer1_outputs(5272) <= not(layer0_outputs(1004));
    layer1_outputs(5273) <= not(layer0_outputs(9083));
    layer1_outputs(5274) <= not(layer0_outputs(9883));
    layer1_outputs(5275) <= (layer0_outputs(5464)) and (layer0_outputs(1050));
    layer1_outputs(5276) <= (layer0_outputs(4771)) and not (layer0_outputs(8291));
    layer1_outputs(5277) <= (layer0_outputs(6295)) and not (layer0_outputs(8118));
    layer1_outputs(5278) <= (layer0_outputs(2658)) and not (layer0_outputs(468));
    layer1_outputs(5279) <= (layer0_outputs(6334)) xor (layer0_outputs(8018));
    layer1_outputs(5280) <= layer0_outputs(5255);
    layer1_outputs(5281) <= '0';
    layer1_outputs(5282) <= not(layer0_outputs(6755));
    layer1_outputs(5283) <= not(layer0_outputs(3714)) or (layer0_outputs(9114));
    layer1_outputs(5284) <= (layer0_outputs(3577)) and (layer0_outputs(9992));
    layer1_outputs(5285) <= layer0_outputs(2036);
    layer1_outputs(5286) <= not((layer0_outputs(5837)) or (layer0_outputs(7621)));
    layer1_outputs(5287) <= not(layer0_outputs(7882));
    layer1_outputs(5288) <= not(layer0_outputs(3438));
    layer1_outputs(5289) <= (layer0_outputs(9328)) and not (layer0_outputs(6709));
    layer1_outputs(5290) <= layer0_outputs(760);
    layer1_outputs(5291) <= not((layer0_outputs(10129)) or (layer0_outputs(5410)));
    layer1_outputs(5292) <= not((layer0_outputs(8550)) or (layer0_outputs(6097)));
    layer1_outputs(5293) <= not(layer0_outputs(6628));
    layer1_outputs(5294) <= layer0_outputs(5139);
    layer1_outputs(5295) <= layer0_outputs(5117);
    layer1_outputs(5296) <= (layer0_outputs(6628)) and (layer0_outputs(3957));
    layer1_outputs(5297) <= (layer0_outputs(2543)) and not (layer0_outputs(9527));
    layer1_outputs(5298) <= not((layer0_outputs(3373)) and (layer0_outputs(10114)));
    layer1_outputs(5299) <= not(layer0_outputs(3631));
    layer1_outputs(5300) <= not(layer0_outputs(3341)) or (layer0_outputs(8966));
    layer1_outputs(5301) <= not(layer0_outputs(1966));
    layer1_outputs(5302) <= not((layer0_outputs(7338)) xor (layer0_outputs(6924)));
    layer1_outputs(5303) <= (layer0_outputs(3856)) or (layer0_outputs(4198));
    layer1_outputs(5304) <= not(layer0_outputs(7406));
    layer1_outputs(5305) <= not(layer0_outputs(4489)) or (layer0_outputs(8587));
    layer1_outputs(5306) <= not((layer0_outputs(8437)) xor (layer0_outputs(3921)));
    layer1_outputs(5307) <= not((layer0_outputs(564)) xor (layer0_outputs(8693)));
    layer1_outputs(5308) <= layer0_outputs(4358);
    layer1_outputs(5309) <= (layer0_outputs(9546)) and not (layer0_outputs(8224));
    layer1_outputs(5310) <= layer0_outputs(3941);
    layer1_outputs(5311) <= (layer0_outputs(6585)) and not (layer0_outputs(9494));
    layer1_outputs(5312) <= not(layer0_outputs(6703));
    layer1_outputs(5313) <= (layer0_outputs(3164)) or (layer0_outputs(7651));
    layer1_outputs(5314) <= not((layer0_outputs(8641)) xor (layer0_outputs(4911)));
    layer1_outputs(5315) <= (layer0_outputs(6031)) and not (layer0_outputs(8890));
    layer1_outputs(5316) <= not((layer0_outputs(3362)) and (layer0_outputs(9277)));
    layer1_outputs(5317) <= (layer0_outputs(9074)) and (layer0_outputs(1399));
    layer1_outputs(5318) <= '0';
    layer1_outputs(5319) <= (layer0_outputs(4558)) or (layer0_outputs(1068));
    layer1_outputs(5320) <= not(layer0_outputs(4920));
    layer1_outputs(5321) <= (layer0_outputs(5435)) and (layer0_outputs(6725));
    layer1_outputs(5322) <= (layer0_outputs(7074)) and not (layer0_outputs(2450));
    layer1_outputs(5323) <= not(layer0_outputs(5532)) or (layer0_outputs(8061));
    layer1_outputs(5324) <= layer0_outputs(1297);
    layer1_outputs(5325) <= (layer0_outputs(3762)) and not (layer0_outputs(3042));
    layer1_outputs(5326) <= (layer0_outputs(6723)) xor (layer0_outputs(1929));
    layer1_outputs(5327) <= not(layer0_outputs(7532));
    layer1_outputs(5328) <= not(layer0_outputs(184)) or (layer0_outputs(3514));
    layer1_outputs(5329) <= not(layer0_outputs(4946));
    layer1_outputs(5330) <= layer0_outputs(1640);
    layer1_outputs(5331) <= not((layer0_outputs(2279)) and (layer0_outputs(1578)));
    layer1_outputs(5332) <= (layer0_outputs(1192)) and not (layer0_outputs(188));
    layer1_outputs(5333) <= (layer0_outputs(2179)) or (layer0_outputs(3955));
    layer1_outputs(5334) <= layer0_outputs(7912);
    layer1_outputs(5335) <= not(layer0_outputs(5542)) or (layer0_outputs(10014));
    layer1_outputs(5336) <= layer0_outputs(2767);
    layer1_outputs(5337) <= layer0_outputs(7528);
    layer1_outputs(5338) <= (layer0_outputs(8436)) and not (layer0_outputs(4586));
    layer1_outputs(5339) <= '1';
    layer1_outputs(5340) <= not(layer0_outputs(19));
    layer1_outputs(5341) <= not((layer0_outputs(2183)) or (layer0_outputs(767)));
    layer1_outputs(5342) <= not(layer0_outputs(1973));
    layer1_outputs(5343) <= not(layer0_outputs(2048)) or (layer0_outputs(7263));
    layer1_outputs(5344) <= layer0_outputs(7240);
    layer1_outputs(5345) <= not(layer0_outputs(860));
    layer1_outputs(5346) <= (layer0_outputs(1786)) and not (layer0_outputs(9673));
    layer1_outputs(5347) <= not(layer0_outputs(6589));
    layer1_outputs(5348) <= not(layer0_outputs(1617));
    layer1_outputs(5349) <= not((layer0_outputs(2415)) and (layer0_outputs(215)));
    layer1_outputs(5350) <= not(layer0_outputs(235));
    layer1_outputs(5351) <= not(layer0_outputs(7783)) or (layer0_outputs(1444));
    layer1_outputs(5352) <= (layer0_outputs(993)) or (layer0_outputs(7930));
    layer1_outputs(5353) <= '0';
    layer1_outputs(5354) <= not(layer0_outputs(9193));
    layer1_outputs(5355) <= not(layer0_outputs(1386));
    layer1_outputs(5356) <= layer0_outputs(5852);
    layer1_outputs(5357) <= (layer0_outputs(5261)) or (layer0_outputs(5636));
    layer1_outputs(5358) <= not(layer0_outputs(30));
    layer1_outputs(5359) <= not(layer0_outputs(1704));
    layer1_outputs(5360) <= not((layer0_outputs(8942)) or (layer0_outputs(145)));
    layer1_outputs(5361) <= not(layer0_outputs(7851)) or (layer0_outputs(3515));
    layer1_outputs(5362) <= layer0_outputs(9516);
    layer1_outputs(5363) <= not((layer0_outputs(2167)) xor (layer0_outputs(4250)));
    layer1_outputs(5364) <= not((layer0_outputs(7187)) and (layer0_outputs(7165)));
    layer1_outputs(5365) <= layer0_outputs(93);
    layer1_outputs(5366) <= (layer0_outputs(734)) or (layer0_outputs(4191));
    layer1_outputs(5367) <= not(layer0_outputs(5960));
    layer1_outputs(5368) <= layer0_outputs(5760);
    layer1_outputs(5369) <= not(layer0_outputs(4130)) or (layer0_outputs(1198));
    layer1_outputs(5370) <= not(layer0_outputs(777));
    layer1_outputs(5371) <= not(layer0_outputs(5009));
    layer1_outputs(5372) <= layer0_outputs(4232);
    layer1_outputs(5373) <= layer0_outputs(2772);
    layer1_outputs(5374) <= not((layer0_outputs(3214)) or (layer0_outputs(10178)));
    layer1_outputs(5375) <= layer0_outputs(8825);
    layer1_outputs(5376) <= (layer0_outputs(3998)) and (layer0_outputs(9845));
    layer1_outputs(5377) <= not((layer0_outputs(9719)) and (layer0_outputs(4264)));
    layer1_outputs(5378) <= not(layer0_outputs(4447));
    layer1_outputs(5379) <= (layer0_outputs(661)) or (layer0_outputs(4698));
    layer1_outputs(5380) <= '1';
    layer1_outputs(5381) <= (layer0_outputs(3975)) and (layer0_outputs(5331));
    layer1_outputs(5382) <= not((layer0_outputs(6470)) xor (layer0_outputs(7629)));
    layer1_outputs(5383) <= not(layer0_outputs(4957)) or (layer0_outputs(341));
    layer1_outputs(5384) <= (layer0_outputs(785)) and not (layer0_outputs(9153));
    layer1_outputs(5385) <= not((layer0_outputs(3562)) or (layer0_outputs(8117)));
    layer1_outputs(5386) <= layer0_outputs(5748);
    layer1_outputs(5387) <= not(layer0_outputs(1091));
    layer1_outputs(5388) <= not(layer0_outputs(1165)) or (layer0_outputs(3785));
    layer1_outputs(5389) <= layer0_outputs(2823);
    layer1_outputs(5390) <= not((layer0_outputs(2073)) and (layer0_outputs(9051)));
    layer1_outputs(5391) <= not((layer0_outputs(8849)) or (layer0_outputs(201)));
    layer1_outputs(5392) <= layer0_outputs(8596);
    layer1_outputs(5393) <= not(layer0_outputs(4114));
    layer1_outputs(5394) <= (layer0_outputs(7396)) and not (layer0_outputs(840));
    layer1_outputs(5395) <= not((layer0_outputs(7804)) or (layer0_outputs(5269)));
    layer1_outputs(5396) <= (layer0_outputs(9864)) and (layer0_outputs(915));
    layer1_outputs(5397) <= not((layer0_outputs(7707)) and (layer0_outputs(7489)));
    layer1_outputs(5398) <= (layer0_outputs(8740)) and (layer0_outputs(6911));
    layer1_outputs(5399) <= layer0_outputs(8664);
    layer1_outputs(5400) <= layer0_outputs(7047);
    layer1_outputs(5401) <= not((layer0_outputs(3236)) or (layer0_outputs(3280)));
    layer1_outputs(5402) <= '1';
    layer1_outputs(5403) <= (layer0_outputs(5442)) and not (layer0_outputs(6596));
    layer1_outputs(5404) <= (layer0_outputs(131)) and not (layer0_outputs(7785));
    layer1_outputs(5405) <= layer0_outputs(3314);
    layer1_outputs(5406) <= not((layer0_outputs(6942)) xor (layer0_outputs(5377)));
    layer1_outputs(5407) <= (layer0_outputs(2493)) and not (layer0_outputs(7903));
    layer1_outputs(5408) <= layer0_outputs(7721);
    layer1_outputs(5409) <= not(layer0_outputs(1323));
    layer1_outputs(5410) <= not(layer0_outputs(6506));
    layer1_outputs(5411) <= (layer0_outputs(9743)) and not (layer0_outputs(870));
    layer1_outputs(5412) <= layer0_outputs(7612);
    layer1_outputs(5413) <= not(layer0_outputs(9693)) or (layer0_outputs(10066));
    layer1_outputs(5414) <= (layer0_outputs(8677)) and (layer0_outputs(7878));
    layer1_outputs(5415) <= not((layer0_outputs(9559)) or (layer0_outputs(2871)));
    layer1_outputs(5416) <= layer0_outputs(8249);
    layer1_outputs(5417) <= not((layer0_outputs(269)) or (layer0_outputs(864)));
    layer1_outputs(5418) <= layer0_outputs(7584);
    layer1_outputs(5419) <= not(layer0_outputs(271)) or (layer0_outputs(7951));
    layer1_outputs(5420) <= not(layer0_outputs(4426)) or (layer0_outputs(4146));
    layer1_outputs(5421) <= not(layer0_outputs(9967));
    layer1_outputs(5422) <= not(layer0_outputs(9363));
    layer1_outputs(5423) <= not(layer0_outputs(5731));
    layer1_outputs(5424) <= not(layer0_outputs(5573)) or (layer0_outputs(3923));
    layer1_outputs(5425) <= not((layer0_outputs(1669)) and (layer0_outputs(612)));
    layer1_outputs(5426) <= not(layer0_outputs(4152)) or (layer0_outputs(3715));
    layer1_outputs(5427) <= not((layer0_outputs(6644)) or (layer0_outputs(8246)));
    layer1_outputs(5428) <= not(layer0_outputs(6681)) or (layer0_outputs(1641));
    layer1_outputs(5429) <= not(layer0_outputs(7593));
    layer1_outputs(5430) <= not(layer0_outputs(6569)) or (layer0_outputs(7738));
    layer1_outputs(5431) <= not((layer0_outputs(4122)) xor (layer0_outputs(3548)));
    layer1_outputs(5432) <= not(layer0_outputs(648)) or (layer0_outputs(2695));
    layer1_outputs(5433) <= (layer0_outputs(3326)) or (layer0_outputs(9523));
    layer1_outputs(5434) <= (layer0_outputs(9375)) or (layer0_outputs(7695));
    layer1_outputs(5435) <= '1';
    layer1_outputs(5436) <= (layer0_outputs(10023)) and not (layer0_outputs(1625));
    layer1_outputs(5437) <= (layer0_outputs(1149)) and not (layer0_outputs(7659));
    layer1_outputs(5438) <= layer0_outputs(6270);
    layer1_outputs(5439) <= not(layer0_outputs(2220));
    layer1_outputs(5440) <= '1';
    layer1_outputs(5441) <= not(layer0_outputs(432));
    layer1_outputs(5442) <= (layer0_outputs(3720)) and not (layer0_outputs(540));
    layer1_outputs(5443) <= not(layer0_outputs(2675));
    layer1_outputs(5444) <= not(layer0_outputs(8307));
    layer1_outputs(5445) <= not(layer0_outputs(4972));
    layer1_outputs(5446) <= not(layer0_outputs(6132));
    layer1_outputs(5447) <= not(layer0_outputs(2524)) or (layer0_outputs(5645));
    layer1_outputs(5448) <= layer0_outputs(6828);
    layer1_outputs(5449) <= not(layer0_outputs(4543));
    layer1_outputs(5450) <= not(layer0_outputs(7557));
    layer1_outputs(5451) <= layer0_outputs(5504);
    layer1_outputs(5452) <= layer0_outputs(2569);
    layer1_outputs(5453) <= (layer0_outputs(2416)) xor (layer0_outputs(9079));
    layer1_outputs(5454) <= layer0_outputs(6729);
    layer1_outputs(5455) <= layer0_outputs(4612);
    layer1_outputs(5456) <= not(layer0_outputs(10195));
    layer1_outputs(5457) <= (layer0_outputs(8197)) xor (layer0_outputs(8345));
    layer1_outputs(5458) <= not(layer0_outputs(491)) or (layer0_outputs(4995));
    layer1_outputs(5459) <= (layer0_outputs(6866)) and not (layer0_outputs(9225));
    layer1_outputs(5460) <= layer0_outputs(4216);
    layer1_outputs(5461) <= (layer0_outputs(1610)) and not (layer0_outputs(1773));
    layer1_outputs(5462) <= not(layer0_outputs(9316));
    layer1_outputs(5463) <= not((layer0_outputs(4725)) and (layer0_outputs(5183)));
    layer1_outputs(5464) <= (layer0_outputs(3417)) and not (layer0_outputs(3991));
    layer1_outputs(5465) <= layer0_outputs(1767);
    layer1_outputs(5466) <= (layer0_outputs(5874)) or (layer0_outputs(1384));
    layer1_outputs(5467) <= not(layer0_outputs(207));
    layer1_outputs(5468) <= not((layer0_outputs(848)) or (layer0_outputs(3909)));
    layer1_outputs(5469) <= not(layer0_outputs(7446)) or (layer0_outputs(9900));
    layer1_outputs(5470) <= not(layer0_outputs(6321));
    layer1_outputs(5471) <= not(layer0_outputs(6850));
    layer1_outputs(5472) <= (layer0_outputs(2362)) and not (layer0_outputs(4823));
    layer1_outputs(5473) <= not(layer0_outputs(8482));
    layer1_outputs(5474) <= layer0_outputs(4747);
    layer1_outputs(5475) <= not((layer0_outputs(7399)) xor (layer0_outputs(1065)));
    layer1_outputs(5476) <= (layer0_outputs(7144)) and (layer0_outputs(2122));
    layer1_outputs(5477) <= not(layer0_outputs(9836)) or (layer0_outputs(2533));
    layer1_outputs(5478) <= not(layer0_outputs(6250));
    layer1_outputs(5479) <= (layer0_outputs(7489)) xor (layer0_outputs(1914));
    layer1_outputs(5480) <= layer0_outputs(7635);
    layer1_outputs(5481) <= layer0_outputs(7838);
    layer1_outputs(5482) <= '0';
    layer1_outputs(5483) <= not((layer0_outputs(2027)) or (layer0_outputs(1617)));
    layer1_outputs(5484) <= '1';
    layer1_outputs(5485) <= layer0_outputs(4481);
    layer1_outputs(5486) <= (layer0_outputs(5748)) or (layer0_outputs(5690));
    layer1_outputs(5487) <= not(layer0_outputs(3123)) or (layer0_outputs(1648));
    layer1_outputs(5488) <= not((layer0_outputs(6007)) or (layer0_outputs(7867)));
    layer1_outputs(5489) <= not(layer0_outputs(3354)) or (layer0_outputs(3755));
    layer1_outputs(5490) <= '0';
    layer1_outputs(5491) <= (layer0_outputs(1421)) and (layer0_outputs(5447));
    layer1_outputs(5492) <= (layer0_outputs(2690)) and not (layer0_outputs(4633));
    layer1_outputs(5493) <= not(layer0_outputs(5204)) or (layer0_outputs(5220));
    layer1_outputs(5494) <= (layer0_outputs(6561)) or (layer0_outputs(9467));
    layer1_outputs(5495) <= layer0_outputs(6148);
    layer1_outputs(5496) <= not((layer0_outputs(6694)) or (layer0_outputs(8146)));
    layer1_outputs(5497) <= layer0_outputs(7032);
    layer1_outputs(5498) <= layer0_outputs(5085);
    layer1_outputs(5499) <= not((layer0_outputs(5637)) xor (layer0_outputs(2894)));
    layer1_outputs(5500) <= not((layer0_outputs(5923)) or (layer0_outputs(3716)));
    layer1_outputs(5501) <= (layer0_outputs(7826)) or (layer0_outputs(1642));
    layer1_outputs(5502) <= not(layer0_outputs(592));
    layer1_outputs(5503) <= not(layer0_outputs(90)) or (layer0_outputs(1096));
    layer1_outputs(5504) <= not((layer0_outputs(5441)) and (layer0_outputs(9424)));
    layer1_outputs(5505) <= (layer0_outputs(821)) and (layer0_outputs(9432));
    layer1_outputs(5506) <= not(layer0_outputs(4694));
    layer1_outputs(5507) <= layer0_outputs(191);
    layer1_outputs(5508) <= (layer0_outputs(1210)) and (layer0_outputs(3276));
    layer1_outputs(5509) <= not(layer0_outputs(7585)) or (layer0_outputs(1450));
    layer1_outputs(5510) <= layer0_outputs(768);
    layer1_outputs(5511) <= layer0_outputs(9761);
    layer1_outputs(5512) <= not((layer0_outputs(8298)) and (layer0_outputs(1727)));
    layer1_outputs(5513) <= not(layer0_outputs(9875));
    layer1_outputs(5514) <= layer0_outputs(3987);
    layer1_outputs(5515) <= not(layer0_outputs(7766));
    layer1_outputs(5516) <= not(layer0_outputs(7486)) or (layer0_outputs(1798));
    layer1_outputs(5517) <= layer0_outputs(3492);
    layer1_outputs(5518) <= not((layer0_outputs(8875)) and (layer0_outputs(6824)));
    layer1_outputs(5519) <= (layer0_outputs(8641)) and (layer0_outputs(4899));
    layer1_outputs(5520) <= not(layer0_outputs(8632)) or (layer0_outputs(6471));
    layer1_outputs(5521) <= layer0_outputs(3089);
    layer1_outputs(5522) <= (layer0_outputs(6880)) and (layer0_outputs(3660));
    layer1_outputs(5523) <= not((layer0_outputs(4133)) and (layer0_outputs(9048)));
    layer1_outputs(5524) <= (layer0_outputs(5433)) or (layer0_outputs(5691));
    layer1_outputs(5525) <= (layer0_outputs(86)) and not (layer0_outputs(595));
    layer1_outputs(5526) <= not((layer0_outputs(5834)) and (layer0_outputs(2348)));
    layer1_outputs(5527) <= (layer0_outputs(4466)) or (layer0_outputs(4864));
    layer1_outputs(5528) <= not(layer0_outputs(2520));
    layer1_outputs(5529) <= (layer0_outputs(7376)) and not (layer0_outputs(3170));
    layer1_outputs(5530) <= not(layer0_outputs(8385)) or (layer0_outputs(97));
    layer1_outputs(5531) <= (layer0_outputs(10218)) xor (layer0_outputs(1818));
    layer1_outputs(5532) <= layer0_outputs(7963);
    layer1_outputs(5533) <= layer0_outputs(9233);
    layer1_outputs(5534) <= not(layer0_outputs(9256));
    layer1_outputs(5535) <= not((layer0_outputs(1108)) or (layer0_outputs(3200)));
    layer1_outputs(5536) <= layer0_outputs(7591);
    layer1_outputs(5537) <= layer0_outputs(7218);
    layer1_outputs(5538) <= not(layer0_outputs(9435)) or (layer0_outputs(2012));
    layer1_outputs(5539) <= layer0_outputs(9811);
    layer1_outputs(5540) <= layer0_outputs(8518);
    layer1_outputs(5541) <= (layer0_outputs(3310)) and not (layer0_outputs(5378));
    layer1_outputs(5542) <= not(layer0_outputs(3997));
    layer1_outputs(5543) <= (layer0_outputs(4885)) or (layer0_outputs(6414));
    layer1_outputs(5544) <= not(layer0_outputs(3368)) or (layer0_outputs(7653));
    layer1_outputs(5545) <= not(layer0_outputs(4925));
    layer1_outputs(5546) <= not(layer0_outputs(5096));
    layer1_outputs(5547) <= (layer0_outputs(9399)) and not (layer0_outputs(1092));
    layer1_outputs(5548) <= (layer0_outputs(2622)) or (layer0_outputs(6660));
    layer1_outputs(5549) <= '1';
    layer1_outputs(5550) <= layer0_outputs(7456);
    layer1_outputs(5551) <= not(layer0_outputs(172)) or (layer0_outputs(2837));
    layer1_outputs(5552) <= (layer0_outputs(7610)) or (layer0_outputs(5688));
    layer1_outputs(5553) <= not(layer0_outputs(5798)) or (layer0_outputs(5958));
    layer1_outputs(5554) <= not(layer0_outputs(4262));
    layer1_outputs(5555) <= not((layer0_outputs(4295)) or (layer0_outputs(6690)));
    layer1_outputs(5556) <= not(layer0_outputs(1080));
    layer1_outputs(5557) <= layer0_outputs(7678);
    layer1_outputs(5558) <= not(layer0_outputs(5356));
    layer1_outputs(5559) <= layer0_outputs(8531);
    layer1_outputs(5560) <= not(layer0_outputs(4401));
    layer1_outputs(5561) <= (layer0_outputs(3330)) and (layer0_outputs(3713));
    layer1_outputs(5562) <= (layer0_outputs(3428)) and not (layer0_outputs(2174));
    layer1_outputs(5563) <= not(layer0_outputs(9726));
    layer1_outputs(5564) <= not(layer0_outputs(4773));
    layer1_outputs(5565) <= not(layer0_outputs(8405));
    layer1_outputs(5566) <= not(layer0_outputs(5429)) or (layer0_outputs(6282));
    layer1_outputs(5567) <= not(layer0_outputs(9304)) or (layer0_outputs(4388));
    layer1_outputs(5568) <= (layer0_outputs(7084)) or (layer0_outputs(6115));
    layer1_outputs(5569) <= layer0_outputs(8077);
    layer1_outputs(5570) <= not(layer0_outputs(3578));
    layer1_outputs(5571) <= (layer0_outputs(162)) and (layer0_outputs(6448));
    layer1_outputs(5572) <= (layer0_outputs(110)) xor (layer0_outputs(2947));
    layer1_outputs(5573) <= not(layer0_outputs(637)) or (layer0_outputs(8540));
    layer1_outputs(5574) <= (layer0_outputs(5539)) and not (layer0_outputs(593));
    layer1_outputs(5575) <= not(layer0_outputs(1059)) or (layer0_outputs(715));
    layer1_outputs(5576) <= not(layer0_outputs(892)) or (layer0_outputs(9774));
    layer1_outputs(5577) <= (layer0_outputs(698)) xor (layer0_outputs(9044));
    layer1_outputs(5578) <= not(layer0_outputs(1433));
    layer1_outputs(5579) <= layer0_outputs(6555);
    layer1_outputs(5580) <= '1';
    layer1_outputs(5581) <= not(layer0_outputs(4692)) or (layer0_outputs(8000));
    layer1_outputs(5582) <= (layer0_outputs(8678)) and (layer0_outputs(3653));
    layer1_outputs(5583) <= (layer0_outputs(8953)) and not (layer0_outputs(3242));
    layer1_outputs(5584) <= not(layer0_outputs(6034)) or (layer0_outputs(7282));
    layer1_outputs(5585) <= not((layer0_outputs(1293)) or (layer0_outputs(2395)));
    layer1_outputs(5586) <= (layer0_outputs(3297)) xor (layer0_outputs(2224));
    layer1_outputs(5587) <= not(layer0_outputs(101));
    layer1_outputs(5588) <= not(layer0_outputs(7072));
    layer1_outputs(5589) <= '1';
    layer1_outputs(5590) <= layer0_outputs(3033);
    layer1_outputs(5591) <= (layer0_outputs(2578)) xor (layer0_outputs(7806));
    layer1_outputs(5592) <= layer0_outputs(550);
    layer1_outputs(5593) <= layer0_outputs(6531);
    layer1_outputs(5594) <= (layer0_outputs(7975)) and not (layer0_outputs(5606));
    layer1_outputs(5595) <= not(layer0_outputs(4841));
    layer1_outputs(5596) <= not(layer0_outputs(5300)) or (layer0_outputs(7275));
    layer1_outputs(5597) <= not(layer0_outputs(2009));
    layer1_outputs(5598) <= '1';
    layer1_outputs(5599) <= (layer0_outputs(3379)) and not (layer0_outputs(7842));
    layer1_outputs(5600) <= layer0_outputs(5035);
    layer1_outputs(5601) <= not((layer0_outputs(8817)) or (layer0_outputs(414)));
    layer1_outputs(5602) <= (layer0_outputs(2384)) and not (layer0_outputs(4639));
    layer1_outputs(5603) <= (layer0_outputs(2335)) or (layer0_outputs(6879));
    layer1_outputs(5604) <= not(layer0_outputs(2410));
    layer1_outputs(5605) <= not(layer0_outputs(1321));
    layer1_outputs(5606) <= layer0_outputs(10064);
    layer1_outputs(5607) <= not((layer0_outputs(3195)) or (layer0_outputs(1123)));
    layer1_outputs(5608) <= not(layer0_outputs(6817));
    layer1_outputs(5609) <= not(layer0_outputs(6061));
    layer1_outputs(5610) <= '1';
    layer1_outputs(5611) <= not(layer0_outputs(13));
    layer1_outputs(5612) <= not(layer0_outputs(3193));
    layer1_outputs(5613) <= not(layer0_outputs(2170));
    layer1_outputs(5614) <= (layer0_outputs(4918)) xor (layer0_outputs(2704));
    layer1_outputs(5615) <= '0';
    layer1_outputs(5616) <= not(layer0_outputs(3117));
    layer1_outputs(5617) <= not(layer0_outputs(10120));
    layer1_outputs(5618) <= not(layer0_outputs(5847));
    layer1_outputs(5619) <= (layer0_outputs(443)) and not (layer0_outputs(4566));
    layer1_outputs(5620) <= layer0_outputs(10028);
    layer1_outputs(5621) <= layer0_outputs(73);
    layer1_outputs(5622) <= layer0_outputs(9978);
    layer1_outputs(5623) <= not(layer0_outputs(200)) or (layer0_outputs(5502));
    layer1_outputs(5624) <= not(layer0_outputs(5988));
    layer1_outputs(5625) <= not(layer0_outputs(7831));
    layer1_outputs(5626) <= layer0_outputs(9695);
    layer1_outputs(5627) <= layer0_outputs(6062);
    layer1_outputs(5628) <= '1';
    layer1_outputs(5629) <= not(layer0_outputs(6008));
    layer1_outputs(5630) <= not(layer0_outputs(1634)) or (layer0_outputs(9521));
    layer1_outputs(5631) <= (layer0_outputs(617)) xor (layer0_outputs(5457));
    layer1_outputs(5632) <= not(layer0_outputs(4752)) or (layer0_outputs(827));
    layer1_outputs(5633) <= not(layer0_outputs(3893));
    layer1_outputs(5634) <= layer0_outputs(6359);
    layer1_outputs(5635) <= layer0_outputs(9602);
    layer1_outputs(5636) <= not(layer0_outputs(7213));
    layer1_outputs(5637) <= not((layer0_outputs(7665)) or (layer0_outputs(6276)));
    layer1_outputs(5638) <= not(layer0_outputs(6991));
    layer1_outputs(5639) <= (layer0_outputs(4437)) and not (layer0_outputs(2607));
    layer1_outputs(5640) <= not(layer0_outputs(5508));
    layer1_outputs(5641) <= (layer0_outputs(5852)) and (layer0_outputs(6244));
    layer1_outputs(5642) <= (layer0_outputs(3922)) or (layer0_outputs(3331));
    layer1_outputs(5643) <= '0';
    layer1_outputs(5644) <= not(layer0_outputs(6045));
    layer1_outputs(5645) <= layer0_outputs(8452);
    layer1_outputs(5646) <= not(layer0_outputs(5056));
    layer1_outputs(5647) <= not((layer0_outputs(6885)) and (layer0_outputs(8194)));
    layer1_outputs(5648) <= not((layer0_outputs(9215)) xor (layer0_outputs(5917)));
    layer1_outputs(5649) <= not(layer0_outputs(4605));
    layer1_outputs(5650) <= not(layer0_outputs(762));
    layer1_outputs(5651) <= layer0_outputs(5795);
    layer1_outputs(5652) <= not(layer0_outputs(4661));
    layer1_outputs(5653) <= (layer0_outputs(5276)) and (layer0_outputs(10173));
    layer1_outputs(5654) <= not((layer0_outputs(6618)) and (layer0_outputs(7699)));
    layer1_outputs(5655) <= '0';
    layer1_outputs(5656) <= not((layer0_outputs(3030)) or (layer0_outputs(1186)));
    layer1_outputs(5657) <= not(layer0_outputs(2908)) or (layer0_outputs(4425));
    layer1_outputs(5658) <= not((layer0_outputs(9697)) and (layer0_outputs(843)));
    layer1_outputs(5659) <= not(layer0_outputs(8967));
    layer1_outputs(5660) <= layer0_outputs(5888);
    layer1_outputs(5661) <= layer0_outputs(8480);
    layer1_outputs(5662) <= (layer0_outputs(3959)) or (layer0_outputs(9386));
    layer1_outputs(5663) <= (layer0_outputs(2300)) or (layer0_outputs(1741));
    layer1_outputs(5664) <= not(layer0_outputs(9361));
    layer1_outputs(5665) <= not((layer0_outputs(6304)) xor (layer0_outputs(773)));
    layer1_outputs(5666) <= layer0_outputs(2893);
    layer1_outputs(5667) <= not(layer0_outputs(6859)) or (layer0_outputs(6419));
    layer1_outputs(5668) <= not((layer0_outputs(6049)) or (layer0_outputs(678)));
    layer1_outputs(5669) <= not(layer0_outputs(7842));
    layer1_outputs(5670) <= layer0_outputs(2433);
    layer1_outputs(5671) <= layer0_outputs(6607);
    layer1_outputs(5672) <= not(layer0_outputs(9859));
    layer1_outputs(5673) <= layer0_outputs(3955);
    layer1_outputs(5674) <= layer0_outputs(1298);
    layer1_outputs(5675) <= not(layer0_outputs(8143)) or (layer0_outputs(3049));
    layer1_outputs(5676) <= not((layer0_outputs(9055)) and (layer0_outputs(7806)));
    layer1_outputs(5677) <= (layer0_outputs(2294)) and not (layer0_outputs(5114));
    layer1_outputs(5678) <= (layer0_outputs(1481)) and not (layer0_outputs(8270));
    layer1_outputs(5679) <= layer0_outputs(5529);
    layer1_outputs(5680) <= layer0_outputs(9441);
    layer1_outputs(5681) <= (layer0_outputs(6337)) or (layer0_outputs(9906));
    layer1_outputs(5682) <= not(layer0_outputs(1178)) or (layer0_outputs(5721));
    layer1_outputs(5683) <= '0';
    layer1_outputs(5684) <= layer0_outputs(3275);
    layer1_outputs(5685) <= (layer0_outputs(5217)) xor (layer0_outputs(79));
    layer1_outputs(5686) <= not((layer0_outputs(5327)) xor (layer0_outputs(1131)));
    layer1_outputs(5687) <= (layer0_outputs(2793)) and not (layer0_outputs(2716));
    layer1_outputs(5688) <= (layer0_outputs(2944)) and not (layer0_outputs(9393));
    layer1_outputs(5689) <= (layer0_outputs(1906)) xor (layer0_outputs(6280));
    layer1_outputs(5690) <= (layer0_outputs(2227)) or (layer0_outputs(724));
    layer1_outputs(5691) <= not(layer0_outputs(6931)) or (layer0_outputs(596));
    layer1_outputs(5692) <= not(layer0_outputs(9564));
    layer1_outputs(5693) <= not((layer0_outputs(8537)) or (layer0_outputs(4877)));
    layer1_outputs(5694) <= layer0_outputs(4795);
    layer1_outputs(5695) <= layer0_outputs(1037);
    layer1_outputs(5696) <= not(layer0_outputs(3457)) or (layer0_outputs(5909));
    layer1_outputs(5697) <= not(layer0_outputs(6819));
    layer1_outputs(5698) <= layer0_outputs(1265);
    layer1_outputs(5699) <= not(layer0_outputs(6070));
    layer1_outputs(5700) <= (layer0_outputs(2445)) and not (layer0_outputs(99));
    layer1_outputs(5701) <= not(layer0_outputs(3561));
    layer1_outputs(5702) <= not(layer0_outputs(5241));
    layer1_outputs(5703) <= (layer0_outputs(3303)) and not (layer0_outputs(9828));
    layer1_outputs(5704) <= '1';
    layer1_outputs(5705) <= (layer0_outputs(7644)) and (layer0_outputs(6278));
    layer1_outputs(5706) <= layer0_outputs(447);
    layer1_outputs(5707) <= not((layer0_outputs(944)) and (layer0_outputs(6197)));
    layer1_outputs(5708) <= layer0_outputs(1668);
    layer1_outputs(5709) <= layer0_outputs(5055);
    layer1_outputs(5710) <= not((layer0_outputs(510)) or (layer0_outputs(2216)));
    layer1_outputs(5711) <= not(layer0_outputs(2240));
    layer1_outputs(5712) <= not(layer0_outputs(627)) or (layer0_outputs(9561));
    layer1_outputs(5713) <= not(layer0_outputs(6470));
    layer1_outputs(5714) <= not((layer0_outputs(535)) or (layer0_outputs(1523)));
    layer1_outputs(5715) <= not(layer0_outputs(4091));
    layer1_outputs(5716) <= layer0_outputs(904);
    layer1_outputs(5717) <= not(layer0_outputs(9322)) or (layer0_outputs(1927));
    layer1_outputs(5718) <= (layer0_outputs(3627)) xor (layer0_outputs(7558));
    layer1_outputs(5719) <= not(layer0_outputs(7268)) or (layer0_outputs(9847));
    layer1_outputs(5720) <= layer0_outputs(7936);
    layer1_outputs(5721) <= not(layer0_outputs(3951));
    layer1_outputs(5722) <= (layer0_outputs(9570)) and not (layer0_outputs(2628));
    layer1_outputs(5723) <= not((layer0_outputs(3609)) or (layer0_outputs(916)));
    layer1_outputs(5724) <= (layer0_outputs(6461)) or (layer0_outputs(4844));
    layer1_outputs(5725) <= not((layer0_outputs(9848)) and (layer0_outputs(5309)));
    layer1_outputs(5726) <= not(layer0_outputs(5134)) or (layer0_outputs(723));
    layer1_outputs(5727) <= not((layer0_outputs(6735)) or (layer0_outputs(5252)));
    layer1_outputs(5728) <= (layer0_outputs(8917)) and (layer0_outputs(1245));
    layer1_outputs(5729) <= not(layer0_outputs(6879));
    layer1_outputs(5730) <= '1';
    layer1_outputs(5731) <= not((layer0_outputs(2146)) and (layer0_outputs(7431)));
    layer1_outputs(5732) <= (layer0_outputs(2352)) and not (layer0_outputs(5403));
    layer1_outputs(5733) <= not(layer0_outputs(8362)) or (layer0_outputs(302));
    layer1_outputs(5734) <= layer0_outputs(1082);
    layer1_outputs(5735) <= not((layer0_outputs(4107)) and (layer0_outputs(3713)));
    layer1_outputs(5736) <= not((layer0_outputs(5129)) and (layer0_outputs(4686)));
    layer1_outputs(5737) <= not(layer0_outputs(2634));
    layer1_outputs(5738) <= layer0_outputs(2411);
    layer1_outputs(5739) <= not(layer0_outputs(2740));
    layer1_outputs(5740) <= layer0_outputs(4105);
    layer1_outputs(5741) <= layer0_outputs(5654);
    layer1_outputs(5742) <= (layer0_outputs(6467)) and not (layer0_outputs(89));
    layer1_outputs(5743) <= not(layer0_outputs(6200));
    layer1_outputs(5744) <= layer0_outputs(9249);
    layer1_outputs(5745) <= layer0_outputs(371);
    layer1_outputs(5746) <= (layer0_outputs(8569)) and (layer0_outputs(4645));
    layer1_outputs(5747) <= layer0_outputs(2723);
    layer1_outputs(5748) <= not(layer0_outputs(1112)) or (layer0_outputs(903));
    layer1_outputs(5749) <= (layer0_outputs(4039)) or (layer0_outputs(7907));
    layer1_outputs(5750) <= '1';
    layer1_outputs(5751) <= (layer0_outputs(6613)) or (layer0_outputs(6322));
    layer1_outputs(5752) <= not(layer0_outputs(10035));
    layer1_outputs(5753) <= not(layer0_outputs(5584)) or (layer0_outputs(6863));
    layer1_outputs(5754) <= not((layer0_outputs(9188)) and (layer0_outputs(4907)));
    layer1_outputs(5755) <= not(layer0_outputs(11));
    layer1_outputs(5756) <= (layer0_outputs(3751)) and (layer0_outputs(6380));
    layer1_outputs(5757) <= (layer0_outputs(6338)) and not (layer0_outputs(8962));
    layer1_outputs(5758) <= layer0_outputs(676);
    layer1_outputs(5759) <= not(layer0_outputs(2337)) or (layer0_outputs(7119));
    layer1_outputs(5760) <= not((layer0_outputs(7654)) xor (layer0_outputs(4789)));
    layer1_outputs(5761) <= '0';
    layer1_outputs(5762) <= (layer0_outputs(3753)) and (layer0_outputs(5386));
    layer1_outputs(5763) <= not(layer0_outputs(7777));
    layer1_outputs(5764) <= not(layer0_outputs(6482));
    layer1_outputs(5765) <= not((layer0_outputs(6643)) xor (layer0_outputs(8942)));
    layer1_outputs(5766) <= layer0_outputs(9236);
    layer1_outputs(5767) <= (layer0_outputs(1541)) and not (layer0_outputs(5968));
    layer1_outputs(5768) <= (layer0_outputs(322)) and (layer0_outputs(6877));
    layer1_outputs(5769) <= not(layer0_outputs(6040));
    layer1_outputs(5770) <= not((layer0_outputs(118)) or (layer0_outputs(9030)));
    layer1_outputs(5771) <= not((layer0_outputs(897)) or (layer0_outputs(4768)));
    layer1_outputs(5772) <= (layer0_outputs(1731)) and not (layer0_outputs(8449));
    layer1_outputs(5773) <= not(layer0_outputs(7381));
    layer1_outputs(5774) <= layer0_outputs(4763);
    layer1_outputs(5775) <= not(layer0_outputs(5296)) or (layer0_outputs(5247));
    layer1_outputs(5776) <= (layer0_outputs(9208)) and not (layer0_outputs(3746));
    layer1_outputs(5777) <= '1';
    layer1_outputs(5778) <= layer0_outputs(8122);
    layer1_outputs(5779) <= (layer0_outputs(7262)) or (layer0_outputs(2254));
    layer1_outputs(5780) <= (layer0_outputs(4864)) or (layer0_outputs(6370));
    layer1_outputs(5781) <= not(layer0_outputs(2522)) or (layer0_outputs(3973));
    layer1_outputs(5782) <= not(layer0_outputs(1319));
    layer1_outputs(5783) <= (layer0_outputs(9940)) xor (layer0_outputs(684));
    layer1_outputs(5784) <= (layer0_outputs(6389)) and not (layer0_outputs(1107));
    layer1_outputs(5785) <= (layer0_outputs(9092)) and (layer0_outputs(180));
    layer1_outputs(5786) <= not(layer0_outputs(2014)) or (layer0_outputs(3099));
    layer1_outputs(5787) <= (layer0_outputs(3398)) and not (layer0_outputs(7939));
    layer1_outputs(5788) <= not((layer0_outputs(9844)) or (layer0_outputs(10172)));
    layer1_outputs(5789) <= layer0_outputs(9027);
    layer1_outputs(5790) <= (layer0_outputs(9181)) and not (layer0_outputs(265));
    layer1_outputs(5791) <= not(layer0_outputs(345));
    layer1_outputs(5792) <= layer0_outputs(7694);
    layer1_outputs(5793) <= layer0_outputs(8578);
    layer1_outputs(5794) <= (layer0_outputs(5661)) and not (layer0_outputs(571));
    layer1_outputs(5795) <= layer0_outputs(7716);
    layer1_outputs(5796) <= not(layer0_outputs(5242));
    layer1_outputs(5797) <= not(layer0_outputs(5533));
    layer1_outputs(5798) <= not(layer0_outputs(382));
    layer1_outputs(5799) <= (layer0_outputs(6141)) xor (layer0_outputs(6260));
    layer1_outputs(5800) <= not(layer0_outputs(9996));
    layer1_outputs(5801) <= layer0_outputs(4740);
    layer1_outputs(5802) <= not(layer0_outputs(2313)) or (layer0_outputs(5630));
    layer1_outputs(5803) <= layer0_outputs(3043);
    layer1_outputs(5804) <= (layer0_outputs(7077)) or (layer0_outputs(9330));
    layer1_outputs(5805) <= (layer0_outputs(1060)) xor (layer0_outputs(10163));
    layer1_outputs(5806) <= not((layer0_outputs(6258)) or (layer0_outputs(4615)));
    layer1_outputs(5807) <= layer0_outputs(899);
    layer1_outputs(5808) <= (layer0_outputs(8255)) and not (layer0_outputs(3822));
    layer1_outputs(5809) <= not(layer0_outputs(8565)) or (layer0_outputs(2348));
    layer1_outputs(5810) <= (layer0_outputs(256)) and not (layer0_outputs(6102));
    layer1_outputs(5811) <= (layer0_outputs(3416)) xor (layer0_outputs(2853));
    layer1_outputs(5812) <= not(layer0_outputs(5051));
    layer1_outputs(5813) <= not(layer0_outputs(6274));
    layer1_outputs(5814) <= not(layer0_outputs(6433)) or (layer0_outputs(8282));
    layer1_outputs(5815) <= (layer0_outputs(3325)) or (layer0_outputs(772));
    layer1_outputs(5816) <= not((layer0_outputs(2312)) and (layer0_outputs(2835)));
    layer1_outputs(5817) <= not(layer0_outputs(8257));
    layer1_outputs(5818) <= not(layer0_outputs(3650));
    layer1_outputs(5819) <= not(layer0_outputs(1696));
    layer1_outputs(5820) <= (layer0_outputs(372)) xor (layer0_outputs(7993));
    layer1_outputs(5821) <= (layer0_outputs(7743)) and not (layer0_outputs(2467));
    layer1_outputs(5822) <= (layer0_outputs(9124)) and not (layer0_outputs(8131));
    layer1_outputs(5823) <= not(layer0_outputs(3772));
    layer1_outputs(5824) <= not(layer0_outputs(8141));
    layer1_outputs(5825) <= layer0_outputs(867);
    layer1_outputs(5826) <= (layer0_outputs(927)) or (layer0_outputs(5398));
    layer1_outputs(5827) <= layer0_outputs(3593);
    layer1_outputs(5828) <= (layer0_outputs(3041)) or (layer0_outputs(3336));
    layer1_outputs(5829) <= '0';
    layer1_outputs(5830) <= (layer0_outputs(3093)) and not (layer0_outputs(5178));
    layer1_outputs(5831) <= not(layer0_outputs(5869));
    layer1_outputs(5832) <= not(layer0_outputs(483));
    layer1_outputs(5833) <= not(layer0_outputs(7724));
    layer1_outputs(5834) <= (layer0_outputs(5518)) and not (layer0_outputs(1556));
    layer1_outputs(5835) <= layer0_outputs(292);
    layer1_outputs(5836) <= (layer0_outputs(6697)) and (layer0_outputs(5547));
    layer1_outputs(5837) <= layer0_outputs(2512);
    layer1_outputs(5838) <= (layer0_outputs(8219)) and not (layer0_outputs(4415));
    layer1_outputs(5839) <= layer0_outputs(1008);
    layer1_outputs(5840) <= layer0_outputs(793);
    layer1_outputs(5841) <= not(layer0_outputs(3945)) or (layer0_outputs(1591));
    layer1_outputs(5842) <= (layer0_outputs(785)) or (layer0_outputs(8784));
    layer1_outputs(5843) <= not((layer0_outputs(1810)) or (layer0_outputs(9146)));
    layer1_outputs(5844) <= (layer0_outputs(1560)) xor (layer0_outputs(1639));
    layer1_outputs(5845) <= not((layer0_outputs(9076)) and (layer0_outputs(7972)));
    layer1_outputs(5846) <= not(layer0_outputs(7675)) or (layer0_outputs(4813));
    layer1_outputs(5847) <= not(layer0_outputs(9186)) or (layer0_outputs(9749));
    layer1_outputs(5848) <= layer0_outputs(2378);
    layer1_outputs(5849) <= not(layer0_outputs(9387));
    layer1_outputs(5850) <= layer0_outputs(3455);
    layer1_outputs(5851) <= layer0_outputs(6896);
    layer1_outputs(5852) <= layer0_outputs(4833);
    layer1_outputs(5853) <= layer0_outputs(8837);
    layer1_outputs(5854) <= not(layer0_outputs(147));
    layer1_outputs(5855) <= not((layer0_outputs(3933)) and (layer0_outputs(5552)));
    layer1_outputs(5856) <= layer0_outputs(5288);
    layer1_outputs(5857) <= '0';
    layer1_outputs(5858) <= not(layer0_outputs(2010));
    layer1_outputs(5859) <= not(layer0_outputs(3632));
    layer1_outputs(5860) <= not(layer0_outputs(2937)) or (layer0_outputs(9588));
    layer1_outputs(5861) <= (layer0_outputs(1215)) and not (layer0_outputs(3863));
    layer1_outputs(5862) <= not(layer0_outputs(2978)) or (layer0_outputs(6163));
    layer1_outputs(5863) <= not(layer0_outputs(1580));
    layer1_outputs(5864) <= not((layer0_outputs(9583)) or (layer0_outputs(2005)));
    layer1_outputs(5865) <= not((layer0_outputs(6998)) or (layer0_outputs(6319)));
    layer1_outputs(5866) <= layer0_outputs(2247);
    layer1_outputs(5867) <= not(layer0_outputs(8306)) or (layer0_outputs(6511));
    layer1_outputs(5868) <= not(layer0_outputs(5098)) or (layer0_outputs(4507));
    layer1_outputs(5869) <= not((layer0_outputs(7656)) and (layer0_outputs(6726)));
    layer1_outputs(5870) <= not(layer0_outputs(8049)) or (layer0_outputs(1497));
    layer1_outputs(5871) <= not(layer0_outputs(5030));
    layer1_outputs(5872) <= (layer0_outputs(3267)) or (layer0_outputs(852));
    layer1_outputs(5873) <= not(layer0_outputs(6893));
    layer1_outputs(5874) <= not(layer0_outputs(9698));
    layer1_outputs(5875) <= not((layer0_outputs(6328)) or (layer0_outputs(3221)));
    layer1_outputs(5876) <= (layer0_outputs(8965)) or (layer0_outputs(3906));
    layer1_outputs(5877) <= not(layer0_outputs(8494)) or (layer0_outputs(8805));
    layer1_outputs(5878) <= not(layer0_outputs(8663));
    layer1_outputs(5879) <= layer0_outputs(7397);
    layer1_outputs(5880) <= layer0_outputs(4000);
    layer1_outputs(5881) <= (layer0_outputs(4309)) and not (layer0_outputs(5382));
    layer1_outputs(5882) <= not((layer0_outputs(7965)) or (layer0_outputs(2404)));
    layer1_outputs(5883) <= not((layer0_outputs(1420)) and (layer0_outputs(5577)));
    layer1_outputs(5884) <= layer0_outputs(626);
    layer1_outputs(5885) <= not((layer0_outputs(5608)) or (layer0_outputs(2318)));
    layer1_outputs(5886) <= not(layer0_outputs(7520));
    layer1_outputs(5887) <= layer0_outputs(3370);
    layer1_outputs(5888) <= not((layer0_outputs(7743)) or (layer0_outputs(9276)));
    layer1_outputs(5889) <= not(layer0_outputs(5383));
    layer1_outputs(5890) <= not((layer0_outputs(7161)) and (layer0_outputs(5262)));
    layer1_outputs(5891) <= (layer0_outputs(3639)) or (layer0_outputs(7264));
    layer1_outputs(5892) <= not(layer0_outputs(7397));
    layer1_outputs(5893) <= not((layer0_outputs(224)) or (layer0_outputs(4971)));
    layer1_outputs(5894) <= not(layer0_outputs(7535));
    layer1_outputs(5895) <= (layer0_outputs(5353)) and not (layer0_outputs(8038));
    layer1_outputs(5896) <= not(layer0_outputs(6513));
    layer1_outputs(5897) <= layer0_outputs(9281);
    layer1_outputs(5898) <= (layer0_outputs(6368)) and (layer0_outputs(3888));
    layer1_outputs(5899) <= layer0_outputs(10052);
    layer1_outputs(5900) <= (layer0_outputs(9947)) and (layer0_outputs(3817));
    layer1_outputs(5901) <= not(layer0_outputs(1535)) or (layer0_outputs(7908));
    layer1_outputs(5902) <= not((layer0_outputs(7156)) or (layer0_outputs(8226)));
    layer1_outputs(5903) <= (layer0_outputs(286)) xor (layer0_outputs(4239));
    layer1_outputs(5904) <= (layer0_outputs(5475)) or (layer0_outputs(6202));
    layer1_outputs(5905) <= not(layer0_outputs(7787)) or (layer0_outputs(10067));
    layer1_outputs(5906) <= not(layer0_outputs(7071));
    layer1_outputs(5907) <= layer0_outputs(1655);
    layer1_outputs(5908) <= layer0_outputs(334);
    layer1_outputs(5909) <= not((layer0_outputs(1538)) or (layer0_outputs(3942)));
    layer1_outputs(5910) <= not(layer0_outputs(2941)) or (layer0_outputs(9558));
    layer1_outputs(5911) <= (layer0_outputs(5874)) and not (layer0_outputs(758));
    layer1_outputs(5912) <= '1';
    layer1_outputs(5913) <= layer0_outputs(8506);
    layer1_outputs(5914) <= not(layer0_outputs(6039));
    layer1_outputs(5915) <= (layer0_outputs(384)) and (layer0_outputs(6006));
    layer1_outputs(5916) <= not(layer0_outputs(2601));
    layer1_outputs(5917) <= not((layer0_outputs(8716)) or (layer0_outputs(9426)));
    layer1_outputs(5918) <= layer0_outputs(1440);
    layer1_outputs(5919) <= layer0_outputs(771);
    layer1_outputs(5920) <= (layer0_outputs(5164)) xor (layer0_outputs(9657));
    layer1_outputs(5921) <= not((layer0_outputs(1605)) and (layer0_outputs(7742)));
    layer1_outputs(5922) <= (layer0_outputs(2482)) and not (layer0_outputs(3619));
    layer1_outputs(5923) <= not(layer0_outputs(3406));
    layer1_outputs(5924) <= not((layer0_outputs(4741)) xor (layer0_outputs(7735)));
    layer1_outputs(5925) <= layer0_outputs(1702);
    layer1_outputs(5926) <= layer0_outputs(9435);
    layer1_outputs(5927) <= (layer0_outputs(6829)) and not (layer0_outputs(6134));
    layer1_outputs(5928) <= not(layer0_outputs(153));
    layer1_outputs(5929) <= (layer0_outputs(3031)) and not (layer0_outputs(3230));
    layer1_outputs(5930) <= (layer0_outputs(5553)) and (layer0_outputs(8094));
    layer1_outputs(5931) <= (layer0_outputs(2817)) and not (layer0_outputs(3966));
    layer1_outputs(5932) <= not(layer0_outputs(9135));
    layer1_outputs(5933) <= (layer0_outputs(6862)) and (layer0_outputs(2867));
    layer1_outputs(5934) <= (layer0_outputs(6827)) and not (layer0_outputs(3220));
    layer1_outputs(5935) <= (layer0_outputs(1545)) and not (layer0_outputs(6247));
    layer1_outputs(5936) <= not((layer0_outputs(434)) or (layer0_outputs(2479)));
    layer1_outputs(5937) <= not(layer0_outputs(8521));
    layer1_outputs(5938) <= layer0_outputs(553);
    layer1_outputs(5939) <= (layer0_outputs(3332)) or (layer0_outputs(9380));
    layer1_outputs(5940) <= (layer0_outputs(9472)) xor (layer0_outputs(7159));
    layer1_outputs(5941) <= not(layer0_outputs(531));
    layer1_outputs(5942) <= layer0_outputs(2365);
    layer1_outputs(5943) <= layer0_outputs(2210);
    layer1_outputs(5944) <= (layer0_outputs(938)) and not (layer0_outputs(141));
    layer1_outputs(5945) <= not(layer0_outputs(3434)) or (layer0_outputs(7717));
    layer1_outputs(5946) <= not((layer0_outputs(6821)) and (layer0_outputs(4419)));
    layer1_outputs(5947) <= layer0_outputs(7231);
    layer1_outputs(5948) <= layer0_outputs(145);
    layer1_outputs(5949) <= '1';
    layer1_outputs(5950) <= not(layer0_outputs(9232)) or (layer0_outputs(9053));
    layer1_outputs(5951) <= (layer0_outputs(792)) and not (layer0_outputs(2949));
    layer1_outputs(5952) <= layer0_outputs(5589);
    layer1_outputs(5953) <= (layer0_outputs(2728)) and (layer0_outputs(3159));
    layer1_outputs(5954) <= not((layer0_outputs(3328)) and (layer0_outputs(4529)));
    layer1_outputs(5955) <= not(layer0_outputs(9063));
    layer1_outputs(5956) <= not(layer0_outputs(5193));
    layer1_outputs(5957) <= not((layer0_outputs(6649)) xor (layer0_outputs(9054)));
    layer1_outputs(5958) <= layer0_outputs(9615);
    layer1_outputs(5959) <= layer0_outputs(7015);
    layer1_outputs(5960) <= not(layer0_outputs(4206)) or (layer0_outputs(3073));
    layer1_outputs(5961) <= (layer0_outputs(7850)) and not (layer0_outputs(9509));
    layer1_outputs(5962) <= not(layer0_outputs(8363));
    layer1_outputs(5963) <= layer0_outputs(7713);
    layer1_outputs(5964) <= layer0_outputs(2877);
    layer1_outputs(5965) <= not(layer0_outputs(5940));
    layer1_outputs(5966) <= layer0_outputs(1796);
    layer1_outputs(5967) <= not(layer0_outputs(6693));
    layer1_outputs(5968) <= not(layer0_outputs(10208)) or (layer0_outputs(3120));
    layer1_outputs(5969) <= not(layer0_outputs(8163)) or (layer0_outputs(9004));
    layer1_outputs(5970) <= not((layer0_outputs(9526)) or (layer0_outputs(5570)));
    layer1_outputs(5971) <= '1';
    layer1_outputs(5972) <= (layer0_outputs(7593)) xor (layer0_outputs(875));
    layer1_outputs(5973) <= (layer0_outputs(7710)) and not (layer0_outputs(1496));
    layer1_outputs(5974) <= (layer0_outputs(1846)) or (layer0_outputs(9077));
    layer1_outputs(5975) <= not(layer0_outputs(9630));
    layer1_outputs(5976) <= not(layer0_outputs(7559));
    layer1_outputs(5977) <= not(layer0_outputs(3754)) or (layer0_outputs(1109));
    layer1_outputs(5978) <= layer0_outputs(4218);
    layer1_outputs(5979) <= not((layer0_outputs(6003)) and (layer0_outputs(6626)));
    layer1_outputs(5980) <= '1';
    layer1_outputs(5981) <= (layer0_outputs(7482)) or (layer0_outputs(4304));
    layer1_outputs(5982) <= not(layer0_outputs(7112));
    layer1_outputs(5983) <= layer0_outputs(9524);
    layer1_outputs(5984) <= layer0_outputs(10181);
    layer1_outputs(5985) <= (layer0_outputs(7752)) or (layer0_outputs(7868));
    layer1_outputs(5986) <= not(layer0_outputs(5074));
    layer1_outputs(5987) <= not(layer0_outputs(4079));
    layer1_outputs(5988) <= not((layer0_outputs(6018)) or (layer0_outputs(10157)));
    layer1_outputs(5989) <= not(layer0_outputs(7899)) or (layer0_outputs(2721));
    layer1_outputs(5990) <= layer0_outputs(6738);
    layer1_outputs(5991) <= not((layer0_outputs(8499)) xor (layer0_outputs(7071)));
    layer1_outputs(5992) <= not(layer0_outputs(5231)) or (layer0_outputs(4872));
    layer1_outputs(5993) <= layer0_outputs(7765);
    layer1_outputs(5994) <= not(layer0_outputs(8927)) or (layer0_outputs(8771));
    layer1_outputs(5995) <= not(layer0_outputs(8078)) or (layer0_outputs(1402));
    layer1_outputs(5996) <= not(layer0_outputs(8866)) or (layer0_outputs(55));
    layer1_outputs(5997) <= not(layer0_outputs(4738));
    layer1_outputs(5998) <= (layer0_outputs(1918)) and not (layer0_outputs(8095));
    layer1_outputs(5999) <= not(layer0_outputs(2636));
    layer1_outputs(6000) <= not(layer0_outputs(2739));
    layer1_outputs(6001) <= (layer0_outputs(5535)) or (layer0_outputs(9503));
    layer1_outputs(6002) <= not(layer0_outputs(5753)) or (layer0_outputs(2545));
    layer1_outputs(6003) <= layer0_outputs(4808);
    layer1_outputs(6004) <= (layer0_outputs(9724)) or (layer0_outputs(5057));
    layer1_outputs(6005) <= layer0_outputs(6010);
    layer1_outputs(6006) <= not((layer0_outputs(2565)) xor (layer0_outputs(1551)));
    layer1_outputs(6007) <= not(layer0_outputs(7578)) or (layer0_outputs(9478));
    layer1_outputs(6008) <= (layer0_outputs(3507)) and not (layer0_outputs(3842));
    layer1_outputs(6009) <= not(layer0_outputs(4890)) or (layer0_outputs(1536));
    layer1_outputs(6010) <= layer0_outputs(1089);
    layer1_outputs(6011) <= not(layer0_outputs(3629));
    layer1_outputs(6012) <= not((layer0_outputs(3763)) or (layer0_outputs(2185)));
    layer1_outputs(6013) <= (layer0_outputs(2349)) xor (layer0_outputs(1321));
    layer1_outputs(6014) <= (layer0_outputs(4895)) and not (layer0_outputs(9499));
    layer1_outputs(6015) <= (layer0_outputs(7346)) and not (layer0_outputs(1111));
    layer1_outputs(6016) <= not(layer0_outputs(9527));
    layer1_outputs(6017) <= layer0_outputs(4032);
    layer1_outputs(6018) <= (layer0_outputs(3338)) or (layer0_outputs(8704));
    layer1_outputs(6019) <= layer0_outputs(3903);
    layer1_outputs(6020) <= (layer0_outputs(1651)) or (layer0_outputs(890));
    layer1_outputs(6021) <= not(layer0_outputs(9597));
    layer1_outputs(6022) <= not(layer0_outputs(8486));
    layer1_outputs(6023) <= not(layer0_outputs(2393)) or (layer0_outputs(548));
    layer1_outputs(6024) <= not((layer0_outputs(2177)) xor (layer0_outputs(2049)));
    layer1_outputs(6025) <= not(layer0_outputs(3287));
    layer1_outputs(6026) <= (layer0_outputs(1584)) and not (layer0_outputs(4372));
    layer1_outputs(6027) <= not(layer0_outputs(986)) or (layer0_outputs(6053));
    layer1_outputs(6028) <= not((layer0_outputs(5514)) or (layer0_outputs(671)));
    layer1_outputs(6029) <= not(layer0_outputs(3046)) or (layer0_outputs(371));
    layer1_outputs(6030) <= not(layer0_outputs(1105));
    layer1_outputs(6031) <= layer0_outputs(6542);
    layer1_outputs(6032) <= (layer0_outputs(1624)) and not (layer0_outputs(3658));
    layer1_outputs(6033) <= (layer0_outputs(5033)) and not (layer0_outputs(9508));
    layer1_outputs(6034) <= (layer0_outputs(3181)) xor (layer0_outputs(3407));
    layer1_outputs(6035) <= (layer0_outputs(7097)) and not (layer0_outputs(7571));
    layer1_outputs(6036) <= layer0_outputs(8767);
    layer1_outputs(6037) <= not(layer0_outputs(1652));
    layer1_outputs(6038) <= layer0_outputs(3325);
    layer1_outputs(6039) <= layer0_outputs(10232);
    layer1_outputs(6040) <= (layer0_outputs(7623)) or (layer0_outputs(156));
    layer1_outputs(6041) <= (layer0_outputs(2570)) and not (layer0_outputs(8351));
    layer1_outputs(6042) <= (layer0_outputs(8760)) and not (layer0_outputs(2597));
    layer1_outputs(6043) <= not(layer0_outputs(8907));
    layer1_outputs(6044) <= not(layer0_outputs(4148)) or (layer0_outputs(155));
    layer1_outputs(6045) <= layer0_outputs(6970);
    layer1_outputs(6046) <= not(layer0_outputs(3348));
    layer1_outputs(6047) <= not(layer0_outputs(3793));
    layer1_outputs(6048) <= not(layer0_outputs(7594));
    layer1_outputs(6049) <= not(layer0_outputs(606));
    layer1_outputs(6050) <= (layer0_outputs(5904)) or (layer0_outputs(2556));
    layer1_outputs(6051) <= layer0_outputs(690);
    layer1_outputs(6052) <= layer0_outputs(3601);
    layer1_outputs(6053) <= not(layer0_outputs(791));
    layer1_outputs(6054) <= (layer0_outputs(9094)) and not (layer0_outputs(1193));
    layer1_outputs(6055) <= layer0_outputs(8253);
    layer1_outputs(6056) <= layer0_outputs(5203);
    layer1_outputs(6057) <= '0';
    layer1_outputs(6058) <= layer0_outputs(1012);
    layer1_outputs(6059) <= (layer0_outputs(1307)) or (layer0_outputs(7290));
    layer1_outputs(6060) <= not((layer0_outputs(427)) and (layer0_outputs(5510)));
    layer1_outputs(6061) <= not((layer0_outputs(5455)) xor (layer0_outputs(6017)));
    layer1_outputs(6062) <= not(layer0_outputs(7488));
    layer1_outputs(6063) <= layer0_outputs(1062);
    layer1_outputs(6064) <= not((layer0_outputs(10107)) or (layer0_outputs(6092)));
    layer1_outputs(6065) <= (layer0_outputs(2645)) and (layer0_outputs(4696));
    layer1_outputs(6066) <= '1';
    layer1_outputs(6067) <= not(layer0_outputs(2314));
    layer1_outputs(6068) <= (layer0_outputs(2598)) and not (layer0_outputs(9313));
    layer1_outputs(6069) <= not(layer0_outputs(4821));
    layer1_outputs(6070) <= not(layer0_outputs(4132)) or (layer0_outputs(4966));
    layer1_outputs(6071) <= not(layer0_outputs(395));
    layer1_outputs(6072) <= not(layer0_outputs(3388)) or (layer0_outputs(6542));
    layer1_outputs(6073) <= not((layer0_outputs(6696)) or (layer0_outputs(5916)));
    layer1_outputs(6074) <= layer0_outputs(7537);
    layer1_outputs(6075) <= not(layer0_outputs(7727)) or (layer0_outputs(3531));
    layer1_outputs(6076) <= (layer0_outputs(1300)) and not (layer0_outputs(2008));
    layer1_outputs(6077) <= layer0_outputs(8134);
    layer1_outputs(6078) <= layer0_outputs(6274);
    layer1_outputs(6079) <= (layer0_outputs(1881)) or (layer0_outputs(4201));
    layer1_outputs(6080) <= not(layer0_outputs(6498));
    layer1_outputs(6081) <= (layer0_outputs(542)) or (layer0_outputs(3878));
    layer1_outputs(6082) <= not(layer0_outputs(3048));
    layer1_outputs(6083) <= layer0_outputs(1202);
    layer1_outputs(6084) <= (layer0_outputs(9939)) and (layer0_outputs(9359));
    layer1_outputs(6085) <= (layer0_outputs(2539)) and not (layer0_outputs(8221));
    layer1_outputs(6086) <= not(layer0_outputs(4687)) or (layer0_outputs(4103));
    layer1_outputs(6087) <= layer0_outputs(9137);
    layer1_outputs(6088) <= not(layer0_outputs(4600));
    layer1_outputs(6089) <= (layer0_outputs(8262)) and not (layer0_outputs(6960));
    layer1_outputs(6090) <= (layer0_outputs(4169)) or (layer0_outputs(4784));
    layer1_outputs(6091) <= (layer0_outputs(7327)) and not (layer0_outputs(8873));
    layer1_outputs(6092) <= (layer0_outputs(3067)) and not (layer0_outputs(3421));
    layer1_outputs(6093) <= layer0_outputs(2429);
    layer1_outputs(6094) <= layer0_outputs(248);
    layer1_outputs(6095) <= not(layer0_outputs(9022));
    layer1_outputs(6096) <= not(layer0_outputs(8376)) or (layer0_outputs(7558));
    layer1_outputs(6097) <= (layer0_outputs(7599)) and not (layer0_outputs(5830));
    layer1_outputs(6098) <= layer0_outputs(3534);
    layer1_outputs(6099) <= not((layer0_outputs(8382)) or (layer0_outputs(4764)));
    layer1_outputs(6100) <= layer0_outputs(3813);
    layer1_outputs(6101) <= not(layer0_outputs(2904));
    layer1_outputs(6102) <= not(layer0_outputs(8779)) or (layer0_outputs(1815));
    layer1_outputs(6103) <= not((layer0_outputs(8469)) or (layer0_outputs(6071)));
    layer1_outputs(6104) <= not(layer0_outputs(6652)) or (layer0_outputs(8047));
    layer1_outputs(6105) <= not(layer0_outputs(9036));
    layer1_outputs(6106) <= layer0_outputs(4448);
    layer1_outputs(6107) <= not(layer0_outputs(2621));
    layer1_outputs(6108) <= (layer0_outputs(2413)) and not (layer0_outputs(910));
    layer1_outputs(6109) <= layer0_outputs(7850);
    layer1_outputs(6110) <= not(layer0_outputs(6001));
    layer1_outputs(6111) <= not(layer0_outputs(7459)) or (layer0_outputs(1706));
    layer1_outputs(6112) <= not(layer0_outputs(8863)) or (layer0_outputs(3492));
    layer1_outputs(6113) <= (layer0_outputs(5147)) xor (layer0_outputs(2892));
    layer1_outputs(6114) <= (layer0_outputs(8101)) or (layer0_outputs(1707));
    layer1_outputs(6115) <= '1';
    layer1_outputs(6116) <= not((layer0_outputs(381)) or (layer0_outputs(2290)));
    layer1_outputs(6117) <= not(layer0_outputs(3131)) or (layer0_outputs(4798));
    layer1_outputs(6118) <= not(layer0_outputs(9272));
    layer1_outputs(6119) <= (layer0_outputs(5523)) and (layer0_outputs(4707));
    layer1_outputs(6120) <= (layer0_outputs(6876)) and (layer0_outputs(7220));
    layer1_outputs(6121) <= not(layer0_outputs(6427));
    layer1_outputs(6122) <= not(layer0_outputs(6243));
    layer1_outputs(6123) <= not(layer0_outputs(5103));
    layer1_outputs(6124) <= not(layer0_outputs(2594));
    layer1_outputs(6125) <= (layer0_outputs(3853)) or (layer0_outputs(6676));
    layer1_outputs(6126) <= layer0_outputs(9565);
    layer1_outputs(6127) <= not((layer0_outputs(7465)) or (layer0_outputs(441)));
    layer1_outputs(6128) <= (layer0_outputs(10149)) and not (layer0_outputs(4654));
    layer1_outputs(6129) <= layer0_outputs(7770);
    layer1_outputs(6130) <= (layer0_outputs(9006)) or (layer0_outputs(4810));
    layer1_outputs(6131) <= not(layer0_outputs(3335)) or (layer0_outputs(4711));
    layer1_outputs(6132) <= not((layer0_outputs(10131)) and (layer0_outputs(4171)));
    layer1_outputs(6133) <= (layer0_outputs(2914)) and not (layer0_outputs(4444));
    layer1_outputs(6134) <= not((layer0_outputs(2970)) and (layer0_outputs(8989)));
    layer1_outputs(6135) <= not(layer0_outputs(57));
    layer1_outputs(6136) <= not(layer0_outputs(9783));
    layer1_outputs(6137) <= not(layer0_outputs(9555));
    layer1_outputs(6138) <= not(layer0_outputs(3126)) or (layer0_outputs(4240));
    layer1_outputs(6139) <= (layer0_outputs(7242)) xor (layer0_outputs(7747));
    layer1_outputs(6140) <= not(layer0_outputs(8157));
    layer1_outputs(6141) <= not(layer0_outputs(3360));
    layer1_outputs(6142) <= not(layer0_outputs(5978));
    layer1_outputs(6143) <= not(layer0_outputs(4131));
    layer1_outputs(6144) <= layer0_outputs(7214);
    layer1_outputs(6145) <= not(layer0_outputs(4514)) or (layer0_outputs(9438));
    layer1_outputs(6146) <= (layer0_outputs(6890)) and not (layer0_outputs(5426));
    layer1_outputs(6147) <= not(layer0_outputs(9776));
    layer1_outputs(6148) <= not(layer0_outputs(5028)) or (layer0_outputs(985));
    layer1_outputs(6149) <= not((layer0_outputs(9124)) and (layer0_outputs(3195)));
    layer1_outputs(6150) <= (layer0_outputs(4247)) and not (layer0_outputs(10156));
    layer1_outputs(6151) <= (layer0_outputs(7663)) and not (layer0_outputs(4436));
    layer1_outputs(6152) <= not(layer0_outputs(1616)) or (layer0_outputs(9986));
    layer1_outputs(6153) <= (layer0_outputs(8177)) xor (layer0_outputs(8645));
    layer1_outputs(6154) <= not(layer0_outputs(5299));
    layer1_outputs(6155) <= not(layer0_outputs(4152));
    layer1_outputs(6156) <= not((layer0_outputs(9882)) and (layer0_outputs(5407)));
    layer1_outputs(6157) <= '0';
    layer1_outputs(6158) <= not(layer0_outputs(10046));
    layer1_outputs(6159) <= (layer0_outputs(2955)) or (layer0_outputs(998));
    layer1_outputs(6160) <= not(layer0_outputs(4731));
    layer1_outputs(6161) <= layer0_outputs(7100);
    layer1_outputs(6162) <= (layer0_outputs(9343)) and (layer0_outputs(8357));
    layer1_outputs(6163) <= layer0_outputs(285);
    layer1_outputs(6164) <= (layer0_outputs(3176)) and not (layer0_outputs(495));
    layer1_outputs(6165) <= layer0_outputs(8951);
    layer1_outputs(6166) <= not(layer0_outputs(3387));
    layer1_outputs(6167) <= not((layer0_outputs(978)) and (layer0_outputs(10199)));
    layer1_outputs(6168) <= not((layer0_outputs(2239)) xor (layer0_outputs(3006)));
    layer1_outputs(6169) <= not((layer0_outputs(7770)) and (layer0_outputs(8093)));
    layer1_outputs(6170) <= not((layer0_outputs(1063)) or (layer0_outputs(736)));
    layer1_outputs(6171) <= not(layer0_outputs(3488)) or (layer0_outputs(5550));
    layer1_outputs(6172) <= layer0_outputs(3452);
    layer1_outputs(6173) <= (layer0_outputs(2628)) and (layer0_outputs(8312));
    layer1_outputs(6174) <= not((layer0_outputs(8671)) or (layer0_outputs(7361)));
    layer1_outputs(6175) <= not(layer0_outputs(2274)) or (layer0_outputs(7819));
    layer1_outputs(6176) <= (layer0_outputs(4533)) and not (layer0_outputs(9415));
    layer1_outputs(6177) <= not((layer0_outputs(4228)) and (layer0_outputs(847)));
    layer1_outputs(6178) <= not(layer0_outputs(5623)) or (layer0_outputs(8837));
    layer1_outputs(6179) <= not(layer0_outputs(4227));
    layer1_outputs(6180) <= not(layer0_outputs(5049)) or (layer0_outputs(8631));
    layer1_outputs(6181) <= not(layer0_outputs(1102)) or (layer0_outputs(1207));
    layer1_outputs(6182) <= '1';
    layer1_outputs(6183) <= not(layer0_outputs(3815));
    layer1_outputs(6184) <= not(layer0_outputs(7916));
    layer1_outputs(6185) <= not(layer0_outputs(2408));
    layer1_outputs(6186) <= not(layer0_outputs(8782));
    layer1_outputs(6187) <= not((layer0_outputs(4245)) and (layer0_outputs(6979)));
    layer1_outputs(6188) <= not(layer0_outputs(7113));
    layer1_outputs(6189) <= not(layer0_outputs(5871));
    layer1_outputs(6190) <= not(layer0_outputs(5925)) or (layer0_outputs(2051));
    layer1_outputs(6191) <= not(layer0_outputs(3041)) or (layer0_outputs(1126));
    layer1_outputs(6192) <= not(layer0_outputs(9779)) or (layer0_outputs(3259));
    layer1_outputs(6193) <= layer0_outputs(5746);
    layer1_outputs(6194) <= not((layer0_outputs(613)) or (layer0_outputs(7780)));
    layer1_outputs(6195) <= not((layer0_outputs(6855)) or (layer0_outputs(3198)));
    layer1_outputs(6196) <= not((layer0_outputs(7564)) or (layer0_outputs(1973)));
    layer1_outputs(6197) <= not(layer0_outputs(7741));
    layer1_outputs(6198) <= (layer0_outputs(5863)) and (layer0_outputs(2921));
    layer1_outputs(6199) <= not(layer0_outputs(692));
    layer1_outputs(6200) <= layer0_outputs(7757);
    layer1_outputs(6201) <= (layer0_outputs(2266)) or (layer0_outputs(4405));
    layer1_outputs(6202) <= (layer0_outputs(7541)) and not (layer0_outputs(8444));
    layer1_outputs(6203) <= not(layer0_outputs(3296));
    layer1_outputs(6204) <= not(layer0_outputs(9245));
    layer1_outputs(6205) <= layer0_outputs(2272);
    layer1_outputs(6206) <= (layer0_outputs(9009)) and not (layer0_outputs(3761));
    layer1_outputs(6207) <= not(layer0_outputs(4681));
    layer1_outputs(6208) <= not((layer0_outputs(1662)) or (layer0_outputs(9203)));
    layer1_outputs(6209) <= not(layer0_outputs(8847));
    layer1_outputs(6210) <= not((layer0_outputs(4066)) and (layer0_outputs(8182)));
    layer1_outputs(6211) <= (layer0_outputs(2622)) and (layer0_outputs(4409));
    layer1_outputs(6212) <= (layer0_outputs(8475)) xor (layer0_outputs(5335));
    layer1_outputs(6213) <= not(layer0_outputs(7866));
    layer1_outputs(6214) <= not(layer0_outputs(7190)) or (layer0_outputs(5206));
    layer1_outputs(6215) <= (layer0_outputs(8042)) or (layer0_outputs(4985));
    layer1_outputs(6216) <= not((layer0_outputs(1910)) or (layer0_outputs(2211)));
    layer1_outputs(6217) <= (layer0_outputs(6837)) and not (layer0_outputs(2786));
    layer1_outputs(6218) <= (layer0_outputs(9969)) or (layer0_outputs(7366));
    layer1_outputs(6219) <= not((layer0_outputs(455)) or (layer0_outputs(9814)));
    layer1_outputs(6220) <= not(layer0_outputs(6744)) or (layer0_outputs(5289));
    layer1_outputs(6221) <= layer0_outputs(2635);
    layer1_outputs(6222) <= layer0_outputs(7370);
    layer1_outputs(6223) <= not(layer0_outputs(1007));
    layer1_outputs(6224) <= not(layer0_outputs(3943));
    layer1_outputs(6225) <= (layer0_outputs(6195)) and not (layer0_outputs(2760));
    layer1_outputs(6226) <= layer0_outputs(8876);
    layer1_outputs(6227) <= not((layer0_outputs(2377)) and (layer0_outputs(8485)));
    layer1_outputs(6228) <= not(layer0_outputs(6574)) or (layer0_outputs(3441));
    layer1_outputs(6229) <= '0';
    layer1_outputs(6230) <= (layer0_outputs(9700)) xor (layer0_outputs(144));
    layer1_outputs(6231) <= layer0_outputs(7486);
    layer1_outputs(6232) <= layer0_outputs(2339);
    layer1_outputs(6233) <= not((layer0_outputs(9273)) and (layer0_outputs(2734)));
    layer1_outputs(6234) <= layer0_outputs(6563);
    layer1_outputs(6235) <= '0';
    layer1_outputs(6236) <= not(layer0_outputs(137));
    layer1_outputs(6237) <= not(layer0_outputs(8247));
    layer1_outputs(6238) <= not(layer0_outputs(3232)) or (layer0_outputs(7143));
    layer1_outputs(6239) <= (layer0_outputs(6043)) xor (layer0_outputs(7417));
    layer1_outputs(6240) <= not((layer0_outputs(5475)) or (layer0_outputs(8174)));
    layer1_outputs(6241) <= (layer0_outputs(211)) and not (layer0_outputs(7311));
    layer1_outputs(6242) <= not((layer0_outputs(9147)) and (layer0_outputs(9873)));
    layer1_outputs(6243) <= (layer0_outputs(1197)) or (layer0_outputs(4754));
    layer1_outputs(6244) <= (layer0_outputs(2511)) and not (layer0_outputs(3360));
    layer1_outputs(6245) <= not((layer0_outputs(1754)) and (layer0_outputs(2447)));
    layer1_outputs(6246) <= '1';
    layer1_outputs(6247) <= layer0_outputs(5801);
    layer1_outputs(6248) <= (layer0_outputs(8145)) and (layer0_outputs(5111));
    layer1_outputs(6249) <= not((layer0_outputs(9311)) and (layer0_outputs(315)));
    layer1_outputs(6250) <= layer0_outputs(2783);
    layer1_outputs(6251) <= (layer0_outputs(6547)) xor (layer0_outputs(5116));
    layer1_outputs(6252) <= layer0_outputs(2604);
    layer1_outputs(6253) <= (layer0_outputs(4291)) xor (layer0_outputs(6275));
    layer1_outputs(6254) <= (layer0_outputs(6944)) xor (layer0_outputs(696));
    layer1_outputs(6255) <= layer0_outputs(3679);
    layer1_outputs(6256) <= not(layer0_outputs(5646));
    layer1_outputs(6257) <= (layer0_outputs(8827)) xor (layer0_outputs(5612));
    layer1_outputs(6258) <= layer0_outputs(3809);
    layer1_outputs(6259) <= (layer0_outputs(471)) and not (layer0_outputs(2255));
    layer1_outputs(6260) <= not(layer0_outputs(8051));
    layer1_outputs(6261) <= (layer0_outputs(2362)) and not (layer0_outputs(3137));
    layer1_outputs(6262) <= not(layer0_outputs(10000)) or (layer0_outputs(2221));
    layer1_outputs(6263) <= (layer0_outputs(1368)) xor (layer0_outputs(1915));
    layer1_outputs(6264) <= not(layer0_outputs(9130));
    layer1_outputs(6265) <= (layer0_outputs(3947)) or (layer0_outputs(5089));
    layer1_outputs(6266) <= not(layer0_outputs(5983)) or (layer0_outputs(8195));
    layer1_outputs(6267) <= not(layer0_outputs(3915)) or (layer0_outputs(4207));
    layer1_outputs(6268) <= not((layer0_outputs(7244)) and (layer0_outputs(5695)));
    layer1_outputs(6269) <= (layer0_outputs(9270)) and not (layer0_outputs(7633));
    layer1_outputs(6270) <= layer0_outputs(6746);
    layer1_outputs(6271) <= layer0_outputs(7340);
    layer1_outputs(6272) <= '1';
    layer1_outputs(6273) <= (layer0_outputs(9095)) and not (layer0_outputs(9069));
    layer1_outputs(6274) <= '1';
    layer1_outputs(6275) <= (layer0_outputs(3533)) xor (layer0_outputs(8592));
    layer1_outputs(6276) <= layer0_outputs(1139);
    layer1_outputs(6277) <= not(layer0_outputs(7086));
    layer1_outputs(6278) <= (layer0_outputs(7857)) xor (layer0_outputs(1056));
    layer1_outputs(6279) <= not(layer0_outputs(2986));
    layer1_outputs(6280) <= not(layer0_outputs(6429)) or (layer0_outputs(4769));
    layer1_outputs(6281) <= not((layer0_outputs(4194)) or (layer0_outputs(683)));
    layer1_outputs(6282) <= layer0_outputs(5068);
    layer1_outputs(6283) <= not((layer0_outputs(4347)) or (layer0_outputs(6356)));
    layer1_outputs(6284) <= not(layer0_outputs(2847));
    layer1_outputs(6285) <= not(layer0_outputs(5505)) or (layer0_outputs(1167));
    layer1_outputs(6286) <= not(layer0_outputs(1416)) or (layer0_outputs(3944));
    layer1_outputs(6287) <= (layer0_outputs(6502)) and not (layer0_outputs(3485));
    layer1_outputs(6288) <= layer0_outputs(7647);
    layer1_outputs(6289) <= not(layer0_outputs(4239)) or (layer0_outputs(7764));
    layer1_outputs(6290) <= (layer0_outputs(4251)) and not (layer0_outputs(1836));
    layer1_outputs(6291) <= layer0_outputs(43);
    layer1_outputs(6292) <= (layer0_outputs(8327)) and not (layer0_outputs(3967));
    layer1_outputs(6293) <= (layer0_outputs(9228)) or (layer0_outputs(3677));
    layer1_outputs(6294) <= not((layer0_outputs(5068)) and (layer0_outputs(6638)));
    layer1_outputs(6295) <= (layer0_outputs(6680)) and (layer0_outputs(2350));
    layer1_outputs(6296) <= '0';
    layer1_outputs(6297) <= not(layer0_outputs(2237));
    layer1_outputs(6298) <= (layer0_outputs(7692)) or (layer0_outputs(949));
    layer1_outputs(6299) <= (layer0_outputs(9725)) xor (layer0_outputs(9751));
    layer1_outputs(6300) <= (layer0_outputs(4596)) and (layer0_outputs(4576));
    layer1_outputs(6301) <= not((layer0_outputs(8552)) xor (layer0_outputs(4970)));
    layer1_outputs(6302) <= (layer0_outputs(2365)) and not (layer0_outputs(4880));
    layer1_outputs(6303) <= not((layer0_outputs(1082)) and (layer0_outputs(5274)));
    layer1_outputs(6304) <= not((layer0_outputs(260)) or (layer0_outputs(4323)));
    layer1_outputs(6305) <= layer0_outputs(9179);
    layer1_outputs(6306) <= layer0_outputs(4349);
    layer1_outputs(6307) <= not((layer0_outputs(3443)) and (layer0_outputs(6940)));
    layer1_outputs(6308) <= not(layer0_outputs(3764)) or (layer0_outputs(119));
    layer1_outputs(6309) <= (layer0_outputs(9601)) or (layer0_outputs(6129));
    layer1_outputs(6310) <= not((layer0_outputs(5635)) or (layer0_outputs(9390)));
    layer1_outputs(6311) <= not((layer0_outputs(5651)) and (layer0_outputs(278)));
    layer1_outputs(6312) <= not(layer0_outputs(6057));
    layer1_outputs(6313) <= (layer0_outputs(8063)) and not (layer0_outputs(6231));
    layer1_outputs(6314) <= not(layer0_outputs(4284));
    layer1_outputs(6315) <= layer0_outputs(3051);
    layer1_outputs(6316) <= not((layer0_outputs(189)) or (layer0_outputs(5734)));
    layer1_outputs(6317) <= '0';
    layer1_outputs(6318) <= layer0_outputs(10018);
    layer1_outputs(6319) <= layer0_outputs(454);
    layer1_outputs(6320) <= (layer0_outputs(8026)) or (layer0_outputs(1992));
    layer1_outputs(6321) <= layer0_outputs(5674);
    layer1_outputs(6322) <= not(layer0_outputs(9422)) or (layer0_outputs(619));
    layer1_outputs(6323) <= (layer0_outputs(630)) and not (layer0_outputs(2718));
    layer1_outputs(6324) <= (layer0_outputs(8783)) and not (layer0_outputs(7620));
    layer1_outputs(6325) <= (layer0_outputs(1317)) or (layer0_outputs(6584));
    layer1_outputs(6326) <= layer0_outputs(6890);
    layer1_outputs(6327) <= not(layer0_outputs(1079)) or (layer0_outputs(196));
    layer1_outputs(6328) <= layer0_outputs(7895);
    layer1_outputs(6329) <= not((layer0_outputs(4551)) and (layer0_outputs(5233)));
    layer1_outputs(6330) <= (layer0_outputs(6800)) and not (layer0_outputs(7046));
    layer1_outputs(6331) <= (layer0_outputs(3365)) or (layer0_outputs(4909));
    layer1_outputs(6332) <= layer0_outputs(3056);
    layer1_outputs(6333) <= (layer0_outputs(272)) and not (layer0_outputs(5619));
    layer1_outputs(6334) <= not(layer0_outputs(9150));
    layer1_outputs(6335) <= layer0_outputs(6232);
    layer1_outputs(6336) <= not(layer0_outputs(7547)) or (layer0_outputs(6292));
    layer1_outputs(6337) <= not(layer0_outputs(9425));
    layer1_outputs(6338) <= not(layer0_outputs(600));
    layer1_outputs(6339) <= not((layer0_outputs(6254)) xor (layer0_outputs(373)));
    layer1_outputs(6340) <= (layer0_outputs(2596)) xor (layer0_outputs(4033));
    layer1_outputs(6341) <= not(layer0_outputs(1264));
    layer1_outputs(6342) <= not(layer0_outputs(5970));
    layer1_outputs(6343) <= (layer0_outputs(2989)) and (layer0_outputs(9651));
    layer1_outputs(6344) <= not((layer0_outputs(7515)) and (layer0_outputs(3600)));
    layer1_outputs(6345) <= layer0_outputs(9720);
    layer1_outputs(6346) <= (layer0_outputs(9752)) and (layer0_outputs(3296));
    layer1_outputs(6347) <= not(layer0_outputs(6841));
    layer1_outputs(6348) <= '1';
    layer1_outputs(6349) <= not(layer0_outputs(8456)) or (layer0_outputs(6796));
    layer1_outputs(6350) <= layer0_outputs(10146);
    layer1_outputs(6351) <= layer0_outputs(7437);
    layer1_outputs(6352) <= not(layer0_outputs(7636)) or (layer0_outputs(4273));
    layer1_outputs(6353) <= not(layer0_outputs(3996));
    layer1_outputs(6354) <= layer0_outputs(4597);
    layer1_outputs(6355) <= layer0_outputs(2664);
    layer1_outputs(6356) <= layer0_outputs(5927);
    layer1_outputs(6357) <= not(layer0_outputs(1098)) or (layer0_outputs(5593));
    layer1_outputs(6358) <= not((layer0_outputs(0)) and (layer0_outputs(10211)));
    layer1_outputs(6359) <= not(layer0_outputs(4230));
    layer1_outputs(6360) <= '0';
    layer1_outputs(6361) <= layer0_outputs(6098);
    layer1_outputs(6362) <= (layer0_outputs(2574)) and (layer0_outputs(4286));
    layer1_outputs(6363) <= (layer0_outputs(1023)) and not (layer0_outputs(9260));
    layer1_outputs(6364) <= (layer0_outputs(3200)) and not (layer0_outputs(10105));
    layer1_outputs(6365) <= (layer0_outputs(7342)) and not (layer0_outputs(5754));
    layer1_outputs(6366) <= (layer0_outputs(8392)) xor (layer0_outputs(7696));
    layer1_outputs(6367) <= not(layer0_outputs(3400)) or (layer0_outputs(1968));
    layer1_outputs(6368) <= not(layer0_outputs(8670));
    layer1_outputs(6369) <= not(layer0_outputs(555)) or (layer0_outputs(4968));
    layer1_outputs(6370) <= not(layer0_outputs(4373)) or (layer0_outputs(4248));
    layer1_outputs(6371) <= not((layer0_outputs(4709)) and (layer0_outputs(3026)));
    layer1_outputs(6372) <= (layer0_outputs(2638)) or (layer0_outputs(4796));
    layer1_outputs(6373) <= layer0_outputs(9016);
    layer1_outputs(6374) <= (layer0_outputs(7332)) and (layer0_outputs(4989));
    layer1_outputs(6375) <= not(layer0_outputs(5572));
    layer1_outputs(6376) <= not((layer0_outputs(2202)) xor (layer0_outputs(1772)));
    layer1_outputs(6377) <= (layer0_outputs(7869)) and not (layer0_outputs(7551));
    layer1_outputs(6378) <= not(layer0_outputs(9547));
    layer1_outputs(6379) <= layer0_outputs(2870);
    layer1_outputs(6380) <= not(layer0_outputs(9344));
    layer1_outputs(6381) <= layer0_outputs(4515);
    layer1_outputs(6382) <= layer0_outputs(7272);
    layer1_outputs(6383) <= not(layer0_outputs(6919));
    layer1_outputs(6384) <= layer0_outputs(7386);
    layer1_outputs(6385) <= not(layer0_outputs(9495)) or (layer0_outputs(5082));
    layer1_outputs(6386) <= layer0_outputs(8621);
    layer1_outputs(6387) <= layer0_outputs(6785);
    layer1_outputs(6388) <= layer0_outputs(10194);
    layer1_outputs(6389) <= layer0_outputs(7301);
    layer1_outputs(6390) <= not(layer0_outputs(7340));
    layer1_outputs(6391) <= not(layer0_outputs(7300));
    layer1_outputs(6392) <= not(layer0_outputs(1954));
    layer1_outputs(6393) <= not(layer0_outputs(3498));
    layer1_outputs(6394) <= '0';
    layer1_outputs(6395) <= (layer0_outputs(7434)) and (layer0_outputs(831));
    layer1_outputs(6396) <= not(layer0_outputs(3384)) or (layer0_outputs(8176));
    layer1_outputs(6397) <= layer0_outputs(381);
    layer1_outputs(6398) <= (layer0_outputs(6535)) and (layer0_outputs(3740));
    layer1_outputs(6399) <= (layer0_outputs(3450)) and not (layer0_outputs(9463));
    layer1_outputs(6400) <= (layer0_outputs(4613)) and (layer0_outputs(1664));
    layer1_outputs(6401) <= layer0_outputs(113);
    layer1_outputs(6402) <= not((layer0_outputs(4495)) xor (layer0_outputs(7423)));
    layer1_outputs(6403) <= (layer0_outputs(1600)) xor (layer0_outputs(4955));
    layer1_outputs(6404) <= (layer0_outputs(9694)) xor (layer0_outputs(2168));
    layer1_outputs(6405) <= '1';
    layer1_outputs(6406) <= layer0_outputs(7469);
    layer1_outputs(6407) <= not(layer0_outputs(8465)) or (layer0_outputs(4167));
    layer1_outputs(6408) <= not(layer0_outputs(1904));
    layer1_outputs(6409) <= layer0_outputs(8342);
    layer1_outputs(6410) <= not(layer0_outputs(406));
    layer1_outputs(6411) <= not(layer0_outputs(8339)) or (layer0_outputs(7191));
    layer1_outputs(6412) <= (layer0_outputs(7778)) or (layer0_outputs(7881));
    layer1_outputs(6413) <= not((layer0_outputs(6140)) or (layer0_outputs(6807)));
    layer1_outputs(6414) <= not((layer0_outputs(8652)) and (layer0_outputs(2865)));
    layer1_outputs(6415) <= not(layer0_outputs(7005));
    layer1_outputs(6416) <= (layer0_outputs(4128)) and (layer0_outputs(7753));
    layer1_outputs(6417) <= layer0_outputs(9324);
    layer1_outputs(6418) <= not(layer0_outputs(5633));
    layer1_outputs(6419) <= (layer0_outputs(3766)) and not (layer0_outputs(6282));
    layer1_outputs(6420) <= not(layer0_outputs(7289));
    layer1_outputs(6421) <= layer0_outputs(8644);
    layer1_outputs(6422) <= not((layer0_outputs(5075)) and (layer0_outputs(3740)));
    layer1_outputs(6423) <= not(layer0_outputs(8177)) or (layer0_outputs(7412));
    layer1_outputs(6424) <= layer0_outputs(7436);
    layer1_outputs(6425) <= layer0_outputs(6698);
    layer1_outputs(6426) <= (layer0_outputs(4612)) and not (layer0_outputs(1392));
    layer1_outputs(6427) <= (layer0_outputs(4394)) and not (layer0_outputs(6082));
    layer1_outputs(6428) <= layer0_outputs(3165);
    layer1_outputs(6429) <= not((layer0_outputs(9263)) and (layer0_outputs(6947)));
    layer1_outputs(6430) <= not(layer0_outputs(6608));
    layer1_outputs(6431) <= (layer0_outputs(3592)) and not (layer0_outputs(3791));
    layer1_outputs(6432) <= layer0_outputs(6019);
    layer1_outputs(6433) <= not((layer0_outputs(10020)) and (layer0_outputs(9907)));
    layer1_outputs(6434) <= not(layer0_outputs(3658));
    layer1_outputs(6435) <= layer0_outputs(1445);
    layer1_outputs(6436) <= not(layer0_outputs(9559));
    layer1_outputs(6437) <= '1';
    layer1_outputs(6438) <= '1';
    layer1_outputs(6439) <= layer0_outputs(7368);
    layer1_outputs(6440) <= layer0_outputs(491);
    layer1_outputs(6441) <= not(layer0_outputs(6988)) or (layer0_outputs(9892));
    layer1_outputs(6442) <= not(layer0_outputs(6082));
    layer1_outputs(6443) <= (layer0_outputs(868)) and not (layer0_outputs(5543));
    layer1_outputs(6444) <= not((layer0_outputs(2608)) and (layer0_outputs(129)));
    layer1_outputs(6445) <= not((layer0_outputs(1447)) and (layer0_outputs(1114)));
    layer1_outputs(6446) <= (layer0_outputs(3872)) or (layer0_outputs(1186));
    layer1_outputs(6447) <= not((layer0_outputs(2851)) and (layer0_outputs(9374)));
    layer1_outputs(6448) <= not(layer0_outputs(4460)) or (layer0_outputs(8045));
    layer1_outputs(6449) <= not(layer0_outputs(282));
    layer1_outputs(6450) <= not(layer0_outputs(3963)) or (layer0_outputs(4069));
    layer1_outputs(6451) <= layer0_outputs(9105);
    layer1_outputs(6452) <= (layer0_outputs(6586)) and not (layer0_outputs(1551));
    layer1_outputs(6453) <= '0';
    layer1_outputs(6454) <= '0';
    layer1_outputs(6455) <= layer0_outputs(5009);
    layer1_outputs(6456) <= not(layer0_outputs(9347));
    layer1_outputs(6457) <= layer0_outputs(1912);
    layer1_outputs(6458) <= layer0_outputs(1125);
    layer1_outputs(6459) <= layer0_outputs(2408);
    layer1_outputs(6460) <= not((layer0_outputs(1962)) or (layer0_outputs(5276)));
    layer1_outputs(6461) <= (layer0_outputs(161)) or (layer0_outputs(10004));
    layer1_outputs(6462) <= not(layer0_outputs(6596));
    layer1_outputs(6463) <= (layer0_outputs(563)) and not (layer0_outputs(8763));
    layer1_outputs(6464) <= not((layer0_outputs(3156)) and (layer0_outputs(5595)));
    layer1_outputs(6465) <= layer0_outputs(9843);
    layer1_outputs(6466) <= (layer0_outputs(7890)) or (layer0_outputs(8360));
    layer1_outputs(6467) <= not(layer0_outputs(1960)) or (layer0_outputs(3463));
    layer1_outputs(6468) <= not(layer0_outputs(9965));
    layer1_outputs(6469) <= not(layer0_outputs(3440)) or (layer0_outputs(4483));
    layer1_outputs(6470) <= not(layer0_outputs(813)) or (layer0_outputs(3770));
    layer1_outputs(6471) <= not(layer0_outputs(4852));
    layer1_outputs(6472) <= layer0_outputs(5465);
    layer1_outputs(6473) <= layer0_outputs(498);
    layer1_outputs(6474) <= '1';
    layer1_outputs(6475) <= not(layer0_outputs(7344));
    layer1_outputs(6476) <= (layer0_outputs(6393)) and (layer0_outputs(7444));
    layer1_outputs(6477) <= not(layer0_outputs(6245));
    layer1_outputs(6478) <= (layer0_outputs(2946)) xor (layer0_outputs(1557));
    layer1_outputs(6479) <= not(layer0_outputs(9028));
    layer1_outputs(6480) <= (layer0_outputs(3907)) xor (layer0_outputs(5407));
    layer1_outputs(6481) <= not((layer0_outputs(9813)) or (layer0_outputs(4707)));
    layer1_outputs(6482) <= (layer0_outputs(9050)) or (layer0_outputs(1091));
    layer1_outputs(6483) <= not(layer0_outputs(8764));
    layer1_outputs(6484) <= (layer0_outputs(1265)) or (layer0_outputs(8098));
    layer1_outputs(6485) <= not(layer0_outputs(4050)) or (layer0_outputs(7736));
    layer1_outputs(6486) <= layer0_outputs(2265);
    layer1_outputs(6487) <= layer0_outputs(2364);
    layer1_outputs(6488) <= not((layer0_outputs(5438)) or (layer0_outputs(2440)));
    layer1_outputs(6489) <= '1';
    layer1_outputs(6490) <= (layer0_outputs(9790)) xor (layer0_outputs(4079));
    layer1_outputs(6491) <= not(layer0_outputs(8571));
    layer1_outputs(6492) <= (layer0_outputs(5694)) and not (layer0_outputs(756));
    layer1_outputs(6493) <= not(layer0_outputs(1194)) or (layer0_outputs(3432));
    layer1_outputs(6494) <= layer0_outputs(4096);
    layer1_outputs(6495) <= layer0_outputs(147);
    layer1_outputs(6496) <= (layer0_outputs(6373)) and not (layer0_outputs(8872));
    layer1_outputs(6497) <= layer0_outputs(5400);
    layer1_outputs(6498) <= not((layer0_outputs(8721)) xor (layer0_outputs(5800)));
    layer1_outputs(6499) <= layer0_outputs(1862);
    layer1_outputs(6500) <= not((layer0_outputs(2603)) and (layer0_outputs(7908)));
    layer1_outputs(6501) <= not(layer0_outputs(10230));
    layer1_outputs(6502) <= layer0_outputs(9450);
    layer1_outputs(6503) <= '1';
    layer1_outputs(6504) <= layer0_outputs(1582);
    layer1_outputs(6505) <= (layer0_outputs(2381)) and not (layer0_outputs(5629));
    layer1_outputs(6506) <= not(layer0_outputs(4101)) or (layer0_outputs(8248));
    layer1_outputs(6507) <= layer0_outputs(1686);
    layer1_outputs(6508) <= not(layer0_outputs(1785));
    layer1_outputs(6509) <= layer0_outputs(5841);
    layer1_outputs(6510) <= not((layer0_outputs(4906)) or (layer0_outputs(2502)));
    layer1_outputs(6511) <= not(layer0_outputs(3651));
    layer1_outputs(6512) <= not(layer0_outputs(8041));
    layer1_outputs(6513) <= not((layer0_outputs(3613)) and (layer0_outputs(9810)));
    layer1_outputs(6514) <= not(layer0_outputs(3855));
    layer1_outputs(6515) <= not((layer0_outputs(241)) xor (layer0_outputs(3257)));
    layer1_outputs(6516) <= layer0_outputs(8455);
    layer1_outputs(6517) <= not((layer0_outputs(1131)) and (layer0_outputs(6220)));
    layer1_outputs(6518) <= not(layer0_outputs(6095));
    layer1_outputs(6519) <= (layer0_outputs(8564)) xor (layer0_outputs(2843));
    layer1_outputs(6520) <= not((layer0_outputs(4731)) xor (layer0_outputs(9442)));
    layer1_outputs(6521) <= (layer0_outputs(2601)) and (layer0_outputs(543));
    layer1_outputs(6522) <= layer0_outputs(3253);
    layer1_outputs(6523) <= layer0_outputs(1781);
    layer1_outputs(6524) <= (layer0_outputs(8259)) or (layer0_outputs(383));
    layer1_outputs(6525) <= not((layer0_outputs(4174)) and (layer0_outputs(4708)));
    layer1_outputs(6526) <= (layer0_outputs(6856)) and not (layer0_outputs(8051));
    layer1_outputs(6527) <= not(layer0_outputs(2688)) or (layer0_outputs(8004));
    layer1_outputs(6528) <= layer0_outputs(4261);
    layer1_outputs(6529) <= layer0_outputs(6968);
    layer1_outputs(6530) <= not((layer0_outputs(1214)) or (layer0_outputs(7027)));
    layer1_outputs(6531) <= (layer0_outputs(486)) and (layer0_outputs(6149));
    layer1_outputs(6532) <= (layer0_outputs(9776)) and (layer0_outputs(5223));
    layer1_outputs(6533) <= '0';
    layer1_outputs(6534) <= not((layer0_outputs(270)) or (layer0_outputs(8299)));
    layer1_outputs(6535) <= (layer0_outputs(9138)) and not (layer0_outputs(1596));
    layer1_outputs(6536) <= layer0_outputs(2804);
    layer1_outputs(6537) <= not((layer0_outputs(6131)) or (layer0_outputs(6927)));
    layer1_outputs(6538) <= (layer0_outputs(4804)) or (layer0_outputs(3847));
    layer1_outputs(6539) <= layer0_outputs(8551);
    layer1_outputs(6540) <= not(layer0_outputs(2627)) or (layer0_outputs(6089));
    layer1_outputs(6541) <= not(layer0_outputs(9019));
    layer1_outputs(6542) <= layer0_outputs(8722);
    layer1_outputs(6543) <= '0';
    layer1_outputs(6544) <= not(layer0_outputs(2953)) or (layer0_outputs(9286));
    layer1_outputs(6545) <= not(layer0_outputs(7690)) or (layer0_outputs(9609));
    layer1_outputs(6546) <= not(layer0_outputs(3376));
    layer1_outputs(6547) <= layer0_outputs(1552);
    layer1_outputs(6548) <= not(layer0_outputs(5016));
    layer1_outputs(6549) <= not(layer0_outputs(7114));
    layer1_outputs(6550) <= not(layer0_outputs(793));
    layer1_outputs(6551) <= layer0_outputs(1480);
    layer1_outputs(6552) <= (layer0_outputs(7282)) and not (layer0_outputs(4794));
    layer1_outputs(6553) <= (layer0_outputs(3395)) xor (layer0_outputs(1569));
    layer1_outputs(6554) <= not((layer0_outputs(3871)) or (layer0_outputs(3046)));
    layer1_outputs(6555) <= layer0_outputs(7437);
    layer1_outputs(6556) <= (layer0_outputs(6730)) and (layer0_outputs(8436));
    layer1_outputs(6557) <= (layer0_outputs(9358)) or (layer0_outputs(7285));
    layer1_outputs(6558) <= layer0_outputs(4053);
    layer1_outputs(6559) <= (layer0_outputs(6330)) and (layer0_outputs(6344));
    layer1_outputs(6560) <= not(layer0_outputs(8158));
    layer1_outputs(6561) <= not(layer0_outputs(946));
    layer1_outputs(6562) <= not((layer0_outputs(3071)) xor (layer0_outputs(3566)));
    layer1_outputs(6563) <= layer0_outputs(9002);
    layer1_outputs(6564) <= not(layer0_outputs(9678));
    layer1_outputs(6565) <= layer0_outputs(9218);
    layer1_outputs(6566) <= not(layer0_outputs(5061)) or (layer0_outputs(10117));
    layer1_outputs(6567) <= not((layer0_outputs(6592)) and (layer0_outputs(2698)));
    layer1_outputs(6568) <= not((layer0_outputs(1182)) or (layer0_outputs(4629)));
    layer1_outputs(6569) <= not(layer0_outputs(10030));
    layer1_outputs(6570) <= not(layer0_outputs(8591)) or (layer0_outputs(1501));
    layer1_outputs(6571) <= (layer0_outputs(4868)) and not (layer0_outputs(9372));
    layer1_outputs(6572) <= layer0_outputs(1588);
    layer1_outputs(6573) <= not((layer0_outputs(5383)) or (layer0_outputs(4963)));
    layer1_outputs(6574) <= layer0_outputs(594);
    layer1_outputs(6575) <= not((layer0_outputs(4702)) xor (layer0_outputs(5351)));
    layer1_outputs(6576) <= '1';
    layer1_outputs(6577) <= (layer0_outputs(632)) and not (layer0_outputs(6512));
    layer1_outputs(6578) <= (layer0_outputs(3106)) xor (layer0_outputs(10083));
    layer1_outputs(6579) <= (layer0_outputs(9518)) or (layer0_outputs(2096));
    layer1_outputs(6580) <= not(layer0_outputs(7421));
    layer1_outputs(6581) <= not(layer0_outputs(9661)) or (layer0_outputs(8050));
    layer1_outputs(6582) <= (layer0_outputs(3126)) and not (layer0_outputs(7183));
    layer1_outputs(6583) <= layer0_outputs(231);
    layer1_outputs(6584) <= not(layer0_outputs(9298));
    layer1_outputs(6585) <= layer0_outputs(5560);
    layer1_outputs(6586) <= '1';
    layer1_outputs(6587) <= not(layer0_outputs(9686));
    layer1_outputs(6588) <= not(layer0_outputs(6680));
    layer1_outputs(6589) <= (layer0_outputs(8431)) and (layer0_outputs(8319));
    layer1_outputs(6590) <= not(layer0_outputs(1462)) or (layer0_outputs(5906));
    layer1_outputs(6591) <= (layer0_outputs(2057)) xor (layer0_outputs(4275));
    layer1_outputs(6592) <= not(layer0_outputs(2824));
    layer1_outputs(6593) <= not(layer0_outputs(8289));
    layer1_outputs(6594) <= not(layer0_outputs(7810)) or (layer0_outputs(2260));
    layer1_outputs(6595) <= not(layer0_outputs(1561));
    layer1_outputs(6596) <= (layer0_outputs(4472)) or (layer0_outputs(1));
    layer1_outputs(6597) <= (layer0_outputs(4730)) and not (layer0_outputs(8977));
    layer1_outputs(6598) <= not(layer0_outputs(9217)) or (layer0_outputs(2040));
    layer1_outputs(6599) <= (layer0_outputs(6998)) and (layer0_outputs(2855));
    layer1_outputs(6600) <= layer0_outputs(240);
    layer1_outputs(6601) <= not(layer0_outputs(1248)) or (layer0_outputs(2351));
    layer1_outputs(6602) <= '1';
    layer1_outputs(6603) <= not(layer0_outputs(5816));
    layer1_outputs(6604) <= not(layer0_outputs(3970)) or (layer0_outputs(3065));
    layer1_outputs(6605) <= (layer0_outputs(3676)) and not (layer0_outputs(4680));
    layer1_outputs(6606) <= not((layer0_outputs(4562)) or (layer0_outputs(5975)));
    layer1_outputs(6607) <= not((layer0_outputs(8931)) or (layer0_outputs(3386)));
    layer1_outputs(6608) <= not(layer0_outputs(515)) or (layer0_outputs(5122));
    layer1_outputs(6609) <= not(layer0_outputs(6275)) or (layer0_outputs(8085));
    layer1_outputs(6610) <= not(layer0_outputs(3390)) or (layer0_outputs(4947));
    layer1_outputs(6611) <= layer0_outputs(8231);
    layer1_outputs(6612) <= not(layer0_outputs(4219)) or (layer0_outputs(8729));
    layer1_outputs(6613) <= not(layer0_outputs(4487));
    layer1_outputs(6614) <= (layer0_outputs(399)) or (layer0_outputs(1823));
    layer1_outputs(6615) <= layer0_outputs(6318);
    layer1_outputs(6616) <= layer0_outputs(6564);
    layer1_outputs(6617) <= (layer0_outputs(6013)) and not (layer0_outputs(8640));
    layer1_outputs(6618) <= (layer0_outputs(3382)) or (layer0_outputs(3573));
    layer1_outputs(6619) <= not(layer0_outputs(4356)) or (layer0_outputs(2032));
    layer1_outputs(6620) <= not(layer0_outputs(6622)) or (layer0_outputs(9340));
    layer1_outputs(6621) <= not(layer0_outputs(3329)) or (layer0_outputs(5912));
    layer1_outputs(6622) <= (layer0_outputs(8916)) or (layer0_outputs(7642));
    layer1_outputs(6623) <= (layer0_outputs(5675)) and not (layer0_outputs(3141));
    layer1_outputs(6624) <= (layer0_outputs(2831)) xor (layer0_outputs(2651));
    layer1_outputs(6625) <= (layer0_outputs(2138)) and not (layer0_outputs(8121));
    layer1_outputs(6626) <= (layer0_outputs(9515)) and not (layer0_outputs(3434));
    layer1_outputs(6627) <= not((layer0_outputs(3073)) and (layer0_outputs(9078)));
    layer1_outputs(6628) <= not(layer0_outputs(5548));
    layer1_outputs(6629) <= not(layer0_outputs(8772));
    layer1_outputs(6630) <= not(layer0_outputs(3997));
    layer1_outputs(6631) <= not((layer0_outputs(2917)) or (layer0_outputs(6480)));
    layer1_outputs(6632) <= layer0_outputs(2311);
    layer1_outputs(6633) <= (layer0_outputs(648)) or (layer0_outputs(3330));
    layer1_outputs(6634) <= layer0_outputs(8535);
    layer1_outputs(6635) <= (layer0_outputs(6773)) and (layer0_outputs(6012));
    layer1_outputs(6636) <= not(layer0_outputs(2859));
    layer1_outputs(6637) <= not(layer0_outputs(932)) or (layer0_outputs(9330));
    layer1_outputs(6638) <= (layer0_outputs(9910)) or (layer0_outputs(3055));
    layer1_outputs(6639) <= layer0_outputs(1908);
    layer1_outputs(6640) <= not(layer0_outputs(3246));
    layer1_outputs(6641) <= (layer0_outputs(7905)) and not (layer0_outputs(10191));
    layer1_outputs(6642) <= not(layer0_outputs(2072));
    layer1_outputs(6643) <= not(layer0_outputs(8047));
    layer1_outputs(6644) <= not(layer0_outputs(8179));
    layer1_outputs(6645) <= (layer0_outputs(9693)) and not (layer0_outputs(4353));
    layer1_outputs(6646) <= (layer0_outputs(1640)) or (layer0_outputs(10191));
    layer1_outputs(6647) <= layer0_outputs(3818);
    layer1_outputs(6648) <= '1';
    layer1_outputs(6649) <= layer0_outputs(419);
    layer1_outputs(6650) <= (layer0_outputs(2627)) and not (layer0_outputs(6083));
    layer1_outputs(6651) <= (layer0_outputs(5357)) or (layer0_outputs(7292));
    layer1_outputs(6652) <= layer0_outputs(1329);
    layer1_outputs(6653) <= (layer0_outputs(6781)) or (layer0_outputs(3415));
    layer1_outputs(6654) <= layer0_outputs(4633);
    layer1_outputs(6655) <= layer0_outputs(8990);
    layer1_outputs(6656) <= (layer0_outputs(3852)) and not (layer0_outputs(3001));
    layer1_outputs(6657) <= (layer0_outputs(8398)) xor (layer0_outputs(1831));
    layer1_outputs(6658) <= (layer0_outputs(7814)) or (layer0_outputs(1864));
    layer1_outputs(6659) <= not(layer0_outputs(8094));
    layer1_outputs(6660) <= not((layer0_outputs(5311)) and (layer0_outputs(8493)));
    layer1_outputs(6661) <= layer0_outputs(8057);
    layer1_outputs(6662) <= not(layer0_outputs(578));
    layer1_outputs(6663) <= layer0_outputs(7400);
    layer1_outputs(6664) <= not(layer0_outputs(1876));
    layer1_outputs(6665) <= layer0_outputs(9661);
    layer1_outputs(6666) <= not(layer0_outputs(9822)) or (layer0_outputs(4351));
    layer1_outputs(6667) <= (layer0_outputs(4987)) and not (layer0_outputs(9766));
    layer1_outputs(6668) <= layer0_outputs(588);
    layer1_outputs(6669) <= not(layer0_outputs(946));
    layer1_outputs(6670) <= not(layer0_outputs(8073));
    layer1_outputs(6671) <= not((layer0_outputs(806)) xor (layer0_outputs(2345)));
    layer1_outputs(6672) <= (layer0_outputs(3049)) and not (layer0_outputs(6162));
    layer1_outputs(6673) <= not(layer0_outputs(8870)) or (layer0_outputs(1650));
    layer1_outputs(6674) <= not(layer0_outputs(9030));
    layer1_outputs(6675) <= layer0_outputs(9011);
    layer1_outputs(6676) <= '1';
    layer1_outputs(6677) <= not((layer0_outputs(1403)) or (layer0_outputs(4153)));
    layer1_outputs(6678) <= layer0_outputs(9131);
    layer1_outputs(6679) <= (layer0_outputs(3024)) and (layer0_outputs(3934));
    layer1_outputs(6680) <= not((layer0_outputs(1222)) xor (layer0_outputs(8313)));
    layer1_outputs(6681) <= not(layer0_outputs(7273));
    layer1_outputs(6682) <= (layer0_outputs(9616)) or (layer0_outputs(6115));
    layer1_outputs(6683) <= not(layer0_outputs(2149)) or (layer0_outputs(8672));
    layer1_outputs(6684) <= (layer0_outputs(4220)) and not (layer0_outputs(392));
    layer1_outputs(6685) <= (layer0_outputs(3821)) and (layer0_outputs(5416));
    layer1_outputs(6686) <= not(layer0_outputs(7531)) or (layer0_outputs(10153));
    layer1_outputs(6687) <= '1';
    layer1_outputs(6688) <= (layer0_outputs(1505)) or (layer0_outputs(420));
    layer1_outputs(6689) <= not((layer0_outputs(5798)) and (layer0_outputs(7142)));
    layer1_outputs(6690) <= not(layer0_outputs(8384)) or (layer0_outputs(6121));
    layer1_outputs(6691) <= not((layer0_outputs(8397)) and (layer0_outputs(4790)));
    layer1_outputs(6692) <= not(layer0_outputs(2713)) or (layer0_outputs(6915));
    layer1_outputs(6693) <= not(layer0_outputs(8812));
    layer1_outputs(6694) <= not(layer0_outputs(645));
    layer1_outputs(6695) <= not(layer0_outputs(1174));
    layer1_outputs(6696) <= not((layer0_outputs(6875)) and (layer0_outputs(3590)));
    layer1_outputs(6697) <= not((layer0_outputs(8985)) xor (layer0_outputs(3970)));
    layer1_outputs(6698) <= '1';
    layer1_outputs(6699) <= (layer0_outputs(2942)) xor (layer0_outputs(2350));
    layer1_outputs(6700) <= layer0_outputs(8171);
    layer1_outputs(6701) <= (layer0_outputs(150)) or (layer0_outputs(9692));
    layer1_outputs(6702) <= not(layer0_outputs(405)) or (layer0_outputs(8582));
    layer1_outputs(6703) <= layer0_outputs(3020);
    layer1_outputs(6704) <= (layer0_outputs(8654)) or (layer0_outputs(7856));
    layer1_outputs(6705) <= '1';
    layer1_outputs(6706) <= not(layer0_outputs(5638)) or (layer0_outputs(8422));
    layer1_outputs(6707) <= layer0_outputs(4746);
    layer1_outputs(6708) <= layer0_outputs(1880);
    layer1_outputs(6709) <= (layer0_outputs(8828)) and not (layer0_outputs(1298));
    layer1_outputs(6710) <= not(layer0_outputs(9628)) or (layer0_outputs(3541));
    layer1_outputs(6711) <= (layer0_outputs(9085)) and (layer0_outputs(1393));
    layer1_outputs(6712) <= '0';
    layer1_outputs(6713) <= not(layer0_outputs(9491));
    layer1_outputs(6714) <= layer0_outputs(9848);
    layer1_outputs(6715) <= (layer0_outputs(3843)) and (layer0_outputs(9713));
    layer1_outputs(6716) <= (layer0_outputs(9079)) xor (layer0_outputs(7813));
    layer1_outputs(6717) <= not(layer0_outputs(3952)) or (layer0_outputs(7687));
    layer1_outputs(6718) <= not(layer0_outputs(10043));
    layer1_outputs(6719) <= not(layer0_outputs(8550));
    layer1_outputs(6720) <= not(layer0_outputs(6190));
    layer1_outputs(6721) <= (layer0_outputs(2588)) xor (layer0_outputs(7901));
    layer1_outputs(6722) <= (layer0_outputs(1214)) and not (layer0_outputs(1805));
    layer1_outputs(6723) <= not(layer0_outputs(2091));
    layer1_outputs(6724) <= '1';
    layer1_outputs(6725) <= not(layer0_outputs(3252));
    layer1_outputs(6726) <= layer0_outputs(2332);
    layer1_outputs(6727) <= not((layer0_outputs(3956)) or (layer0_outputs(530)));
    layer1_outputs(6728) <= not(layer0_outputs(4438));
    layer1_outputs(6729) <= not(layer0_outputs(50));
    layer1_outputs(6730) <= layer0_outputs(5924);
    layer1_outputs(6731) <= (layer0_outputs(1549)) and not (layer0_outputs(2968));
    layer1_outputs(6732) <= not(layer0_outputs(5233)) or (layer0_outputs(4732));
    layer1_outputs(6733) <= layer0_outputs(4672);
    layer1_outputs(6734) <= layer0_outputs(9211);
    layer1_outputs(6735) <= layer0_outputs(203);
    layer1_outputs(6736) <= not(layer0_outputs(3800));
    layer1_outputs(6737) <= not((layer0_outputs(2454)) and (layer0_outputs(4889)));
    layer1_outputs(6738) <= layer0_outputs(1150);
    layer1_outputs(6739) <= (layer0_outputs(6864)) and not (layer0_outputs(4321));
    layer1_outputs(6740) <= not(layer0_outputs(10135)) or (layer0_outputs(10186));
    layer1_outputs(6741) <= (layer0_outputs(2769)) and not (layer0_outputs(1558));
    layer1_outputs(6742) <= not(layer0_outputs(3233));
    layer1_outputs(6743) <= '0';
    layer1_outputs(6744) <= layer0_outputs(9664);
    layer1_outputs(6745) <= not((layer0_outputs(7148)) and (layer0_outputs(517)));
    layer1_outputs(6746) <= not((layer0_outputs(6218)) and (layer0_outputs(5515)));
    layer1_outputs(6747) <= layer0_outputs(5327);
    layer1_outputs(6748) <= '1';
    layer1_outputs(6749) <= layer0_outputs(5843);
    layer1_outputs(6750) <= layer0_outputs(10007);
    layer1_outputs(6751) <= (layer0_outputs(296)) or (layer0_outputs(2827));
    layer1_outputs(6752) <= not(layer0_outputs(125));
    layer1_outputs(6753) <= not(layer0_outputs(7981));
    layer1_outputs(6754) <= (layer0_outputs(1598)) or (layer0_outputs(5160));
    layer1_outputs(6755) <= (layer0_outputs(2182)) and not (layer0_outputs(5643));
    layer1_outputs(6756) <= not(layer0_outputs(8976));
    layer1_outputs(6757) <= layer0_outputs(5618);
    layer1_outputs(6758) <= not(layer0_outputs(8068)) or (layer0_outputs(845));
    layer1_outputs(6759) <= not(layer0_outputs(1691));
    layer1_outputs(6760) <= not(layer0_outputs(8548)) or (layer0_outputs(6567));
    layer1_outputs(6761) <= not(layer0_outputs(5810));
    layer1_outputs(6762) <= layer0_outputs(3107);
    layer1_outputs(6763) <= not(layer0_outputs(257));
    layer1_outputs(6764) <= (layer0_outputs(3111)) and (layer0_outputs(4157));
    layer1_outputs(6765) <= not(layer0_outputs(3896));
    layer1_outputs(6766) <= layer0_outputs(7480);
    layer1_outputs(6767) <= not((layer0_outputs(5485)) xor (layer0_outputs(5257)));
    layer1_outputs(6768) <= (layer0_outputs(1697)) and not (layer0_outputs(5358));
    layer1_outputs(6769) <= '0';
    layer1_outputs(6770) <= not((layer0_outputs(7024)) xor (layer0_outputs(2391)));
    layer1_outputs(6771) <= not(layer0_outputs(5153));
    layer1_outputs(6772) <= not(layer0_outputs(6209));
    layer1_outputs(6773) <= (layer0_outputs(7345)) and not (layer0_outputs(3791));
    layer1_outputs(6774) <= (layer0_outputs(7206)) and not (layer0_outputs(803));
    layer1_outputs(6775) <= (layer0_outputs(2372)) and (layer0_outputs(9489));
    layer1_outputs(6776) <= (layer0_outputs(3866)) xor (layer0_outputs(1246));
    layer1_outputs(6777) <= not(layer0_outputs(8183));
    layer1_outputs(6778) <= layer0_outputs(908);
    layer1_outputs(6779) <= (layer0_outputs(558)) or (layer0_outputs(3917));
    layer1_outputs(6780) <= not(layer0_outputs(7702)) or (layer0_outputs(85));
    layer1_outputs(6781) <= not((layer0_outputs(7830)) or (layer0_outputs(3405)));
    layer1_outputs(6782) <= not(layer0_outputs(6661)) or (layer0_outputs(2515));
    layer1_outputs(6783) <= not(layer0_outputs(7874));
    layer1_outputs(6784) <= not(layer0_outputs(4713));
    layer1_outputs(6785) <= not(layer0_outputs(1389)) or (layer0_outputs(4940));
    layer1_outputs(6786) <= not(layer0_outputs(824));
    layer1_outputs(6787) <= (layer0_outputs(1514)) or (layer0_outputs(4658));
    layer1_outputs(6788) <= not(layer0_outputs(9366)) or (layer0_outputs(9334));
    layer1_outputs(6789) <= not(layer0_outputs(3962));
    layer1_outputs(6790) <= not(layer0_outputs(8319)) or (layer0_outputs(3634));
    layer1_outputs(6791) <= layer0_outputs(2771);
    layer1_outputs(6792) <= not(layer0_outputs(7684)) or (layer0_outputs(5005));
    layer1_outputs(6793) <= (layer0_outputs(8129)) xor (layer0_outputs(9611));
    layer1_outputs(6794) <= not((layer0_outputs(5344)) or (layer0_outputs(3993)));
    layer1_outputs(6795) <= (layer0_outputs(3895)) and not (layer0_outputs(6337));
    layer1_outputs(6796) <= (layer0_outputs(8774)) or (layer0_outputs(3394));
    layer1_outputs(6797) <= not(layer0_outputs(10115)) or (layer0_outputs(7333));
    layer1_outputs(6798) <= not(layer0_outputs(2389));
    layer1_outputs(6799) <= layer0_outputs(2208);
    layer1_outputs(6800) <= not((layer0_outputs(8906)) xor (layer0_outputs(7740)));
    layer1_outputs(6801) <= not(layer0_outputs(9621)) or (layer0_outputs(5763));
    layer1_outputs(6802) <= not((layer0_outputs(3352)) or (layer0_outputs(729)));
    layer1_outputs(6803) <= not(layer0_outputs(7941));
    layer1_outputs(6804) <= not(layer0_outputs(2274)) or (layer0_outputs(7277));
    layer1_outputs(6805) <= not((layer0_outputs(3202)) and (layer0_outputs(9744)));
    layer1_outputs(6806) <= not((layer0_outputs(2984)) or (layer0_outputs(4269)));
    layer1_outputs(6807) <= not((layer0_outputs(4785)) or (layer0_outputs(5578)));
    layer1_outputs(6808) <= (layer0_outputs(5796)) and not (layer0_outputs(3916));
    layer1_outputs(6809) <= not(layer0_outputs(440));
    layer1_outputs(6810) <= (layer0_outputs(6741)) xor (layer0_outputs(7967));
    layer1_outputs(6811) <= (layer0_outputs(1323)) xor (layer0_outputs(3823));
    layer1_outputs(6812) <= layer0_outputs(3980);
    layer1_outputs(6813) <= not((layer0_outputs(3879)) and (layer0_outputs(10169)));
    layer1_outputs(6814) <= not(layer0_outputs(1217)) or (layer0_outputs(4433));
    layer1_outputs(6815) <= not(layer0_outputs(3651)) or (layer0_outputs(6136));
    layer1_outputs(6816) <= not(layer0_outputs(6870));
    layer1_outputs(6817) <= (layer0_outputs(9380)) xor (layer0_outputs(8136));
    layer1_outputs(6818) <= not(layer0_outputs(2130));
    layer1_outputs(6819) <= not((layer0_outputs(4322)) and (layer0_outputs(953)));
    layer1_outputs(6820) <= not(layer0_outputs(9732));
    layer1_outputs(6821) <= not(layer0_outputs(6091)) or (layer0_outputs(8756));
    layer1_outputs(6822) <= layer0_outputs(5878);
    layer1_outputs(6823) <= not(layer0_outputs(9587)) or (layer0_outputs(571));
    layer1_outputs(6824) <= '0';
    layer1_outputs(6825) <= not(layer0_outputs(3901));
    layer1_outputs(6826) <= (layer0_outputs(805)) and (layer0_outputs(2464));
    layer1_outputs(6827) <= not(layer0_outputs(577));
    layer1_outputs(6828) <= layer0_outputs(3444);
    layer1_outputs(6829) <= not((layer0_outputs(9207)) or (layer0_outputs(4994)));
    layer1_outputs(6830) <= layer0_outputs(9193);
    layer1_outputs(6831) <= layer0_outputs(4616);
    layer1_outputs(6832) <= '1';
    layer1_outputs(6833) <= not(layer0_outputs(7949)) or (layer0_outputs(6373));
    layer1_outputs(6834) <= not((layer0_outputs(8293)) or (layer0_outputs(610)));
    layer1_outputs(6835) <= not(layer0_outputs(5711)) or (layer0_outputs(2089));
    layer1_outputs(6836) <= layer0_outputs(1658);
    layer1_outputs(6837) <= layer0_outputs(7027);
    layer1_outputs(6838) <= not(layer0_outputs(542));
    layer1_outputs(6839) <= layer0_outputs(5546);
    layer1_outputs(6840) <= (layer0_outputs(3123)) xor (layer0_outputs(8682));
    layer1_outputs(6841) <= not((layer0_outputs(7247)) and (layer0_outputs(1808)));
    layer1_outputs(6842) <= not(layer0_outputs(10105));
    layer1_outputs(6843) <= (layer0_outputs(5001)) or (layer0_outputs(7985));
    layer1_outputs(6844) <= not(layer0_outputs(3209)) or (layer0_outputs(2034));
    layer1_outputs(6845) <= not(layer0_outputs(9763));
    layer1_outputs(6846) <= not((layer0_outputs(3978)) and (layer0_outputs(3169)));
    layer1_outputs(6847) <= (layer0_outputs(2595)) or (layer0_outputs(10066));
    layer1_outputs(6848) <= layer0_outputs(5806);
    layer1_outputs(6849) <= (layer0_outputs(2429)) and not (layer0_outputs(796));
    layer1_outputs(6850) <= not((layer0_outputs(7664)) or (layer0_outputs(10162)));
    layer1_outputs(6851) <= not(layer0_outputs(5177));
    layer1_outputs(6852) <= layer0_outputs(3562);
    layer1_outputs(6853) <= not(layer0_outputs(34)) or (layer0_outputs(3214));
    layer1_outputs(6854) <= (layer0_outputs(718)) xor (layer0_outputs(2176));
    layer1_outputs(6855) <= not(layer0_outputs(5151));
    layer1_outputs(6856) <= not((layer0_outputs(4118)) xor (layer0_outputs(7418)));
    layer1_outputs(6857) <= not(layer0_outputs(1347)) or (layer0_outputs(61));
    layer1_outputs(6858) <= layer0_outputs(1269);
    layer1_outputs(6859) <= layer0_outputs(4952);
    layer1_outputs(6860) <= not(layer0_outputs(1264));
    layer1_outputs(6861) <= (layer0_outputs(2619)) and (layer0_outputs(8332));
    layer1_outputs(6862) <= not((layer0_outputs(8463)) or (layer0_outputs(3677)));
    layer1_outputs(6863) <= (layer0_outputs(8107)) and not (layer0_outputs(9348));
    layer1_outputs(6864) <= not(layer0_outputs(7883)) or (layer0_outputs(8575));
    layer1_outputs(6865) <= (layer0_outputs(6728)) and not (layer0_outputs(523));
    layer1_outputs(6866) <= not(layer0_outputs(8491));
    layer1_outputs(6867) <= layer0_outputs(625);
    layer1_outputs(6868) <= layer0_outputs(8946);
    layer1_outputs(6869) <= layer0_outputs(1991);
    layer1_outputs(6870) <= layer0_outputs(234);
    layer1_outputs(6871) <= (layer0_outputs(5879)) and not (layer0_outputs(6418));
    layer1_outputs(6872) <= layer0_outputs(6414);
    layer1_outputs(6873) <= not((layer0_outputs(9904)) xor (layer0_outputs(9178)));
    layer1_outputs(6874) <= (layer0_outputs(9562)) and not (layer0_outputs(10238));
    layer1_outputs(6875) <= not(layer0_outputs(2757));
    layer1_outputs(6876) <= not(layer0_outputs(4382));
    layer1_outputs(6877) <= layer0_outputs(10127);
    layer1_outputs(6878) <= (layer0_outputs(726)) and not (layer0_outputs(5804));
    layer1_outputs(6879) <= layer0_outputs(400);
    layer1_outputs(6880) <= not((layer0_outputs(9632)) and (layer0_outputs(5439)));
    layer1_outputs(6881) <= (layer0_outputs(8347)) and not (layer0_outputs(9447));
    layer1_outputs(6882) <= layer0_outputs(4611);
    layer1_outputs(6883) <= not(layer0_outputs(9898));
    layer1_outputs(6884) <= not(layer0_outputs(671));
    layer1_outputs(6885) <= not(layer0_outputs(5419));
    layer1_outputs(6886) <= layer0_outputs(1052);
    layer1_outputs(6887) <= (layer0_outputs(9092)) and not (layer0_outputs(3888));
    layer1_outputs(6888) <= layer0_outputs(8314);
    layer1_outputs(6889) <= (layer0_outputs(2655)) and not (layer0_outputs(6124));
    layer1_outputs(6890) <= not(layer0_outputs(2608)) or (layer0_outputs(8729));
    layer1_outputs(6891) <= (layer0_outputs(3794)) or (layer0_outputs(4049));
    layer1_outputs(6892) <= not((layer0_outputs(2953)) or (layer0_outputs(5730)));
    layer1_outputs(6893) <= layer0_outputs(1148);
    layer1_outputs(6894) <= not(layer0_outputs(1856));
    layer1_outputs(6895) <= (layer0_outputs(3586)) or (layer0_outputs(1668));
    layer1_outputs(6896) <= not(layer0_outputs(1879));
    layer1_outputs(6897) <= not((layer0_outputs(1052)) or (layer0_outputs(7628)));
    layer1_outputs(6898) <= (layer0_outputs(9273)) and not (layer0_outputs(5429));
    layer1_outputs(6899) <= layer0_outputs(1206);
    layer1_outputs(6900) <= layer0_outputs(9739);
    layer1_outputs(6901) <= (layer0_outputs(5490)) and not (layer0_outputs(9066));
    layer1_outputs(6902) <= (layer0_outputs(2963)) and not (layer0_outputs(860));
    layer1_outputs(6903) <= (layer0_outputs(2025)) and (layer0_outputs(5682));
    layer1_outputs(6904) <= layer0_outputs(7721);
    layer1_outputs(6905) <= not(layer0_outputs(7007)) or (layer0_outputs(745));
    layer1_outputs(6906) <= '0';
    layer1_outputs(6907) <= not(layer0_outputs(2726));
    layer1_outputs(6908) <= not((layer0_outputs(5279)) and (layer0_outputs(3753)));
    layer1_outputs(6909) <= layer0_outputs(6567);
    layer1_outputs(6910) <= not((layer0_outputs(1613)) and (layer0_outputs(2667)));
    layer1_outputs(6911) <= layer0_outputs(9391);
    layer1_outputs(6912) <= layer0_outputs(7931);
    layer1_outputs(6913) <= (layer0_outputs(6263)) and (layer0_outputs(3466));
    layer1_outputs(6914) <= not(layer0_outputs(4846));
    layer1_outputs(6915) <= layer0_outputs(3560);
    layer1_outputs(6916) <= layer0_outputs(2083);
    layer1_outputs(6917) <= not(layer0_outputs(7896));
    layer1_outputs(6918) <= not(layer0_outputs(2962)) or (layer0_outputs(8510));
    layer1_outputs(6919) <= not(layer0_outputs(9101));
    layer1_outputs(6920) <= not(layer0_outputs(4671)) or (layer0_outputs(62));
    layer1_outputs(6921) <= (layer0_outputs(7452)) and not (layer0_outputs(4630));
    layer1_outputs(6922) <= '1';
    layer1_outputs(6923) <= (layer0_outputs(267)) or (layer0_outputs(8546));
    layer1_outputs(6924) <= not((layer0_outputs(59)) and (layer0_outputs(4572)));
    layer1_outputs(6925) <= (layer0_outputs(4473)) or (layer0_outputs(7639));
    layer1_outputs(6926) <= not((layer0_outputs(7818)) and (layer0_outputs(1950)));
    layer1_outputs(6927) <= not(layer0_outputs(9289));
    layer1_outputs(6928) <= not(layer0_outputs(487)) or (layer0_outputs(7566));
    layer1_outputs(6929) <= layer0_outputs(1944);
    layer1_outputs(6930) <= layer0_outputs(6440);
    layer1_outputs(6931) <= not((layer0_outputs(5790)) or (layer0_outputs(9643)));
    layer1_outputs(6932) <= not(layer0_outputs(850));
    layer1_outputs(6933) <= (layer0_outputs(5704)) or (layer0_outputs(3536));
    layer1_outputs(6934) <= not(layer0_outputs(7125));
    layer1_outputs(6935) <= '1';
    layer1_outputs(6936) <= not((layer0_outputs(7984)) xor (layer0_outputs(329)));
    layer1_outputs(6937) <= layer0_outputs(9578);
    layer1_outputs(6938) <= layer0_outputs(6852);
    layer1_outputs(6939) <= not((layer0_outputs(9675)) and (layer0_outputs(140)));
    layer1_outputs(6940) <= not(layer0_outputs(3099));
    layer1_outputs(6941) <= not(layer0_outputs(3089)) or (layer0_outputs(9021));
    layer1_outputs(6942) <= layer0_outputs(8042);
    layer1_outputs(6943) <= not((layer0_outputs(2702)) xor (layer0_outputs(7224)));
    layer1_outputs(6944) <= (layer0_outputs(2002)) and not (layer0_outputs(7559));
    layer1_outputs(6945) <= not(layer0_outputs(1235));
    layer1_outputs(6946) <= not(layer0_outputs(512));
    layer1_outputs(6947) <= layer0_outputs(3069);
    layer1_outputs(6948) <= layer0_outputs(8751);
    layer1_outputs(6949) <= (layer0_outputs(1911)) and not (layer0_outputs(2356));
    layer1_outputs(6950) <= (layer0_outputs(1564)) and not (layer0_outputs(4196));
    layer1_outputs(6951) <= layer0_outputs(8938);
    layer1_outputs(6952) <= not(layer0_outputs(4593));
    layer1_outputs(6953) <= not((layer0_outputs(3726)) xor (layer0_outputs(10121)));
    layer1_outputs(6954) <= not(layer0_outputs(3850));
    layer1_outputs(6955) <= layer0_outputs(6024);
    layer1_outputs(6956) <= not(layer0_outputs(8308)) or (layer0_outputs(1299));
    layer1_outputs(6957) <= (layer0_outputs(5045)) xor (layer0_outputs(4004));
    layer1_outputs(6958) <= not(layer0_outputs(1838));
    layer1_outputs(6959) <= layer0_outputs(4182);
    layer1_outputs(6960) <= (layer0_outputs(2258)) and not (layer0_outputs(721));
    layer1_outputs(6961) <= not((layer0_outputs(8329)) and (layer0_outputs(1240)));
    layer1_outputs(6962) <= layer0_outputs(9006);
    layer1_outputs(6963) <= not((layer0_outputs(6483)) xor (layer0_outputs(1084)));
    layer1_outputs(6964) <= layer0_outputs(660);
    layer1_outputs(6965) <= not((layer0_outputs(4923)) and (layer0_outputs(2525)));
    layer1_outputs(6966) <= not(layer0_outputs(124));
    layer1_outputs(6967) <= (layer0_outputs(6962)) or (layer0_outputs(800));
    layer1_outputs(6968) <= not((layer0_outputs(8048)) or (layer0_outputs(1300)));
    layer1_outputs(6969) <= not(layer0_outputs(14)) or (layer0_outputs(7675));
    layer1_outputs(6970) <= not(layer0_outputs(5282));
    layer1_outputs(6971) <= not(layer0_outputs(5862));
    layer1_outputs(6972) <= (layer0_outputs(4192)) and not (layer0_outputs(8348));
    layer1_outputs(6973) <= not(layer0_outputs(8198)) or (layer0_outputs(4574));
    layer1_outputs(6974) <= '0';
    layer1_outputs(6975) <= (layer0_outputs(5335)) or (layer0_outputs(3583));
    layer1_outputs(6976) <= (layer0_outputs(6215)) and not (layer0_outputs(6928));
    layer1_outputs(6977) <= (layer0_outputs(5176)) and (layer0_outputs(5700));
    layer1_outputs(6978) <= (layer0_outputs(6556)) xor (layer0_outputs(1361));
    layer1_outputs(6979) <= not(layer0_outputs(3927)) or (layer0_outputs(7195));
    layer1_outputs(6980) <= not((layer0_outputs(1051)) xor (layer0_outputs(3320)));
    layer1_outputs(6981) <= not(layer0_outputs(8483));
    layer1_outputs(6982) <= (layer0_outputs(260)) xor (layer0_outputs(1111));
    layer1_outputs(6983) <= (layer0_outputs(6433)) or (layer0_outputs(8440));
    layer1_outputs(6984) <= layer0_outputs(9771);
    layer1_outputs(6985) <= not(layer0_outputs(3695));
    layer1_outputs(6986) <= not(layer0_outputs(2211));
    layer1_outputs(6987) <= layer0_outputs(7312);
    layer1_outputs(6988) <= (layer0_outputs(9547)) and not (layer0_outputs(7854));
    layer1_outputs(6989) <= not(layer0_outputs(7982));
    layer1_outputs(6990) <= not((layer0_outputs(7584)) and (layer0_outputs(9406)));
    layer1_outputs(6991) <= layer0_outputs(4714);
    layer1_outputs(6992) <= not(layer0_outputs(4563)) or (layer0_outputs(3903));
    layer1_outputs(6993) <= (layer0_outputs(7925)) and not (layer0_outputs(344));
    layer1_outputs(6994) <= not(layer0_outputs(5591));
    layer1_outputs(6995) <= (layer0_outputs(8513)) and (layer0_outputs(3183));
    layer1_outputs(6996) <= layer0_outputs(5208);
    layer1_outputs(6997) <= not(layer0_outputs(4593)) or (layer0_outputs(8315));
    layer1_outputs(6998) <= not((layer0_outputs(4493)) and (layer0_outputs(8264)));
    layer1_outputs(6999) <= layer0_outputs(1548);
    layer1_outputs(7000) <= not(layer0_outputs(2022));
    layer1_outputs(7001) <= not((layer0_outputs(2166)) or (layer0_outputs(7529)));
    layer1_outputs(7002) <= '0';
    layer1_outputs(7003) <= not((layer0_outputs(4823)) and (layer0_outputs(3990)));
    layer1_outputs(7004) <= not(layer0_outputs(293)) or (layer0_outputs(5989));
    layer1_outputs(7005) <= not((layer0_outputs(8313)) xor (layer0_outputs(1814)));
    layer1_outputs(7006) <= (layer0_outputs(2193)) and not (layer0_outputs(4111));
    layer1_outputs(7007) <= not(layer0_outputs(5818));
    layer1_outputs(7008) <= (layer0_outputs(7425)) and not (layer0_outputs(6977));
    layer1_outputs(7009) <= not(layer0_outputs(8630)) or (layer0_outputs(6636));
    layer1_outputs(7010) <= (layer0_outputs(2891)) xor (layer0_outputs(7907));
    layer1_outputs(7011) <= not(layer0_outputs(1464));
    layer1_outputs(7012) <= not(layer0_outputs(3028));
    layer1_outputs(7013) <= layer0_outputs(1874);
    layer1_outputs(7014) <= (layer0_outputs(386)) and (layer0_outputs(2585));
    layer1_outputs(7015) <= layer0_outputs(6339);
    layer1_outputs(7016) <= not(layer0_outputs(6100)) or (layer0_outputs(6386));
    layer1_outputs(7017) <= not(layer0_outputs(753));
    layer1_outputs(7018) <= layer0_outputs(2912);
    layer1_outputs(7019) <= not(layer0_outputs(9031));
    layer1_outputs(7020) <= not(layer0_outputs(8210));
    layer1_outputs(7021) <= not(layer0_outputs(4726)) or (layer0_outputs(4551));
    layer1_outputs(7022) <= not(layer0_outputs(8625)) or (layer0_outputs(3871));
    layer1_outputs(7023) <= layer0_outputs(1335);
    layer1_outputs(7024) <= (layer0_outputs(3190)) xor (layer0_outputs(5949));
    layer1_outputs(7025) <= not(layer0_outputs(4262));
    layer1_outputs(7026) <= not(layer0_outputs(7411));
    layer1_outputs(7027) <= not((layer0_outputs(5778)) or (layer0_outputs(4073)));
    layer1_outputs(7028) <= not((layer0_outputs(3990)) or (layer0_outputs(6002)));
    layer1_outputs(7029) <= layer0_outputs(8003);
    layer1_outputs(7030) <= not((layer0_outputs(1369)) xor (layer0_outputs(8889)));
    layer1_outputs(7031) <= not((layer0_outputs(999)) xor (layer0_outputs(8642)));
    layer1_outputs(7032) <= (layer0_outputs(2057)) xor (layer0_outputs(4876));
    layer1_outputs(7033) <= (layer0_outputs(4377)) and (layer0_outputs(5458));
    layer1_outputs(7034) <= layer0_outputs(4670);
    layer1_outputs(7035) <= not((layer0_outputs(31)) or (layer0_outputs(9130)));
    layer1_outputs(7036) <= not((layer0_outputs(7964)) and (layer0_outputs(7595)));
    layer1_outputs(7037) <= (layer0_outputs(1184)) and not (layer0_outputs(7212));
    layer1_outputs(7038) <= not(layer0_outputs(1310));
    layer1_outputs(7039) <= not(layer0_outputs(2903));
    layer1_outputs(7040) <= not(layer0_outputs(1892)) or (layer0_outputs(470));
    layer1_outputs(7041) <= layer0_outputs(7904);
    layer1_outputs(7042) <= not(layer0_outputs(2205));
    layer1_outputs(7043) <= not((layer0_outputs(335)) or (layer0_outputs(7884)));
    layer1_outputs(7044) <= layer0_outputs(9709);
    layer1_outputs(7045) <= not(layer0_outputs(9557));
    layer1_outputs(7046) <= layer0_outputs(1326);
    layer1_outputs(7047) <= (layer0_outputs(2936)) xor (layer0_outputs(2947));
    layer1_outputs(7048) <= not((layer0_outputs(6246)) and (layer0_outputs(7256)));
    layer1_outputs(7049) <= not(layer0_outputs(4574));
    layer1_outputs(7050) <= (layer0_outputs(5937)) and (layer0_outputs(133));
    layer1_outputs(7051) <= not((layer0_outputs(8203)) and (layer0_outputs(4258)));
    layer1_outputs(7052) <= not(layer0_outputs(9964));
    layer1_outputs(7053) <= not(layer0_outputs(8273));
    layer1_outputs(7054) <= not(layer0_outputs(5952));
    layer1_outputs(7055) <= not(layer0_outputs(346));
    layer1_outputs(7056) <= (layer0_outputs(1289)) and not (layer0_outputs(9673));
    layer1_outputs(7057) <= not((layer0_outputs(3606)) and (layer0_outputs(5687)));
    layer1_outputs(7058) <= (layer0_outputs(4316)) xor (layer0_outputs(9319));
    layer1_outputs(7059) <= layer0_outputs(10008);
    layer1_outputs(7060) <= (layer0_outputs(4632)) and not (layer0_outputs(2839));
    layer1_outputs(7061) <= layer0_outputs(1653);
    layer1_outputs(7062) <= layer0_outputs(6925);
    layer1_outputs(7063) <= (layer0_outputs(583)) xor (layer0_outputs(5499));
    layer1_outputs(7064) <= '0';
    layer1_outputs(7065) <= not(layer0_outputs(8162)) or (layer0_outputs(489));
    layer1_outputs(7066) <= not(layer0_outputs(1110)) or (layer0_outputs(788));
    layer1_outputs(7067) <= (layer0_outputs(3724)) xor (layer0_outputs(4549));
    layer1_outputs(7068) <= not(layer0_outputs(1448));
    layer1_outputs(7069) <= not((layer0_outputs(4656)) xor (layer0_outputs(3754)));
    layer1_outputs(7070) <= not(layer0_outputs(9516));
    layer1_outputs(7071) <= (layer0_outputs(961)) or (layer0_outputs(5639));
    layer1_outputs(7072) <= not((layer0_outputs(7227)) or (layer0_outputs(9284)));
    layer1_outputs(7073) <= (layer0_outputs(139)) and not (layer0_outputs(5732));
    layer1_outputs(7074) <= (layer0_outputs(3604)) and not (layer0_outputs(7259));
    layer1_outputs(7075) <= not(layer0_outputs(5771));
    layer1_outputs(7076) <= not(layer0_outputs(7104)) or (layer0_outputs(6588));
    layer1_outputs(7077) <= not(layer0_outputs(3712)) or (layer0_outputs(1930));
    layer1_outputs(7078) <= not(layer0_outputs(1526));
    layer1_outputs(7079) <= not(layer0_outputs(9156));
    layer1_outputs(7080) <= (layer0_outputs(6595)) and not (layer0_outputs(6449));
    layer1_outputs(7081) <= (layer0_outputs(1493)) and not (layer0_outputs(1193));
    layer1_outputs(7082) <= layer0_outputs(8123);
    layer1_outputs(7083) <= (layer0_outputs(909)) xor (layer0_outputs(4777));
    layer1_outputs(7084) <= not(layer0_outputs(9394)) or (layer0_outputs(9620));
    layer1_outputs(7085) <= (layer0_outputs(7357)) and not (layer0_outputs(706));
    layer1_outputs(7086) <= not(layer0_outputs(5985)) or (layer0_outputs(3109));
    layer1_outputs(7087) <= not(layer0_outputs(554));
    layer1_outputs(7088) <= not(layer0_outputs(4762));
    layer1_outputs(7089) <= layer0_outputs(9871);
    layer1_outputs(7090) <= (layer0_outputs(3719)) and not (layer0_outputs(557));
    layer1_outputs(7091) <= (layer0_outputs(4173)) xor (layer0_outputs(7163));
    layer1_outputs(7092) <= (layer0_outputs(1382)) or (layer0_outputs(5660));
    layer1_outputs(7093) <= (layer0_outputs(2292)) and not (layer0_outputs(9343));
    layer1_outputs(7094) <= not(layer0_outputs(9794));
    layer1_outputs(7095) <= '0';
    layer1_outputs(7096) <= layer0_outputs(2282);
    layer1_outputs(7097) <= not(layer0_outputs(7012));
    layer1_outputs(7098) <= layer0_outputs(6424);
    layer1_outputs(7099) <= layer0_outputs(199);
    layer1_outputs(7100) <= layer0_outputs(6205);
    layer1_outputs(7101) <= (layer0_outputs(955)) and (layer0_outputs(9556));
    layer1_outputs(7102) <= not(layer0_outputs(1946));
    layer1_outputs(7103) <= layer0_outputs(2508);
    layer1_outputs(7104) <= layer0_outputs(5058);
    layer1_outputs(7105) <= not(layer0_outputs(4404));
    layer1_outputs(7106) <= '0';
    layer1_outputs(7107) <= not(layer0_outputs(6117)) or (layer0_outputs(5600));
    layer1_outputs(7108) <= layer0_outputs(2334);
    layer1_outputs(7109) <= (layer0_outputs(4608)) and (layer0_outputs(9032));
    layer1_outputs(7110) <= layer0_outputs(4243);
    layer1_outputs(7111) <= (layer0_outputs(497)) and (layer0_outputs(2070));
    layer1_outputs(7112) <= not(layer0_outputs(6482));
    layer1_outputs(7113) <= not(layer0_outputs(2499));
    layer1_outputs(7114) <= (layer0_outputs(1330)) and not (layer0_outputs(5278));
    layer1_outputs(7115) <= (layer0_outputs(4974)) or (layer0_outputs(1356));
    layer1_outputs(7116) <= (layer0_outputs(1041)) or (layer0_outputs(7116));
    layer1_outputs(7117) <= (layer0_outputs(3275)) and (layer0_outputs(4338));
    layer1_outputs(7118) <= layer0_outputs(3982);
    layer1_outputs(7119) <= not((layer0_outputs(8636)) xor (layer0_outputs(8690)));
    layer1_outputs(7120) <= not((layer0_outputs(10103)) or (layer0_outputs(4195)));
    layer1_outputs(7121) <= not(layer0_outputs(2238));
    layer1_outputs(7122) <= layer0_outputs(9364);
    layer1_outputs(7123) <= (layer0_outputs(7995)) and not (layer0_outputs(6159));
    layer1_outputs(7124) <= not((layer0_outputs(6812)) and (layer0_outputs(646)));
    layer1_outputs(7125) <= (layer0_outputs(7080)) and (layer0_outputs(4637));
    layer1_outputs(7126) <= not((layer0_outputs(8613)) and (layer0_outputs(10104)));
    layer1_outputs(7127) <= layer0_outputs(9522);
    layer1_outputs(7128) <= '1';
    layer1_outputs(7129) <= layer0_outputs(7697);
    layer1_outputs(7130) <= not(layer0_outputs(3175));
    layer1_outputs(7131) <= (layer0_outputs(5953)) xor (layer0_outputs(8004));
    layer1_outputs(7132) <= not((layer0_outputs(3500)) and (layer0_outputs(4374)));
    layer1_outputs(7133) <= not((layer0_outputs(10106)) or (layer0_outputs(6941)));
    layer1_outputs(7134) <= layer0_outputs(1270);
    layer1_outputs(7135) <= not(layer0_outputs(5277));
    layer1_outputs(7136) <= layer0_outputs(461);
    layer1_outputs(7137) <= not(layer0_outputs(5116)) or (layer0_outputs(951));
    layer1_outputs(7138) <= '0';
    layer1_outputs(7139) <= (layer0_outputs(2453)) and not (layer0_outputs(4679));
    layer1_outputs(7140) <= (layer0_outputs(6568)) and not (layer0_outputs(1566));
    layer1_outputs(7141) <= not((layer0_outputs(4534)) or (layer0_outputs(9595)));
    layer1_outputs(7142) <= layer0_outputs(8773);
    layer1_outputs(7143) <= (layer0_outputs(1219)) or (layer0_outputs(6457));
    layer1_outputs(7144) <= layer0_outputs(520);
    layer1_outputs(7145) <= not(layer0_outputs(8263)) or (layer0_outputs(3229));
    layer1_outputs(7146) <= not(layer0_outputs(9351)) or (layer0_outputs(6284));
    layer1_outputs(7147) <= not((layer0_outputs(9444)) or (layer0_outputs(5088)));
    layer1_outputs(7148) <= not(layer0_outputs(741)) or (layer0_outputs(2617));
    layer1_outputs(7149) <= not(layer0_outputs(5235));
    layer1_outputs(7150) <= not((layer0_outputs(280)) or (layer0_outputs(7527)));
    layer1_outputs(7151) <= layer0_outputs(5648);
    layer1_outputs(7152) <= not(layer0_outputs(3240)) or (layer0_outputs(6251));
    layer1_outputs(7153) <= (layer0_outputs(1905)) or (layer0_outputs(21));
    layer1_outputs(7154) <= layer0_outputs(4751);
    layer1_outputs(7155) <= not(layer0_outputs(3166));
    layer1_outputs(7156) <= (layer0_outputs(2799)) or (layer0_outputs(7419));
    layer1_outputs(7157) <= (layer0_outputs(5140)) and (layer0_outputs(4881));
    layer1_outputs(7158) <= not(layer0_outputs(1608)) or (layer0_outputs(2134));
    layer1_outputs(7159) <= not((layer0_outputs(388)) or (layer0_outputs(2064)));
    layer1_outputs(7160) <= not((layer0_outputs(6631)) or (layer0_outputs(2133)));
    layer1_outputs(7161) <= layer0_outputs(8159);
    layer1_outputs(7162) <= not(layer0_outputs(9454));
    layer1_outputs(7163) <= not(layer0_outputs(1027)) or (layer0_outputs(4774));
    layer1_outputs(7164) <= not(layer0_outputs(2436)) or (layer0_outputs(2331));
    layer1_outputs(7165) <= layer0_outputs(6365);
    layer1_outputs(7166) <= not(layer0_outputs(4604)) or (layer0_outputs(8589));
    layer1_outputs(7167) <= not((layer0_outputs(3254)) and (layer0_outputs(5144)));
    layer1_outputs(7168) <= (layer0_outputs(4818)) and not (layer0_outputs(8154));
    layer1_outputs(7169) <= layer0_outputs(9431);
    layer1_outputs(7170) <= not(layer0_outputs(6684)) or (layer0_outputs(3159));
    layer1_outputs(7171) <= layer0_outputs(4472);
    layer1_outputs(7172) <= (layer0_outputs(1244)) and (layer0_outputs(7274));
    layer1_outputs(7173) <= layer0_outputs(4700);
    layer1_outputs(7174) <= not(layer0_outputs(3848));
    layer1_outputs(7175) <= layer0_outputs(6495);
    layer1_outputs(7176) <= not(layer0_outputs(9787));
    layer1_outputs(7177) <= not((layer0_outputs(3280)) or (layer0_outputs(2175)));
    layer1_outputs(7178) <= not((layer0_outputs(896)) or (layer0_outputs(7621)));
    layer1_outputs(7179) <= not(layer0_outputs(5681));
    layer1_outputs(7180) <= not(layer0_outputs(111));
    layer1_outputs(7181) <= not(layer0_outputs(2396));
    layer1_outputs(7182) <= not(layer0_outputs(1077)) or (layer0_outputs(3683));
    layer1_outputs(7183) <= layer0_outputs(10022);
    layer1_outputs(7184) <= layer0_outputs(5808);
    layer1_outputs(7185) <= (layer0_outputs(8627)) and not (layer0_outputs(4082));
    layer1_outputs(7186) <= not(layer0_outputs(2506));
    layer1_outputs(7187) <= not(layer0_outputs(8133));
    layer1_outputs(7188) <= layer0_outputs(6859);
    layer1_outputs(7189) <= (layer0_outputs(6026)) and (layer0_outputs(1386));
    layer1_outputs(7190) <= not((layer0_outputs(86)) and (layer0_outputs(745)));
    layer1_outputs(7191) <= (layer0_outputs(1593)) or (layer0_outputs(6549));
    layer1_outputs(7192) <= (layer0_outputs(3160)) and (layer0_outputs(2886));
    layer1_outputs(7193) <= not(layer0_outputs(6504));
    layer1_outputs(7194) <= not((layer0_outputs(2620)) xor (layer0_outputs(7038)));
    layer1_outputs(7195) <= '1';
    layer1_outputs(7196) <= layer0_outputs(6026);
    layer1_outputs(7197) <= layer0_outputs(714);
    layer1_outputs(7198) <= layer0_outputs(5040);
    layer1_outputs(7199) <= layer0_outputs(12);
    layer1_outputs(7200) <= (layer0_outputs(1856)) and not (layer0_outputs(6195));
    layer1_outputs(7201) <= not((layer0_outputs(6664)) and (layer0_outputs(10017)));
    layer1_outputs(7202) <= layer0_outputs(6252);
    layer1_outputs(7203) <= not((layer0_outputs(7409)) and (layer0_outputs(2897)));
    layer1_outputs(7204) <= layer0_outputs(2645);
    layer1_outputs(7205) <= layer0_outputs(5493);
    layer1_outputs(7206) <= not(layer0_outputs(8608));
    layer1_outputs(7207) <= not(layer0_outputs(9874)) or (layer0_outputs(10054));
    layer1_outputs(7208) <= not(layer0_outputs(7473));
    layer1_outputs(7209) <= (layer0_outputs(4928)) xor (layer0_outputs(9379));
    layer1_outputs(7210) <= not(layer0_outputs(842));
    layer1_outputs(7211) <= (layer0_outputs(7065)) and not (layer0_outputs(5583));
    layer1_outputs(7212) <= (layer0_outputs(9984)) xor (layer0_outputs(7005));
    layer1_outputs(7213) <= not(layer0_outputs(9866)) or (layer0_outputs(1121));
    layer1_outputs(7214) <= not(layer0_outputs(10077));
    layer1_outputs(7215) <= (layer0_outputs(7810)) and not (layer0_outputs(532));
    layer1_outputs(7216) <= not((layer0_outputs(5857)) xor (layer0_outputs(7560)));
    layer1_outputs(7217) <= not((layer0_outputs(7657)) or (layer0_outputs(10123)));
    layer1_outputs(7218) <= (layer0_outputs(3491)) and not (layer0_outputs(2880));
    layer1_outputs(7219) <= not((layer0_outputs(8359)) xor (layer0_outputs(2367)));
    layer1_outputs(7220) <= not((layer0_outputs(7718)) xor (layer0_outputs(528)));
    layer1_outputs(7221) <= layer0_outputs(9068);
    layer1_outputs(7222) <= (layer0_outputs(5452)) and not (layer0_outputs(653));
    layer1_outputs(7223) <= '1';
    layer1_outputs(7224) <= layer0_outputs(5302);
    layer1_outputs(7225) <= layer0_outputs(1935);
    layer1_outputs(7226) <= not(layer0_outputs(1537)) or (layer0_outputs(576));
    layer1_outputs(7227) <= layer0_outputs(4130);
    layer1_outputs(7228) <= (layer0_outputs(8522)) and (layer0_outputs(9400));
    layer1_outputs(7229) <= not(layer0_outputs(7035)) or (layer0_outputs(4600));
    layer1_outputs(7230) <= (layer0_outputs(9476)) and (layer0_outputs(3443));
    layer1_outputs(7231) <= not(layer0_outputs(4197));
    layer1_outputs(7232) <= (layer0_outputs(7395)) and (layer0_outputs(6584));
    layer1_outputs(7233) <= not(layer0_outputs(8545)) or (layer0_outputs(7171));
    layer1_outputs(7234) <= layer0_outputs(1278);
    layer1_outputs(7235) <= not((layer0_outputs(4718)) xor (layer0_outputs(6036)));
    layer1_outputs(7236) <= not(layer0_outputs(8724));
    layer1_outputs(7237) <= (layer0_outputs(1783)) and (layer0_outputs(5396));
    layer1_outputs(7238) <= (layer0_outputs(6736)) and not (layer0_outputs(5793));
    layer1_outputs(7239) <= (layer0_outputs(8538)) or (layer0_outputs(7355));
    layer1_outputs(7240) <= layer0_outputs(295);
    layer1_outputs(7241) <= layer0_outputs(3620);
    layer1_outputs(7242) <= (layer0_outputs(6432)) and not (layer0_outputs(7428));
    layer1_outputs(7243) <= not((layer0_outputs(3251)) and (layer0_outputs(8775)));
    layer1_outputs(7244) <= not((layer0_outputs(1639)) or (layer0_outputs(8928)));
    layer1_outputs(7245) <= (layer0_outputs(6235)) and not (layer0_outputs(4381));
    layer1_outputs(7246) <= not((layer0_outputs(2546)) or (layer0_outputs(5117)));
    layer1_outputs(7247) <= not(layer0_outputs(7624));
    layer1_outputs(7248) <= not(layer0_outputs(972));
    layer1_outputs(7249) <= not((layer0_outputs(6720)) xor (layer0_outputs(5272)));
    layer1_outputs(7250) <= layer0_outputs(6152);
    layer1_outputs(7251) <= not(layer0_outputs(2709));
    layer1_outputs(7252) <= (layer0_outputs(7539)) xor (layer0_outputs(3265));
    layer1_outputs(7253) <= not((layer0_outputs(1295)) xor (layer0_outputs(2509)));
    layer1_outputs(7254) <= not(layer0_outputs(930)) or (layer0_outputs(6571));
    layer1_outputs(7255) <= not(layer0_outputs(1406));
    layer1_outputs(7256) <= (layer0_outputs(5666)) and (layer0_outputs(9096));
    layer1_outputs(7257) <= not((layer0_outputs(6139)) or (layer0_outputs(4157)));
    layer1_outputs(7258) <= layer0_outputs(6772);
    layer1_outputs(7259) <= not(layer0_outputs(2970));
    layer1_outputs(7260) <= not(layer0_outputs(2095)) or (layer0_outputs(8687));
    layer1_outputs(7261) <= not(layer0_outputs(1650));
    layer1_outputs(7262) <= layer0_outputs(4290);
    layer1_outputs(7263) <= (layer0_outputs(3491)) and (layer0_outputs(6926));
    layer1_outputs(7264) <= not(layer0_outputs(1751));
    layer1_outputs(7265) <= not((layer0_outputs(9718)) and (layer0_outputs(7230)));
    layer1_outputs(7266) <= not(layer0_outputs(8767));
    layer1_outputs(7267) <= (layer0_outputs(7172)) and not (layer0_outputs(3953));
    layer1_outputs(7268) <= (layer0_outputs(7001)) or (layer0_outputs(2829));
    layer1_outputs(7269) <= (layer0_outputs(1333)) and not (layer0_outputs(8126));
    layer1_outputs(7270) <= '0';
    layer1_outputs(7271) <= layer0_outputs(765);
    layer1_outputs(7272) <= (layer0_outputs(7002)) or (layer0_outputs(9162));
    layer1_outputs(7273) <= layer0_outputs(5537);
    layer1_outputs(7274) <= '0';
    layer1_outputs(7275) <= (layer0_outputs(9721)) or (layer0_outputs(3310));
    layer1_outputs(7276) <= not(layer0_outputs(80));
    layer1_outputs(7277) <= not((layer0_outputs(9388)) and (layer0_outputs(4784)));
    layer1_outputs(7278) <= '0';
    layer1_outputs(7279) <= (layer0_outputs(1159)) and (layer0_outputs(3247));
    layer1_outputs(7280) <= not(layer0_outputs(9525)) or (layer0_outputs(8480));
    layer1_outputs(7281) <= (layer0_outputs(8075)) and not (layer0_outputs(7519));
    layer1_outputs(7282) <= layer0_outputs(2060);
    layer1_outputs(7283) <= '0';
    layer1_outputs(7284) <= not(layer0_outputs(4)) or (layer0_outputs(6500));
    layer1_outputs(7285) <= not((layer0_outputs(2964)) and (layer0_outputs(5945)));
    layer1_outputs(7286) <= not(layer0_outputs(6175)) or (layer0_outputs(3795));
    layer1_outputs(7287) <= not(layer0_outputs(4695)) or (layer0_outputs(3832));
    layer1_outputs(7288) <= not((layer0_outputs(2120)) and (layer0_outputs(8112)));
    layer1_outputs(7289) <= (layer0_outputs(8619)) xor (layer0_outputs(5725));
    layer1_outputs(7290) <= not((layer0_outputs(4006)) or (layer0_outputs(5244)));
    layer1_outputs(7291) <= not(layer0_outputs(620)) or (layer0_outputs(4913));
    layer1_outputs(7292) <= not(layer0_outputs(4684));
    layer1_outputs(7293) <= not(layer0_outputs(9921));
    layer1_outputs(7294) <= '0';
    layer1_outputs(7295) <= layer0_outputs(8614);
    layer1_outputs(7296) <= not((layer0_outputs(8937)) xor (layer0_outputs(4389)));
    layer1_outputs(7297) <= not((layer0_outputs(7625)) xor (layer0_outputs(270)));
    layer1_outputs(7298) <= not(layer0_outputs(2468));
    layer1_outputs(7299) <= (layer0_outputs(5214)) and (layer0_outputs(7127));
    layer1_outputs(7300) <= not((layer0_outputs(3756)) or (layer0_outputs(7102)));
    layer1_outputs(7301) <= not(layer0_outputs(240));
    layer1_outputs(7302) <= (layer0_outputs(8245)) and (layer0_outputs(3551));
    layer1_outputs(7303) <= layer0_outputs(8965);
    layer1_outputs(7304) <= (layer0_outputs(7937)) and (layer0_outputs(2158));
    layer1_outputs(7305) <= not(layer0_outputs(7782)) or (layer0_outputs(5812));
    layer1_outputs(7306) <= not(layer0_outputs(469));
    layer1_outputs(7307) <= (layer0_outputs(7473)) or (layer0_outputs(5427));
    layer1_outputs(7308) <= layer0_outputs(492);
    layer1_outputs(7309) <= not(layer0_outputs(920)) or (layer0_outputs(2045));
    layer1_outputs(7310) <= (layer0_outputs(981)) and not (layer0_outputs(2813));
    layer1_outputs(7311) <= not(layer0_outputs(9536)) or (layer0_outputs(2178));
    layer1_outputs(7312) <= not((layer0_outputs(4420)) and (layer0_outputs(2749)));
    layer1_outputs(7313) <= not((layer0_outputs(8230)) and (layer0_outputs(9722)));
    layer1_outputs(7314) <= not(layer0_outputs(10091));
    layer1_outputs(7315) <= (layer0_outputs(7973)) and not (layer0_outputs(2416));
    layer1_outputs(7316) <= (layer0_outputs(4752)) and (layer0_outputs(10044));
    layer1_outputs(7317) <= not((layer0_outputs(3531)) and (layer0_outputs(7048)));
    layer1_outputs(7318) <= not(layer0_outputs(5665));
    layer1_outputs(7319) <= not(layer0_outputs(188)) or (layer0_outputs(1945));
    layer1_outputs(7320) <= not((layer0_outputs(631)) or (layer0_outputs(1267)));
    layer1_outputs(7321) <= (layer0_outputs(1793)) and not (layer0_outputs(9938));
    layer1_outputs(7322) <= '1';
    layer1_outputs(7323) <= not(layer0_outputs(9836));
    layer1_outputs(7324) <= not((layer0_outputs(3393)) xor (layer0_outputs(306)));
    layer1_outputs(7325) <= (layer0_outputs(9706)) and (layer0_outputs(2303));
    layer1_outputs(7326) <= not(layer0_outputs(1224)) or (layer0_outputs(2527));
    layer1_outputs(7327) <= layer0_outputs(9819);
    layer1_outputs(7328) <= not(layer0_outputs(4392));
    layer1_outputs(7329) <= not(layer0_outputs(5317)) or (layer0_outputs(2423));
    layer1_outputs(7330) <= (layer0_outputs(9065)) and not (layer0_outputs(3890));
    layer1_outputs(7331) <= not((layer0_outputs(9238)) or (layer0_outputs(9413)));
    layer1_outputs(7332) <= not((layer0_outputs(2437)) xor (layer0_outputs(1922)));
    layer1_outputs(7333) <= not(layer0_outputs(5155));
    layer1_outputs(7334) <= (layer0_outputs(6457)) and not (layer0_outputs(7075));
    layer1_outputs(7335) <= not((layer0_outputs(3086)) or (layer0_outputs(409)));
    layer1_outputs(7336) <= not(layer0_outputs(4780)) or (layer0_outputs(1658));
    layer1_outputs(7337) <= not(layer0_outputs(3423)) or (layer0_outputs(7210));
    layer1_outputs(7338) <= (layer0_outputs(9451)) and not (layer0_outputs(1977));
    layer1_outputs(7339) <= not(layer0_outputs(2641)) or (layer0_outputs(7303));
    layer1_outputs(7340) <= layer0_outputs(3015);
    layer1_outputs(7341) <= not(layer0_outputs(1837));
    layer1_outputs(7342) <= not(layer0_outputs(852));
    layer1_outputs(7343) <= not((layer0_outputs(10048)) or (layer0_outputs(1963)));
    layer1_outputs(7344) <= not(layer0_outputs(8968));
    layer1_outputs(7345) <= (layer0_outputs(8149)) and not (layer0_outputs(5777));
    layer1_outputs(7346) <= not(layer0_outputs(8216));
    layer1_outputs(7347) <= not((layer0_outputs(8891)) or (layer0_outputs(5669)));
    layer1_outputs(7348) <= not(layer0_outputs(7875)) or (layer0_outputs(1344));
    layer1_outputs(7349) <= layer0_outputs(4376);
    layer1_outputs(7350) <= not(layer0_outputs(2567));
    layer1_outputs(7351) <= not(layer0_outputs(1349));
    layer1_outputs(7352) <= (layer0_outputs(354)) and not (layer0_outputs(3475));
    layer1_outputs(7353) <= (layer0_outputs(7461)) and not (layer0_outputs(5363));
    layer1_outputs(7354) <= not(layer0_outputs(6855)) or (layer0_outputs(5981));
    layer1_outputs(7355) <= not(layer0_outputs(3983));
    layer1_outputs(7356) <= (layer0_outputs(6575)) and (layer0_outputs(10157));
    layer1_outputs(7357) <= not(layer0_outputs(2691));
    layer1_outputs(7358) <= layer0_outputs(3456);
    layer1_outputs(7359) <= (layer0_outputs(3758)) and (layer0_outputs(2927));
    layer1_outputs(7360) <= not(layer0_outputs(3644));
    layer1_outputs(7361) <= (layer0_outputs(687)) and not (layer0_outputs(10120));
    layer1_outputs(7362) <= (layer0_outputs(467)) and not (layer0_outputs(249));
    layer1_outputs(7363) <= not((layer0_outputs(1254)) and (layer0_outputs(8748)));
    layer1_outputs(7364) <= not((layer0_outputs(9543)) and (layer0_outputs(9605)));
    layer1_outputs(7365) <= not(layer0_outputs(2760)) or (layer0_outputs(964));
    layer1_outputs(7366) <= (layer0_outputs(1197)) and not (layer0_outputs(1515));
    layer1_outputs(7367) <= not((layer0_outputs(1297)) or (layer0_outputs(816)));
    layer1_outputs(7368) <= not(layer0_outputs(7853)) or (layer0_outputs(10000));
    layer1_outputs(7369) <= (layer0_outputs(424)) and not (layer0_outputs(9785));
    layer1_outputs(7370) <= (layer0_outputs(6006)) and (layer0_outputs(9005));
    layer1_outputs(7371) <= (layer0_outputs(1652)) and not (layer0_outputs(2189));
    layer1_outputs(7372) <= (layer0_outputs(9857)) and not (layer0_outputs(6120));
    layer1_outputs(7373) <= not((layer0_outputs(8323)) xor (layer0_outputs(880)));
    layer1_outputs(7374) <= not(layer0_outputs(8035)) or (layer0_outputs(2333));
    layer1_outputs(7375) <= layer0_outputs(7457);
    layer1_outputs(7376) <= layer0_outputs(6953);
    layer1_outputs(7377) <= not(layer0_outputs(3946)) or (layer0_outputs(4477));
    layer1_outputs(7378) <= layer0_outputs(9754);
    layer1_outputs(7379) <= '1';
    layer1_outputs(7380) <= not(layer0_outputs(6874));
    layer1_outputs(7381) <= not(layer0_outputs(8707));
    layer1_outputs(7382) <= (layer0_outputs(4900)) or (layer0_outputs(573));
    layer1_outputs(7383) <= (layer0_outputs(7128)) and not (layer0_outputs(7728));
    layer1_outputs(7384) <= (layer0_outputs(8777)) and not (layer0_outputs(3751));
    layer1_outputs(7385) <= (layer0_outputs(67)) and not (layer0_outputs(8516));
    layer1_outputs(7386) <= (layer0_outputs(3660)) and (layer0_outputs(2736));
    layer1_outputs(7387) <= not(layer0_outputs(9432));
    layer1_outputs(7388) <= '1';
    layer1_outputs(7389) <= not((layer0_outputs(1908)) and (layer0_outputs(5728)));
    layer1_outputs(7390) <= not(layer0_outputs(7605));
    layer1_outputs(7391) <= (layer0_outputs(7569)) and not (layer0_outputs(2843));
    layer1_outputs(7392) <= (layer0_outputs(5938)) and not (layer0_outputs(8009));
    layer1_outputs(7393) <= (layer0_outputs(3312)) and not (layer0_outputs(984));
    layer1_outputs(7394) <= layer0_outputs(9253);
    layer1_outputs(7395) <= '0';
    layer1_outputs(7396) <= (layer0_outputs(5049)) and not (layer0_outputs(5093));
    layer1_outputs(7397) <= not((layer0_outputs(3284)) and (layer0_outputs(5823)));
    layer1_outputs(7398) <= layer0_outputs(4910);
    layer1_outputs(7399) <= (layer0_outputs(7479)) and not (layer0_outputs(3908));
    layer1_outputs(7400) <= not(layer0_outputs(305)) or (layer0_outputs(7754));
    layer1_outputs(7401) <= layer0_outputs(4681);
    layer1_outputs(7402) <= not(layer0_outputs(6551)) or (layer0_outputs(9596));
    layer1_outputs(7403) <= layer0_outputs(1135);
    layer1_outputs(7404) <= not(layer0_outputs(7367));
    layer1_outputs(7405) <= (layer0_outputs(5114)) and (layer0_outputs(7405));
    layer1_outputs(7406) <= layer0_outputs(8890);
    layer1_outputs(7407) <= (layer0_outputs(4580)) and not (layer0_outputs(5840));
    layer1_outputs(7408) <= layer0_outputs(33);
    layer1_outputs(7409) <= not(layer0_outputs(8355)) or (layer0_outputs(1287));
    layer1_outputs(7410) <= layer0_outputs(4975);
    layer1_outputs(7411) <= (layer0_outputs(1795)) and (layer0_outputs(5715));
    layer1_outputs(7412) <= (layer0_outputs(2992)) or (layer0_outputs(948));
    layer1_outputs(7413) <= not(layer0_outputs(9221));
    layer1_outputs(7414) <= '1';
    layer1_outputs(7415) <= (layer0_outputs(906)) xor (layer0_outputs(2854));
    layer1_outputs(7416) <= not(layer0_outputs(4537)) or (layer0_outputs(4117));
    layer1_outputs(7417) <= (layer0_outputs(6383)) and not (layer0_outputs(6111));
    layer1_outputs(7418) <= '0';
    layer1_outputs(7419) <= not(layer0_outputs(218));
    layer1_outputs(7420) <= not(layer0_outputs(1102)) or (layer0_outputs(6005));
    layer1_outputs(7421) <= not(layer0_outputs(5959));
    layer1_outputs(7422) <= layer0_outputs(2553);
    layer1_outputs(7423) <= not(layer0_outputs(9416));
    layer1_outputs(7424) <= layer0_outputs(1012);
    layer1_outputs(7425) <= not(layer0_outputs(3720)) or (layer0_outputs(4009));
    layer1_outputs(7426) <= not(layer0_outputs(3692)) or (layer0_outputs(9224));
    layer1_outputs(7427) <= not(layer0_outputs(6639)) or (layer0_outputs(4954));
    layer1_outputs(7428) <= not((layer0_outputs(5191)) and (layer0_outputs(6570)));
    layer1_outputs(7429) <= not(layer0_outputs(2884));
    layer1_outputs(7430) <= not((layer0_outputs(6312)) or (layer0_outputs(3039)));
    layer1_outputs(7431) <= not((layer0_outputs(2446)) or (layer0_outputs(3790)));
    layer1_outputs(7432) <= not(layer0_outputs(430));
    layer1_outputs(7433) <= layer0_outputs(801);
    layer1_outputs(7434) <= not(layer0_outputs(9807));
    layer1_outputs(7435) <= not(layer0_outputs(55));
    layer1_outputs(7436) <= not((layer0_outputs(5974)) and (layer0_outputs(4061)));
    layer1_outputs(7437) <= not((layer0_outputs(1428)) and (layer0_outputs(1322)));
    layer1_outputs(7438) <= layer0_outputs(8399);
    layer1_outputs(7439) <= layer0_outputs(2720);
    layer1_outputs(7440) <= not(layer0_outputs(8749)) or (layer0_outputs(6447));
    layer1_outputs(7441) <= (layer0_outputs(6932)) and (layer0_outputs(5677));
    layer1_outputs(7442) <= not(layer0_outputs(4062));
    layer1_outputs(7443) <= not(layer0_outputs(1791));
    layer1_outputs(7444) <= not(layer0_outputs(4898));
    layer1_outputs(7445) <= (layer0_outputs(4695)) and (layer0_outputs(2054));
    layer1_outputs(7446) <= not(layer0_outputs(7741)) or (layer0_outputs(7448));
    layer1_outputs(7447) <= layer0_outputs(1992);
    layer1_outputs(7448) <= not(layer0_outputs(502));
    layer1_outputs(7449) <= layer0_outputs(1200);
    layer1_outputs(7450) <= not(layer0_outputs(7512)) or (layer0_outputs(5793));
    layer1_outputs(7451) <= (layer0_outputs(9243)) and (layer0_outputs(3685));
    layer1_outputs(7452) <= not((layer0_outputs(9853)) or (layer0_outputs(7689)));
    layer1_outputs(7453) <= layer0_outputs(4280);
    layer1_outputs(7454) <= not(layer0_outputs(4005)) or (layer0_outputs(5812));
    layer1_outputs(7455) <= '1';
    layer1_outputs(7456) <= not(layer0_outputs(1365));
    layer1_outputs(7457) <= not(layer0_outputs(5110)) or (layer0_outputs(9493));
    layer1_outputs(7458) <= layer0_outputs(7798);
    layer1_outputs(7459) <= not((layer0_outputs(2744)) xor (layer0_outputs(414)));
    layer1_outputs(7460) <= '1';
    layer1_outputs(7461) <= not(layer0_outputs(5911));
    layer1_outputs(7462) <= not(layer0_outputs(8143));
    layer1_outputs(7463) <= not(layer0_outputs(7982)) or (layer0_outputs(8785));
    layer1_outputs(7464) <= (layer0_outputs(1448)) and (layer0_outputs(1408));
    layer1_outputs(7465) <= layer0_outputs(346);
    layer1_outputs(7466) <= (layer0_outputs(1215)) and not (layer0_outputs(9302));
    layer1_outputs(7467) <= not(layer0_outputs(5005)) or (layer0_outputs(3984));
    layer1_outputs(7468) <= not(layer0_outputs(716));
    layer1_outputs(7469) <= (layer0_outputs(5097)) and (layer0_outputs(1070));
    layer1_outputs(7470) <= not(layer0_outputs(5318));
    layer1_outputs(7471) <= layer0_outputs(8378);
    layer1_outputs(7472) <= layer0_outputs(9029);
    layer1_outputs(7473) <= (layer0_outputs(323)) and not (layer0_outputs(8852));
    layer1_outputs(7474) <= layer0_outputs(2344);
    layer1_outputs(7475) <= not(layer0_outputs(3680)) or (layer0_outputs(1421));
    layer1_outputs(7476) <= not(layer0_outputs(991));
    layer1_outputs(7477) <= layer0_outputs(2659);
    layer1_outputs(7478) <= (layer0_outputs(9468)) and not (layer0_outputs(1095));
    layer1_outputs(7479) <= layer0_outputs(2914);
    layer1_outputs(7480) <= not(layer0_outputs(7996));
    layer1_outputs(7481) <= layer0_outputs(3070);
    layer1_outputs(7482) <= (layer0_outputs(8269)) and (layer0_outputs(5093));
    layer1_outputs(7483) <= not(layer0_outputs(7882)) or (layer0_outputs(1457));
    layer1_outputs(7484) <= (layer0_outputs(447)) or (layer0_outputs(8142));
    layer1_outputs(7485) <= not(layer0_outputs(8338));
    layer1_outputs(7486) <= layer0_outputs(8499);
    layer1_outputs(7487) <= not(layer0_outputs(6743));
    layer1_outputs(7488) <= not((layer0_outputs(5773)) xor (layer0_outputs(2648)));
    layer1_outputs(7489) <= not(layer0_outputs(9116));
    layer1_outputs(7490) <= not(layer0_outputs(69));
    layer1_outputs(7491) <= (layer0_outputs(6987)) and not (layer0_outputs(3557));
    layer1_outputs(7492) <= (layer0_outputs(9471)) or (layer0_outputs(1771));
    layer1_outputs(7493) <= (layer0_outputs(4943)) and (layer0_outputs(9191));
    layer1_outputs(7494) <= not((layer0_outputs(10168)) and (layer0_outputs(9685)));
    layer1_outputs(7495) <= not((layer0_outputs(3016)) or (layer0_outputs(881)));
    layer1_outputs(7496) <= not(layer0_outputs(289));
    layer1_outputs(7497) <= layer0_outputs(3710);
    layer1_outputs(7498) <= (layer0_outputs(9177)) and not (layer0_outputs(6392));
    layer1_outputs(7499) <= (layer0_outputs(2636)) xor (layer0_outputs(237));
    layer1_outputs(7500) <= (layer0_outputs(5866)) and not (layer0_outputs(6113));
    layer1_outputs(7501) <= layer0_outputs(9399);
    layer1_outputs(7502) <= (layer0_outputs(4505)) and (layer0_outputs(597));
    layer1_outputs(7503) <= not(layer0_outputs(6788));
    layer1_outputs(7504) <= layer0_outputs(3205);
    layer1_outputs(7505) <= not(layer0_outputs(9441));
    layer1_outputs(7506) <= layer0_outputs(6248);
    layer1_outputs(7507) <= (layer0_outputs(8439)) xor (layer0_outputs(6776));
    layer1_outputs(7508) <= not(layer0_outputs(10216)) or (layer0_outputs(1178));
    layer1_outputs(7509) <= not((layer0_outputs(5501)) xor (layer0_outputs(6489)));
    layer1_outputs(7510) <= not(layer0_outputs(4276)) or (layer0_outputs(889));
    layer1_outputs(7511) <= not(layer0_outputs(7927)) or (layer0_outputs(7149));
    layer1_outputs(7512) <= layer0_outputs(6011);
    layer1_outputs(7513) <= not(layer0_outputs(2743)) or (layer0_outputs(7846));
    layer1_outputs(7514) <= not((layer0_outputs(8947)) or (layer0_outputs(8685)));
    layer1_outputs(7515) <= (layer0_outputs(877)) or (layer0_outputs(7649));
    layer1_outputs(7516) <= not(layer0_outputs(224));
    layer1_outputs(7517) <= not(layer0_outputs(7947)) or (layer0_outputs(3287));
    layer1_outputs(7518) <= '0';
    layer1_outputs(7519) <= not(layer0_outputs(9948));
    layer1_outputs(7520) <= not((layer0_outputs(8974)) xor (layer0_outputs(7736)));
    layer1_outputs(7521) <= (layer0_outputs(4352)) or (layer0_outputs(7576));
    layer1_outputs(7522) <= not((layer0_outputs(5749)) xor (layer0_outputs(3215)));
    layer1_outputs(7523) <= not(layer0_outputs(5605));
    layer1_outputs(7524) <= not(layer0_outputs(360));
    layer1_outputs(7525) <= (layer0_outputs(4647)) and (layer0_outputs(7427));
    layer1_outputs(7526) <= (layer0_outputs(3575)) and not (layer0_outputs(9797));
    layer1_outputs(7527) <= (layer0_outputs(1574)) and not (layer0_outputs(2637));
    layer1_outputs(7528) <= layer0_outputs(3594);
    layer1_outputs(7529) <= not(layer0_outputs(6277)) or (layer0_outputs(3288));
    layer1_outputs(7530) <= not(layer0_outputs(5017)) or (layer0_outputs(6048));
    layer1_outputs(7531) <= not((layer0_outputs(9285)) and (layer0_outputs(4662)));
    layer1_outputs(7532) <= not(layer0_outputs(1671)) or (layer0_outputs(9045));
    layer1_outputs(7533) <= not(layer0_outputs(4628));
    layer1_outputs(7534) <= layer0_outputs(7534);
    layer1_outputs(7535) <= not(layer0_outputs(10001)) or (layer0_outputs(2840));
    layer1_outputs(7536) <= not((layer0_outputs(250)) or (layer0_outputs(2929)));
    layer1_outputs(7537) <= (layer0_outputs(210)) and not (layer0_outputs(7524));
    layer1_outputs(7538) <= layer0_outputs(5522);
    layer1_outputs(7539) <= (layer0_outputs(1334)) or (layer0_outputs(4129));
    layer1_outputs(7540) <= not(layer0_outputs(7625));
    layer1_outputs(7541) <= not((layer0_outputs(2614)) xor (layer0_outputs(8261)));
    layer1_outputs(7542) <= (layer0_outputs(3184)) xor (layer0_outputs(730));
    layer1_outputs(7543) <= layer0_outputs(4089);
    layer1_outputs(7544) <= (layer0_outputs(3104)) and (layer0_outputs(8036));
    layer1_outputs(7545) <= layer0_outputs(259);
    layer1_outputs(7546) <= not((layer0_outputs(1718)) or (layer0_outputs(6790)));
    layer1_outputs(7547) <= not(layer0_outputs(1662));
    layer1_outputs(7548) <= (layer0_outputs(8807)) and (layer0_outputs(7606));
    layer1_outputs(7549) <= not(layer0_outputs(5054));
    layer1_outputs(7550) <= not(layer0_outputs(6157));
    layer1_outputs(7551) <= not((layer0_outputs(3101)) or (layer0_outputs(5596)));
    layer1_outputs(7552) <= '1';
    layer1_outputs(7553) <= (layer0_outputs(9585)) xor (layer0_outputs(2457));
    layer1_outputs(7554) <= (layer0_outputs(1735)) and (layer0_outputs(1154));
    layer1_outputs(7555) <= (layer0_outputs(232)) xor (layer0_outputs(1414));
    layer1_outputs(7556) <= not((layer0_outputs(4801)) and (layer0_outputs(2172)));
    layer1_outputs(7557) <= not((layer0_outputs(8044)) or (layer0_outputs(6079)));
    layer1_outputs(7558) <= (layer0_outputs(5148)) and not (layer0_outputs(911));
    layer1_outputs(7559) <= layer0_outputs(3063);
    layer1_outputs(7560) <= layer0_outputs(3745);
    layer1_outputs(7561) <= layer0_outputs(5133);
    layer1_outputs(7562) <= (layer0_outputs(7824)) xor (layer0_outputs(4439));
    layer1_outputs(7563) <= layer0_outputs(2353);
    layer1_outputs(7564) <= (layer0_outputs(9700)) and (layer0_outputs(3741));
    layer1_outputs(7565) <= (layer0_outputs(9569)) and not (layer0_outputs(1453));
    layer1_outputs(7566) <= (layer0_outputs(8605)) or (layer0_outputs(5087));
    layer1_outputs(7567) <= not((layer0_outputs(6342)) xor (layer0_outputs(4124)));
    layer1_outputs(7568) <= not((layer0_outputs(5655)) or (layer0_outputs(8466)));
    layer1_outputs(7569) <= (layer0_outputs(8969)) and not (layer0_outputs(3262));
    layer1_outputs(7570) <= not((layer0_outputs(2116)) or (layer0_outputs(2697)));
    layer1_outputs(7571) <= layer0_outputs(5489);
    layer1_outputs(7572) <= not(layer0_outputs(2848)) or (layer0_outputs(9749));
    layer1_outputs(7573) <= layer0_outputs(2125);
    layer1_outputs(7574) <= layer0_outputs(1266);
    layer1_outputs(7575) <= not((layer0_outputs(9779)) or (layer0_outputs(307)));
    layer1_outputs(7576) <= not(layer0_outputs(6372)) or (layer0_outputs(2907));
    layer1_outputs(7577) <= (layer0_outputs(9248)) and not (layer0_outputs(454));
    layer1_outputs(7578) <= not((layer0_outputs(2717)) and (layer0_outputs(9594)));
    layer1_outputs(7579) <= layer0_outputs(9815);
    layer1_outputs(7580) <= not(layer0_outputs(2222));
    layer1_outputs(7581) <= not(layer0_outputs(4465)) or (layer0_outputs(7492));
    layer1_outputs(7582) <= (layer0_outputs(10201)) or (layer0_outputs(9656));
    layer1_outputs(7583) <= not(layer0_outputs(7377));
    layer1_outputs(7584) <= (layer0_outputs(7078)) or (layer0_outputs(693));
    layer1_outputs(7585) <= (layer0_outputs(829)) and not (layer0_outputs(2277));
    layer1_outputs(7586) <= not((layer0_outputs(8018)) and (layer0_outputs(2414)));
    layer1_outputs(7587) <= not(layer0_outputs(6406));
    layer1_outputs(7588) <= not(layer0_outputs(3311));
    layer1_outputs(7589) <= not((layer0_outputs(4384)) and (layer0_outputs(7746)));
    layer1_outputs(7590) <= (layer0_outputs(2769)) and not (layer0_outputs(10197));
    layer1_outputs(7591) <= not(layer0_outputs(2574)) or (layer0_outputs(1752));
    layer1_outputs(7592) <= layer0_outputs(928);
    layer1_outputs(7593) <= (layer0_outputs(7055)) and (layer0_outputs(4098));
    layer1_outputs(7594) <= not((layer0_outputs(3640)) and (layer0_outputs(5404)));
    layer1_outputs(7595) <= not((layer0_outputs(8332)) xor (layer0_outputs(8620)));
    layer1_outputs(7596) <= not(layer0_outputs(2277)) or (layer0_outputs(2871));
    layer1_outputs(7597) <= not((layer0_outputs(6662)) and (layer0_outputs(3655)));
    layer1_outputs(7598) <= not((layer0_outputs(2755)) or (layer0_outputs(8185)));
    layer1_outputs(7599) <= '0';
    layer1_outputs(7600) <= layer0_outputs(2217);
    layer1_outputs(7601) <= layer0_outputs(8196);
    layer1_outputs(7602) <= (layer0_outputs(2641)) and not (layer0_outputs(7096));
    layer1_outputs(7603) <= layer0_outputs(9958);
    layer1_outputs(7604) <= '0';
    layer1_outputs(7605) <= (layer0_outputs(2242)) or (layer0_outputs(10056));
    layer1_outputs(7606) <= not(layer0_outputs(105));
    layer1_outputs(7607) <= layer0_outputs(3859);
    layer1_outputs(7608) <= layer0_outputs(7294);
    layer1_outputs(7609) <= (layer0_outputs(3378)) or (layer0_outputs(8040));
    layer1_outputs(7610) <= '1';
    layer1_outputs(7611) <= not(layer0_outputs(7662));
    layer1_outputs(7612) <= (layer0_outputs(403)) or (layer0_outputs(6679));
    layer1_outputs(7613) <= not(layer0_outputs(2787));
    layer1_outputs(7614) <= not(layer0_outputs(2144)) or (layer0_outputs(8461));
    layer1_outputs(7615) <= not((layer0_outputs(6167)) xor (layer0_outputs(7707)));
    layer1_outputs(7616) <= not(layer0_outputs(3442));
    layer1_outputs(7617) <= '0';
    layer1_outputs(7618) <= layer0_outputs(420);
    layer1_outputs(7619) <= not(layer0_outputs(9465)) or (layer0_outputs(3464));
    layer1_outputs(7620) <= (layer0_outputs(6598)) xor (layer0_outputs(1654));
    layer1_outputs(7621) <= not(layer0_outputs(6909));
    layer1_outputs(7622) <= (layer0_outputs(618)) or (layer0_outputs(5329));
    layer1_outputs(7623) <= '0';
    layer1_outputs(7624) <= not(layer0_outputs(4069));
    layer1_outputs(7625) <= (layer0_outputs(3721)) xor (layer0_outputs(7014));
    layer1_outputs(7626) <= not((layer0_outputs(1638)) or (layer0_outputs(5372)));
    layer1_outputs(7627) <= not(layer0_outputs(8445)) or (layer0_outputs(9320));
    layer1_outputs(7628) <= (layer0_outputs(82)) and not (layer0_outputs(3543));
    layer1_outputs(7629) <= '1';
    layer1_outputs(7630) <= layer0_outputs(8529);
    layer1_outputs(7631) <= (layer0_outputs(8892)) or (layer0_outputs(1211));
    layer1_outputs(7632) <= (layer0_outputs(4522)) xor (layer0_outputs(2498));
    layer1_outputs(7633) <= (layer0_outputs(71)) and not (layer0_outputs(10063));
    layer1_outputs(7634) <= not(layer0_outputs(4047));
    layer1_outputs(7635) <= not((layer0_outputs(342)) and (layer0_outputs(7749)));
    layer1_outputs(7636) <= layer0_outputs(888);
    layer1_outputs(7637) <= not(layer0_outputs(7052));
    layer1_outputs(7638) <= not((layer0_outputs(4910)) xor (layer0_outputs(1390)));
    layer1_outputs(7639) <= not((layer0_outputs(4853)) and (layer0_outputs(704)));
    layer1_outputs(7640) <= layer0_outputs(1072);
    layer1_outputs(7641) <= layer0_outputs(4988);
    layer1_outputs(7642) <= (layer0_outputs(9325)) and not (layer0_outputs(2553));
    layer1_outputs(7643) <= (layer0_outputs(7233)) and (layer0_outputs(5742));
    layer1_outputs(7644) <= not(layer0_outputs(3786)) or (layer0_outputs(3539));
    layer1_outputs(7645) <= (layer0_outputs(8269)) and (layer0_outputs(4887));
    layer1_outputs(7646) <= not(layer0_outputs(10060));
    layer1_outputs(7647) <= layer0_outputs(1840);
    layer1_outputs(7648) <= not(layer0_outputs(1196));
    layer1_outputs(7649) <= '1';
    layer1_outputs(7650) <= not((layer0_outputs(9975)) and (layer0_outputs(7069)));
    layer1_outputs(7651) <= (layer0_outputs(4476)) or (layer0_outputs(3502));
    layer1_outputs(7652) <= not(layer0_outputs(3352)) or (layer0_outputs(3812));
    layer1_outputs(7653) <= not(layer0_outputs(6406)) or (layer0_outputs(6725));
    layer1_outputs(7654) <= not(layer0_outputs(7628));
    layer1_outputs(7655) <= (layer0_outputs(5554)) and not (layer0_outputs(5803));
    layer1_outputs(7656) <= layer0_outputs(1316);
    layer1_outputs(7657) <= (layer0_outputs(2915)) and not (layer0_outputs(755));
    layer1_outputs(7658) <= layer0_outputs(7795);
    layer1_outputs(7659) <= not(layer0_outputs(8369)) or (layer0_outputs(3659));
    layer1_outputs(7660) <= not(layer0_outputs(1802));
    layer1_outputs(7661) <= layer0_outputs(8518);
    layer1_outputs(7662) <= not(layer0_outputs(6794)) or (layer0_outputs(4625));
    layer1_outputs(7663) <= layer0_outputs(9505);
    layer1_outputs(7664) <= (layer0_outputs(396)) and not (layer0_outputs(8699));
    layer1_outputs(7665) <= not(layer0_outputs(5887));
    layer1_outputs(7666) <= not((layer0_outputs(2470)) and (layer0_outputs(8842)));
    layer1_outputs(7667) <= not(layer0_outputs(6501)) or (layer0_outputs(8811));
    layer1_outputs(7668) <= (layer0_outputs(7011)) or (layer0_outputs(7077));
    layer1_outputs(7669) <= not(layer0_outputs(569));
    layer1_outputs(7670) <= not((layer0_outputs(2495)) or (layer0_outputs(4110)));
    layer1_outputs(7671) <= layer0_outputs(1535);
    layer1_outputs(7672) <= (layer0_outputs(4648)) and (layer0_outputs(2249));
    layer1_outputs(7673) <= (layer0_outputs(7900)) and not (layer0_outputs(7825));
    layer1_outputs(7674) <= not(layer0_outputs(5253));
    layer1_outputs(7675) <= (layer0_outputs(7513)) or (layer0_outputs(6629));
    layer1_outputs(7676) <= not(layer0_outputs(5170)) or (layer0_outputs(9101));
    layer1_outputs(7677) <= layer0_outputs(4206);
    layer1_outputs(7678) <= layer0_outputs(7454);
    layer1_outputs(7679) <= layer0_outputs(3403);
    layer1_outputs(7680) <= not((layer0_outputs(8883)) xor (layer0_outputs(5935)));
    layer1_outputs(7681) <= layer0_outputs(1290);
    layer1_outputs(7682) <= not(layer0_outputs(2314));
    layer1_outputs(7683) <= not(layer0_outputs(3143));
    layer1_outputs(7684) <= (layer0_outputs(7072)) or (layer0_outputs(194));
    layer1_outputs(7685) <= (layer0_outputs(8036)) and not (layer0_outputs(6046));
    layer1_outputs(7686) <= not(layer0_outputs(1104));
    layer1_outputs(7687) <= not((layer0_outputs(7223)) and (layer0_outputs(6918)));
    layer1_outputs(7688) <= not(layer0_outputs(5319));
    layer1_outputs(7689) <= layer0_outputs(8881);
    layer1_outputs(7690) <= (layer0_outputs(8602)) or (layer0_outputs(7645));
    layer1_outputs(7691) <= not((layer0_outputs(1995)) and (layer0_outputs(6898)));
    layer1_outputs(7692) <= (layer0_outputs(8888)) or (layer0_outputs(6775));
    layer1_outputs(7693) <= not((layer0_outputs(6779)) and (layer0_outputs(4847)));
    layer1_outputs(7694) <= (layer0_outputs(1525)) and not (layer0_outputs(2059));
    layer1_outputs(7695) <= not(layer0_outputs(1488)) or (layer0_outputs(5404));
    layer1_outputs(7696) <= (layer0_outputs(10099)) and not (layer0_outputs(10227));
    layer1_outputs(7697) <= not((layer0_outputs(6952)) xor (layer0_outputs(3881)));
    layer1_outputs(7698) <= (layer0_outputs(8019)) and not (layer0_outputs(4678));
    layer1_outputs(7699) <= layer0_outputs(8507);
    layer1_outputs(7700) <= layer0_outputs(4875);
    layer1_outputs(7701) <= not((layer0_outputs(2134)) or (layer0_outputs(8222)));
    layer1_outputs(7702) <= not((layer0_outputs(851)) xor (layer0_outputs(1187)));
    layer1_outputs(7703) <= (layer0_outputs(6213)) and (layer0_outputs(5974));
    layer1_outputs(7704) <= layer0_outputs(6841);
    layer1_outputs(7705) <= not((layer0_outputs(5811)) or (layer0_outputs(7976)));
    layer1_outputs(7706) <= not(layer0_outputs(4232)) or (layer0_outputs(3203));
    layer1_outputs(7707) <= layer0_outputs(5687);
    layer1_outputs(7708) <= layer0_outputs(9660);
    layer1_outputs(7709) <= not(layer0_outputs(7109));
    layer1_outputs(7710) <= not((layer0_outputs(9672)) xor (layer0_outputs(7164)));
    layer1_outputs(7711) <= (layer0_outputs(8215)) and (layer0_outputs(4690));
    layer1_outputs(7712) <= not(layer0_outputs(1222));
    layer1_outputs(7713) <= not(layer0_outputs(2960));
    layer1_outputs(7714) <= layer0_outputs(1627);
    layer1_outputs(7715) <= not((layer0_outputs(1204)) xor (layer0_outputs(3519)));
    layer1_outputs(7716) <= (layer0_outputs(9427)) and (layer0_outputs(5638));
    layer1_outputs(7717) <= '1';
    layer1_outputs(7718) <= not((layer0_outputs(7950)) and (layer0_outputs(8937)));
    layer1_outputs(7719) <= not(layer0_outputs(2624));
    layer1_outputs(7720) <= (layer0_outputs(2835)) and (layer0_outputs(9573));
    layer1_outputs(7721) <= not((layer0_outputs(4000)) xor (layer0_outputs(100)));
    layer1_outputs(7722) <= not((layer0_outputs(4685)) and (layer0_outputs(9125)));
    layer1_outputs(7723) <= not(layer0_outputs(8324)) or (layer0_outputs(3886));
    layer1_outputs(7724) <= (layer0_outputs(8544)) xor (layer0_outputs(6064));
    layer1_outputs(7725) <= (layer0_outputs(8797)) and not (layer0_outputs(4984));
    layer1_outputs(7726) <= (layer0_outputs(8388)) and not (layer0_outputs(8554));
    layer1_outputs(7727) <= not(layer0_outputs(6036));
    layer1_outputs(7728) <= not(layer0_outputs(10193));
    layer1_outputs(7729) <= layer0_outputs(6630);
    layer1_outputs(7730) <= not((layer0_outputs(1348)) or (layer0_outputs(3684)));
    layer1_outputs(7731) <= not((layer0_outputs(2858)) xor (layer0_outputs(8776)));
    layer1_outputs(7732) <= layer0_outputs(4402);
    layer1_outputs(7733) <= not(layer0_outputs(1146)) or (layer0_outputs(2537));
    layer1_outputs(7734) <= (layer0_outputs(3535)) and (layer0_outputs(769));
    layer1_outputs(7735) <= not((layer0_outputs(10200)) and (layer0_outputs(5342)));
    layer1_outputs(7736) <= layer0_outputs(3923);
    layer1_outputs(7737) <= (layer0_outputs(1903)) or (layer0_outputs(889));
    layer1_outputs(7738) <= not((layer0_outputs(9908)) and (layer0_outputs(84)));
    layer1_outputs(7739) <= not((layer0_outputs(5789)) and (layer0_outputs(9286)));
    layer1_outputs(7740) <= layer0_outputs(169);
    layer1_outputs(7741) <= not(layer0_outputs(2801));
    layer1_outputs(7742) <= not(layer0_outputs(8915));
    layer1_outputs(7743) <= not((layer0_outputs(5838)) xor (layer0_outputs(3309)));
    layer1_outputs(7744) <= (layer0_outputs(4306)) and not (layer0_outputs(9676));
    layer1_outputs(7745) <= not(layer0_outputs(755)) or (layer0_outputs(1676));
    layer1_outputs(7746) <= (layer0_outputs(7334)) or (layer0_outputs(2877));
    layer1_outputs(7747) <= (layer0_outputs(5193)) and not (layer0_outputs(9793));
    layer1_outputs(7748) <= not(layer0_outputs(8193));
    layer1_outputs(7749) <= (layer0_outputs(4649)) and not (layer0_outputs(3204));
    layer1_outputs(7750) <= layer0_outputs(6588);
    layer1_outputs(7751) <= not(layer0_outputs(7507)) or (layer0_outputs(9546));
    layer1_outputs(7752) <= not(layer0_outputs(4055)) or (layer0_outputs(8144));
    layer1_outputs(7753) <= layer0_outputs(2371);
    layer1_outputs(7754) <= layer0_outputs(7127);
    layer1_outputs(7755) <= not((layer0_outputs(7262)) xor (layer0_outputs(3306)));
    layer1_outputs(7756) <= (layer0_outputs(719)) and (layer0_outputs(3989));
    layer1_outputs(7757) <= not((layer0_outputs(9446)) or (layer0_outputs(585)));
    layer1_outputs(7758) <= not((layer0_outputs(10204)) or (layer0_outputs(3224)));
    layer1_outputs(7759) <= not(layer0_outputs(1198));
    layer1_outputs(7760) <= (layer0_outputs(190)) and (layer0_outputs(6370));
    layer1_outputs(7761) <= not((layer0_outputs(6340)) and (layer0_outputs(1384)));
    layer1_outputs(7762) <= layer0_outputs(7120);
    layer1_outputs(7763) <= layer0_outputs(6738);
    layer1_outputs(7764) <= not(layer0_outputs(5767));
    layer1_outputs(7765) <= layer0_outputs(6991);
    layer1_outputs(7766) <= not((layer0_outputs(10003)) xor (layer0_outputs(3904)));
    layer1_outputs(7767) <= '1';
    layer1_outputs(7768) <= not((layer0_outputs(7433)) xor (layer0_outputs(3205)));
    layer1_outputs(7769) <= (layer0_outputs(670)) and (layer0_outputs(7577));
    layer1_outputs(7770) <= (layer0_outputs(5729)) and (layer0_outputs(8766));
    layer1_outputs(7771) <= not((layer0_outputs(466)) or (layer0_outputs(4313)));
    layer1_outputs(7772) <= (layer0_outputs(5834)) and not (layer0_outputs(6418));
    layer1_outputs(7773) <= (layer0_outputs(8140)) and (layer0_outputs(4845));
    layer1_outputs(7774) <= '0';
    layer1_outputs(7775) <= not(layer0_outputs(7006)) or (layer0_outputs(7885));
    layer1_outputs(7776) <= (layer0_outputs(8206)) xor (layer0_outputs(6280));
    layer1_outputs(7777) <= layer0_outputs(7141);
    layer1_outputs(7778) <= not(layer0_outputs(428));
    layer1_outputs(7779) <= layer0_outputs(893);
    layer1_outputs(7780) <= layer0_outputs(1953);
    layer1_outputs(7781) <= layer0_outputs(2814);
    layer1_outputs(7782) <= layer0_outputs(3425);
    layer1_outputs(7783) <= not((layer0_outputs(8827)) or (layer0_outputs(1870)));
    layer1_outputs(7784) <= layer0_outputs(5271);
    layer1_outputs(7785) <= (layer0_outputs(1616)) and not (layer0_outputs(7709));
    layer1_outputs(7786) <= (layer0_outputs(3783)) xor (layer0_outputs(4642));
    layer1_outputs(7787) <= not((layer0_outputs(8743)) xor (layer0_outputs(682)));
    layer1_outputs(7788) <= not(layer0_outputs(6070)) or (layer0_outputs(3665));
    layer1_outputs(7789) <= not(layer0_outputs(6677));
    layer1_outputs(7790) <= '1';
    layer1_outputs(7791) <= (layer0_outputs(51)) and not (layer0_outputs(5480));
    layer1_outputs(7792) <= (layer0_outputs(5992)) xor (layer0_outputs(5876));
    layer1_outputs(7793) <= not((layer0_outputs(5249)) or (layer0_outputs(3323)));
    layer1_outputs(7794) <= (layer0_outputs(6907)) and not (layer0_outputs(971));
    layer1_outputs(7795) <= layer0_outputs(476);
    layer1_outputs(7796) <= not(layer0_outputs(8622)) or (layer0_outputs(2341));
    layer1_outputs(7797) <= layer0_outputs(1158);
    layer1_outputs(7798) <= not((layer0_outputs(4723)) and (layer0_outputs(2449)));
    layer1_outputs(7799) <= not((layer0_outputs(8945)) and (layer0_outputs(1792)));
    layer1_outputs(7800) <= layer0_outputs(585);
    layer1_outputs(7801) <= (layer0_outputs(7940)) and (layer0_outputs(6253));
    layer1_outputs(7802) <= layer0_outputs(2025);
    layer1_outputs(7803) <= (layer0_outputs(2752)) and (layer0_outputs(5829));
    layer1_outputs(7804) <= (layer0_outputs(947)) or (layer0_outputs(3811));
    layer1_outputs(7805) <= not(layer0_outputs(5603));
    layer1_outputs(7806) <= (layer0_outputs(9536)) and not (layer0_outputs(8501));
    layer1_outputs(7807) <= not(layer0_outputs(6009));
    layer1_outputs(7808) <= not(layer0_outputs(9777)) or (layer0_outputs(8852));
    layer1_outputs(7809) <= layer0_outputs(4949);
    layer1_outputs(7810) <= not(layer0_outputs(6363)) or (layer0_outputs(7053));
    layer1_outputs(7811) <= not((layer0_outputs(1790)) or (layer0_outputs(5073)));
    layer1_outputs(7812) <= not(layer0_outputs(830));
    layer1_outputs(7813) <= not((layer0_outputs(639)) and (layer0_outputs(2763)));
    layer1_outputs(7814) <= not(layer0_outputs(5551)) or (layer0_outputs(9760));
    layer1_outputs(7815) <= (layer0_outputs(7028)) or (layer0_outputs(8278));
    layer1_outputs(7816) <= layer0_outputs(9375);
    layer1_outputs(7817) <= layer0_outputs(4137);
    layer1_outputs(7818) <= layer0_outputs(6699);
    layer1_outputs(7819) <= (layer0_outputs(1826)) and not (layer0_outputs(2637));
    layer1_outputs(7820) <= not(layer0_outputs(2003)) or (layer0_outputs(10119));
    layer1_outputs(7821) <= not((layer0_outputs(9759)) xor (layer0_outputs(3230)));
    layer1_outputs(7822) <= layer0_outputs(2884);
    layer1_outputs(7823) <= not(layer0_outputs(2905));
    layer1_outputs(7824) <= (layer0_outputs(8559)) and not (layer0_outputs(9755));
    layer1_outputs(7825) <= (layer0_outputs(264)) and not (layer0_outputs(7008));
    layer1_outputs(7826) <= '0';
    layer1_outputs(7827) <= not(layer0_outputs(1889)) or (layer0_outputs(7898));
    layer1_outputs(7828) <= not((layer0_outputs(1132)) xor (layer0_outputs(6892)));
    layer1_outputs(7829) <= layer0_outputs(9462);
    layer1_outputs(7830) <= not(layer0_outputs(1341)) or (layer0_outputs(3706));
    layer1_outputs(7831) <= not(layer0_outputs(5013)) or (layer0_outputs(5058));
    layer1_outputs(7832) <= '0';
    layer1_outputs(7833) <= not((layer0_outputs(48)) xor (layer0_outputs(3532)));
    layer1_outputs(7834) <= layer0_outputs(7705);
    layer1_outputs(7835) <= not(layer0_outputs(5346));
    layer1_outputs(7836) <= (layer0_outputs(10140)) and not (layer0_outputs(9429));
    layer1_outputs(7837) <= (layer0_outputs(5427)) or (layer0_outputs(8000));
    layer1_outputs(7838) <= (layer0_outputs(2017)) and not (layer0_outputs(6657));
    layer1_outputs(7839) <= not((layer0_outputs(315)) or (layer0_outputs(3533)));
    layer1_outputs(7840) <= not(layer0_outputs(2697)) or (layer0_outputs(9266));
    layer1_outputs(7841) <= not((layer0_outputs(4550)) or (layer0_outputs(8207)));
    layer1_outputs(7842) <= (layer0_outputs(7927)) and not (layer0_outputs(3462));
    layer1_outputs(7843) <= (layer0_outputs(1951)) and not (layer0_outputs(841));
    layer1_outputs(7844) <= not(layer0_outputs(3227));
    layer1_outputs(7845) <= not(layer0_outputs(2308));
    layer1_outputs(7846) <= (layer0_outputs(3940)) xor (layer0_outputs(4052));
    layer1_outputs(7847) <= not((layer0_outputs(2915)) or (layer0_outputs(5672)));
    layer1_outputs(7848) <= (layer0_outputs(9061)) and not (layer0_outputs(287));
    layer1_outputs(7849) <= not((layer0_outputs(4391)) and (layer0_outputs(7047)));
    layer1_outputs(7850) <= not(layer0_outputs(7976));
    layer1_outputs(7851) <= not(layer0_outputs(5290)) or (layer0_outputs(422));
    layer1_outputs(7852) <= layer0_outputs(1279);
    layer1_outputs(7853) <= not((layer0_outputs(986)) or (layer0_outputs(8462)));
    layer1_outputs(7854) <= layer0_outputs(8229);
    layer1_outputs(7855) <= layer0_outputs(3683);
    layer1_outputs(7856) <= not(layer0_outputs(4986)) or (layer0_outputs(1278));
    layer1_outputs(7857) <= not((layer0_outputs(9198)) or (layer0_outputs(1768)));
    layer1_outputs(7858) <= layer0_outputs(940);
    layer1_outputs(7859) <= '0';
    layer1_outputs(7860) <= not(layer0_outputs(3342)) or (layer0_outputs(5608));
    layer1_outputs(7861) <= (layer0_outputs(4043)) and not (layer0_outputs(5993));
    layer1_outputs(7862) <= layer0_outputs(4902);
    layer1_outputs(7863) <= layer0_outputs(652);
    layer1_outputs(7864) <= not((layer0_outputs(9153)) or (layer0_outputs(3978)));
    layer1_outputs(7865) <= '0';
    layer1_outputs(7866) <= (layer0_outputs(8016)) and not (layer0_outputs(8917));
    layer1_outputs(7867) <= not(layer0_outputs(7032));
    layer1_outputs(7868) <= (layer0_outputs(4618)) and not (layer0_outputs(3333));
    layer1_outputs(7869) <= (layer0_outputs(4431)) and not (layer0_outputs(356));
    layer1_outputs(7870) <= not((layer0_outputs(7748)) or (layer0_outputs(3988)));
    layer1_outputs(7871) <= not(layer0_outputs(5579));
    layer1_outputs(7872) <= '1';
    layer1_outputs(7873) <= layer0_outputs(6930);
    layer1_outputs(7874) <= (layer0_outputs(7453)) or (layer0_outputs(7110));
    layer1_outputs(7875) <= not(layer0_outputs(1221)) or (layer0_outputs(6564));
    layer1_outputs(7876) <= (layer0_outputs(5880)) or (layer0_outputs(8982));
    layer1_outputs(7877) <= layer0_outputs(6010);
    layer1_outputs(7878) <= not(layer0_outputs(6783));
    layer1_outputs(7879) <= not((layer0_outputs(7812)) xor (layer0_outputs(3868)));
    layer1_outputs(7880) <= layer0_outputs(1759);
    layer1_outputs(7881) <= not(layer0_outputs(7739));
    layer1_outputs(7882) <= not(layer0_outputs(2944));
    layer1_outputs(7883) <= (layer0_outputs(8882)) or (layer0_outputs(1172));
    layer1_outputs(7884) <= not(layer0_outputs(9728)) or (layer0_outputs(8861));
    layer1_outputs(7885) <= not(layer0_outputs(7399));
    layer1_outputs(7886) <= not(layer0_outputs(7421));
    layer1_outputs(7887) <= not(layer0_outputs(711));
    layer1_outputs(7888) <= layer0_outputs(5275);
    layer1_outputs(7889) <= not(layer0_outputs(2999));
    layer1_outputs(7890) <= not(layer0_outputs(7587)) or (layer0_outputs(7708));
    layer1_outputs(7891) <= (layer0_outputs(7602)) or (layer0_outputs(817));
    layer1_outputs(7892) <= not((layer0_outputs(1049)) or (layer0_outputs(1911)));
    layer1_outputs(7893) <= '1';
    layer1_outputs(7894) <= not(layer0_outputs(4918)) or (layer0_outputs(2399));
    layer1_outputs(7895) <= not(layer0_outputs(5334));
    layer1_outputs(7896) <= not(layer0_outputs(4035));
    layer1_outputs(7897) <= (layer0_outputs(8543)) xor (layer0_outputs(8524));
    layer1_outputs(7898) <= not((layer0_outputs(9579)) and (layer0_outputs(6840)));
    layer1_outputs(7899) <= not(layer0_outputs(5818));
    layer1_outputs(7900) <= layer0_outputs(6758);
    layer1_outputs(7901) <= (layer0_outputs(516)) and (layer0_outputs(5057));
    layer1_outputs(7902) <= (layer0_outputs(2931)) and not (layer0_outputs(7797));
    layer1_outputs(7903) <= not((layer0_outputs(4093)) or (layer0_outputs(5520)));
    layer1_outputs(7904) <= (layer0_outputs(8892)) xor (layer0_outputs(7786));
    layer1_outputs(7905) <= not((layer0_outputs(7554)) xor (layer0_outputs(1026)));
    layer1_outputs(7906) <= not((layer0_outputs(5197)) and (layer0_outputs(8041)));
    layer1_outputs(7907) <= (layer0_outputs(3375)) or (layer0_outputs(5954));
    layer1_outputs(7908) <= (layer0_outputs(1374)) or (layer0_outputs(3894));
    layer1_outputs(7909) <= '0';
    layer1_outputs(7910) <= layer0_outputs(7232);
    layer1_outputs(7911) <= not(layer0_outputs(8612)) or (layer0_outputs(886));
    layer1_outputs(7912) <= not(layer0_outputs(3478)) or (layer0_outputs(5175));
    layer1_outputs(7913) <= '0';
    layer1_outputs(7914) <= not(layer0_outputs(8178)) or (layer0_outputs(4378));
    layer1_outputs(7915) <= '1';
    layer1_outputs(7916) <= (layer0_outputs(8161)) and not (layer0_outputs(2269));
    layer1_outputs(7917) <= (layer0_outputs(3643)) xor (layer0_outputs(8394));
    layer1_outputs(7918) <= not(layer0_outputs(941));
    layer1_outputs(7919) <= not(layer0_outputs(7359));
    layer1_outputs(7920) <= (layer0_outputs(5689)) or (layer0_outputs(9340));
    layer1_outputs(7921) <= not(layer0_outputs(6472));
    layer1_outputs(7922) <= not((layer0_outputs(4977)) and (layer0_outputs(5227)));
    layer1_outputs(7923) <= layer0_outputs(7089);
    layer1_outputs(7924) <= not(layer0_outputs(7651));
    layer1_outputs(7925) <= layer0_outputs(5527);
    layer1_outputs(7926) <= (layer0_outputs(2492)) and not (layer0_outputs(1035));
    layer1_outputs(7927) <= (layer0_outputs(5677)) xor (layer0_outputs(4561));
    layer1_outputs(7928) <= not((layer0_outputs(4715)) or (layer0_outputs(9742)));
    layer1_outputs(7929) <= (layer0_outputs(10220)) and not (layer0_outputs(3700));
    layer1_outputs(7930) <= (layer0_outputs(9226)) and not (layer0_outputs(4313));
    layer1_outputs(7931) <= (layer0_outputs(3023)) xor (layer0_outputs(7424));
    layer1_outputs(7932) <= (layer0_outputs(2298)) and not (layer0_outputs(5513));
    layer1_outputs(7933) <= (layer0_outputs(6501)) or (layer0_outputs(5873));
    layer1_outputs(7934) <= (layer0_outputs(3686)) or (layer0_outputs(9406));
    layer1_outputs(7935) <= (layer0_outputs(140)) or (layer0_outputs(4520));
    layer1_outputs(7936) <= not(layer0_outputs(1463));
    layer1_outputs(7937) <= layer0_outputs(5921);
    layer1_outputs(7938) <= layer0_outputs(2438);
    layer1_outputs(7939) <= not(layer0_outputs(8743));
    layer1_outputs(7940) <= (layer0_outputs(560)) and not (layer0_outputs(8929));
    layer1_outputs(7941) <= not((layer0_outputs(10192)) and (layer0_outputs(957)));
    layer1_outputs(7942) <= (layer0_outputs(4216)) and not (layer0_outputs(6600));
    layer1_outputs(7943) <= '1';
    layer1_outputs(7944) <= layer0_outputs(9371);
    layer1_outputs(7945) <= not(layer0_outputs(6214));
    layer1_outputs(7946) <= (layer0_outputs(937)) or (layer0_outputs(9936));
    layer1_outputs(7947) <= not(layer0_outputs(2741)) or (layer0_outputs(5002));
    layer1_outputs(7948) <= not(layer0_outputs(8129));
    layer1_outputs(7949) <= not(layer0_outputs(8250));
    layer1_outputs(7950) <= layer0_outputs(7727);
    layer1_outputs(7951) <= layer0_outputs(9386);
    layer1_outputs(7952) <= not(layer0_outputs(5792));
    layer1_outputs(7953) <= layer0_outputs(8476);
    layer1_outputs(7954) <= not((layer0_outputs(5997)) and (layer0_outputs(3605)));
    layer1_outputs(7955) <= layer0_outputs(6124);
    layer1_outputs(7956) <= not(layer0_outputs(1187));
    layer1_outputs(7957) <= not(layer0_outputs(8301));
    layer1_outputs(7958) <= not((layer0_outputs(7209)) xor (layer0_outputs(1320)));
    layer1_outputs(7959) <= (layer0_outputs(1739)) or (layer0_outputs(1708));
    layer1_outputs(7960) <= (layer0_outputs(9090)) and not (layer0_outputs(763));
    layer1_outputs(7961) <= (layer0_outputs(1001)) or (layer0_outputs(4455));
    layer1_outputs(7962) <= not((layer0_outputs(8790)) or (layer0_outputs(5195)));
    layer1_outputs(7963) <= (layer0_outputs(4351)) or (layer0_outputs(786));
    layer1_outputs(7964) <= (layer0_outputs(6236)) and (layer0_outputs(2791));
    layer1_outputs(7965) <= not((layer0_outputs(776)) or (layer0_outputs(7136)));
    layer1_outputs(7966) <= (layer0_outputs(5362)) xor (layer0_outputs(5757));
    layer1_outputs(7967) <= not(layer0_outputs(3077));
    layer1_outputs(7968) <= not((layer0_outputs(1775)) xor (layer0_outputs(9944)));
    layer1_outputs(7969) <= not(layer0_outputs(9772));
    layer1_outputs(7970) <= '1';
    layer1_outputs(7971) <= not((layer0_outputs(1273)) and (layer0_outputs(3045)));
    layer1_outputs(7972) <= not(layer0_outputs(2263)) or (layer0_outputs(130));
    layer1_outputs(7973) <= not(layer0_outputs(2303));
    layer1_outputs(7974) <= not(layer0_outputs(5788));
    layer1_outputs(7975) <= not(layer0_outputs(8672)) or (layer0_outputs(3779));
    layer1_outputs(7976) <= (layer0_outputs(2793)) xor (layer0_outputs(6532));
    layer1_outputs(7977) <= layer0_outputs(2595);
    layer1_outputs(7978) <= (layer0_outputs(3554)) and not (layer0_outputs(1418));
    layer1_outputs(7979) <= layer0_outputs(4736);
    layer1_outputs(7980) <= layer0_outputs(9165);
    layer1_outputs(7981) <= (layer0_outputs(5928)) and not (layer0_outputs(1158));
    layer1_outputs(7982) <= not((layer0_outputs(1657)) or (layer0_outputs(4626)));
    layer1_outputs(7983) <= not((layer0_outputs(2263)) xor (layer0_outputs(7242)));
    layer1_outputs(7984) <= (layer0_outputs(4607)) xor (layer0_outputs(4861));
    layer1_outputs(7985) <= (layer0_outputs(519)) and not (layer0_outputs(7588));
    layer1_outputs(7986) <= (layer0_outputs(2366)) and not (layer0_outputs(5048));
    layer1_outputs(7987) <= not((layer0_outputs(8725)) xor (layer0_outputs(3130)));
    layer1_outputs(7988) <= not((layer0_outputs(9465)) and (layer0_outputs(8511)));
    layer1_outputs(7989) <= (layer0_outputs(8141)) and not (layer0_outputs(1924));
    layer1_outputs(7990) <= not(layer0_outputs(2388));
    layer1_outputs(7991) <= layer0_outputs(2463);
    layer1_outputs(7992) <= not(layer0_outputs(4485));
    layer1_outputs(7993) <= not(layer0_outputs(6222)) or (layer0_outputs(9681));
    layer1_outputs(7994) <= not((layer0_outputs(5422)) or (layer0_outputs(5557)));
    layer1_outputs(7995) <= layer0_outputs(1404);
    layer1_outputs(7996) <= (layer0_outputs(8155)) and not (layer0_outputs(310));
    layer1_outputs(7997) <= not(layer0_outputs(3243));
    layer1_outputs(7998) <= not(layer0_outputs(6119));
    layer1_outputs(7999) <= layer0_outputs(5942);
    layer1_outputs(8000) <= '1';
    layer1_outputs(8001) <= layer0_outputs(2505);
    layer1_outputs(8002) <= layer0_outputs(3106);
    layer1_outputs(8003) <= not(layer0_outputs(1440));
    layer1_outputs(8004) <= (layer0_outputs(4829)) or (layer0_outputs(5094));
    layer1_outputs(8005) <= layer0_outputs(8801);
    layer1_outputs(8006) <= not((layer0_outputs(6324)) and (layer0_outputs(1611)));
    layer1_outputs(8007) <= (layer0_outputs(4872)) and not (layer0_outputs(3010));
    layer1_outputs(8008) <= not((layer0_outputs(8166)) xor (layer0_outputs(7818)));
    layer1_outputs(8009) <= (layer0_outputs(2752)) and not (layer0_outputs(8099));
    layer1_outputs(8010) <= not(layer0_outputs(6675));
    layer1_outputs(8011) <= not(layer0_outputs(1933)) or (layer0_outputs(6631));
    layer1_outputs(8012) <= layer0_outputs(2562);
    layer1_outputs(8013) <= not(layer0_outputs(2156));
    layer1_outputs(8014) <= not(layer0_outputs(3567));
    layer1_outputs(8015) <= (layer0_outputs(3675)) and (layer0_outputs(2463));
    layer1_outputs(8016) <= not(layer0_outputs(7880));
    layer1_outputs(8017) <= not((layer0_outputs(7760)) or (layer0_outputs(5764)));
    layer1_outputs(8018) <= not(layer0_outputs(2320));
    layer1_outputs(8019) <= not(layer0_outputs(3321)) or (layer0_outputs(4721));
    layer1_outputs(8020) <= layer0_outputs(5944);
    layer1_outputs(8021) <= not(layer0_outputs(2800)) or (layer0_outputs(3324));
    layer1_outputs(8022) <= not(layer0_outputs(4669)) or (layer0_outputs(4883));
    layer1_outputs(8023) <= not(layer0_outputs(3782)) or (layer0_outputs(6873));
    layer1_outputs(8024) <= not(layer0_outputs(2120));
    layer1_outputs(8025) <= not(layer0_outputs(967));
    layer1_outputs(8026) <= not(layer0_outputs(5894));
    layer1_outputs(8027) <= not(layer0_outputs(9838));
    layer1_outputs(8028) <= layer0_outputs(6950);
    layer1_outputs(8029) <= not(layer0_outputs(2116));
    layer1_outputs(8030) <= not((layer0_outputs(9199)) or (layer0_outputs(1097)));
    layer1_outputs(8031) <= '0';
    layer1_outputs(8032) <= not((layer0_outputs(7292)) and (layer0_outputs(3518)));
    layer1_outputs(8033) <= layer0_outputs(8692);
    layer1_outputs(8034) <= (layer0_outputs(7619)) or (layer0_outputs(6904));
    layer1_outputs(8035) <= not(layer0_outputs(3767)) or (layer0_outputs(9655));
    layer1_outputs(8036) <= not(layer0_outputs(1087));
    layer1_outputs(8037) <= layer0_outputs(8371);
    layer1_outputs(8038) <= '1';
    layer1_outputs(8039) <= not(layer0_outputs(7364)) or (layer0_outputs(9672));
    layer1_outputs(8040) <= not(layer0_outputs(10006)) or (layer0_outputs(6943));
    layer1_outputs(8041) <= '1';
    layer1_outputs(8042) <= not((layer0_outputs(4345)) and (layer0_outputs(3958)));
    layer1_outputs(8043) <= layer0_outputs(2139);
    layer1_outputs(8044) <= layer0_outputs(2239);
    layer1_outputs(8045) <= (layer0_outputs(2106)) and (layer0_outputs(42));
    layer1_outputs(8046) <= not(layer0_outputs(7233));
    layer1_outputs(8047) <= '1';
    layer1_outputs(8048) <= layer0_outputs(8562);
    layer1_outputs(8049) <= not(layer0_outputs(8176));
    layer1_outputs(8050) <= not(layer0_outputs(2074));
    layer1_outputs(8051) <= layer0_outputs(1179);
    layer1_outputs(8052) <= (layer0_outputs(1604)) or (layer0_outputs(9430));
    layer1_outputs(8053) <= not((layer0_outputs(4182)) or (layer0_outputs(9035)));
    layer1_outputs(8054) <= not(layer0_outputs(1171));
    layer1_outputs(8055) <= not((layer0_outputs(5719)) and (layer0_outputs(9903)));
    layer1_outputs(8056) <= layer0_outputs(1135);
    layer1_outputs(8057) <= not(layer0_outputs(9418)) or (layer0_outputs(4222));
    layer1_outputs(8058) <= not(layer0_outputs(2531));
    layer1_outputs(8059) <= not(layer0_outputs(3655)) or (layer0_outputs(667));
    layer1_outputs(8060) <= layer0_outputs(49);
    layer1_outputs(8061) <= not(layer0_outputs(8243));
    layer1_outputs(8062) <= not(layer0_outputs(6911));
    layer1_outputs(8063) <= layer0_outputs(1843);
    layer1_outputs(8064) <= not((layer0_outputs(7466)) and (layer0_outputs(8997)));
    layer1_outputs(8065) <= not((layer0_outputs(914)) and (layer0_outputs(5239)));
    layer1_outputs(8066) <= (layer0_outputs(3039)) and not (layer0_outputs(8477));
    layer1_outputs(8067) <= not(layer0_outputs(4122)) or (layer0_outputs(9247));
    layer1_outputs(8068) <= (layer0_outputs(3045)) and (layer0_outputs(5752));
    layer1_outputs(8069) <= not(layer0_outputs(5707)) or (layer0_outputs(4307));
    layer1_outputs(8070) <= not(layer0_outputs(1572));
    layer1_outputs(8071) <= layer0_outputs(2103);
    layer1_outputs(8072) <= not(layer0_outputs(5963));
    layer1_outputs(8073) <= not(layer0_outputs(5906));
    layer1_outputs(8074) <= not(layer0_outputs(1999)) or (layer0_outputs(10173));
    layer1_outputs(8075) <= not((layer0_outputs(6611)) or (layer0_outputs(9202)));
    layer1_outputs(8076) <= (layer0_outputs(8806)) and not (layer0_outputs(3914));
    layer1_outputs(8077) <= layer0_outputs(7353);
    layer1_outputs(8078) <= not(layer0_outputs(7660)) or (layer0_outputs(6740));
    layer1_outputs(8079) <= not(layer0_outputs(6487));
    layer1_outputs(8080) <= not((layer0_outputs(7695)) and (layer0_outputs(9830)));
    layer1_outputs(8081) <= layer0_outputs(415);
    layer1_outputs(8082) <= not(layer0_outputs(10206)) or (layer0_outputs(2207));
    layer1_outputs(8083) <= (layer0_outputs(5927)) xor (layer0_outputs(2150));
    layer1_outputs(8084) <= not((layer0_outputs(665)) and (layer0_outputs(7902)));
    layer1_outputs(8085) <= layer0_outputs(5703);
    layer1_outputs(8086) <= not((layer0_outputs(10215)) and (layer0_outputs(9072)));
    layer1_outputs(8087) <= not((layer0_outputs(582)) or (layer0_outputs(5907)));
    layer1_outputs(8088) <= not((layer0_outputs(5412)) or (layer0_outputs(8426)));
    layer1_outputs(8089) <= not(layer0_outputs(2815)) or (layer0_outputs(10205));
    layer1_outputs(8090) <= layer0_outputs(7174);
    layer1_outputs(8091) <= layer0_outputs(823);
    layer1_outputs(8092) <= not(layer0_outputs(4748));
    layer1_outputs(8093) <= layer0_outputs(4391);
    layer1_outputs(8094) <= not(layer0_outputs(5202)) or (layer0_outputs(3315));
    layer1_outputs(8095) <= (layer0_outputs(4003)) and not (layer0_outputs(7775));
    layer1_outputs(8096) <= not(layer0_outputs(210));
    layer1_outputs(8097) <= (layer0_outputs(5882)) or (layer0_outputs(1660));
    layer1_outputs(8098) <= not((layer0_outputs(7611)) xor (layer0_outputs(7860)));
    layer1_outputs(8099) <= layer0_outputs(2651);
    layer1_outputs(8100) <= layer0_outputs(3028);
    layer1_outputs(8101) <= not(layer0_outputs(6411));
    layer1_outputs(8102) <= (layer0_outputs(6969)) and not (layer0_outputs(9000));
    layer1_outputs(8103) <= (layer0_outputs(5905)) and (layer0_outputs(1829));
    layer1_outputs(8104) <= not(layer0_outputs(1414)) or (layer0_outputs(9479));
    layer1_outputs(8105) <= not(layer0_outputs(4663)) or (layer0_outputs(7223));
    layer1_outputs(8106) <= layer0_outputs(7948);
    layer1_outputs(8107) <= not((layer0_outputs(301)) and (layer0_outputs(9275)));
    layer1_outputs(8108) <= not(layer0_outputs(4583)) or (layer0_outputs(8290));
    layer1_outputs(8109) <= not(layer0_outputs(8960));
    layer1_outputs(8110) <= not(layer0_outputs(2790));
    layer1_outputs(8111) <= not(layer0_outputs(5893));
    layer1_outputs(8112) <= layer0_outputs(4095);
    layer1_outputs(8113) <= layer0_outputs(2465);
    layer1_outputs(8114) <= (layer0_outputs(8903)) xor (layer0_outputs(2082));
    layer1_outputs(8115) <= layer0_outputs(9935);
    layer1_outputs(8116) <= (layer0_outputs(5168)) and (layer0_outputs(2200));
    layer1_outputs(8117) <= (layer0_outputs(95)) xor (layer0_outputs(3535));
    layer1_outputs(8118) <= not(layer0_outputs(1553)) or (layer0_outputs(9936));
    layer1_outputs(8119) <= not(layer0_outputs(3121));
    layer1_outputs(8120) <= not(layer0_outputs(61));
    layer1_outputs(8121) <= not(layer0_outputs(6051));
    layer1_outputs(8122) <= not((layer0_outputs(5326)) or (layer0_outputs(8662)));
    layer1_outputs(8123) <= (layer0_outputs(9575)) or (layer0_outputs(9210));
    layer1_outputs(8124) <= not((layer0_outputs(7674)) or (layer0_outputs(9382)));
    layer1_outputs(8125) <= (layer0_outputs(6439)) and (layer0_outputs(2550));
    layer1_outputs(8126) <= not(layer0_outputs(514));
    layer1_outputs(8127) <= not((layer0_outputs(5826)) or (layer0_outputs(3277)));
    layer1_outputs(8128) <= not(layer0_outputs(7123));
    layer1_outputs(8129) <= (layer0_outputs(6308)) xor (layer0_outputs(8346));
    layer1_outputs(8130) <= '0';
    layer1_outputs(8131) <= not(layer0_outputs(7583)) or (layer0_outputs(1575));
    layer1_outputs(8132) <= layer0_outputs(2965);
    layer1_outputs(8133) <= (layer0_outputs(10145)) xor (layer0_outputs(2638));
    layer1_outputs(8134) <= (layer0_outputs(994)) or (layer0_outputs(5466));
    layer1_outputs(8135) <= layer0_outputs(8568);
    layer1_outputs(8136) <= not(layer0_outputs(8020));
    layer1_outputs(8137) <= not((layer0_outputs(6851)) and (layer0_outputs(1863)));
    layer1_outputs(8138) <= not(layer0_outputs(1731));
    layer1_outputs(8139) <= (layer0_outputs(8653)) xor (layer0_outputs(1670));
    layer1_outputs(8140) <= layer0_outputs(3290);
    layer1_outputs(8141) <= layer0_outputs(8317);
    layer1_outputs(8142) <= (layer0_outputs(2900)) or (layer0_outputs(9747));
    layer1_outputs(8143) <= not((layer0_outputs(7400)) or (layer0_outputs(340)));
    layer1_outputs(8144) <= (layer0_outputs(5229)) or (layer0_outputs(6298));
    layer1_outputs(8145) <= (layer0_outputs(9709)) and not (layer0_outputs(4591));
    layer1_outputs(8146) <= not(layer0_outputs(4219));
    layer1_outputs(8147) <= not((layer0_outputs(1274)) xor (layer0_outputs(8040)));
    layer1_outputs(8148) <= '1';
    layer1_outputs(8149) <= layer0_outputs(7163);
    layer1_outputs(8150) <= (layer0_outputs(740)) and (layer0_outputs(1983));
    layer1_outputs(8151) <= not((layer0_outputs(7170)) xor (layer0_outputs(674)));
    layer1_outputs(8152) <= not((layer0_outputs(10036)) and (layer0_outputs(442)));
    layer1_outputs(8153) <= not((layer0_outputs(4587)) and (layer0_outputs(3981)));
    layer1_outputs(8154) <= not((layer0_outputs(8234)) and (layer0_outputs(2039)));
    layer1_outputs(8155) <= (layer0_outputs(1101)) xor (layer0_outputs(5196));
    layer1_outputs(8156) <= not(layer0_outputs(3829)) or (layer0_outputs(5341));
    layer1_outputs(8157) <= not(layer0_outputs(4562));
    layer1_outputs(8158) <= layer0_outputs(2240);
    layer1_outputs(8159) <= layer0_outputs(4883);
    layer1_outputs(8160) <= layer0_outputs(8003);
    layer1_outputs(8161) <= not(layer0_outputs(9486));
    layer1_outputs(8162) <= layer0_outputs(7519);
    layer1_outputs(8163) <= layer0_outputs(7309);
    layer1_outputs(8164) <= (layer0_outputs(8923)) and not (layer0_outputs(4343));
    layer1_outputs(8165) <= (layer0_outputs(3711)) and not (layer0_outputs(2767));
    layer1_outputs(8166) <= not(layer0_outputs(750));
    layer1_outputs(8167) <= not(layer0_outputs(10088));
    layer1_outputs(8168) <= (layer0_outputs(1614)) and not (layer0_outputs(3504));
    layer1_outputs(8169) <= not((layer0_outputs(8532)) xor (layer0_outputs(8710)));
    layer1_outputs(8170) <= '0';
    layer1_outputs(8171) <= not((layer0_outputs(5377)) and (layer0_outputs(180)));
    layer1_outputs(8172) <= not(layer0_outputs(6330)) or (layer0_outputs(3932));
    layer1_outputs(8173) <= not((layer0_outputs(2909)) or (layer0_outputs(9746)));
    layer1_outputs(8174) <= not((layer0_outputs(9707)) or (layer0_outputs(8001)));
    layer1_outputs(8175) <= (layer0_outputs(5997)) and not (layer0_outputs(4202));
    layer1_outputs(8176) <= not(layer0_outputs(4084));
    layer1_outputs(8177) <= not(layer0_outputs(2623));
    layer1_outputs(8178) <= layer0_outputs(3191);
    layer1_outputs(8179) <= not(layer0_outputs(6264)) or (layer0_outputs(9853));
    layer1_outputs(8180) <= not((layer0_outputs(5826)) and (layer0_outputs(7199)));
    layer1_outputs(8181) <= (layer0_outputs(2754)) and not (layer0_outputs(7552));
    layer1_outputs(8182) <= layer0_outputs(4851);
    layer1_outputs(8183) <= not(layer0_outputs(5560));
    layer1_outputs(8184) <= not(layer0_outputs(3339));
    layer1_outputs(8185) <= not(layer0_outputs(3676)) or (layer0_outputs(8752));
    layer1_outputs(8186) <= not(layer0_outputs(6166)) or (layer0_outputs(3727));
    layer1_outputs(8187) <= not(layer0_outputs(3825));
    layer1_outputs(8188) <= not(layer0_outputs(7764));
    layer1_outputs(8189) <= layer0_outputs(4114);
    layer1_outputs(8190) <= (layer0_outputs(2280)) or (layer0_outputs(10217));
    layer1_outputs(8191) <= not((layer0_outputs(9103)) or (layer0_outputs(9355)));
    layer1_outputs(8192) <= not(layer0_outputs(1957));
    layer1_outputs(8193) <= (layer0_outputs(9687)) and not (layer0_outputs(5349));
    layer1_outputs(8194) <= not(layer0_outputs(2883));
    layer1_outputs(8195) <= not(layer0_outputs(97)) or (layer0_outputs(6556));
    layer1_outputs(8196) <= (layer0_outputs(8330)) or (layer0_outputs(6743));
    layer1_outputs(8197) <= not((layer0_outputs(6032)) xor (layer0_outputs(423)));
    layer1_outputs(8198) <= not(layer0_outputs(2812)) or (layer0_outputs(7384));
    layer1_outputs(8199) <= (layer0_outputs(997)) and not (layer0_outputs(6059));
    layer1_outputs(8200) <= not((layer0_outputs(110)) and (layer0_outputs(9735)));
    layer1_outputs(8201) <= not(layer0_outputs(4838));
    layer1_outputs(8202) <= not(layer0_outputs(3393));
    layer1_outputs(8203) <= layer0_outputs(2510);
    layer1_outputs(8204) <= (layer0_outputs(2451)) and not (layer0_outputs(6797));
    layer1_outputs(8205) <= not(layer0_outputs(9803));
    layer1_outputs(8206) <= (layer0_outputs(2681)) and not (layer0_outputs(98));
    layer1_outputs(8207) <= (layer0_outputs(7302)) and (layer0_outputs(6294));
    layer1_outputs(8208) <= not((layer0_outputs(78)) xor (layer0_outputs(6772)));
    layer1_outputs(8209) <= layer0_outputs(6917);
    layer1_outputs(8210) <= (layer0_outputs(4880)) and not (layer0_outputs(2714));
    layer1_outputs(8211) <= (layer0_outputs(7781)) and (layer0_outputs(485));
    layer1_outputs(8212) <= layer0_outputs(2982);
    layer1_outputs(8213) <= (layer0_outputs(9548)) and not (layer0_outputs(905));
    layer1_outputs(8214) <= not((layer0_outputs(9876)) xor (layer0_outputs(5582)));
    layer1_outputs(8215) <= layer0_outputs(5883);
    layer1_outputs(8216) <= not(layer0_outputs(8747));
    layer1_outputs(8217) <= not(layer0_outputs(6502));
    layer1_outputs(8218) <= layer0_outputs(4078);
    layer1_outputs(8219) <= layer0_outputs(9299);
    layer1_outputs(8220) <= layer0_outputs(2026);
    layer1_outputs(8221) <= not(layer0_outputs(2840));
    layer1_outputs(8222) <= layer0_outputs(9207);
    layer1_outputs(8223) <= layer0_outputs(2918);
    layer1_outputs(8224) <= layer0_outputs(8665);
    layer1_outputs(8225) <= (layer0_outputs(3081)) and not (layer0_outputs(5387));
    layer1_outputs(8226) <= not((layer0_outputs(2810)) xor (layer0_outputs(6380)));
    layer1_outputs(8227) <= (layer0_outputs(158)) and not (layer0_outputs(6891));
    layer1_outputs(8228) <= layer0_outputs(4277);
    layer1_outputs(8229) <= layer0_outputs(5204);
    layer1_outputs(8230) <= (layer0_outputs(3789)) or (layer0_outputs(8315));
    layer1_outputs(8231) <= not((layer0_outputs(5708)) and (layer0_outputs(1561)));
    layer1_outputs(8232) <= layer0_outputs(6385);
    layer1_outputs(8233) <= (layer0_outputs(628)) and not (layer0_outputs(8733));
    layer1_outputs(8234) <= not((layer0_outputs(7832)) xor (layer0_outputs(1589)));
    layer1_outputs(8235) <= not(layer0_outputs(4162)) or (layer0_outputs(8244));
    layer1_outputs(8236) <= not(layer0_outputs(361));
    layer1_outputs(8237) <= not(layer0_outputs(2261));
    layer1_outputs(8238) <= not(layer0_outputs(7101));
    layer1_outputs(8239) <= not(layer0_outputs(6210));
    layer1_outputs(8240) <= layer0_outputs(6523);
    layer1_outputs(8241) <= (layer0_outputs(7693)) or (layer0_outputs(9995));
    layer1_outputs(8242) <= '0';
    layer1_outputs(8243) <= not(layer0_outputs(9024)) or (layer0_outputs(5674));
    layer1_outputs(8244) <= not((layer0_outputs(4452)) or (layer0_outputs(8002)));
    layer1_outputs(8245) <= (layer0_outputs(8181)) or (layer0_outputs(4329));
    layer1_outputs(8246) <= layer0_outputs(5275);
    layer1_outputs(8247) <= layer0_outputs(8568);
    layer1_outputs(8248) <= (layer0_outputs(753)) or (layer0_outputs(515));
    layer1_outputs(8249) <= not(layer0_outputs(7623));
    layer1_outputs(8250) <= not(layer0_outputs(1813));
    layer1_outputs(8251) <= layer0_outputs(9674);
    layer1_outputs(8252) <= not(layer0_outputs(1208));
    layer1_outputs(8253) <= layer0_outputs(2534);
    layer1_outputs(8254) <= (layer0_outputs(3679)) and not (layer0_outputs(5503));
    layer1_outputs(8255) <= not(layer0_outputs(8228)) or (layer0_outputs(6691));
    layer1_outputs(8256) <= layer0_outputs(8015);
    layer1_outputs(8257) <= layer0_outputs(4960);
    layer1_outputs(8258) <= not(layer0_outputs(9778));
    layer1_outputs(8259) <= not(layer0_outputs(7537));
    layer1_outputs(8260) <= '0';
    layer1_outputs(8261) <= '1';
    layer1_outputs(8262) <= not((layer0_outputs(3389)) and (layer0_outputs(2462)));
    layer1_outputs(8263) <= not((layer0_outputs(1350)) and (layer0_outputs(1698)));
    layer1_outputs(8264) <= not((layer0_outputs(2564)) or (layer0_outputs(4934)));
    layer1_outputs(8265) <= not(layer0_outputs(6465)) or (layer0_outputs(9271));
    layer1_outputs(8266) <= (layer0_outputs(783)) xor (layer0_outputs(29));
    layer1_outputs(8267) <= not(layer0_outputs(10));
    layer1_outputs(8268) <= (layer0_outputs(63)) or (layer0_outputs(7540));
    layer1_outputs(8269) <= not(layer0_outputs(8333));
    layer1_outputs(8270) <= layer0_outputs(8649);
    layer1_outputs(8271) <= not(layer0_outputs(3116));
    layer1_outputs(8272) <= (layer0_outputs(6720)) and not (layer0_outputs(1851));
    layer1_outputs(8273) <= not(layer0_outputs(7955));
    layer1_outputs(8274) <= (layer0_outputs(4374)) and (layer0_outputs(5889));
    layer1_outputs(8275) <= not(layer0_outputs(5107));
    layer1_outputs(8276) <= layer0_outputs(10037);
    layer1_outputs(8277) <= not(layer0_outputs(5822));
    layer1_outputs(8278) <= not(layer0_outputs(6268));
    layer1_outputs(8279) <= not(layer0_outputs(8936));
    layer1_outputs(8280) <= not(layer0_outputs(2380)) or (layer0_outputs(8872));
    layer1_outputs(8281) <= layer0_outputs(5394);
    layer1_outputs(8282) <= layer0_outputs(3098);
    layer1_outputs(8283) <= not((layer0_outputs(814)) xor (layer0_outputs(4475)));
    layer1_outputs(8284) <= layer0_outputs(8800);
    layer1_outputs(8285) <= not((layer0_outputs(8655)) xor (layer0_outputs(7590)));
    layer1_outputs(8286) <= (layer0_outputs(2507)) and (layer0_outputs(6419));
    layer1_outputs(8287) <= (layer0_outputs(3661)) and not (layer0_outputs(4750));
    layer1_outputs(8288) <= not((layer0_outputs(591)) and (layer0_outputs(1145)));
    layer1_outputs(8289) <= not(layer0_outputs(3079));
    layer1_outputs(8290) <= not(layer0_outputs(3549)) or (layer0_outputs(2591));
    layer1_outputs(8291) <= (layer0_outputs(4294)) and not (layer0_outputs(6316));
    layer1_outputs(8292) <= layer0_outputs(6539);
    layer1_outputs(8293) <= (layer0_outputs(9257)) or (layer0_outputs(4412));
    layer1_outputs(8294) <= (layer0_outputs(9891)) and not (layer0_outputs(4964));
    layer1_outputs(8295) <= '0';
    layer1_outputs(8296) <= (layer0_outputs(854)) and not (layer0_outputs(7495));
    layer1_outputs(8297) <= layer0_outputs(9979);
    layer1_outputs(8298) <= (layer0_outputs(7566)) and not (layer0_outputs(6816));
    layer1_outputs(8299) <= not(layer0_outputs(4621));
    layer1_outputs(8300) <= not(layer0_outputs(3253));
    layer1_outputs(8301) <= (layer0_outputs(10148)) or (layer0_outputs(6055));
    layer1_outputs(8302) <= not((layer0_outputs(892)) or (layer0_outputs(5125)));
    layer1_outputs(8303) <= not(layer0_outputs(5702));
    layer1_outputs(8304) <= (layer0_outputs(3265)) and not (layer0_outputs(4860));
    layer1_outputs(8305) <= (layer0_outputs(6300)) and (layer0_outputs(7855));
    layer1_outputs(8306) <= not(layer0_outputs(7180));
    layer1_outputs(8307) <= not(layer0_outputs(9341));
    layer1_outputs(8308) <= not((layer0_outputs(9412)) xor (layer0_outputs(7148)));
    layer1_outputs(8309) <= not(layer0_outputs(808));
    layer1_outputs(8310) <= (layer0_outputs(5172)) and not (layer0_outputs(1249));
    layer1_outputs(8311) <= layer0_outputs(8993);
    layer1_outputs(8312) <= (layer0_outputs(1572)) or (layer0_outputs(10016));
    layer1_outputs(8313) <= not((layer0_outputs(3090)) or (layer0_outputs(5788)));
    layer1_outputs(8314) <= layer0_outputs(1690);
    layer1_outputs(8315) <= not(layer0_outputs(5356));
    layer1_outputs(8316) <= not(layer0_outputs(4770));
    layer1_outputs(8317) <= not(layer0_outputs(2872));
    layer1_outputs(8318) <= (layer0_outputs(8574)) or (layer0_outputs(8241));
    layer1_outputs(8319) <= not(layer0_outputs(3313)) or (layer0_outputs(1061));
    layer1_outputs(8320) <= not((layer0_outputs(5833)) or (layer0_outputs(4788)));
    layer1_outputs(8321) <= not(layer0_outputs(8645));
    layer1_outputs(8322) <= not(layer0_outputs(455));
    layer1_outputs(8323) <= (layer0_outputs(9299)) and not (layer0_outputs(2449));
    layer1_outputs(8324) <= (layer0_outputs(6540)) or (layer0_outputs(5202));
    layer1_outputs(8325) <= not((layer0_outputs(602)) and (layer0_outputs(1517)));
    layer1_outputs(8326) <= not((layer0_outputs(588)) and (layer0_outputs(1442)));
    layer1_outputs(8327) <= layer0_outputs(3128);
    layer1_outputs(8328) <= (layer0_outputs(8275)) and not (layer0_outputs(9179));
    layer1_outputs(8329) <= not(layer0_outputs(4058)) or (layer0_outputs(1397));
    layer1_outputs(8330) <= not((layer0_outputs(3093)) and (layer0_outputs(7328)));
    layer1_outputs(8331) <= layer0_outputs(5806);
    layer1_outputs(8332) <= (layer0_outputs(4254)) or (layer0_outputs(3294));
    layer1_outputs(8333) <= not(layer0_outputs(5578));
    layer1_outputs(8334) <= layer0_outputs(104);
    layer1_outputs(8335) <= (layer0_outputs(9115)) or (layer0_outputs(472));
    layer1_outputs(8336) <= '1';
    layer1_outputs(8337) <= (layer0_outputs(4067)) or (layer0_outputs(7574));
    layer1_outputs(8338) <= (layer0_outputs(5174)) xor (layer0_outputs(1492));
    layer1_outputs(8339) <= (layer0_outputs(6409)) and not (layer0_outputs(6689));
    layer1_outputs(8340) <= layer0_outputs(1388);
    layer1_outputs(8341) <= (layer0_outputs(7952)) and not (layer0_outputs(1622));
    layer1_outputs(8342) <= layer0_outputs(1789);
    layer1_outputs(8343) <= not(layer0_outputs(7576));
    layer1_outputs(8344) <= not(layer0_outputs(844));
    layer1_outputs(8345) <= not(layer0_outputs(3127));
    layer1_outputs(8346) <= not(layer0_outputs(2492));
    layer1_outputs(8347) <= not(layer0_outputs(8809));
    layer1_outputs(8348) <= not(layer0_outputs(5844)) or (layer0_outputs(8472));
    layer1_outputs(8349) <= not(layer0_outputs(6391));
    layer1_outputs(8350) <= not(layer0_outputs(5353)) or (layer0_outputs(3630));
    layer1_outputs(8351) <= (layer0_outputs(2890)) and (layer0_outputs(479));
    layer1_outputs(8352) <= (layer0_outputs(2267)) and not (layer0_outputs(2045));
    layer1_outputs(8353) <= '1';
    layer1_outputs(8354) <= not(layer0_outputs(2696));
    layer1_outputs(8355) <= not((layer0_outputs(2330)) and (layer0_outputs(7427)));
    layer1_outputs(8356) <= (layer0_outputs(1211)) and (layer0_outputs(6469));
    layer1_outputs(8357) <= (layer0_outputs(4139)) or (layer0_outputs(6402));
    layer1_outputs(8358) <= not(layer0_outputs(5698));
    layer1_outputs(8359) <= layer0_outputs(5105);
    layer1_outputs(8360) <= layer0_outputs(7903);
    layer1_outputs(8361) <= not(layer0_outputs(10069));
    layer1_outputs(8362) <= (layer0_outputs(3211)) and not (layer0_outputs(8522));
    layer1_outputs(8363) <= not(layer0_outputs(2742));
    layer1_outputs(8364) <= not(layer0_outputs(3872));
    layer1_outputs(8365) <= (layer0_outputs(5069)) and (layer0_outputs(9445));
    layer1_outputs(8366) <= not(layer0_outputs(10065)) or (layer0_outputs(1003));
    layer1_outputs(8367) <= not(layer0_outputs(5784));
    layer1_outputs(8368) <= not(layer0_outputs(9745));
    layer1_outputs(8369) <= not(layer0_outputs(4179));
    layer1_outputs(8370) <= (layer0_outputs(5679)) or (layer0_outputs(9102));
    layer1_outputs(8371) <= not((layer0_outputs(3020)) xor (layer0_outputs(4261)));
    layer1_outputs(8372) <= not(layer0_outputs(9913));
    layer1_outputs(8373) <= not(layer0_outputs(9968)) or (layer0_outputs(8432));
    layer1_outputs(8374) <= (layer0_outputs(2788)) and not (layer0_outputs(6745));
    layer1_outputs(8375) <= (layer0_outputs(9577)) and (layer0_outputs(695));
    layer1_outputs(8376) <= layer0_outputs(10188);
    layer1_outputs(8377) <= layer0_outputs(7971);
    layer1_outputs(8378) <= not((layer0_outputs(2737)) xor (layer0_outputs(10023)));
    layer1_outputs(8379) <= (layer0_outputs(3362)) and not (layer0_outputs(7828));
    layer1_outputs(8380) <= layer0_outputs(6529);
    layer1_outputs(8381) <= '1';
    layer1_outputs(8382) <= (layer0_outputs(5161)) and not (layer0_outputs(8161));
    layer1_outputs(8383) <= not(layer0_outputs(10064));
    layer1_outputs(8384) <= not((layer0_outputs(352)) and (layer0_outputs(3044)));
    layer1_outputs(8385) <= layer0_outputs(4170);
    layer1_outputs(8386) <= layer0_outputs(7522);
    layer1_outputs(8387) <= '1';
    layer1_outputs(8388) <= layer0_outputs(10174);
    layer1_outputs(8389) <= layer0_outputs(8458);
    layer1_outputs(8390) <= not(layer0_outputs(8733));
    layer1_outputs(8391) <= '0';
    layer1_outputs(8392) <= not((layer0_outputs(9711)) or (layer0_outputs(8070)));
    layer1_outputs(8393) <= not(layer0_outputs(7934));
    layer1_outputs(8394) <= (layer0_outputs(525)) xor (layer0_outputs(82));
    layer1_outputs(8395) <= not((layer0_outputs(8275)) xor (layer0_outputs(694)));
    layer1_outputs(8396) <= (layer0_outputs(2024)) or (layer0_outputs(3185));
    layer1_outputs(8397) <= not(layer0_outputs(1315)) or (layer0_outputs(2511));
    layer1_outputs(8398) <= not((layer0_outputs(2118)) or (layer0_outputs(4638)));
    layer1_outputs(8399) <= not(layer0_outputs(9748));
    layer1_outputs(8400) <= not((layer0_outputs(9882)) and (layer0_outputs(1577)));
    layer1_outputs(8401) <= not(layer0_outputs(663));
    layer1_outputs(8402) <= layer0_outputs(3954);
    layer1_outputs(8403) <= not(layer0_outputs(5176)) or (layer0_outputs(4234));
    layer1_outputs(8404) <= not((layer0_outputs(7571)) or (layer0_outputs(4434)));
    layer1_outputs(8405) <= layer0_outputs(2212);
    layer1_outputs(8406) <= (layer0_outputs(4685)) and not (layer0_outputs(8146));
    layer1_outputs(8407) <= not((layer0_outputs(190)) xor (layer0_outputs(9902)));
    layer1_outputs(8408) <= not(layer0_outputs(8901));
    layer1_outputs(8409) <= (layer0_outputs(4691)) or (layer0_outputs(10010));
    layer1_outputs(8410) <= (layer0_outputs(4914)) or (layer0_outputs(6434));
    layer1_outputs(8411) <= (layer0_outputs(4790)) and (layer0_outputs(6789));
    layer1_outputs(8412) <= (layer0_outputs(712)) or (layer0_outputs(7169));
    layer1_outputs(8413) <= not(layer0_outputs(9806));
    layer1_outputs(8414) <= (layer0_outputs(8385)) and not (layer0_outputs(6982));
    layer1_outputs(8415) <= not(layer0_outputs(6847));
    layer1_outputs(8416) <= layer0_outputs(2084);
    layer1_outputs(8417) <= (layer0_outputs(23)) or (layer0_outputs(5648));
    layer1_outputs(8418) <= (layer0_outputs(53)) and not (layer0_outputs(3101));
    layer1_outputs(8419) <= not(layer0_outputs(5945)) or (layer0_outputs(8633));
    layer1_outputs(8420) <= '1';
    layer1_outputs(8421) <= (layer0_outputs(7824)) xor (layer0_outputs(5042));
    layer1_outputs(8422) <= not((layer0_outputs(4927)) or (layer0_outputs(1999)));
    layer1_outputs(8423) <= not(layer0_outputs(5036));
    layer1_outputs(8424) <= (layer0_outputs(4922)) and not (layer0_outputs(1542));
    layer1_outputs(8425) <= layer0_outputs(9135);
    layer1_outputs(8426) <= not((layer0_outputs(1173)) xor (layer0_outputs(5536)));
    layer1_outputs(8427) <= not(layer0_outputs(1317));
    layer1_outputs(8428) <= (layer0_outputs(2049)) and not (layer0_outputs(2624));
    layer1_outputs(8429) <= layer0_outputs(8578);
    layer1_outputs(8430) <= not(layer0_outputs(4312));
    layer1_outputs(8431) <= (layer0_outputs(331)) xor (layer0_outputs(1894));
    layer1_outputs(8432) <= layer0_outputs(6127);
    layer1_outputs(8433) <= not((layer0_outputs(5918)) xor (layer0_outputs(5412)));
    layer1_outputs(8434) <= not((layer0_outputs(2538)) or (layer0_outputs(3366)));
    layer1_outputs(8435) <= (layer0_outputs(5000)) or (layer0_outputs(8752));
    layer1_outputs(8436) <= not(layer0_outputs(7803));
    layer1_outputs(8437) <= (layer0_outputs(9213)) or (layer0_outputs(1439));
    layer1_outputs(8438) <= (layer0_outputs(1863)) or (layer0_outputs(5283));
    layer1_outputs(8439) <= not((layer0_outputs(9296)) and (layer0_outputs(6553)));
    layer1_outputs(8440) <= layer0_outputs(6305);
    layer1_outputs(8441) <= '1';
    layer1_outputs(8442) <= not(layer0_outputs(3110));
    layer1_outputs(8443) <= not(layer0_outputs(2516));
    layer1_outputs(8444) <= (layer0_outputs(8801)) or (layer0_outputs(837));
    layer1_outputs(8445) <= not(layer0_outputs(8139));
    layer1_outputs(8446) <= not(layer0_outputs(7470));
    layer1_outputs(8447) <= not(layer0_outputs(6355)) or (layer0_outputs(8142));
    layer1_outputs(8448) <= not(layer0_outputs(1459));
    layer1_outputs(8449) <= not(layer0_outputs(6143));
    layer1_outputs(8450) <= not(layer0_outputs(3977)) or (layer0_outputs(6848));
    layer1_outputs(8451) <= not(layer0_outputs(1019));
    layer1_outputs(8452) <= layer0_outputs(2036);
    layer1_outputs(8453) <= (layer0_outputs(3152)) or (layer0_outputs(1943));
    layer1_outputs(8454) <= layer0_outputs(8109);
    layer1_outputs(8455) <= not(layer0_outputs(8705)) or (layer0_outputs(2891));
    layer1_outputs(8456) <= not(layer0_outputs(2518)) or (layer0_outputs(5312));
    layer1_outputs(8457) <= not(layer0_outputs(7211)) or (layer0_outputs(6343));
    layer1_outputs(8458) <= not((layer0_outputs(2900)) xor (layer0_outputs(7015)));
    layer1_outputs(8459) <= not((layer0_outputs(3640)) and (layer0_outputs(9729)));
    layer1_outputs(8460) <= (layer0_outputs(5386)) and not (layer0_outputs(24));
    layer1_outputs(8461) <= not((layer0_outputs(2759)) xor (layer0_outputs(8510)));
    layer1_outputs(8462) <= not((layer0_outputs(40)) and (layer0_outputs(6106)));
    layer1_outputs(8463) <= layer0_outputs(704);
    layer1_outputs(8464) <= not(layer0_outputs(2091));
    layer1_outputs(8465) <= layer0_outputs(8697);
    layer1_outputs(8466) <= layer0_outputs(6456);
    layer1_outputs(8467) <= not(layer0_outputs(9091));
    layer1_outputs(8468) <= '1';
    layer1_outputs(8469) <= (layer0_outputs(9680)) or (layer0_outputs(3840));
    layer1_outputs(8470) <= layer0_outputs(3972);
    layer1_outputs(8471) <= layer0_outputs(4978);
    layer1_outputs(8472) <= not(layer0_outputs(1272));
    layer1_outputs(8473) <= not(layer0_outputs(6787));
    layer1_outputs(8474) <= layer0_outputs(1474);
    layer1_outputs(8475) <= (layer0_outputs(3574)) xor (layer0_outputs(9062));
    layer1_outputs(8476) <= not(layer0_outputs(2855)) or (layer0_outputs(654));
    layer1_outputs(8477) <= layer0_outputs(624);
    layer1_outputs(8478) <= (layer0_outputs(1822)) and not (layer0_outputs(1733));
    layer1_outputs(8479) <= not(layer0_outputs(1954));
    layer1_outputs(8480) <= layer0_outputs(3482);
    layer1_outputs(8481) <= layer0_outputs(9502);
    layer1_outputs(8482) <= (layer0_outputs(5031)) and not (layer0_outputs(1528));
    layer1_outputs(8483) <= not(layer0_outputs(941));
    layer1_outputs(8484) <= not((layer0_outputs(9462)) and (layer0_outputs(3128)));
    layer1_outputs(8485) <= (layer0_outputs(5365)) xor (layer0_outputs(244));
    layer1_outputs(8486) <= (layer0_outputs(2280)) or (layer0_outputs(5956));
    layer1_outputs(8487) <= (layer0_outputs(6181)) and not (layer0_outputs(5929));
    layer1_outputs(8488) <= layer0_outputs(8778);
    layer1_outputs(8489) <= not(layer0_outputs(8276)) or (layer0_outputs(8439));
    layer1_outputs(8490) <= not(layer0_outputs(9580)) or (layer0_outputs(2346));
    layer1_outputs(8491) <= (layer0_outputs(6681)) or (layer0_outputs(2162));
    layer1_outputs(8492) <= not((layer0_outputs(7668)) or (layer0_outputs(2347)));
    layer1_outputs(8493) <= layer0_outputs(5642);
    layer1_outputs(8494) <= not(layer0_outputs(6877)) or (layer0_outputs(6940));
    layer1_outputs(8495) <= '1';
    layer1_outputs(8496) <= not(layer0_outputs(2857));
    layer1_outputs(8497) <= layer0_outputs(7205);
    layer1_outputs(8498) <= not((layer0_outputs(501)) or (layer0_outputs(5270)));
    layer1_outputs(8499) <= not((layer0_outputs(622)) and (layer0_outputs(4700)));
    layer1_outputs(8500) <= '1';
    layer1_outputs(8501) <= not((layer0_outputs(8403)) xor (layer0_outputs(1000)));
    layer1_outputs(8502) <= not((layer0_outputs(9195)) xor (layer0_outputs(3179)));
    layer1_outputs(8503) <= not(layer0_outputs(8606)) or (layer0_outputs(8440));
    layer1_outputs(8504) <= (layer0_outputs(8389)) and not (layer0_outputs(304));
    layer1_outputs(8505) <= not(layer0_outputs(4178));
    layer1_outputs(8506) <= not(layer0_outputs(7812));
    layer1_outputs(8507) <= (layer0_outputs(245)) and not (layer0_outputs(3652));
    layer1_outputs(8508) <= layer0_outputs(2053);
    layer1_outputs(8509) <= not((layer0_outputs(5255)) and (layer0_outputs(7703)));
    layer1_outputs(8510) <= not(layer0_outputs(6325)) or (layer0_outputs(2938));
    layer1_outputs(8511) <= not(layer0_outputs(7139));
    layer1_outputs(8512) <= (layer0_outputs(4582)) and not (layer0_outputs(9416));
    layer1_outputs(8513) <= layer0_outputs(7807);
    layer1_outputs(8514) <= not((layer0_outputs(3259)) and (layer0_outputs(2731)));
    layer1_outputs(8515) <= (layer0_outputs(673)) and not (layer0_outputs(1743));
    layer1_outputs(8516) <= not((layer0_outputs(3440)) xor (layer0_outputs(5845)));
    layer1_outputs(8517) <= layer0_outputs(3102);
    layer1_outputs(8518) <= layer0_outputs(4602);
    layer1_outputs(8519) <= not((layer0_outputs(7483)) and (layer0_outputs(9076)));
    layer1_outputs(8520) <= (layer0_outputs(2038)) and not (layer0_outputs(3088));
    layer1_outputs(8521) <= (layer0_outputs(3144)) and not (layer0_outputs(6937));
    layer1_outputs(8522) <= not(layer0_outputs(6545));
    layer1_outputs(8523) <= not(layer0_outputs(6670));
    layer1_outputs(8524) <= not(layer0_outputs(7986));
    layer1_outputs(8525) <= not(layer0_outputs(1014));
    layer1_outputs(8526) <= not((layer0_outputs(950)) xor (layer0_outputs(5864)));
    layer1_outputs(8527) <= not(layer0_outputs(4025));
    layer1_outputs(8528) <= layer0_outputs(2202);
    layer1_outputs(8529) <= not(layer0_outputs(7080)) or (layer0_outputs(464));
    layer1_outputs(8530) <= (layer0_outputs(968)) or (layer0_outputs(5733));
    layer1_outputs(8531) <= (layer0_outputs(6559)) and not (layer0_outputs(3669));
    layer1_outputs(8532) <= layer0_outputs(7564);
    layer1_outputs(8533) <= layer0_outputs(8110);
    layer1_outputs(8534) <= not(layer0_outputs(7836));
    layer1_outputs(8535) <= not(layer0_outputs(2199));
    layer1_outputs(8536) <= layer0_outputs(9747);
    layer1_outputs(8537) <= not((layer0_outputs(5787)) and (layer0_outputs(3460)));
    layer1_outputs(8538) <= (layer0_outputs(9304)) and not (layer0_outputs(9993));
    layer1_outputs(8539) <= not((layer0_outputs(4158)) xor (layer0_outputs(9686)));
    layer1_outputs(8540) <= '1';
    layer1_outputs(8541) <= not(layer0_outputs(182));
    layer1_outputs(8542) <= not(layer0_outputs(9461)) or (layer0_outputs(3228));
    layer1_outputs(8543) <= not(layer0_outputs(7657));
    layer1_outputs(8544) <= not((layer0_outputs(10161)) xor (layer0_outputs(2062)));
    layer1_outputs(8545) <= not(layer0_outputs(7654)) or (layer0_outputs(8751));
    layer1_outputs(8546) <= (layer0_outputs(2406)) or (layer0_outputs(5378));
    layer1_outputs(8547) <= (layer0_outputs(2484)) and not (layer0_outputs(1126));
    layer1_outputs(8548) <= not(layer0_outputs(4197));
    layer1_outputs(8549) <= '1';
    layer1_outputs(8550) <= not(layer0_outputs(4702));
    layer1_outputs(8551) <= not(layer0_outputs(7582));
    layer1_outputs(8552) <= not((layer0_outputs(5720)) xor (layer0_outputs(9098)));
    layer1_outputs(8553) <= (layer0_outputs(5171)) and not (layer0_outputs(5942));
    layer1_outputs(8554) <= not(layer0_outputs(9251));
    layer1_outputs(8555) <= not(layer0_outputs(3956)) or (layer0_outputs(10143));
    layer1_outputs(8556) <= (layer0_outputs(7895)) and not (layer0_outputs(8768));
    layer1_outputs(8557) <= (layer0_outputs(6375)) and (layer0_outputs(1034));
    layer1_outputs(8558) <= not(layer0_outputs(2517));
    layer1_outputs(8559) <= '0';
    layer1_outputs(8560) <= not(layer0_outputs(5838));
    layer1_outputs(8561) <= (layer0_outputs(4693)) and not (layer0_outputs(8453));
    layer1_outputs(8562) <= not(layer0_outputs(178)) or (layer0_outputs(5074));
    layer1_outputs(8563) <= '0';
    layer1_outputs(8564) <= not(layer0_outputs(1469));
    layer1_outputs(8565) <= (layer0_outputs(3983)) or (layer0_outputs(1148));
    layer1_outputs(8566) <= layer0_outputs(5142);
    layer1_outputs(8567) <= not(layer0_outputs(4111));
    layer1_outputs(8568) <= not(layer0_outputs(3279)) or (layer0_outputs(8940));
    layer1_outputs(8569) <= layer0_outputs(7474);
    layer1_outputs(8570) <= (layer0_outputs(8914)) and not (layer0_outputs(2609));
    layer1_outputs(8571) <= layer0_outputs(4462);
    layer1_outputs(8572) <= not((layer0_outputs(4705)) or (layer0_outputs(3415)));
    layer1_outputs(8573) <= not(layer0_outputs(7095));
    layer1_outputs(8574) <= not(layer0_outputs(8542));
    layer1_outputs(8575) <= not(layer0_outputs(7269)) or (layer0_outputs(3657));
    layer1_outputs(8576) <= not((layer0_outputs(2250)) and (layer0_outputs(2484)));
    layer1_outputs(8577) <= not(layer0_outputs(4084));
    layer1_outputs(8578) <= layer0_outputs(4027);
    layer1_outputs(8579) <= not((layer0_outputs(5900)) and (layer0_outputs(10227)));
    layer1_outputs(8580) <= (layer0_outputs(229)) or (layer0_outputs(8780));
    layer1_outputs(8581) <= (layer0_outputs(6875)) or (layer0_outputs(6733));
    layer1_outputs(8582) <= (layer0_outputs(4568)) and (layer0_outputs(5738));
    layer1_outputs(8583) <= not(layer0_outputs(6171)) or (layer0_outputs(6217));
    layer1_outputs(8584) <= not(layer0_outputs(1853));
    layer1_outputs(8585) <= (layer0_outputs(8389)) and not (layer0_outputs(2558));
    layer1_outputs(8586) <= not(layer0_outputs(6354)) or (layer0_outputs(6884));
    layer1_outputs(8587) <= not((layer0_outputs(1140)) and (layer0_outputs(6785)));
    layer1_outputs(8588) <= (layer0_outputs(1567)) and (layer0_outputs(7118));
    layer1_outputs(8589) <= not(layer0_outputs(2296));
    layer1_outputs(8590) <= (layer0_outputs(1268)) and not (layer0_outputs(8454));
    layer1_outputs(8591) <= (layer0_outputs(6302)) and not (layer0_outputs(1369));
    layer1_outputs(8592) <= (layer0_outputs(935)) or (layer0_outputs(526));
    layer1_outputs(8593) <= layer0_outputs(8314);
    layer1_outputs(8594) <= '1';
    layer1_outputs(8595) <= (layer0_outputs(2826)) and (layer0_outputs(8905));
    layer1_outputs(8596) <= (layer0_outputs(4531)) and not (layer0_outputs(5060));
    layer1_outputs(8597) <= layer0_outputs(7624);
    layer1_outputs(8598) <= not(layer0_outputs(4879));
    layer1_outputs(8599) <= (layer0_outputs(266)) and not (layer0_outputs(7472));
    layer1_outputs(8600) <= not(layer0_outputs(1452));
    layer1_outputs(8601) <= not(layer0_outputs(7093));
    layer1_outputs(8602) <= not((layer0_outputs(3749)) and (layer0_outputs(8209)));
    layer1_outputs(8603) <= layer0_outputs(10019);
    layer1_outputs(8604) <= not(layer0_outputs(7952)) or (layer0_outputs(998));
    layer1_outputs(8605) <= '0';
    layer1_outputs(8606) <= (layer0_outputs(7514)) and (layer0_outputs(9570));
    layer1_outputs(8607) <= (layer0_outputs(4031)) xor (layer0_outputs(4065));
    layer1_outputs(8608) <= not(layer0_outputs(5870));
    layer1_outputs(8609) <= (layer0_outputs(3692)) and (layer0_outputs(5724));
    layer1_outputs(8610) <= layer0_outputs(4510);
    layer1_outputs(8611) <= not(layer0_outputs(9800)) or (layer0_outputs(9290));
    layer1_outputs(8612) <= (layer0_outputs(7295)) and not (layer0_outputs(377));
    layer1_outputs(8613) <= layer0_outputs(10015);
    layer1_outputs(8614) <= not(layer0_outputs(4470));
    layer1_outputs(8615) <= not((layer0_outputs(4229)) and (layer0_outputs(2015)));
    layer1_outputs(8616) <= not(layer0_outputs(3723));
    layer1_outputs(8617) <= (layer0_outputs(1981)) and not (layer0_outputs(5132));
    layer1_outputs(8618) <= not(layer0_outputs(2100));
    layer1_outputs(8619) <= not(layer0_outputs(6481)) or (layer0_outputs(8665));
    layer1_outputs(8620) <= layer0_outputs(8585);
    layer1_outputs(8621) <= not((layer0_outputs(7237)) or (layer0_outputs(1679)));
    layer1_outputs(8622) <= not(layer0_outputs(4199));
    layer1_outputs(8623) <= not((layer0_outputs(8239)) or (layer0_outputs(285)));
    layer1_outputs(8624) <= not(layer0_outputs(7203));
    layer1_outputs(8625) <= layer0_outputs(9866);
    layer1_outputs(8626) <= '1';
    layer1_outputs(8627) <= not((layer0_outputs(1941)) and (layer0_outputs(9517)));
    layer1_outputs(8628) <= not(layer0_outputs(6849));
    layer1_outputs(8629) <= layer0_outputs(2423);
    layer1_outputs(8630) <= not(layer0_outputs(2451));
    layer1_outputs(8631) <= not((layer0_outputs(9104)) xor (layer0_outputs(7147)));
    layer1_outputs(8632) <= not((layer0_outputs(3762)) and (layer0_outputs(4622)));
    layer1_outputs(8633) <= not(layer0_outputs(10209));
    layer1_outputs(8634) <= not(layer0_outputs(5095));
    layer1_outputs(8635) <= layer0_outputs(6390);
    layer1_outputs(8636) <= not(layer0_outputs(7222));
    layer1_outputs(8637) <= not(layer0_outputs(9805));
    layer1_outputs(8638) <= not(layer0_outputs(1333)) or (layer0_outputs(4108));
    layer1_outputs(8639) <= not(layer0_outputs(5500)) or (layer0_outputs(844));
    layer1_outputs(8640) <= not(layer0_outputs(5248));
    layer1_outputs(8641) <= layer0_outputs(9243);
    layer1_outputs(8642) <= '0';
    layer1_outputs(8643) <= not(layer0_outputs(3805)) or (layer0_outputs(4636));
    layer1_outputs(8644) <= (layer0_outputs(4447)) and (layer0_outputs(5652));
    layer1_outputs(8645) <= layer0_outputs(9051);
    layer1_outputs(8646) <= (layer0_outputs(1627)) and (layer0_outputs(2367));
    layer1_outputs(8647) <= (layer0_outputs(6016)) or (layer0_outputs(6317));
    layer1_outputs(8648) <= not((layer0_outputs(8029)) or (layer0_outputs(3475)));
    layer1_outputs(8649) <= (layer0_outputs(6087)) and not (layer0_outputs(888));
    layer1_outputs(8650) <= (layer0_outputs(5990)) xor (layer0_outputs(6587));
    layer1_outputs(8651) <= not(layer0_outputs(5536));
    layer1_outputs(8652) <= (layer0_outputs(2275)) or (layer0_outputs(8834));
    layer1_outputs(8653) <= not(layer0_outputs(9539));
    layer1_outputs(8654) <= (layer0_outputs(10219)) and not (layer0_outputs(10222));
    layer1_outputs(8655) <= (layer0_outputs(4022)) and not (layer0_outputs(9449));
    layer1_outputs(8656) <= layer0_outputs(8116);
    layer1_outputs(8657) <= (layer0_outputs(9143)) and not (layer0_outputs(9535));
    layer1_outputs(8658) <= not(layer0_outputs(1044));
    layer1_outputs(8659) <= (layer0_outputs(5651)) and not (layer0_outputs(2579));
    layer1_outputs(8660) <= not(layer0_outputs(243)) or (layer0_outputs(7113));
    layer1_outputs(8661) <= (layer0_outputs(6404)) and not (layer0_outputs(7968));
    layer1_outputs(8662) <= (layer0_outputs(9501)) and (layer0_outputs(2085));
    layer1_outputs(8663) <= not((layer0_outputs(5331)) and (layer0_outputs(9410)));
    layer1_outputs(8664) <= (layer0_outputs(9524)) and not (layer0_outputs(495));
    layer1_outputs(8665) <= layer0_outputs(4704);
    layer1_outputs(8666) <= not((layer0_outputs(556)) or (layer0_outputs(2582)));
    layer1_outputs(8667) <= not(layer0_outputs(2552));
    layer1_outputs(8668) <= layer0_outputs(1931);
    layer1_outputs(8669) <= '1';
    layer1_outputs(8670) <= layer0_outputs(154);
    layer1_outputs(8671) <= not(layer0_outputs(9071)) or (layer0_outputs(6706));
    layer1_outputs(8672) <= (layer0_outputs(5079)) or (layer0_outputs(1257));
    layer1_outputs(8673) <= layer0_outputs(4613);
    layer1_outputs(8674) <= not((layer0_outputs(1586)) and (layer0_outputs(7547)));
    layer1_outputs(8675) <= layer0_outputs(2745);
    layer1_outputs(8676) <= layer0_outputs(2630);
    layer1_outputs(8677) <= (layer0_outputs(9488)) and not (layer0_outputs(6336));
    layer1_outputs(8678) <= (layer0_outputs(6566)) xor (layer0_outputs(4829));
    layer1_outputs(8679) <= (layer0_outputs(2205)) xor (layer0_outputs(1100));
    layer1_outputs(8680) <= not(layer0_outputs(4490));
    layer1_outputs(8681) <= not(layer0_outputs(4023));
    layer1_outputs(8682) <= layer0_outputs(1234);
    layer1_outputs(8683) <= not((layer0_outputs(4223)) xor (layer0_outputs(10166)));
    layer1_outputs(8684) <= (layer0_outputs(4894)) and (layer0_outputs(1718));
    layer1_outputs(8685) <= not(layer0_outputs(575));
    layer1_outputs(8686) <= not((layer0_outputs(385)) or (layer0_outputs(5003)));
    layer1_outputs(8687) <= (layer0_outputs(7490)) and not (layer0_outputs(6746));
    layer1_outputs(8688) <= (layer0_outputs(10069)) and not (layer0_outputs(4903));
    layer1_outputs(8689) <= not((layer0_outputs(7994)) xor (layer0_outputs(2184)));
    layer1_outputs(8690) <= (layer0_outputs(6710)) and not (layer0_outputs(9367));
    layer1_outputs(8691) <= (layer0_outputs(7422)) and not (layer0_outputs(1047));
    layer1_outputs(8692) <= (layer0_outputs(4404)) or (layer0_outputs(594));
    layer1_outputs(8693) <= not(layer0_outputs(2153));
    layer1_outputs(8694) <= (layer0_outputs(2521)) or (layer0_outputs(1956));
    layer1_outputs(8695) <= not(layer0_outputs(4693));
    layer1_outputs(8696) <= layer0_outputs(8818);
    layer1_outputs(8697) <= not(layer0_outputs(6078));
    layer1_outputs(8698) <= '0';
    layer1_outputs(8699) <= layer0_outputs(4282);
    layer1_outputs(8700) <= not((layer0_outputs(3318)) xor (layer0_outputs(5580)));
    layer1_outputs(8701) <= not(layer0_outputs(2774));
    layer1_outputs(8702) <= not((layer0_outputs(4402)) and (layer0_outputs(6818)));
    layer1_outputs(8703) <= not(layer0_outputs(6978)) or (layer0_outputs(5443));
    layer1_outputs(8704) <= not(layer0_outputs(8831));
    layer1_outputs(8705) <= not(layer0_outputs(8031));
    layer1_outputs(8706) <= not(layer0_outputs(7488));
    layer1_outputs(8707) <= (layer0_outputs(3066)) and (layer0_outputs(1739));
    layer1_outputs(8708) <= layer0_outputs(4231);
    layer1_outputs(8709) <= (layer0_outputs(4163)) and (layer0_outputs(968));
    layer1_outputs(8710) <= not(layer0_outputs(3698));
    layer1_outputs(8711) <= '0';
    layer1_outputs(8712) <= (layer0_outputs(8922)) and not (layer0_outputs(4950));
    layer1_outputs(8713) <= layer0_outputs(4638);
    layer1_outputs(8714) <= layer0_outputs(1031);
    layer1_outputs(8715) <= not(layer0_outputs(2195));
    layer1_outputs(8716) <= not(layer0_outputs(2725)) or (layer0_outputs(8213));
    layer1_outputs(8717) <= layer0_outputs(581);
    layer1_outputs(8718) <= not((layer0_outputs(8988)) or (layer0_outputs(7533)));
    layer1_outputs(8719) <= (layer0_outputs(1031)) and not (layer0_outputs(3837));
    layer1_outputs(8720) <= layer0_outputs(2717);
    layer1_outputs(8721) <= not(layer0_outputs(5696));
    layer1_outputs(8722) <= not(layer0_outputs(6347));
    layer1_outputs(8723) <= (layer0_outputs(5985)) and (layer0_outputs(1784));
    layer1_outputs(8724) <= not(layer0_outputs(3905));
    layer1_outputs(8725) <= not(layer0_outputs(7966));
    layer1_outputs(8726) <= '1';
    layer1_outputs(8727) <= not(layer0_outputs(7435));
    layer1_outputs(8728) <= (layer0_outputs(3005)) or (layer0_outputs(1056));
    layer1_outputs(8729) <= not(layer0_outputs(5314));
    layer1_outputs(8730) <= not(layer0_outputs(9639));
    layer1_outputs(8731) <= not(layer0_outputs(9336));
    layer1_outputs(8732) <= not((layer0_outputs(8465)) or (layer0_outputs(3391)));
    layer1_outputs(8733) <= (layer0_outputs(1723)) and not (layer0_outputs(6935));
    layer1_outputs(8734) <= not(layer0_outputs(4545));
    layer1_outputs(8735) <= not(layer0_outputs(1365));
    layer1_outputs(8736) <= not(layer0_outputs(9953));
    layer1_outputs(8737) <= not(layer0_outputs(2726));
    layer1_outputs(8738) <= not((layer0_outputs(7257)) and (layer0_outputs(9089)));
    layer1_outputs(8739) <= layer0_outputs(5181);
    layer1_outputs(8740) <= (layer0_outputs(4912)) or (layer0_outputs(7216));
    layer1_outputs(8741) <= not(layer0_outputs(887)) or (layer0_outputs(661));
    layer1_outputs(8742) <= (layer0_outputs(5459)) and not (layer0_outputs(1481));
    layer1_outputs(8743) <= not((layer0_outputs(4314)) or (layer0_outputs(6938)));
    layer1_outputs(8744) <= not(layer0_outputs(1261));
    layer1_outputs(8745) <= not((layer0_outputs(3057)) and (layer0_outputs(3717)));
    layer1_outputs(8746) <= (layer0_outputs(1938)) xor (layer0_outputs(3575));
    layer1_outputs(8747) <= not(layer0_outputs(7390));
    layer1_outputs(8748) <= layer0_outputs(5673);
    layer1_outputs(8749) <= not(layer0_outputs(6574));
    layer1_outputs(8750) <= layer0_outputs(2393);
    layer1_outputs(8751) <= (layer0_outputs(8500)) and not (layer0_outputs(2489));
    layer1_outputs(8752) <= not(layer0_outputs(7239)) or (layer0_outputs(2943));
    layer1_outputs(8753) <= not((layer0_outputs(8331)) or (layer0_outputs(4396)));
    layer1_outputs(8754) <= (layer0_outputs(4166)) and not (layer0_outputs(2678));
    layer1_outputs(8755) <= layer0_outputs(5092);
    layer1_outputs(8756) <= layer0_outputs(3709);
    layer1_outputs(8757) <= not((layer0_outputs(1208)) xor (layer0_outputs(8010)));
    layer1_outputs(8758) <= not(layer0_outputs(1532));
    layer1_outputs(8759) <= not((layer0_outputs(7568)) xor (layer0_outputs(4185)));
    layer1_outputs(8760) <= not((layer0_outputs(3536)) or (layer0_outputs(780)));
    layer1_outputs(8761) <= not(layer0_outputs(1981)) or (layer0_outputs(2593));
    layer1_outputs(8762) <= not(layer0_outputs(1978));
    layer1_outputs(8763) <= not(layer0_outputs(9663));
    layer1_outputs(8764) <= (layer0_outputs(822)) and not (layer0_outputs(1513));
    layer1_outputs(8765) <= layer0_outputs(2875);
    layer1_outputs(8766) <= not((layer0_outputs(871)) or (layer0_outputs(5024)));
    layer1_outputs(8767) <= layer0_outputs(6173);
    layer1_outputs(8768) <= not(layer0_outputs(6573)) or (layer0_outputs(2971));
    layer1_outputs(8769) <= not((layer0_outputs(5667)) xor (layer0_outputs(6065)));
    layer1_outputs(8770) <= (layer0_outputs(4414)) xor (layer0_outputs(9031));
    layer1_outputs(8771) <= layer0_outputs(3611);
    layer1_outputs(8772) <= not((layer0_outputs(1828)) xor (layer0_outputs(8235)));
    layer1_outputs(8773) <= not(layer0_outputs(8327)) or (layer0_outputs(9647));
    layer1_outputs(8774) <= '1';
    layer1_outputs(8775) <= not(layer0_outputs(4729));
    layer1_outputs(8776) <= not(layer0_outputs(7890));
    layer1_outputs(8777) <= not(layer0_outputs(2518));
    layer1_outputs(8778) <= (layer0_outputs(8080)) and not (layer0_outputs(8631));
    layer1_outputs(8779) <= layer0_outputs(886);
    layer1_outputs(8780) <= layer0_outputs(5604);
    layer1_outputs(8781) <= not(layer0_outputs(3277)) or (layer0_outputs(9577));
    layer1_outputs(8782) <= not((layer0_outputs(2566)) xor (layer0_outputs(2681)));
    layer1_outputs(8783) <= (layer0_outputs(8368)) or (layer0_outputs(3064));
    layer1_outputs(8784) <= not((layer0_outputs(10143)) and (layer0_outputs(5859)));
    layer1_outputs(8785) <= not(layer0_outputs(3617));
    layer1_outputs(8786) <= layer0_outputs(4664);
    layer1_outputs(8787) <= not(layer0_outputs(7145));
    layer1_outputs(8788) <= not((layer0_outputs(2435)) and (layer0_outputs(556)));
    layer1_outputs(8789) <= not((layer0_outputs(2219)) or (layer0_outputs(7254)));
    layer1_outputs(8790) <= (layer0_outputs(7439)) xor (layer0_outputs(5598));
    layer1_outputs(8791) <= not((layer0_outputs(8318)) and (layer0_outputs(6883)));
    layer1_outputs(8792) <= not(layer0_outputs(799));
    layer1_outputs(8793) <= '0';
    layer1_outputs(8794) <= (layer0_outputs(4710)) and not (layer0_outputs(9957));
    layer1_outputs(8795) <= not((layer0_outputs(5768)) or (layer0_outputs(6410)));
    layer1_outputs(8796) <= layer0_outputs(7545);
    layer1_outputs(8797) <= layer0_outputs(4225);
    layer1_outputs(8798) <= not(layer0_outputs(8971));
    layer1_outputs(8799) <= not(layer0_outputs(8717));
    layer1_outputs(8800) <= not((layer0_outputs(159)) and (layer0_outputs(3376)));
    layer1_outputs(8801) <= not((layer0_outputs(9284)) xor (layer0_outputs(7485)));
    layer1_outputs(8802) <= not((layer0_outputs(3079)) and (layer0_outputs(4814)));
    layer1_outputs(8803) <= (layer0_outputs(5775)) or (layer0_outputs(6163));
    layer1_outputs(8804) <= not(layer0_outputs(369)) or (layer0_outputs(3875));
    layer1_outputs(8805) <= (layer0_outputs(1096)) and (layer0_outputs(8604));
    layer1_outputs(8806) <= not(layer0_outputs(1260));
    layer1_outputs(8807) <= not((layer0_outputs(8366)) xor (layer0_outputs(9428)));
    layer1_outputs(8808) <= not(layer0_outputs(6238)) or (layer0_outputs(6517));
    layer1_outputs(8809) <= layer0_outputs(3979);
    layer1_outputs(8810) <= layer0_outputs(5423);
    layer1_outputs(8811) <= layer0_outputs(3920);
    layer1_outputs(8812) <= not(layer0_outputs(7265));
    layer1_outputs(8813) <= (layer0_outputs(9704)) and (layer0_outputs(1737));
    layer1_outputs(8814) <= layer0_outputs(8450);
    layer1_outputs(8815) <= layer0_outputs(1569);
    layer1_outputs(8816) <= (layer0_outputs(5503)) and not (layer0_outputs(9086));
    layer1_outputs(8817) <= (layer0_outputs(4198)) and not (layer0_outputs(9369));
    layer1_outputs(8818) <= not((layer0_outputs(451)) and (layer0_outputs(5624)));
    layer1_outputs(8819) <= layer0_outputs(5264);
    layer1_outputs(8820) <= layer0_outputs(2691);
    layer1_outputs(8821) <= layer0_outputs(6682);
    layer1_outputs(8822) <= (layer0_outputs(9561)) and (layer0_outputs(5544));
    layer1_outputs(8823) <= not(layer0_outputs(6371)) or (layer0_outputs(7548));
    layer1_outputs(8824) <= not(layer0_outputs(6765));
    layer1_outputs(8825) <= layer0_outputs(7552);
    layer1_outputs(8826) <= (layer0_outputs(3379)) xor (layer0_outputs(9021));
    layer1_outputs(8827) <= (layer0_outputs(345)) or (layer0_outputs(3019));
    layer1_outputs(8828) <= (layer0_outputs(3163)) and not (layer0_outputs(481));
    layer1_outputs(8829) <= not(layer0_outputs(650)) or (layer0_outputs(5271));
    layer1_outputs(8830) <= (layer0_outputs(173)) and not (layer0_outputs(6889));
    layer1_outputs(8831) <= layer0_outputs(5223);
    layer1_outputs(8832) <= (layer0_outputs(4769)) or (layer0_outputs(1438));
    layer1_outputs(8833) <= layer0_outputs(4841);
    layer1_outputs(8834) <= not((layer0_outputs(5639)) or (layer0_outputs(9118)));
    layer1_outputs(8835) <= not((layer0_outputs(4103)) or (layer0_outputs(7827)));
    layer1_outputs(8836) <= not(layer0_outputs(8122));
    layer1_outputs(8837) <= not((layer0_outputs(9950)) xor (layer0_outputs(1765)));
    layer1_outputs(8838) <= not((layer0_outputs(7258)) and (layer0_outputs(2417)));
    layer1_outputs(8839) <= (layer0_outputs(4843)) or (layer0_outputs(2097));
    layer1_outputs(8840) <= not(layer0_outputs(1894));
    layer1_outputs(8841) <= layer0_outputs(3647);
    layer1_outputs(8842) <= not((layer0_outputs(6422)) and (layer0_outputs(1051)));
    layer1_outputs(8843) <= not((layer0_outputs(4793)) and (layer0_outputs(1842)));
    layer1_outputs(8844) <= (layer0_outputs(5516)) and not (layer0_outputs(7979));
    layer1_outputs(8845) <= not(layer0_outputs(9139));
    layer1_outputs(8846) <= not(layer0_outputs(7129));
    layer1_outputs(8847) <= (layer0_outputs(1446)) and not (layer0_outputs(5891));
    layer1_outputs(8848) <= not((layer0_outputs(5745)) and (layer0_outputs(4040)));
    layer1_outputs(8849) <= (layer0_outputs(403)) and not (layer0_outputs(5346));
    layer1_outputs(8850) <= not(layer0_outputs(4010)) or (layer0_outputs(10061));
    layer1_outputs(8851) <= layer0_outputs(308);
    layer1_outputs(8852) <= not((layer0_outputs(6279)) xor (layer0_outputs(5448)));
    layer1_outputs(8853) <= not(layer0_outputs(8119));
    layer1_outputs(8854) <= not((layer0_outputs(9909)) and (layer0_outputs(2267)));
    layer1_outputs(8855) <= (layer0_outputs(9082)) and (layer0_outputs(6037));
    layer1_outputs(8856) <= not(layer0_outputs(5470)) or (layer0_outputs(2676));
    layer1_outputs(8857) <= '0';
    layer1_outputs(8858) <= not((layer0_outputs(1536)) or (layer0_outputs(3429)));
    layer1_outputs(8859) <= not((layer0_outputs(7381)) or (layer0_outputs(5098)));
    layer1_outputs(8860) <= not((layer0_outputs(8087)) and (layer0_outputs(6919)));
    layer1_outputs(8861) <= layer0_outputs(2876);
    layer1_outputs(8862) <= not((layer0_outputs(4532)) and (layer0_outputs(10037)));
    layer1_outputs(8863) <= not(layer0_outputs(3484));
    layer1_outputs(8864) <= not(layer0_outputs(9016)) or (layer0_outputs(6023));
    layer1_outputs(8865) <= (layer0_outputs(641)) or (layer0_outputs(1262));
    layer1_outputs(8866) <= layer0_outputs(5739);
    layer1_outputs(8867) <= not((layer0_outputs(2692)) xor (layer0_outputs(5273)));
    layer1_outputs(8868) <= layer0_outputs(3964);
    layer1_outputs(8869) <= (layer0_outputs(6247)) or (layer0_outputs(8153));
    layer1_outputs(8870) <= not(layer0_outputs(5885));
    layer1_outputs(8871) <= not(layer0_outputs(3098)) or (layer0_outputs(8727));
    layer1_outputs(8872) <= (layer0_outputs(7535)) and (layer0_outputs(4160));
    layer1_outputs(8873) <= not(layer0_outputs(2268)) or (layer0_outputs(1457));
    layer1_outputs(8874) <= (layer0_outputs(2028)) or (layer0_outputs(2258));
    layer1_outputs(8875) <= not((layer0_outputs(6293)) or (layer0_outputs(408)));
    layer1_outputs(8876) <= not((layer0_outputs(9239)) or (layer0_outputs(3892)));
    layer1_outputs(8877) <= layer0_outputs(4417);
    layer1_outputs(8878) <= not(layer0_outputs(9912));
    layer1_outputs(8879) <= layer0_outputs(854);
    layer1_outputs(8880) <= not(layer0_outputs(1397));
    layer1_outputs(8881) <= not(layer0_outputs(1885));
    layer1_outputs(8882) <= not(layer0_outputs(4255));
    layer1_outputs(8883) <= layer0_outputs(3914);
    layer1_outputs(8884) <= not((layer0_outputs(6759)) xor (layer0_outputs(9811)));
    layer1_outputs(8885) <= not(layer0_outputs(522));
    layer1_outputs(8886) <= (layer0_outputs(9163)) and not (layer0_outputs(10202));
    layer1_outputs(8887) <= not(layer0_outputs(7114)) or (layer0_outputs(8120));
    layer1_outputs(8888) <= layer0_outputs(5753);
    layer1_outputs(8889) <= not((layer0_outputs(4087)) and (layer0_outputs(3096)));
    layer1_outputs(8890) <= (layer0_outputs(2159)) or (layer0_outputs(3500));
    layer1_outputs(8891) <= (layer0_outputs(3461)) or (layer0_outputs(5850));
    layer1_outputs(8892) <= layer0_outputs(8525);
    layer1_outputs(8893) <= not((layer0_outputs(3381)) and (layer0_outputs(9484)));
    layer1_outputs(8894) <= not(layer0_outputs(7022)) or (layer0_outputs(2503));
    layer1_outputs(8895) <= layer0_outputs(1522);
    layer1_outputs(8896) <= not(layer0_outputs(7439));
    layer1_outputs(8897) <= (layer0_outputs(9327)) and (layer0_outputs(2128));
    layer1_outputs(8898) <= '0';
    layer1_outputs(8899) <= (layer0_outputs(3407)) and not (layer0_outputs(1231));
    layer1_outputs(8900) <= not(layer0_outputs(5022));
    layer1_outputs(8901) <= layer0_outputs(6329);
    layer1_outputs(8902) <= layer0_outputs(6668);
    layer1_outputs(8903) <= not(layer0_outputs(8520)) or (layer0_outputs(4684));
    layer1_outputs(8904) <= (layer0_outputs(8794)) and not (layer0_outputs(6325));
    layer1_outputs(8905) <= not((layer0_outputs(6910)) and (layer0_outputs(7049)));
    layer1_outputs(8906) <= not(layer0_outputs(5167));
    layer1_outputs(8907) <= layer0_outputs(8723);
    layer1_outputs(8908) <= (layer0_outputs(3995)) and not (layer0_outputs(9980));
    layer1_outputs(8909) <= layer0_outputs(7518);
    layer1_outputs(8910) <= not(layer0_outputs(4148));
    layer1_outputs(8911) <= not(layer0_outputs(2361));
    layer1_outputs(8912) <= (layer0_outputs(5453)) and (layer0_outputs(7402));
    layer1_outputs(8913) <= not((layer0_outputs(7589)) and (layer0_outputs(956)));
    layer1_outputs(8914) <= '0';
    layer1_outputs(8915) <= not(layer0_outputs(10042));
    layer1_outputs(8916) <= not(layer0_outputs(8850)) or (layer0_outputs(3767));
    layer1_outputs(8917) <= (layer0_outputs(4735)) or (layer0_outputs(7858));
    layer1_outputs(8918) <= layer0_outputs(7297);
    layer1_outputs(8919) <= layer0_outputs(199);
    layer1_outputs(8920) <= not(layer0_outputs(5322));
    layer1_outputs(8921) <= not(layer0_outputs(5532));
    layer1_outputs(8922) <= not((layer0_outputs(1394)) or (layer0_outputs(6449)));
    layer1_outputs(8923) <= not(layer0_outputs(5234));
    layer1_outputs(8924) <= not(layer0_outputs(6224));
    layer1_outputs(8925) <= layer0_outputs(1106);
    layer1_outputs(8926) <= layer0_outputs(1839);
    layer1_outputs(8927) <= not((layer0_outputs(5224)) or (layer0_outputs(6672)));
    layer1_outputs(8928) <= not(layer0_outputs(1205));
    layer1_outputs(8929) <= layer0_outputs(8860);
    layer1_outputs(8930) <= not(layer0_outputs(7339));
    layer1_outputs(8931) <= not((layer0_outputs(2235)) or (layer0_outputs(5214)));
    layer1_outputs(8932) <= not(layer0_outputs(3158));
    layer1_outputs(8933) <= '1';
    layer1_outputs(8934) <= not(layer0_outputs(1710));
    layer1_outputs(8935) <= not(layer0_outputs(7774));
    layer1_outputs(8936) <= '0';
    layer1_outputs(8937) <= not(layer0_outputs(8113));
    layer1_outputs(8938) <= not((layer0_outputs(5931)) or (layer0_outputs(4204)));
    layer1_outputs(8939) <= (layer0_outputs(3882)) and not (layer0_outputs(1709));
    layer1_outputs(8940) <= not(layer0_outputs(1661));
    layer1_outputs(8941) <= not(layer0_outputs(9353));
    layer1_outputs(8942) <= (layer0_outputs(4671)) or (layer0_outputs(9637));
    layer1_outputs(8943) <= (layer0_outputs(1237)) and not (layer0_outputs(6747));
    layer1_outputs(8944) <= not(layer0_outputs(9154));
    layer1_outputs(8945) <= not(layer0_outputs(5783)) or (layer0_outputs(4089));
    layer1_outputs(8946) <= not(layer0_outputs(4363));
    layer1_outputs(8947) <= not((layer0_outputs(3632)) or (layer0_outputs(5794)));
    layer1_outputs(8948) <= layer0_outputs(2154);
    layer1_outputs(8949) <= layer0_outputs(3469);
    layer1_outputs(8950) <= not(layer0_outputs(2490));
    layer1_outputs(8951) <= (layer0_outputs(1271)) or (layer0_outputs(9826));
    layer1_outputs(8952) <= (layer0_outputs(10199)) or (layer0_outputs(3823));
    layer1_outputs(8953) <= not(layer0_outputs(1420)) or (layer0_outputs(9097));
    layer1_outputs(8954) <= not(layer0_outputs(8623)) or (layer0_outputs(8312));
    layer1_outputs(8955) <= not(layer0_outputs(2751)) or (layer0_outputs(3083));
    layer1_outputs(8956) <= '0';
    layer1_outputs(8957) <= not((layer0_outputs(10085)) or (layer0_outputs(9890)));
    layer1_outputs(8958) <= (layer0_outputs(8577)) and (layer0_outputs(2565));
    layer1_outputs(8959) <= layer0_outputs(1695);
    layer1_outputs(8960) <= layer0_outputs(5872);
    layer1_outputs(8961) <= (layer0_outputs(2551)) and (layer0_outputs(204));
    layer1_outputs(8962) <= (layer0_outputs(3281)) xor (layer0_outputs(1521));
    layer1_outputs(8963) <= not((layer0_outputs(5286)) xor (layer0_outputs(296)));
    layer1_outputs(8964) <= not((layer0_outputs(9235)) xor (layer0_outputs(1328)));
    layer1_outputs(8965) <= not(layer0_outputs(4475));
    layer1_outputs(8966) <= not(layer0_outputs(1313));
    layer1_outputs(8967) <= layer0_outputs(904);
    layer1_outputs(8968) <= '0';
    layer1_outputs(8969) <= layer0_outputs(5900);
    layer1_outputs(8970) <= (layer0_outputs(9781)) and (layer0_outputs(4268));
    layer1_outputs(8971) <= '0';
    layer1_outputs(8972) <= layer0_outputs(9761);
    layer1_outputs(8973) <= not(layer0_outputs(4592));
    layer1_outputs(8974) <= not(layer0_outputs(7051));
    layer1_outputs(8975) <= layer0_outputs(3945);
    layer1_outputs(8976) <= not(layer0_outputs(6481));
    layer1_outputs(8977) <= layer0_outputs(2747);
    layer1_outputs(8978) <= '1';
    layer1_outputs(8979) <= (layer0_outputs(8532)) and (layer0_outputs(4821));
    layer1_outputs(8980) <= layer0_outputs(1985);
    layer1_outputs(8981) <= (layer0_outputs(3684)) and not (layer0_outputs(1039));
    layer1_outputs(8982) <= not(layer0_outputs(8063));
    layer1_outputs(8983) <= not(layer0_outputs(2676));
    layer1_outputs(8984) <= layer0_outputs(614);
    layer1_outputs(8985) <= (layer0_outputs(1654)) or (layer0_outputs(8604));
    layer1_outputs(8986) <= (layer0_outputs(10063)) xor (layer0_outputs(4370));
    layer1_outputs(8987) <= not(layer0_outputs(6722)) or (layer0_outputs(10126));
    layer1_outputs(8988) <= layer0_outputs(7379);
    layer1_outputs(8989) <= not(layer0_outputs(4965));
    layer1_outputs(8990) <= not(layer0_outputs(7000)) or (layer0_outputs(5219));
    layer1_outputs(8991) <= not(layer0_outputs(3886)) or (layer0_outputs(1822));
    layer1_outputs(8992) <= '0';
    layer1_outputs(8993) <= not(layer0_outputs(5268)) or (layer0_outputs(10212));
    layer1_outputs(8994) <= (layer0_outputs(5170)) and not (layer0_outputs(357));
    layer1_outputs(8995) <= not(layer0_outputs(3924));
    layer1_outputs(8996) <= layer0_outputs(7768);
    layer1_outputs(8997) <= '0';
    layer1_outputs(8998) <= layer0_outputs(8688);
    layer1_outputs(8999) <= layer0_outputs(4456);
    layer1_outputs(9000) <= layer0_outputs(7673);
    layer1_outputs(9001) <= (layer0_outputs(5779)) or (layer0_outputs(5206));
    layer1_outputs(9002) <= not(layer0_outputs(9185));
    layer1_outputs(9003) <= (layer0_outputs(3999)) and (layer0_outputs(3052));
    layer1_outputs(9004) <= not((layer0_outputs(453)) or (layer0_outputs(9754)));
    layer1_outputs(9005) <= not(layer0_outputs(8457));
    layer1_outputs(9006) <= not(layer0_outputs(1760)) or (layer0_outputs(1348));
    layer1_outputs(9007) <= layer0_outputs(540);
    layer1_outputs(9008) <= (layer0_outputs(8858)) and not (layer0_outputs(3235));
    layer1_outputs(9009) <= (layer0_outputs(1473)) and not (layer0_outputs(7281));
    layer1_outputs(9010) <= layer0_outputs(3453);
    layer1_outputs(9011) <= layer0_outputs(9812);
    layer1_outputs(9012) <= not(layer0_outputs(8867));
    layer1_outputs(9013) <= layer0_outputs(8791);
    layer1_outputs(9014) <= not(layer0_outputs(83)) or (layer0_outputs(9282));
    layer1_outputs(9015) <= not((layer0_outputs(10124)) or (layer0_outputs(682)));
    layer1_outputs(9016) <= layer0_outputs(7183);
    layer1_outputs(9017) <= not(layer0_outputs(6039));
    layer1_outputs(9018) <= not(layer0_outputs(3481));
    layer1_outputs(9019) <= not(layer0_outputs(6190)) or (layer0_outputs(1790));
    layer1_outputs(9020) <= layer0_outputs(3638);
    layer1_outputs(9021) <= (layer0_outputs(5371)) or (layer0_outputs(8259));
    layer1_outputs(9022) <= not(layer0_outputs(4030)) or (layer0_outputs(2110));
    layer1_outputs(9023) <= (layer0_outputs(4015)) or (layer0_outputs(8448));
    layer1_outputs(9024) <= (layer0_outputs(7958)) or (layer0_outputs(1122));
    layer1_outputs(9025) <= not((layer0_outputs(4354)) and (layer0_outputs(7861)));
    layer1_outputs(9026) <= not(layer0_outputs(9617));
    layer1_outputs(9027) <= layer0_outputs(7457);
    layer1_outputs(9028) <= not(layer0_outputs(5943));
    layer1_outputs(9029) <= not((layer0_outputs(1276)) xor (layer0_outputs(4176)));
    layer1_outputs(9030) <= (layer0_outputs(6752)) and not (layer0_outputs(8074));
    layer1_outputs(9031) <= not(layer0_outputs(9691));
    layer1_outputs(9032) <= (layer0_outputs(6027)) and (layer0_outputs(6576));
    layer1_outputs(9033) <= (layer0_outputs(3182)) or (layer0_outputs(9103));
    layer1_outputs(9034) <= (layer0_outputs(7250)) or (layer0_outputs(2685));
    layer1_outputs(9035) <= not(layer0_outputs(1853)) or (layer0_outputs(9437));
    layer1_outputs(9036) <= not(layer0_outputs(5027));
    layer1_outputs(9037) <= '1';
    layer1_outputs(9038) <= (layer0_outputs(4426)) or (layer0_outputs(3775));
    layer1_outputs(9039) <= not(layer0_outputs(4543));
    layer1_outputs(9040) <= not((layer0_outputs(3256)) or (layer0_outputs(2236)));
    layer1_outputs(9041) <= (layer0_outputs(1683)) and (layer0_outputs(387));
    layer1_outputs(9042) <= not(layer0_outputs(3339));
    layer1_outputs(9043) <= not((layer0_outputs(4125)) xor (layer0_outputs(6485)));
    layer1_outputs(9044) <= not((layer0_outputs(9628)) and (layer0_outputs(6451)));
    layer1_outputs(9045) <= not((layer0_outputs(9347)) or (layer0_outputs(5265)));
    layer1_outputs(9046) <= (layer0_outputs(9843)) and not (layer0_outputs(4494));
    layer1_outputs(9047) <= not((layer0_outputs(6509)) xor (layer0_outputs(3648)));
    layer1_outputs(9048) <= layer0_outputs(410);
    layer1_outputs(9049) <= layer0_outputs(8560);
    layer1_outputs(9050) <= (layer0_outputs(5966)) and (layer0_outputs(6464));
    layer1_outputs(9051) <= layer0_outputs(6796);
    layer1_outputs(9052) <= not(layer0_outputs(4099));
    layer1_outputs(9053) <= (layer0_outputs(8408)) and not (layer0_outputs(2509));
    layer1_outputs(9054) <= not(layer0_outputs(1895));
    layer1_outputs(9055) <= not(layer0_outputs(6487)) or (layer0_outputs(1720));
    layer1_outputs(9056) <= not(layer0_outputs(1067));
    layer1_outputs(9057) <= layer0_outputs(4413);
    layer1_outputs(9058) <= (layer0_outputs(1522)) and not (layer0_outputs(1748));
    layer1_outputs(9059) <= (layer0_outputs(314)) and not (layer0_outputs(547));
    layer1_outputs(9060) <= (layer0_outputs(4759)) and (layer0_outputs(365));
    layer1_outputs(9061) <= not(layer0_outputs(2389));
    layer1_outputs(9062) <= (layer0_outputs(9968)) and not (layer0_outputs(5817));
    layer1_outputs(9063) <= layer0_outputs(7490);
    layer1_outputs(9064) <= not((layer0_outputs(3234)) or (layer0_outputs(3836)));
    layer1_outputs(9065) <= layer0_outputs(3412);
    layer1_outputs(9066) <= not(layer0_outputs(7061));
    layer1_outputs(9067) <= (layer0_outputs(3257)) and not (layer0_outputs(7451));
    layer1_outputs(9068) <= '0';
    layer1_outputs(9069) <= not(layer0_outputs(3202)) or (layer0_outputs(6973));
    layer1_outputs(9070) <= (layer0_outputs(7)) or (layer0_outputs(6352));
    layer1_outputs(9071) <= not(layer0_outputs(3895));
    layer1_outputs(9072) <= not(layer0_outputs(1898)) or (layer0_outputs(7299));
    layer1_outputs(9073) <= (layer0_outputs(3809)) and (layer0_outputs(9949));
    layer1_outputs(9074) <= layer0_outputs(3496);
    layer1_outputs(9075) <= (layer0_outputs(962)) and not (layer0_outputs(8802));
    layer1_outputs(9076) <= layer0_outputs(373);
    layer1_outputs(9077) <= not(layer0_outputs(7250)) or (layer0_outputs(6392));
    layer1_outputs(9078) <= not((layer0_outputs(5099)) xor (layer0_outputs(4364)));
    layer1_outputs(9079) <= not(layer0_outputs(2557)) or (layer0_outputs(9638));
    layer1_outputs(9080) <= not(layer0_outputs(2495));
    layer1_outputs(9081) <= not(layer0_outputs(8072));
    layer1_outputs(9082) <= (layer0_outputs(8274)) and (layer0_outputs(3861));
    layer1_outputs(9083) <= (layer0_outputs(4400)) and (layer0_outputs(608));
    layer1_outputs(9084) <= not(layer0_outputs(8996));
    layer1_outputs(9085) <= not(layer0_outputs(9790));
    layer1_outputs(9086) <= not((layer0_outputs(5090)) or (layer0_outputs(5)));
    layer1_outputs(9087) <= layer0_outputs(6255);
    layer1_outputs(9088) <= (layer0_outputs(655)) and not (layer0_outputs(4443));
    layer1_outputs(9089) <= not(layer0_outputs(1221));
    layer1_outputs(9090) <= not(layer0_outputs(2475));
    layer1_outputs(9091) <= (layer0_outputs(9895)) and not (layer0_outputs(3219));
    layer1_outputs(9092) <= not((layer0_outputs(4240)) and (layer0_outputs(1847)));
    layer1_outputs(9093) <= not(layer0_outputs(7000));
    layer1_outputs(9094) <= (layer0_outputs(6962)) and not (layer0_outputs(8656));
    layer1_outputs(9095) <= layer0_outputs(2657);
    layer1_outputs(9096) <= not(layer0_outputs(6774));
    layer1_outputs(9097) <= '0';
    layer1_outputs(9098) <= '0';
    layer1_outputs(9099) <= '1';
    layer1_outputs(9100) <= not(layer0_outputs(3611));
    layer1_outputs(9101) <= not((layer0_outputs(4863)) and (layer0_outputs(770)));
    layer1_outputs(9102) <= not(layer0_outputs(10114)) or (layer0_outputs(3612));
    layer1_outputs(9103) <= (layer0_outputs(9675)) and (layer0_outputs(5293));
    layer1_outputs(9104) <= (layer0_outputs(9224)) xor (layer0_outputs(2246));
    layer1_outputs(9105) <= not(layer0_outputs(5070));
    layer1_outputs(9106) <= not((layer0_outputs(1720)) or (layer0_outputs(2112)));
    layer1_outputs(9107) <= not((layer0_outputs(3426)) or (layer0_outputs(10179)));
    layer1_outputs(9108) <= (layer0_outputs(1914)) xor (layer0_outputs(314));
    layer1_outputs(9109) <= layer0_outputs(7420);
    layer1_outputs(9110) <= (layer0_outputs(10126)) and not (layer0_outputs(7891));
    layer1_outputs(9111) <= not(layer0_outputs(6468));
    layer1_outputs(9112) <= layer0_outputs(2528);
    layer1_outputs(9113) <= (layer0_outputs(4275)) and not (layer0_outputs(143));
    layer1_outputs(9114) <= not(layer0_outputs(7176));
    layer1_outputs(9115) <= not((layer0_outputs(1969)) xor (layer0_outputs(5106)));
    layer1_outputs(9116) <= (layer0_outputs(7215)) or (layer0_outputs(8714));
    layer1_outputs(9117) <= (layer0_outputs(3418)) xor (layer0_outputs(2482));
    layer1_outputs(9118) <= '1';
    layer1_outputs(9119) <= (layer0_outputs(5081)) or (layer0_outputs(3235));
    layer1_outputs(9120) <= (layer0_outputs(9542)) and (layer0_outputs(5474));
    layer1_outputs(9121) <= (layer0_outputs(8915)) or (layer0_outputs(1376));
    layer1_outputs(9122) <= '0';
    layer1_outputs(9123) <= not(layer0_outputs(4274));
    layer1_outputs(9124) <= (layer0_outputs(2293)) xor (layer0_outputs(8163));
    layer1_outputs(9125) <= not(layer0_outputs(8731));
    layer1_outputs(9126) <= not(layer0_outputs(5736));
    layer1_outputs(9127) <= not(layer0_outputs(9654)) or (layer0_outputs(9823));
    layer1_outputs(9128) <= layer0_outputs(3670);
    layer1_outputs(9129) <= not(layer0_outputs(9329));
    layer1_outputs(9130) <= layer0_outputs(1248);
    layer1_outputs(9131) <= not(layer0_outputs(9629));
    layer1_outputs(9132) <= '1';
    layer1_outputs(9133) <= (layer0_outputs(6646)) and (layer0_outputs(3355));
    layer1_outputs(9134) <= not(layer0_outputs(7841));
    layer1_outputs(9135) <= (layer0_outputs(5813)) and (layer0_outputs(1177));
    layer1_outputs(9136) <= not(layer0_outputs(2576)) or (layer0_outputs(5135));
    layer1_outputs(9137) <= layer0_outputs(737);
    layer1_outputs(9138) <= not((layer0_outputs(7658)) or (layer0_outputs(8119)));
    layer1_outputs(9139) <= not(layer0_outputs(7112));
    layer1_outputs(9140) <= not((layer0_outputs(5228)) and (layer0_outputs(42)));
    layer1_outputs(9141) <= layer0_outputs(4191);
    layer1_outputs(9142) <= (layer0_outputs(3685)) and not (layer0_outputs(1989));
    layer1_outputs(9143) <= not((layer0_outputs(2360)) xor (layer0_outputs(957)));
    layer1_outputs(9144) <= not(layer0_outputs(9783));
    layer1_outputs(9145) <= not(layer0_outputs(2922));
    layer1_outputs(9146) <= not(layer0_outputs(6074));
    layer1_outputs(9147) <= (layer0_outputs(5094)) and (layer0_outputs(4051));
    layer1_outputs(9148) <= (layer0_outputs(841)) or (layer0_outputs(3604));
    layer1_outputs(9149) <= (layer0_outputs(2787)) and (layer0_outputs(7162));
    layer1_outputs(9150) <= not(layer0_outputs(6719)) or (layer0_outputs(9552));
    layer1_outputs(9151) <= not(layer0_outputs(6017));
    layer1_outputs(9152) <= not(layer0_outputs(909)) or (layer0_outputs(156));
    layer1_outputs(9153) <= layer0_outputs(9040);
    layer1_outputs(9154) <= (layer0_outputs(6978)) and (layer0_outputs(667));
    layer1_outputs(9155) <= (layer0_outputs(9396)) and not (layer0_outputs(6916));
    layer1_outputs(9156) <= not(layer0_outputs(589)) or (layer0_outputs(5840));
    layer1_outputs(9157) <= not(layer0_outputs(1740));
    layer1_outputs(9158) <= (layer0_outputs(6516)) xor (layer0_outputs(8973));
    layer1_outputs(9159) <= layer0_outputs(6295);
    layer1_outputs(9160) <= not((layer0_outputs(655)) or (layer0_outputs(4350)));
    layer1_outputs(9161) <= not(layer0_outputs(5967));
    layer1_outputs(9162) <= not(layer0_outputs(5421));
    layer1_outputs(9163) <= (layer0_outputs(1433)) and not (layer0_outputs(6897));
    layer1_outputs(9164) <= '1';
    layer1_outputs(9165) <= not(layer0_outputs(6985)) or (layer0_outputs(2223));
    layer1_outputs(9166) <= layer0_outputs(4464);
    layer1_outputs(9167) <= '1';
    layer1_outputs(9168) <= (layer0_outputs(8243)) and (layer0_outputs(5897));
    layer1_outputs(9169) <= (layer0_outputs(2317)) xor (layer0_outputs(6020));
    layer1_outputs(9170) <= (layer0_outputs(3618)) or (layer0_outputs(1425));
    layer1_outputs(9171) <= not(layer0_outputs(2301)) or (layer0_outputs(3494));
    layer1_outputs(9172) <= (layer0_outputs(5724)) and not (layer0_outputs(8792));
    layer1_outputs(9173) <= not((layer0_outputs(4703)) or (layer0_outputs(2983)));
    layer1_outputs(9174) <= not((layer0_outputs(6120)) or (layer0_outputs(1680)));
    layer1_outputs(9175) <= layer0_outputs(5911);
    layer1_outputs(9176) <= not(layer0_outputs(4757));
    layer1_outputs(9177) <= not((layer0_outputs(1516)) and (layer0_outputs(10052)));
    layer1_outputs(9178) <= not(layer0_outputs(5139));
    layer1_outputs(9179) <= not(layer0_outputs(7724)) or (layer0_outputs(4720));
    layer1_outputs(9180) <= '1';
    layer1_outputs(9181) <= layer0_outputs(8150);
    layer1_outputs(9182) <= layer0_outputs(634);
    layer1_outputs(9183) <= not(layer0_outputs(2845)) or (layer0_outputs(9525));
    layer1_outputs(9184) <= not(layer0_outputs(975)) or (layer0_outputs(8544));
    layer1_outputs(9185) <= (layer0_outputs(9878)) and not (layer0_outputs(5868));
    layer1_outputs(9186) <= not(layer0_outputs(737));
    layer1_outputs(9187) <= (layer0_outputs(5288)) and not (layer0_outputs(7734));
    layer1_outputs(9188) <= (layer0_outputs(4307)) and (layer0_outputs(391));
    layer1_outputs(9189) <= (layer0_outputs(9269)) and not (layer0_outputs(4204));
    layer1_outputs(9190) <= not(layer0_outputs(321)) or (layer0_outputs(5707));
    layer1_outputs(9191) <= (layer0_outputs(7054)) or (layer0_outputs(2229));
    layer1_outputs(9192) <= not((layer0_outputs(3851)) or (layer0_outputs(256)));
    layer1_outputs(9193) <= layer0_outputs(7567);
    layer1_outputs(9194) <= not((layer0_outputs(4002)) and (layer0_outputs(7973)));
    layer1_outputs(9195) <= not(layer0_outputs(7749));
    layer1_outputs(9196) <= layer0_outputs(5984);
    layer1_outputs(9197) <= (layer0_outputs(2132)) xor (layer0_outputs(4085));
    layer1_outputs(9198) <= layer0_outputs(7324);
    layer1_outputs(9199) <= layer0_outputs(6624);
    layer1_outputs(9200) <= not(layer0_outputs(8489));
    layer1_outputs(9201) <= (layer0_outputs(8173)) xor (layer0_outputs(7217));
    layer1_outputs(9202) <= not(layer0_outputs(916)) or (layer0_outputs(4721));
    layer1_outputs(9203) <= not(layer0_outputs(8806)) or (layer0_outputs(5385));
    layer1_outputs(9204) <= layer0_outputs(1596);
    layer1_outputs(9205) <= not(layer0_outputs(6809)) or (layer0_outputs(164));
    layer1_outputs(9206) <= not(layer0_outputs(2029)) or (layer0_outputs(9479));
    layer1_outputs(9207) <= not(layer0_outputs(1997));
    layer1_outputs(9208) <= layer0_outputs(3645);
    layer1_outputs(9209) <= (layer0_outputs(4900)) and not (layer0_outputs(6381));
    layer1_outputs(9210) <= not(layer0_outputs(9346));
    layer1_outputs(9211) <= (layer0_outputs(8071)) or (layer0_outputs(7897));
    layer1_outputs(9212) <= layer0_outputs(65);
    layer1_outputs(9213) <= layer0_outputs(3304);
    layer1_outputs(9214) <= not(layer0_outputs(8972));
    layer1_outputs(9215) <= '1';
    layer1_outputs(9216) <= layer0_outputs(3131);
    layer1_outputs(9217) <= not((layer0_outputs(5158)) xor (layer0_outputs(2130)));
    layer1_outputs(9218) <= (layer0_outputs(4882)) or (layer0_outputs(8049));
    layer1_outputs(9219) <= '1';
    layer1_outputs(9220) <= not(layer0_outputs(4930)) or (layer0_outputs(5631));
    layer1_outputs(9221) <= (layer0_outputs(7161)) and not (layer0_outputs(251));
    layer1_outputs(9222) <= (layer0_outputs(2099)) and not (layer0_outputs(2735));
    layer1_outputs(9223) <= (layer0_outputs(7167)) and not (layer0_outputs(6934));
    layer1_outputs(9224) <= not(layer0_outputs(9470)) or (layer0_outputs(7455));
    layer1_outputs(9225) <= layer0_outputs(4577);
    layer1_outputs(9226) <= layer0_outputs(9907);
    layer1_outputs(9227) <= not(layer0_outputs(8781)) or (layer0_outputs(3329));
    layer1_outputs(9228) <= not((layer0_outputs(2305)) or (layer0_outputs(8362)));
    layer1_outputs(9229) <= not((layer0_outputs(4333)) and (layer0_outputs(1971)));
    layer1_outputs(9230) <= not((layer0_outputs(5660)) and (layer0_outputs(8098)));
    layer1_outputs(9231) <= (layer0_outputs(2190)) and (layer0_outputs(9974));
    layer1_outputs(9232) <= (layer0_outputs(9642)) and not (layer0_outputs(1399));
    layer1_outputs(9233) <= (layer0_outputs(1283)) and not (layer0_outputs(4398));
    layer1_outputs(9234) <= (layer0_outputs(4917)) and (layer0_outputs(3802));
    layer1_outputs(9235) <= (layer0_outputs(5445)) or (layer0_outputs(7100));
    layer1_outputs(9236) <= not(layer0_outputs(4873));
    layer1_outputs(9237) <= (layer0_outputs(3507)) and not (layer0_outputs(1411));
    layer1_outputs(9238) <= '1';
    layer1_outputs(9239) <= layer0_outputs(8686);
    layer1_outputs(9240) <= not(layer0_outputs(8895));
    layer1_outputs(9241) <= '1';
    layer1_outputs(9242) <= not((layer0_outputs(3196)) or (layer0_outputs(9795)));
    layer1_outputs(9243) <= (layer0_outputs(4569)) and not (layer0_outputs(3196));
    layer1_outputs(9244) <= not(layer0_outputs(5272));
    layer1_outputs(9245) <= not((layer0_outputs(8438)) and (layer0_outputs(1119)));
    layer1_outputs(9246) <= layer0_outputs(7117);
    layer1_outputs(9247) <= layer0_outputs(3300);
    layer1_outputs(9248) <= (layer0_outputs(4573)) and not (layer0_outputs(6381));
    layer1_outputs(9249) <= not(layer0_outputs(9987)) or (layer0_outputs(1090));
    layer1_outputs(9250) <= not(layer0_outputs(5218));
    layer1_outputs(9251) <= (layer0_outputs(7031)) and (layer0_outputs(9625));
    layer1_outputs(9252) <= (layer0_outputs(9338)) xor (layer0_outputs(6219));
    layer1_outputs(9253) <= not(layer0_outputs(9833));
    layer1_outputs(9254) <= not(layer0_outputs(6371));
    layer1_outputs(9255) <= '1';
    layer1_outputs(9256) <= not(layer0_outputs(3804));
    layer1_outputs(9257) <= layer0_outputs(9317);
    layer1_outputs(9258) <= layer0_outputs(4220);
    layer1_outputs(9259) <= layer0_outputs(3932);
    layer1_outputs(9260) <= not(layer0_outputs(3588));
    layer1_outputs(9261) <= not(layer0_outputs(2809)) or (layer0_outputs(20));
    layer1_outputs(9262) <= (layer0_outputs(8574)) or (layer0_outputs(757));
    layer1_outputs(9263) <= not(layer0_outputs(6952));
    layer1_outputs(9264) <= layer0_outputs(9000);
    layer1_outputs(9265) <= layer0_outputs(2034);
    layer1_outputs(9266) <= not((layer0_outputs(637)) xor (layer0_outputs(523)));
    layer1_outputs(9267) <= not(layer0_outputs(2911)) or (layer0_outputs(7019));
    layer1_outputs(9268) <= not(layer0_outputs(4557));
    layer1_outputs(9269) <= not((layer0_outputs(7360)) or (layer0_outputs(518)));
    layer1_outputs(9270) <= layer0_outputs(8437);
    layer1_outputs(9271) <= not(layer0_outputs(1055)) or (layer0_outputs(1761));
    layer1_outputs(9272) <= not((layer0_outputs(10018)) or (layer0_outputs(10065)));
    layer1_outputs(9273) <= not(layer0_outputs(5994));
    layer1_outputs(9274) <= (layer0_outputs(3705)) and not (layer0_outputs(4916));
    layer1_outputs(9275) <= not(layer0_outputs(5856));
    layer1_outputs(9276) <= not(layer0_outputs(5199)) or (layer0_outputs(9508));
    layer1_outputs(9277) <= '1';
    layer1_outputs(9278) <= layer0_outputs(8866);
    layer1_outputs(9279) <= not(layer0_outputs(102));
    layer1_outputs(9280) <= (layer0_outputs(8139)) or (layer0_outputs(1934));
    layer1_outputs(9281) <= (layer0_outputs(2693)) and not (layer0_outputs(9397));
    layer1_outputs(9282) <= layer0_outputs(697);
    layer1_outputs(9283) <= not(layer0_outputs(8720));
    layer1_outputs(9284) <= (layer0_outputs(7371)) xor (layer0_outputs(8871));
    layer1_outputs(9285) <= not((layer0_outputs(8239)) or (layer0_outputs(1707)));
    layer1_outputs(9286) <= (layer0_outputs(4983)) and (layer0_outputs(9945));
    layer1_outputs(9287) <= (layer0_outputs(9183)) xor (layer0_outputs(2747));
    layer1_outputs(9288) <= not(layer0_outputs(1917));
    layer1_outputs(9289) <= (layer0_outputs(8472)) and not (layer0_outputs(9719));
    layer1_outputs(9290) <= layer0_outputs(4522);
    layer1_outputs(9291) <= (layer0_outputs(6095)) and not (layer0_outputs(16));
    layer1_outputs(9292) <= not(layer0_outputs(8735));
    layer1_outputs(9293) <= not(layer0_outputs(9922));
    layer1_outputs(9294) <= not(layer0_outputs(4991));
    layer1_outputs(9295) <= not(layer0_outputs(9158)) or (layer0_outputs(9295));
    layer1_outputs(9296) <= not((layer0_outputs(677)) xor (layer0_outputs(9842)));
    layer1_outputs(9297) <= not(layer0_outputs(1336));
    layer1_outputs(9298) <= not(layer0_outputs(8739));
    layer1_outputs(9299) <= (layer0_outputs(5234)) and (layer0_outputs(9162));
    layer1_outputs(9300) <= (layer0_outputs(1257)) or (layer0_outputs(8829));
    layer1_outputs(9301) <= (layer0_outputs(6971)) and not (layer0_outputs(1103));
    layer1_outputs(9302) <= (layer0_outputs(758)) xor (layer0_outputs(9241));
    layer1_outputs(9303) <= not((layer0_outputs(8762)) xor (layer0_outputs(2913)));
    layer1_outputs(9304) <= not((layer0_outputs(170)) and (layer0_outputs(2774)));
    layer1_outputs(9305) <= not((layer0_outputs(954)) and (layer0_outputs(9727)));
    layer1_outputs(9306) <= '0';
    layer1_outputs(9307) <= (layer0_outputs(9944)) xor (layer0_outputs(2554));
    layer1_outputs(9308) <= (layer0_outputs(8715)) and (layer0_outputs(3304));
    layer1_outputs(9309) <= (layer0_outputs(7323)) xor (layer0_outputs(7505));
    layer1_outputs(9310) <= '1';
    layer1_outputs(9311) <= not((layer0_outputs(3773)) or (layer0_outputs(496)));
    layer1_outputs(9312) <= not(layer0_outputs(5696));
    layer1_outputs(9313) <= layer0_outputs(8101);
    layer1_outputs(9314) <= not((layer0_outputs(936)) or (layer0_outputs(3012)));
    layer1_outputs(9315) <= not((layer0_outputs(3742)) xor (layer0_outputs(3472)));
    layer1_outputs(9316) <= layer0_outputs(1398);
    layer1_outputs(9317) <= layer0_outputs(5559);
    layer1_outputs(9318) <= not(layer0_outputs(869));
    layer1_outputs(9319) <= (layer0_outputs(5295)) and not (layer0_outputs(7108));
    layer1_outputs(9320) <= not(layer0_outputs(511));
    layer1_outputs(9321) <= not((layer0_outputs(2206)) and (layer0_outputs(8294)));
    layer1_outputs(9322) <= layer0_outputs(221);
    layer1_outputs(9323) <= not((layer0_outputs(9218)) or (layer0_outputs(4478)));
    layer1_outputs(9324) <= not(layer0_outputs(3004));
    layer1_outputs(9325) <= not(layer0_outputs(4010)) or (layer0_outputs(8116));
    layer1_outputs(9326) <= not((layer0_outputs(2951)) xor (layer0_outputs(3704)));
    layer1_outputs(9327) <= not(layer0_outputs(9095)) or (layer0_outputs(1391));
    layer1_outputs(9328) <= (layer0_outputs(663)) xor (layer0_outputs(3054));
    layer1_outputs(9329) <= (layer0_outputs(2093)) and (layer0_outputs(3829));
    layer1_outputs(9330) <= layer0_outputs(1443);
    layer1_outputs(9331) <= (layer0_outputs(10122)) and (layer0_outputs(6101));
    layer1_outputs(9332) <= not(layer0_outputs(1239)) or (layer0_outputs(9493));
    layer1_outputs(9333) <= layer0_outputs(3308);
    layer1_outputs(9334) <= layer0_outputs(8816);
    layer1_outputs(9335) <= layer0_outputs(8675);
    layer1_outputs(9336) <= not((layer0_outputs(2233)) or (layer0_outputs(5451)));
    layer1_outputs(9337) <= not(layer0_outputs(9919)) or (layer0_outputs(7275));
    layer1_outputs(9338) <= (layer0_outputs(9532)) and (layer0_outputs(1922));
    layer1_outputs(9339) <= layer0_outputs(4483);
    layer1_outputs(9340) <= not((layer0_outputs(6399)) and (layer0_outputs(5574)));
    layer1_outputs(9341) <= layer0_outputs(10005);
    layer1_outputs(9342) <= (layer0_outputs(812)) and not (layer0_outputs(6249));
    layer1_outputs(9343) <= (layer0_outputs(364)) and not (layer0_outputs(3320));
    layer1_outputs(9344) <= layer0_outputs(6715);
    layer1_outputs(9345) <= not(layer0_outputs(7782));
    layer1_outputs(9346) <= not(layer0_outputs(6301)) or (layer0_outputs(5615));
    layer1_outputs(9347) <= layer0_outputs(4465);
    layer1_outputs(9348) <= not((layer0_outputs(423)) xor (layer0_outputs(1861)));
    layer1_outputs(9349) <= layer0_outputs(8053);
    layer1_outputs(9350) <= not(layer0_outputs(3104));
    layer1_outputs(9351) <= (layer0_outputs(5779)) or (layer0_outputs(9777));
    layer1_outputs(9352) <= (layer0_outputs(1802)) and (layer0_outputs(8200));
    layer1_outputs(9353) <= (layer0_outputs(3585)) xor (layer0_outputs(7798));
    layer1_outputs(9354) <= layer0_outputs(4648);
    layer1_outputs(9355) <= layer0_outputs(7873);
    layer1_outputs(9356) <= '0';
    layer1_outputs(9357) <= layer0_outputs(8328);
    layer1_outputs(9358) <= layer0_outputs(5977);
    layer1_outputs(9359) <= not(layer0_outputs(6528)) or (layer0_outputs(7500));
    layer1_outputs(9360) <= (layer0_outputs(6544)) or (layer0_outputs(1859));
    layer1_outputs(9361) <= '0';
    layer1_outputs(9362) <= '0';
    layer1_outputs(9363) <= layer0_outputs(2810);
    layer1_outputs(9364) <= '0';
    layer1_outputs(9365) <= not(layer0_outputs(8147));
    layer1_outputs(9366) <= (layer0_outputs(2169)) or (layer0_outputs(7056));
    layer1_outputs(9367) <= (layer0_outputs(8212)) and not (layer0_outputs(10098));
    layer1_outputs(9368) <= not(layer0_outputs(2464));
    layer1_outputs(9369) <= layer0_outputs(5518);
    layer1_outputs(9370) <= (layer0_outputs(4531)) and not (layer0_outputs(3493));
    layer1_outputs(9371) <= '0';
    layer1_outputs(9372) <= not(layer0_outputs(7364)) or (layer0_outputs(6156));
    layer1_outputs(9373) <= not((layer0_outputs(5508)) or (layer0_outputs(4705)));
    layer1_outputs(9374) <= (layer0_outputs(9354)) xor (layer0_outputs(8788));
    layer1_outputs(9375) <= not((layer0_outputs(689)) xor (layer0_outputs(9685)));
    layer1_outputs(9376) <= (layer0_outputs(8346)) and not (layer0_outputs(635));
    layer1_outputs(9377) <= (layer0_outputs(1719)) and not (layer0_outputs(18));
    layer1_outputs(9378) <= not((layer0_outputs(8202)) or (layer0_outputs(2869)));
    layer1_outputs(9379) <= not(layer0_outputs(2244));
    layer1_outputs(9380) <= not(layer0_outputs(5041)) or (layer0_outputs(7900));
    layer1_outputs(9381) <= (layer0_outputs(5481)) and not (layer0_outputs(6982));
    layer1_outputs(9382) <= not(layer0_outputs(136));
    layer1_outputs(9383) <= (layer0_outputs(471)) and (layer0_outputs(5418));
    layer1_outputs(9384) <= not((layer0_outputs(7948)) or (layer0_outputs(3984)));
    layer1_outputs(9385) <= not((layer0_outputs(865)) and (layer0_outputs(658)));
    layer1_outputs(9386) <= not(layer0_outputs(1637)) or (layer0_outputs(9718));
    layer1_outputs(9387) <= (layer0_outputs(2078)) and not (layer0_outputs(437));
    layer1_outputs(9388) <= not(layer0_outputs(9244));
    layer1_outputs(9389) <= (layer0_outputs(2584)) and (layer0_outputs(6298));
    layer1_outputs(9390) <= not(layer0_outputs(2409)) or (layer0_outputs(8894));
    layer1_outputs(9391) <= not(layer0_outputs(501));
    layer1_outputs(9392) <= layer0_outputs(3417);
    layer1_outputs(9393) <= not(layer0_outputs(10145));
    layer1_outputs(9394) <= (layer0_outputs(2374)) and not (layer0_outputs(438));
    layer1_outputs(9395) <= layer0_outputs(475);
    layer1_outputs(9396) <= not((layer0_outputs(6981)) xor (layer0_outputs(545)));
    layer1_outputs(9397) <= not(layer0_outputs(5015));
    layer1_outputs(9398) <= not((layer0_outputs(8062)) or (layer0_outputs(3874)));
    layer1_outputs(9399) <= not(layer0_outputs(8017));
    layer1_outputs(9400) <= layer0_outputs(5990);
    layer1_outputs(9401) <= not(layer0_outputs(2668));
    layer1_outputs(9402) <= (layer0_outputs(10032)) and not (layer0_outputs(6790));
    layer1_outputs(9403) <= not((layer0_outputs(4657)) or (layer0_outputs(3430)));
    layer1_outputs(9404) <= (layer0_outputs(8862)) or (layer0_outputs(10053));
    layer1_outputs(9405) <= not((layer0_outputs(8336)) and (layer0_outputs(9548)));
    layer1_outputs(9406) <= layer0_outputs(6486);
    layer1_outputs(9407) <= not(layer0_outputs(1622));
    layer1_outputs(9408) <= not(layer0_outputs(6186));
    layer1_outputs(9409) <= not(layer0_outputs(7090));
    layer1_outputs(9410) <= not(layer0_outputs(838)) or (layer0_outputs(5090));
    layer1_outputs(9411) <= not(layer0_outputs(10024));
    layer1_outputs(9412) <= (layer0_outputs(4258)) and (layer0_outputs(5196));
    layer1_outputs(9413) <= layer0_outputs(5825);
    layer1_outputs(9414) <= not((layer0_outputs(1890)) and (layer0_outputs(445)));
    layer1_outputs(9415) <= '1';
    layer1_outputs(9416) <= '1';
    layer1_outputs(9417) <= not(layer0_outputs(8317));
    layer1_outputs(9418) <= not((layer0_outputs(8302)) and (layer0_outputs(4945)));
    layer1_outputs(9419) <= not((layer0_outputs(3172)) or (layer0_outputs(1815)));
    layer1_outputs(9420) <= not(layer0_outputs(2589));
    layer1_outputs(9421) <= layer0_outputs(4302);
    layer1_outputs(9422) <= not(layer0_outputs(10097));
    layer1_outputs(9423) <= (layer0_outputs(72)) and not (layer0_outputs(7115));
    layer1_outputs(9424) <= not(layer0_outputs(3095));
    layer1_outputs(9425) <= not(layer0_outputs(9156));
    layer1_outputs(9426) <= (layer0_outputs(9825)) and (layer0_outputs(7070));
    layer1_outputs(9427) <= not(layer0_outputs(2656)) or (layer0_outputs(7109));
    layer1_outputs(9428) <= (layer0_outputs(7990)) and not (layer0_outputs(1976));
    layer1_outputs(9429) <= not(layer0_outputs(5052));
    layer1_outputs(9430) <= layer0_outputs(6417);
    layer1_outputs(9431) <= not((layer0_outputs(2613)) and (layer0_outputs(5855)));
    layer1_outputs(9432) <= layer0_outputs(1983);
    layer1_outputs(9433) <= not((layer0_outputs(5180)) and (layer0_outputs(9824)));
    layer1_outputs(9434) <= not(layer0_outputs(1229));
    layer1_outputs(9435) <= not(layer0_outputs(10014));
    layer1_outputs(9436) <= not(layer0_outputs(1476));
    layer1_outputs(9437) <= (layer0_outputs(679)) and not (layer0_outputs(6666));
    layer1_outputs(9438) <= not(layer0_outputs(5841));
    layer1_outputs(9439) <= layer0_outputs(2032);
    layer1_outputs(9440) <= not(layer0_outputs(685));
    layer1_outputs(9441) <= (layer0_outputs(4969)) and (layer0_outputs(213));
    layer1_outputs(9442) <= (layer0_outputs(5292)) and not (layer0_outputs(10136));
    layer1_outputs(9443) <= (layer0_outputs(617)) and not (layer0_outputs(8175));
    layer1_outputs(9444) <= not(layer0_outputs(6401));
    layer1_outputs(9445) <= not(layer0_outputs(8477)) or (layer0_outputs(4923));
    layer1_outputs(9446) <= not(layer0_outputs(3266));
    layer1_outputs(9447) <= not((layer0_outputs(3438)) and (layer0_outputs(6223)));
    layer1_outputs(9448) <= (layer0_outputs(6932)) xor (layer0_outputs(7415));
    layer1_outputs(9449) <= (layer0_outputs(2111)) and not (layer0_outputs(6145));
    layer1_outputs(9450) <= not(layer0_outputs(3316)) or (layer0_outputs(5935));
    layer1_outputs(9451) <= layer0_outputs(9213);
    layer1_outputs(9452) <= layer0_outputs(3595);
    layer1_outputs(9453) <= layer0_outputs(1855);
    layer1_outputs(9454) <= not(layer0_outputs(9060));
    layer1_outputs(9455) <= layer0_outputs(1934);
    layer1_outputs(9456) <= layer0_outputs(8131);
    layer1_outputs(9457) <= not(layer0_outputs(912)) or (layer0_outputs(908));
    layer1_outputs(9458) <= not((layer0_outputs(2265)) xor (layer0_outputs(9499)));
    layer1_outputs(9459) <= not(layer0_outputs(2911)) or (layer0_outputs(4021));
    layer1_outputs(9460) <= not(layer0_outputs(7627));
    layer1_outputs(9461) <= layer0_outputs(1418);
    layer1_outputs(9462) <= not(layer0_outputs(3278));
    layer1_outputs(9463) <= (layer0_outputs(2587)) or (layer0_outputs(8619));
    layer1_outputs(9464) <= not((layer0_outputs(5712)) or (layer0_outputs(1811)));
    layer1_outputs(9465) <= not((layer0_outputs(4908)) and (layer0_outputs(3112)));
    layer1_outputs(9466) <= '1';
    layer1_outputs(9467) <= not(layer0_outputs(1020));
    layer1_outputs(9468) <= not(layer0_outputs(6066));
    layer1_outputs(9469) <= not(layer0_outputs(7834));
    layer1_outputs(9470) <= layer0_outputs(2715);
    layer1_outputs(9471) <= (layer0_outputs(456)) and not (layer0_outputs(301));
    layer1_outputs(9472) <= '0';
    layer1_outputs(9473) <= layer0_outputs(1405);
    layer1_outputs(9474) <= '0';
    layer1_outputs(9475) <= (layer0_outputs(379)) xor (layer0_outputs(9041));
    layer1_outputs(9476) <= not(layer0_outputs(408));
    layer1_outputs(9477) <= (layer0_outputs(279)) xor (layer0_outputs(4436));
    layer1_outputs(9478) <= layer0_outputs(7429);
    layer1_outputs(9479) <= not(layer0_outputs(7974)) or (layer0_outputs(8681));
    layer1_outputs(9480) <= '0';
    layer1_outputs(9481) <= layer0_outputs(4732);
    layer1_outputs(9482) <= not((layer0_outputs(6687)) or (layer0_outputs(6931)));
    layer1_outputs(9483) <= layer0_outputs(4761);
    layer1_outputs(9484) <= not(layer0_outputs(2391)) or (layer0_outputs(3071));
    layer1_outputs(9485) <= not(layer0_outputs(1368));
    layer1_outputs(9486) <= (layer0_outputs(6678)) and (layer0_outputs(8736));
    layer1_outputs(9487) <= not(layer0_outputs(6331));
    layer1_outputs(9488) <= not(layer0_outputs(8864));
    layer1_outputs(9489) <= (layer0_outputs(3345)) and (layer0_outputs(5739));
    layer1_outputs(9490) <= not(layer0_outputs(6146)) or (layer0_outputs(4113));
    layer1_outputs(9491) <= layer0_outputs(9710);
    layer1_outputs(9492) <= (layer0_outputs(9602)) and not (layer0_outputs(3197));
    layer1_outputs(9493) <= layer0_outputs(8054);
    layer1_outputs(9494) <= (layer0_outputs(2778)) xor (layer0_outputs(6020));
    layer1_outputs(9495) <= layer0_outputs(7767);
    layer1_outputs(9496) <= (layer0_outputs(3643)) xor (layer0_outputs(7813));
    layer1_outputs(9497) <= not((layer0_outputs(2693)) xor (layer0_outputs(4990)));
    layer1_outputs(9498) <= layer0_outputs(4340);
    layer1_outputs(9499) <= '1';
    layer1_outputs(9500) <= layer0_outputs(3347);
    layer1_outputs(9501) <= (layer0_outputs(9987)) or (layer0_outputs(10005));
    layer1_outputs(9502) <= (layer0_outputs(8414)) xor (layer0_outputs(8646));
    layer1_outputs(9503) <= (layer0_outputs(10214)) xor (layer0_outputs(3837));
    layer1_outputs(9504) <= (layer0_outputs(6541)) and not (layer0_outputs(9839));
    layer1_outputs(9505) <= layer0_outputs(1565);
    layer1_outputs(9506) <= '0';
    layer1_outputs(9507) <= (layer0_outputs(6346)) or (layer0_outputs(7957));
    layer1_outputs(9508) <= (layer0_outputs(4594)) and not (layer0_outputs(1085));
    layer1_outputs(9509) <= (layer0_outputs(5565)) and not (layer0_outputs(3298));
    layer1_outputs(9510) <= not((layer0_outputs(2326)) or (layer0_outputs(2748)));
    layer1_outputs(9511) <= not((layer0_outputs(1249)) and (layer0_outputs(7918)));
    layer1_outputs(9512) <= layer0_outputs(6871);
    layer1_outputs(9513) <= layer0_outputs(9323);
    layer1_outputs(9514) <= not(layer0_outputs(5887)) or (layer0_outputs(2712));
    layer1_outputs(9515) <= not(layer0_outputs(5286)) or (layer0_outputs(2398));
    layer1_outputs(9516) <= not(layer0_outputs(4730)) or (layer0_outputs(1064));
    layer1_outputs(9517) <= layer0_outputs(10176);
    layer1_outputs(9518) <= not((layer0_outputs(63)) xor (layer0_outputs(9258)));
    layer1_outputs(9519) <= layer0_outputs(7835);
    layer1_outputs(9520) <= (layer0_outputs(9838)) and (layer0_outputs(7510));
    layer1_outputs(9521) <= (layer0_outputs(3697)) xor (layer0_outputs(3892));
    layer1_outputs(9522) <= (layer0_outputs(8878)) and (layer0_outputs(3210));
    layer1_outputs(9523) <= layer0_outputs(58);
    layer1_outputs(9524) <= layer0_outputs(1694);
    layer1_outputs(9525) <= layer0_outputs(9640);
    layer1_outputs(9526) <= not(layer0_outputs(160)) or (layer0_outputs(7371));
    layer1_outputs(9527) <= (layer0_outputs(5858)) and not (layer0_outputs(10115));
    layer1_outputs(9528) <= (layer0_outputs(2228)) and not (layer0_outputs(5460));
    layer1_outputs(9529) <= not(layer0_outputs(5359)) or (layer0_outputs(5121));
    layer1_outputs(9530) <= layer0_outputs(5610);
    layer1_outputs(9531) <= layer0_outputs(7811);
    layer1_outputs(9532) <= (layer0_outputs(1379)) and not (layer0_outputs(4517));
    layer1_outputs(9533) <= not(layer0_outputs(4951));
    layer1_outputs(9534) <= (layer0_outputs(4159)) and not (layer0_outputs(1066));
    layer1_outputs(9535) <= not(layer0_outputs(5705));
    layer1_outputs(9536) <= not(layer0_outputs(6467)) or (layer0_outputs(6356));
    layer1_outputs(9537) <= (layer0_outputs(5693)) and (layer0_outputs(620));
    layer1_outputs(9538) <= not(layer0_outputs(6309));
    layer1_outputs(9539) <= '1';
    layer1_outputs(9540) <= not((layer0_outputs(193)) and (layer0_outputs(10095)));
    layer1_outputs(9541) <= (layer0_outputs(3845)) or (layer0_outputs(2895));
    layer1_outputs(9542) <= (layer0_outputs(4858)) and not (layer0_outputs(127));
    layer1_outputs(9543) <= '1';
    layer1_outputs(9544) <= (layer0_outputs(4181)) and not (layer0_outputs(7523));
    layer1_outputs(9545) <= (layer0_outputs(75)) and (layer0_outputs(7310));
    layer1_outputs(9546) <= (layer0_outputs(9433)) and not (layer0_outputs(8277));
    layer1_outputs(9547) <= not(layer0_outputs(8333)) or (layer0_outputs(6011));
    layer1_outputs(9548) <= layer0_outputs(9039);
    layer1_outputs(9549) <= not(layer0_outputs(7311));
    layer1_outputs(9550) <= not(layer0_outputs(6583));
    layer1_outputs(9551) <= not((layer0_outputs(4331)) or (layer0_outputs(7932)));
    layer1_outputs(9552) <= (layer0_outputs(6349)) and not (layer0_outputs(552));
    layer1_outputs(9553) <= not((layer0_outputs(4568)) and (layer0_outputs(9934)));
    layer1_outputs(9554) <= layer0_outputs(2684);
    layer1_outputs(9555) <= (layer0_outputs(6771)) xor (layer0_outputs(8079));
    layer1_outputs(9556) <= '1';
    layer1_outputs(9557) <= layer0_outputs(5744);
    layer1_outputs(9558) <= not(layer0_outputs(7463)) or (layer0_outputs(7703));
    layer1_outputs(9559) <= (layer0_outputs(6825)) or (layer0_outputs(6748));
    layer1_outputs(9560) <= not((layer0_outputs(6285)) or (layer0_outputs(135)));
    layer1_outputs(9561) <= layer0_outputs(3723);
    layer1_outputs(9562) <= (layer0_outputs(9485)) and (layer0_outputs(1223));
    layer1_outputs(9563) <= not((layer0_outputs(7826)) xor (layer0_outputs(5994)));
    layer1_outputs(9564) <= not(layer0_outputs(7481));
    layer1_outputs(9565) <= (layer0_outputs(8433)) xor (layer0_outputs(8258));
    layer1_outputs(9566) <= (layer0_outputs(9)) and not (layer0_outputs(2781));
    layer1_outputs(9567) <= not(layer0_outputs(1301)) or (layer0_outputs(567));
    layer1_outputs(9568) <= (layer0_outputs(6413)) and (layer0_outputs(2513));
    layer1_outputs(9569) <= (layer0_outputs(9293)) and not (layer0_outputs(1852));
    layer1_outputs(9570) <= '1';
    layer1_outputs(9571) <= not(layer0_outputs(3711));
    layer1_outputs(9572) <= layer0_outputs(1779);
    layer1_outputs(9573) <= layer0_outputs(5585);
    layer1_outputs(9574) <= (layer0_outputs(1824)) and (layer0_outputs(5211));
    layer1_outputs(9575) <= not(layer0_outputs(298));
    layer1_outputs(9576) <= not(layer0_outputs(4279)) or (layer0_outputs(8409));
    layer1_outputs(9577) <= (layer0_outputs(9358)) and not (layer0_outputs(10057));
    layer1_outputs(9578) <= (layer0_outputs(6901)) and not (layer0_outputs(3272));
    layer1_outputs(9579) <= (layer0_outputs(10142)) and not (layer0_outputs(6206));
    layer1_outputs(9580) <= (layer0_outputs(3309)) or (layer0_outputs(7719));
    layer1_outputs(9581) <= layer0_outputs(142);
    layer1_outputs(9582) <= not(layer0_outputs(9205));
    layer1_outputs(9583) <= not(layer0_outputs(2573));
    layer1_outputs(9584) <= layer0_outputs(2602);
    layer1_outputs(9585) <= not(layer0_outputs(1028));
    layer1_outputs(9586) <= (layer0_outputs(3441)) and not (layer0_outputs(1141));
    layer1_outputs(9587) <= not((layer0_outputs(7520)) xor (layer0_outputs(603)));
    layer1_outputs(9588) <= (layer0_outputs(8364)) or (layer0_outputs(6454));
    layer1_outputs(9589) <= not(layer0_outputs(8815)) or (layer0_outputs(7336));
    layer1_outputs(9590) <= not(layer0_outputs(10185)) or (layer0_outputs(918));
    layer1_outputs(9591) <= layer0_outputs(9879);
    layer1_outputs(9592) <= (layer0_outputs(622)) and not (layer0_outputs(8624));
    layer1_outputs(9593) <= layer0_outputs(7248);
    layer1_outputs(9594) <= not(layer0_outputs(6972));
    layer1_outputs(9595) <= not(layer0_outputs(1095));
    layer1_outputs(9596) <= (layer0_outputs(3731)) and not (layer0_outputs(9997));
    layer1_outputs(9597) <= (layer0_outputs(5100)) and (layer0_outputs(8171));
    layer1_outputs(9598) <= not(layer0_outputs(1465));
    layer1_outputs(9599) <= layer0_outputs(219);
    layer1_outputs(9600) <= not(layer0_outputs(948)) or (layer0_outputs(2218));
    layer1_outputs(9601) <= not(layer0_outputs(1957));
    layer1_outputs(9602) <= not((layer0_outputs(2816)) and (layer0_outputs(1177)));
    layer1_outputs(9603) <= not(layer0_outputs(9093));
    layer1_outputs(9604) <= (layer0_outputs(3447)) and (layer0_outputs(7453));
    layer1_outputs(9605) <= not(layer0_outputs(3733));
    layer1_outputs(9606) <= layer0_outputs(1722);
    layer1_outputs(9607) <= '0';
    layer1_outputs(9608) <= not(layer0_outputs(10025));
    layer1_outputs(9609) <= not((layer0_outputs(7572)) xor (layer0_outputs(5337)));
    layer1_outputs(9610) <= not(layer0_outputs(106)) or (layer0_outputs(70));
    layer1_outputs(9611) <= not(layer0_outputs(8818)) or (layer0_outputs(4996));
    layer1_outputs(9612) <= not(layer0_outputs(3661)) or (layer0_outputs(6526));
    layer1_outputs(9613) <= (layer0_outputs(3636)) and (layer0_outputs(9504));
    layer1_outputs(9614) <= not(layer0_outputs(2426));
    layer1_outputs(9615) <= not((layer0_outputs(7682)) and (layer0_outputs(9985)));
    layer1_outputs(9616) <= (layer0_outputs(767)) xor (layer0_outputs(393));
    layer1_outputs(9617) <= not(layer0_outputs(7237)) or (layer0_outputs(9448));
    layer1_outputs(9618) <= not((layer0_outputs(8086)) and (layer0_outputs(5141)));
    layer1_outputs(9619) <= not(layer0_outputs(3454)) or (layer0_outputs(8435));
    layer1_outputs(9620) <= layer0_outputs(2055);
    layer1_outputs(9621) <= (layer0_outputs(2477)) and not (layer0_outputs(3085));
    layer1_outputs(9622) <= not((layer0_outputs(9679)) or (layer0_outputs(8043)));
    layer1_outputs(9623) <= not((layer0_outputs(4226)) and (layer0_outputs(6829)));
    layer1_outputs(9624) <= (layer0_outputs(8588)) and not (layer0_outputs(1262));
    layer1_outputs(9625) <= not((layer0_outputs(800)) and (layer0_outputs(6377)));
    layer1_outputs(9626) <= layer0_outputs(1086);
    layer1_outputs(9627) <= not((layer0_outputs(7406)) or (layer0_outputs(8930)));
    layer1_outputs(9628) <= layer0_outputs(6562);
    layer1_outputs(9629) <= (layer0_outputs(2694)) xor (layer0_outputs(8416));
    layer1_outputs(9630) <= (layer0_outputs(9860)) and not (layer0_outputs(2306));
    layer1_outputs(9631) <= not(layer0_outputs(8697));
    layer1_outputs(9632) <= (layer0_outputs(10085)) and (layer0_outputs(2738));
    layer1_outputs(9633) <= (layer0_outputs(166)) and not (layer0_outputs(4251));
    layer1_outputs(9634) <= (layer0_outputs(8939)) and (layer0_outputs(1680));
    layer1_outputs(9635) <= not(layer0_outputs(6084)) or (layer0_outputs(9496));
    layer1_outputs(9636) <= (layer0_outputs(5044)) and not (layer0_outputs(7229));
    layer1_outputs(9637) <= layer0_outputs(6168);
    layer1_outputs(9638) <= (layer0_outputs(7058)) xor (layer0_outputs(5488));
    layer1_outputs(9639) <= not(layer0_outputs(272));
    layer1_outputs(9640) <= not(layer0_outputs(6355));
    layer1_outputs(9641) <= not((layer0_outputs(242)) and (layer0_outputs(2417)));
    layer1_outputs(9642) <= not((layer0_outputs(7175)) or (layer0_outputs(3351)));
    layer1_outputs(9643) <= '0';
    layer1_outputs(9644) <= '1';
    layer1_outputs(9645) <= not((layer0_outputs(5418)) or (layer0_outputs(1451)));
    layer1_outputs(9646) <= (layer0_outputs(6656)) and not (layer0_outputs(1728));
    layer1_outputs(9647) <= layer0_outputs(1638);
    layer1_outputs(9648) <= layer0_outputs(10031);
    layer1_outputs(9649) <= not(layer0_outputs(7362));
    layer1_outputs(9650) <= (layer0_outputs(1227)) xor (layer0_outputs(6921));
    layer1_outputs(9651) <= not(layer0_outputs(3340));
    layer1_outputs(9652) <= not(layer0_outputs(3034));
    layer1_outputs(9653) <= (layer0_outputs(2254)) xor (layer0_outputs(8934));
    layer1_outputs(9654) <= not(layer0_outputs(4961));
    layer1_outputs(9655) <= (layer0_outputs(5899)) and not (layer0_outputs(5219));
    layer1_outputs(9656) <= layer0_outputs(5516);
    layer1_outputs(9657) <= not(layer0_outputs(6384));
    layer1_outputs(9658) <= layer0_outputs(5307);
    layer1_outputs(9659) <= not(layer0_outputs(6054));
    layer1_outputs(9660) <= not(layer0_outputs(6929));
    layer1_outputs(9661) <= not(layer0_outputs(5438));
    layer1_outputs(9662) <= not(layer0_outputs(3840));
    layer1_outputs(9663) <= not(layer0_outputs(3327)) or (layer0_outputs(4396));
    layer1_outputs(9664) <= (layer0_outputs(4946)) and not (layer0_outputs(1747));
    layer1_outputs(9665) <= layer0_outputs(2424);
    layer1_outputs(9666) <= layer0_outputs(5482);
    layer1_outputs(9667) <= layer0_outputs(136);
    layer1_outputs(9668) <= not(layer0_outputs(597));
    layer1_outputs(9669) <= not((layer0_outputs(7041)) and (layer0_outputs(9483)));
    layer1_outputs(9670) <= not((layer0_outputs(8037)) xor (layer0_outputs(6602)));
    layer1_outputs(9671) <= (layer0_outputs(65)) or (layer0_outputs(5367));
    layer1_outputs(9672) <= (layer0_outputs(7825)) and not (layer0_outputs(7779));
    layer1_outputs(9673) <= not(layer0_outputs(9566));
    layer1_outputs(9674) <= not((layer0_outputs(6551)) and (layer0_outputs(3766)));
    layer1_outputs(9675) <= not(layer0_outputs(5235)) or (layer0_outputs(3078));
    layer1_outputs(9676) <= not(layer0_outputs(8479)) or (layer0_outputs(2369));
    layer1_outputs(9677) <= (layer0_outputs(7060)) and (layer0_outputs(9943));
    layer1_outputs(9678) <= layer0_outputs(4558);
    layer1_outputs(9679) <= layer0_outputs(8661);
    layer1_outputs(9680) <= (layer0_outputs(6903)) xor (layer0_outputs(5311));
    layer1_outputs(9681) <= '1';
    layer1_outputs(9682) <= not(layer0_outputs(7698));
    layer1_outputs(9683) <= not(layer0_outputs(9928)) or (layer0_outputs(1108));
    layer1_outputs(9684) <= layer0_outputs(6453);
    layer1_outputs(9685) <= layer0_outputs(9801);
    layer1_outputs(9686) <= layer0_outputs(2621);
    layer1_outputs(9687) <= layer0_outputs(300);
    layer1_outputs(9688) <= '0';
    layer1_outputs(9689) <= layer0_outputs(5273);
    layer1_outputs(9690) <= (layer0_outputs(7416)) and not (layer0_outputs(4092));
    layer1_outputs(9691) <= not(layer0_outputs(10149));
    layer1_outputs(9692) <= (layer0_outputs(1311)) xor (layer0_outputs(228));
    layer1_outputs(9693) <= not((layer0_outputs(8096)) xor (layer0_outputs(6078)));
    layer1_outputs(9694) <= not(layer0_outputs(5309));
    layer1_outputs(9695) <= not(layer0_outputs(5940));
    layer1_outputs(9696) <= not(layer0_outputs(4860));
    layer1_outputs(9697) <= layer0_outputs(8608);
    layer1_outputs(9698) <= not(layer0_outputs(9690));
    layer1_outputs(9699) <= not(layer0_outputs(7688));
    layer1_outputs(9700) <= not(layer0_outputs(7830));
    layer1_outputs(9701) <= not(layer0_outputs(9262)) or (layer0_outputs(4458));
    layer1_outputs(9702) <= (layer0_outputs(3794)) and not (layer0_outputs(4045));
    layer1_outputs(9703) <= not(layer0_outputs(6846));
    layer1_outputs(9704) <= not(layer0_outputs(8646));
    layer1_outputs(9705) <= not(layer0_outputs(9616));
    layer1_outputs(9706) <= not((layer0_outputs(9088)) and (layer0_outputs(4511)));
    layer1_outputs(9707) <= not(layer0_outputs(3355));
    layer1_outputs(9708) <= layer0_outputs(2849);
    layer1_outputs(9709) <= (layer0_outputs(6949)) or (layer0_outputs(2129));
    layer1_outputs(9710) <= (layer0_outputs(8664)) and (layer0_outputs(101));
    layer1_outputs(9711) <= not((layer0_outputs(6644)) or (layer0_outputs(1347)));
    layer1_outputs(9712) <= layer0_outputs(4226);
    layer1_outputs(9713) <= (layer0_outputs(4799)) and (layer0_outputs(6416));
    layer1_outputs(9714) <= not(layer0_outputs(5909));
    layer1_outputs(9715) <= not(layer0_outputs(4500));
    layer1_outputs(9716) <= not(layer0_outputs(7525));
    layer1_outputs(9717) <= not(layer0_outputs(1967));
    layer1_outputs(9718) <= layer0_outputs(8104);
    layer1_outputs(9719) <= not((layer0_outputs(7620)) or (layer0_outputs(5477)));
    layer1_outputs(9720) <= not(layer0_outputs(7569)) or (layer0_outputs(8643));
    layer1_outputs(9721) <= '0';
    layer1_outputs(9722) <= layer0_outputs(7996);
    layer1_outputs(9723) <= not((layer0_outputs(1182)) or (layer0_outputs(1854)));
    layer1_outputs(9724) <= not((layer0_outputs(2209)) xor (layer0_outputs(6208)));
    layer1_outputs(9725) <= layer0_outputs(6920);
    layer1_outputs(9726) <= (layer0_outputs(8793)) and not (layer0_outputs(3916));
    layer1_outputs(9727) <= layer0_outputs(6620);
    layer1_outputs(9728) <= (layer0_outputs(6518)) and not (layer0_outputs(924));
    layer1_outputs(9729) <= (layer0_outputs(6000)) xor (layer0_outputs(7494));
    layer1_outputs(9730) <= not(layer0_outputs(7338)) or (layer0_outputs(2478));
    layer1_outputs(9731) <= not(layer0_outputs(9305)) or (layer0_outputs(2930));
    layer1_outputs(9732) <= not(layer0_outputs(4878)) or (layer0_outputs(2906));
    layer1_outputs(9733) <= not(layer0_outputs(2452)) or (layer0_outputs(402));
    layer1_outputs(9734) <= not(layer0_outputs(320));
    layer1_outputs(9735) <= not(layer0_outputs(3291));
    layer1_outputs(9736) <= layer0_outputs(7067);
    layer1_outputs(9737) <= (layer0_outputs(5507)) and not (layer0_outputs(1328));
    layer1_outputs(9738) <= not(layer0_outputs(6179));
    layer1_outputs(9739) <= (layer0_outputs(2146)) and not (layer0_outputs(119));
    layer1_outputs(9740) <= (layer0_outputs(9498)) or (layer0_outputs(8899));
    layer1_outputs(9741) <= layer0_outputs(4230);
    layer1_outputs(9742) <= layer0_outputs(7065);
    layer1_outputs(9743) <= (layer0_outputs(7252)) and not (layer0_outputs(8750));
    layer1_outputs(9744) <= not(layer0_outputs(9959)) or (layer0_outputs(4361));
    layer1_outputs(9745) <= not(layer0_outputs(280)) or (layer0_outputs(1304));
    layer1_outputs(9746) <= not(layer0_outputs(7089)) or (layer0_outputs(9900));
    layer1_outputs(9747) <= not(layer0_outputs(2147)) or (layer0_outputs(6204));
    layer1_outputs(9748) <= layer0_outputs(4063);
    layer1_outputs(9749) <= (layer0_outputs(853)) and not (layer0_outputs(8279));
    layer1_outputs(9750) <= not((layer0_outputs(2297)) xor (layer0_outputs(5034)));
    layer1_outputs(9751) <= (layer0_outputs(3964)) and (layer0_outputs(4469));
    layer1_outputs(9752) <= not(layer0_outputs(4333));
    layer1_outputs(9753) <= layer0_outputs(8958);
    layer1_outputs(9754) <= layer0_outputs(4658);
    layer1_outputs(9755) <= not(layer0_outputs(6437));
    layer1_outputs(9756) <= layer0_outputs(7125);
    layer1_outputs(9757) <= not((layer0_outputs(3591)) and (layer0_outputs(5760)));
    layer1_outputs(9758) <= not(layer0_outputs(2635)) or (layer0_outputs(8167));
    layer1_outputs(9759) <= layer0_outputs(2771);
    layer1_outputs(9760) <= (layer0_outputs(5112)) and not (layer0_outputs(818));
    layer1_outputs(9761) <= '1';
    layer1_outputs(9762) <= not((layer0_outputs(7094)) xor (layer0_outputs(9799)));
    layer1_outputs(9763) <= not(layer0_outputs(9654));
    layer1_outputs(9764) <= (layer0_outputs(627)) and not (layer0_outputs(4809));
    layer1_outputs(9765) <= (layer0_outputs(560)) and not (layer0_outputs(5348));
    layer1_outputs(9766) <= not(layer0_outputs(4030)) or (layer0_outputs(3910));
    layer1_outputs(9767) <= not((layer0_outputs(10159)) or (layer0_outputs(4954)));
    layer1_outputs(9768) <= layer0_outputs(539);
    layer1_outputs(9769) <= not(layer0_outputs(7697));
    layer1_outputs(9770) <= layer0_outputs(2317);
    layer1_outputs(9771) <= layer0_outputs(9543);
    layer1_outputs(9772) <= (layer0_outputs(9038)) and (layer0_outputs(5108));
    layer1_outputs(9773) <= not((layer0_outputs(6233)) and (layer0_outputs(1470)));
    layer1_outputs(9774) <= not((layer0_outputs(1538)) or (layer0_outputs(802)));
    layer1_outputs(9775) <= not((layer0_outputs(7792)) xor (layer0_outputs(4577)));
    layer1_outputs(9776) <= layer0_outputs(5848);
    layer1_outputs(9777) <= not(layer0_outputs(3348));
    layer1_outputs(9778) <= not(layer0_outputs(2291)) or (layer0_outputs(5076));
    layer1_outputs(9779) <= layer0_outputs(8261);
    layer1_outputs(9780) <= not(layer0_outputs(7772));
    layer1_outputs(9781) <= not((layer0_outputs(4033)) and (layer0_outputs(7201)));
    layer1_outputs(9782) <= not(layer0_outputs(2526)) or (layer0_outputs(2287));
    layer1_outputs(9783) <= (layer0_outputs(842)) and not (layer0_outputs(4964));
    layer1_outputs(9784) <= not(layer0_outputs(8484));
    layer1_outputs(9785) <= (layer0_outputs(181)) or (layer0_outputs(1068));
    layer1_outputs(9786) <= not(layer0_outputs(3850));
    layer1_outputs(9787) <= layer0_outputs(6289);
    layer1_outputs(9788) <= layer0_outputs(7353);
    layer1_outputs(9789) <= not((layer0_outputs(6056)) xor (layer0_outputs(8361)));
    layer1_outputs(9790) <= not(layer0_outputs(6346));
    layer1_outputs(9791) <= layer0_outputs(2879);
    layer1_outputs(9792) <= not((layer0_outputs(9433)) xor (layer0_outputs(4776)));
    layer1_outputs(9793) <= not(layer0_outputs(2614));
    layer1_outputs(9794) <= (layer0_outputs(8238)) and (layer0_outputs(292));
    layer1_outputs(9795) <= (layer0_outputs(10060)) and not (layer0_outputs(7500));
    layer1_outputs(9796) <= not((layer0_outputs(1777)) and (layer0_outputs(6905)));
    layer1_outputs(9797) <= not(layer0_outputs(6591)) or (layer0_outputs(6965));
    layer1_outputs(9798) <= (layer0_outputs(8953)) or (layer0_outputs(3462));
    layer1_outputs(9799) <= not(layer0_outputs(5726));
    layer1_outputs(9800) <= not(layer0_outputs(154));
    layer1_outputs(9801) <= not(layer0_outputs(2443));
    layer1_outputs(9802) <= not(layer0_outputs(2887));
    layer1_outputs(9803) <= not(layer0_outputs(4487));
    layer1_outputs(9804) <= (layer0_outputs(5070)) and not (layer0_outputs(5381));
    layer1_outputs(9805) <= not((layer0_outputs(6533)) and (layer0_outputs(8285)));
    layer1_outputs(9806) <= not((layer0_outputs(6524)) or (layer0_outputs(2201)));
    layer1_outputs(9807) <= not(layer0_outputs(4046)) or (layer0_outputs(3845));
    layer1_outputs(9808) <= (layer0_outputs(6309)) or (layer0_outputs(8396));
    layer1_outputs(9809) <= not(layer0_outputs(461)) or (layer0_outputs(7897));
    layer1_outputs(9810) <= (layer0_outputs(1763)) and not (layer0_outputs(7026));
    layer1_outputs(9811) <= layer0_outputs(3367);
    layer1_outputs(9812) <= (layer0_outputs(4354)) and not (layer0_outputs(2142));
    layer1_outputs(9813) <= layer0_outputs(8180);
    layer1_outputs(9814) <= not((layer0_outputs(8778)) or (layer0_outputs(1625)));
    layer1_outputs(9815) <= layer0_outputs(9439);
    layer1_outputs(9816) <= not(layer0_outputs(6473));
    layer1_outputs(9817) <= layer0_outputs(6603);
    layer1_outputs(9818) <= not((layer0_outputs(6895)) or (layer0_outputs(3029)));
    layer1_outputs(9819) <= not(layer0_outputs(8008));
    layer1_outputs(9820) <= layer0_outputs(4664);
    layer1_outputs(9821) <= not(layer0_outputs(3372)) or (layer0_outputs(1460));
    layer1_outputs(9822) <= (layer0_outputs(2632)) or (layer0_outputs(4070));
    layer1_outputs(9823) <= not((layer0_outputs(8407)) and (layer0_outputs(5750)));
    layer1_outputs(9824) <= not(layer0_outputs(5292)) or (layer0_outputs(8959));
    layer1_outputs(9825) <= not(layer0_outputs(8666));
    layer1_outputs(9826) <= (layer0_outputs(9384)) or (layer0_outputs(2));
    layer1_outputs(9827) <= not(layer0_outputs(6529));
    layer1_outputs(9828) <= not(layer0_outputs(5355));
    layer1_outputs(9829) <= (layer0_outputs(9053)) and not (layer0_outputs(6187));
    layer1_outputs(9830) <= not(layer0_outputs(359)) or (layer0_outputs(3830));
    layer1_outputs(9831) <= layer0_outputs(9140);
    layer1_outputs(9832) <= layer0_outputs(4099);
    layer1_outputs(9833) <= layer0_outputs(5232);
    layer1_outputs(9834) <= not(layer0_outputs(7985));
    layer1_outputs(9835) <= not((layer0_outputs(7129)) or (layer0_outputs(1504)));
    layer1_outputs(9836) <= not(layer0_outputs(5962));
    layer1_outputs(9837) <= not((layer0_outputs(563)) xor (layer0_outputs(310)));
    layer1_outputs(9838) <= not(layer0_outputs(7497)) or (layer0_outputs(9278));
    layer1_outputs(9839) <= not((layer0_outputs(7575)) and (layer0_outputs(9402)));
    layer1_outputs(9840) <= not(layer0_outputs(5487));
    layer1_outputs(9841) <= not((layer0_outputs(6777)) and (layer0_outputs(9237)));
    layer1_outputs(9842) <= '0';
    layer1_outputs(9843) <= (layer0_outputs(7491)) and not (layer0_outputs(5153));
    layer1_outputs(9844) <= not((layer0_outputs(8145)) and (layer0_outputs(6894)));
    layer1_outputs(9845) <= not(layer0_outputs(1872));
    layer1_outputs(9846) <= layer0_outputs(8512);
    layer1_outputs(9847) <= not(layer0_outputs(1169)) or (layer0_outputs(827));
    layer1_outputs(9848) <= not(layer0_outputs(5795)) or (layer0_outputs(2307));
    layer1_outputs(9849) <= not(layer0_outputs(8747));
    layer1_outputs(9850) <= not(layer0_outputs(2126));
    layer1_outputs(9851) <= layer0_outputs(3612);
    layer1_outputs(9852) <= (layer0_outputs(5337)) and not (layer0_outputs(8182));
    layer1_outputs(9853) <= (layer0_outputs(5721)) xor (layer0_outputs(4742));
    layer1_outputs(9854) <= (layer0_outputs(2206)) and (layer0_outputs(1537));
    layer1_outputs(9855) <= (layer0_outputs(5414)) and (layer0_outputs(10125));
    layer1_outputs(9856) <= not(layer0_outputs(972)) or (layer0_outputs(3789));
    layer1_outputs(9857) <= layer0_outputs(13);
    layer1_outputs(9858) <= not(layer0_outputs(9008));
    layer1_outputs(9859) <= not(layer0_outputs(1383));
    layer1_outputs(9860) <= not((layer0_outputs(2472)) and (layer0_outputs(2979)));
    layer1_outputs(9861) <= layer0_outputs(1909);
    layer1_outputs(9862) <= not((layer0_outputs(6999)) and (layer0_outputs(8811)));
    layer1_outputs(9863) <= (layer0_outputs(4448)) and not (layer0_outputs(5815));
    layer1_outputs(9864) <= not(layer0_outputs(8187));
    layer1_outputs(9865) <= (layer0_outputs(1230)) and (layer0_outputs(2158));
    layer1_outputs(9866) <= not(layer0_outputs(5723)) or (layer0_outputs(5307));
    layer1_outputs(9867) <= '1';
    layer1_outputs(9868) <= not(layer0_outputs(9834));
    layer1_outputs(9869) <= not((layer0_outputs(8656)) or (layer0_outputs(8443)));
    layer1_outputs(9870) <= '0';
    layer1_outputs(9871) <= not((layer0_outputs(2048)) and (layer0_outputs(1745)));
    layer1_outputs(9872) <= not((layer0_outputs(5600)) and (layer0_outputs(9195)));
    layer1_outputs(9873) <= (layer0_outputs(10073)) and not (layer0_outputs(8793));
    layer1_outputs(9874) <= not(layer0_outputs(1530)) or (layer0_outputs(1820));
    layer1_outputs(9875) <= (layer0_outputs(7009)) and not (layer0_outputs(1559));
    layer1_outputs(9876) <= not(layer0_outputs(7321));
    layer1_outputs(9877) <= (layer0_outputs(318)) or (layer0_outputs(2214));
    layer1_outputs(9878) <= layer0_outputs(8304);
    layer1_outputs(9879) <= not(layer0_outputs(4556)) or (layer0_outputs(7778));
    layer1_outputs(9880) <= not((layer0_outputs(2873)) xor (layer0_outputs(5209)));
    layer1_outputs(9881) <= not(layer0_outputs(4576));
    layer1_outputs(9882) <= (layer0_outputs(9782)) and (layer0_outputs(5713));
    layer1_outputs(9883) <= not(layer0_outputs(9845)) or (layer0_outputs(326));
    layer1_outputs(9884) <= layer0_outputs(6778);
    layer1_outputs(9885) <= (layer0_outputs(8217)) xor (layer0_outputs(8341));
    layer1_outputs(9886) <= not((layer0_outputs(4036)) and (layer0_outputs(9850)));
    layer1_outputs(9887) <= not(layer0_outputs(355));
    layer1_outputs(9888) <= layer0_outputs(8055);
    layer1_outputs(9889) <= layer0_outputs(866);
    layer1_outputs(9890) <= not(layer0_outputs(8077)) or (layer0_outputs(9868));
    layer1_outputs(9891) <= not(layer0_outputs(3056));
    layer1_outputs(9892) <= not(layer0_outputs(6030)) or (layer0_outputs(1285));
    layer1_outputs(9893) <= not((layer0_outputs(4463)) or (layer0_outputs(399)));
    layer1_outputs(9894) <= not(layer0_outputs(3323));
    layer1_outputs(9895) <= (layer0_outputs(8156)) or (layer0_outputs(3835));
    layer1_outputs(9896) <= (layer0_outputs(9863)) or (layer0_outputs(3620));
    layer1_outputs(9897) <= not((layer0_outputs(929)) or (layer0_outputs(6623)));
    layer1_outputs(9898) <= layer0_outputs(4940);
    layer1_outputs(9899) <= not(layer0_outputs(2523));
    layer1_outputs(9900) <= not(layer0_outputs(8364)) or (layer0_outputs(9975));
    layer1_outputs(9901) <= (layer0_outputs(7801)) xor (layer0_outputs(2519));
    layer1_outputs(9902) <= not(layer0_outputs(8523));
    layer1_outputs(9903) <= (layer0_outputs(9252)) and not (layer0_outputs(1932));
    layer1_outputs(9904) <= not((layer0_outputs(4490)) and (layer0_outputs(2499)));
    layer1_outputs(9905) <= not(layer0_outputs(6265)) or (layer0_outputs(2187));
    layer1_outputs(9906) <= not(layer0_outputs(5)) or (layer0_outputs(2259));
    layer1_outputs(9907) <= not(layer0_outputs(567)) or (layer0_outputs(9134));
    layer1_outputs(9908) <= (layer0_outputs(7832)) and (layer0_outputs(5053));
    layer1_outputs(9909) <= not(layer0_outputs(3810));
    layer1_outputs(9910) <= (layer0_outputs(3322)) and not (layer0_outputs(5778));
    layer1_outputs(9911) <= (layer0_outputs(3621)) or (layer0_outputs(6953));
    layer1_outputs(9912) <= layer0_outputs(9139);
    layer1_outputs(9913) <= (layer0_outputs(3800)) and not (layer0_outputs(9808));
    layer1_outputs(9914) <= (layer0_outputs(21)) and not (layer0_outputs(2674));
    layer1_outputs(9915) <= not(layer0_outputs(5487));
    layer1_outputs(9916) <= layer0_outputs(8375);
    layer1_outputs(9917) <= layer0_outputs(2758);
    layer1_outputs(9918) <= layer0_outputs(8564);
    layer1_outputs(9919) <= not(layer0_outputs(247));
    layer1_outputs(9920) <= layer0_outputs(2813);
    layer1_outputs(9921) <= layer0_outputs(5362);
    layer1_outputs(9922) <= layer0_outputs(564);
    layer1_outputs(9923) <= not((layer0_outputs(8509)) or (layer0_outputs(1598)));
    layer1_outputs(9924) <= not(layer0_outputs(4656));
    layer1_outputs(9925) <= layer0_outputs(7020);
    layer1_outputs(9926) <= (layer0_outputs(5198)) and not (layer0_outputs(1256));
    layer1_outputs(9927) <= '0';
    layer1_outputs(9928) <= (layer0_outputs(451)) or (layer0_outputs(2164));
    layer1_outputs(9929) <= (layer0_outputs(8048)) and not (layer0_outputs(4001));
    layer1_outputs(9930) <= not((layer0_outputs(212)) or (layer0_outputs(5827)));
    layer1_outputs(9931) <= not((layer0_outputs(8553)) or (layer0_outputs(6187)));
    layer1_outputs(9932) <= not(layer0_outputs(4505)) or (layer0_outputs(7133));
    layer1_outputs(9933) <= (layer0_outputs(6379)) xor (layer0_outputs(7320));
    layer1_outputs(9934) <= (layer0_outputs(7549)) and (layer0_outputs(1721));
    layer1_outputs(9935) <= layer0_outputs(7230);
    layer1_outputs(9936) <= (layer0_outputs(5709)) or (layer0_outputs(9557));
    layer1_outputs(9937) <= not(layer0_outputs(6794));
    layer1_outputs(9938) <= (layer0_outputs(8591)) or (layer0_outputs(1693));
    layer1_outputs(9939) <= not(layer0_outputs(10003));
    layer1_outputs(9940) <= '0';
    layer1_outputs(9941) <= not(layer0_outputs(9128));
    layer1_outputs(9942) <= layer0_outputs(6658);
    layer1_outputs(9943) <= not(layer0_outputs(6184)) or (layer0_outputs(952));
    layer1_outputs(9944) <= not(layer0_outputs(6883)) or (layer0_outputs(3558));
    layer1_outputs(9945) <= not((layer0_outputs(3732)) xor (layer0_outputs(6077)));
    layer1_outputs(9946) <= not(layer0_outputs(1531)) or (layer0_outputs(5919));
    layer1_outputs(9947) <= not(layer0_outputs(5649)) or (layer0_outputs(1603));
    layer1_outputs(9948) <= (layer0_outputs(8707)) and not (layer0_outputs(4247));
    layer1_outputs(9949) <= (layer0_outputs(7356)) xor (layer0_outputs(347));
    layer1_outputs(9950) <= not((layer0_outputs(2670)) and (layer0_outputs(8173)));
    layer1_outputs(9951) <= (layer0_outputs(1001)) and (layer0_outputs(9306));
    layer1_outputs(9952) <= (layer0_outputs(837)) or (layer0_outputs(9974));
    layer1_outputs(9953) <= layer0_outputs(10237);
    layer1_outputs(9954) <= layer0_outputs(7198);
    layer1_outputs(9955) <= layer0_outputs(1621);
    layer1_outputs(9956) <= not(layer0_outputs(1493));
    layer1_outputs(9957) <= not(layer0_outputs(931)) or (layer0_outputs(1351));
    layer1_outputs(9958) <= layer0_outputs(8921);
    layer1_outputs(9959) <= (layer0_outputs(2527)) and not (layer0_outputs(3819));
    layer1_outputs(9960) <= not(layer0_outputs(2010)) or (layer0_outputs(4800));
    layer1_outputs(9961) <= layer0_outputs(2119);
    layer1_outputs(9962) <= '1';
    layer1_outputs(9963) <= not(layer0_outputs(4075));
    layer1_outputs(9964) <= not(layer0_outputs(3605));
    layer1_outputs(9965) <= not(layer0_outputs(876));
    layer1_outputs(9966) <= not(layer0_outputs(2740));
    layer1_outputs(9967) <= not((layer0_outputs(1528)) xor (layer0_outputs(923)));
    layer1_outputs(9968) <= (layer0_outputs(3146)) and not (layer0_outputs(3971));
    layer1_outputs(9969) <= not(layer0_outputs(259));
    layer1_outputs(9970) <= layer0_outputs(1062);
    layer1_outputs(9971) <= not(layer0_outputs(3482));
    layer1_outputs(9972) <= (layer0_outputs(5890)) and (layer0_outputs(10161));
    layer1_outputs(9973) <= not((layer0_outputs(9142)) and (layer0_outputs(5512)));
    layer1_outputs(9974) <= '1';
    layer1_outputs(9975) <= (layer0_outputs(449)) xor (layer0_outputs(9897));
    layer1_outputs(9976) <= not((layer0_outputs(9328)) and (layer0_outputs(4758)));
    layer1_outputs(9977) <= not(layer0_outputs(8978)) or (layer0_outputs(882));
    layer1_outputs(9978) <= (layer0_outputs(8587)) and not (layer0_outputs(1136));
    layer1_outputs(9979) <= not(layer0_outputs(3890));
    layer1_outputs(9980) <= not(layer0_outputs(9899)) or (layer0_outputs(6128));
    layer1_outputs(9981) <= not(layer0_outputs(5944)) or (layer0_outputs(1022));
    layer1_outputs(9982) <= layer0_outputs(2755);
    layer1_outputs(9983) <= (layer0_outputs(4601)) or (layer0_outputs(4091));
    layer1_outputs(9984) <= not(layer0_outputs(4107)) or (layer0_outputs(6873));
    layer1_outputs(9985) <= (layer0_outputs(4440)) and not (layer0_outputs(9007));
    layer1_outputs(9986) <= not((layer0_outputs(5354)) and (layer0_outputs(7616)));
    layer1_outputs(9987) <= (layer0_outputs(7301)) xor (layer0_outputs(743));
    layer1_outputs(9988) <= (layer0_outputs(1533)) and not (layer0_outputs(8135));
    layer1_outputs(9989) <= (layer0_outputs(7107)) or (layer0_outputs(5751));
    layer1_outputs(9990) <= (layer0_outputs(8092)) and not (layer0_outputs(2496));
    layer1_outputs(9991) <= not(layer0_outputs(3134)) or (layer0_outputs(3498));
    layer1_outputs(9992) <= not(layer0_outputs(9415));
    layer1_outputs(9993) <= (layer0_outputs(2799)) and not (layer0_outputs(9457));
    layer1_outputs(9994) <= '1';
    layer1_outputs(9995) <= not(layer0_outputs(3258)) or (layer0_outputs(175));
    layer1_outputs(9996) <= layer0_outputs(3298);
    layer1_outputs(9997) <= not(layer0_outputs(7312));
    layer1_outputs(9998) <= not(layer0_outputs(6437));
    layer1_outputs(9999) <= layer0_outputs(3483);
    layer1_outputs(10000) <= not((layer0_outputs(3506)) and (layer0_outputs(5804)));
    layer1_outputs(10001) <= not((layer0_outputs(7226)) and (layer0_outputs(5428)));
    layer1_outputs(10002) <= layer0_outputs(8726);
    layer1_outputs(10003) <= not(layer0_outputs(6388));
    layer1_outputs(10004) <= (layer0_outputs(1938)) and not (layer0_outputs(9314));
    layer1_outputs(10005) <= not((layer0_outputs(3574)) or (layer0_outputs(8571)));
    layer1_outputs(10006) <= layer0_outputs(2095);
    layer1_outputs(10007) <= (layer0_outputs(8403)) xor (layer0_outputs(1717));
    layer1_outputs(10008) <= not((layer0_outputs(8201)) or (layer0_outputs(8237)));
    layer1_outputs(10009) <= layer0_outputs(2023);
    layer1_outputs(10010) <= not((layer0_outputs(5080)) xor (layer0_outputs(4507)));
    layer1_outputs(10011) <= layer0_outputs(8486);
    layer1_outputs(10012) <= (layer0_outputs(6566)) and not (layer0_outputs(3537));
    layer1_outputs(10013) <= '0';
    layer1_outputs(10014) <= (layer0_outputs(303)) and (layer0_outputs(1469));
    layer1_outputs(10015) <= not(layer0_outputs(4334));
    layer1_outputs(10016) <= not(layer0_outputs(3876));
    layer1_outputs(10017) <= not((layer0_outputs(2962)) and (layer0_outputs(1290)));
    layer1_outputs(10018) <= not(layer0_outputs(6068)) or (layer0_outputs(2384));
    layer1_outputs(10019) <= not((layer0_outputs(4967)) xor (layer0_outputs(6659)));
    layer1_outputs(10020) <= layer0_outputs(7681);
    layer1_outputs(10021) <= not((layer0_outputs(5396)) or (layer0_outputs(2487)));
    layer1_outputs(10022) <= layer0_outputs(5259);
    layer1_outputs(10023) <= (layer0_outputs(6714)) or (layer0_outputs(4295));
    layer1_outputs(10024) <= layer0_outputs(1884);
    layer1_outputs(10025) <= '0';
    layer1_outputs(10026) <= not(layer0_outputs(6792)) or (layer0_outputs(4250));
    layer1_outputs(10027) <= not(layer0_outputs(1921));
    layer1_outputs(10028) <= (layer0_outputs(2401)) and (layer0_outputs(4073));
    layer1_outputs(10029) <= not((layer0_outputs(4449)) and (layer0_outputs(7601)));
    layer1_outputs(10030) <= (layer0_outputs(4160)) or (layer0_outputs(7470));
    layer1_outputs(10031) <= not(layer0_outputs(9036));
    layer1_outputs(10032) <= layer0_outputs(6077);
    layer1_outputs(10033) <= not(layer0_outputs(3686));
    layer1_outputs(10034) <= layer0_outputs(9152);
    layer1_outputs(10035) <= not(layer0_outputs(2916));
    layer1_outputs(10036) <= layer0_outputs(351);
    layer1_outputs(10037) <= not(layer0_outputs(3674));
    layer1_outputs(10038) <= (layer0_outputs(7561)) and not (layer0_outputs(9447));
    layer1_outputs(10039) <= not(layer0_outputs(5577)) or (layer0_outputs(6086));
    layer1_outputs(10040) <= not((layer0_outputs(4596)) and (layer0_outputs(9970)));
    layer1_outputs(10041) <= '0';
    layer1_outputs(10042) <= not(layer0_outputs(8861)) or (layer0_outputs(8132));
    layer1_outputs(10043) <= (layer0_outputs(7745)) and not (layer0_outputs(9977));
    layer1_outputs(10044) <= not((layer0_outputs(1919)) or (layer0_outputs(505)));
    layer1_outputs(10045) <= (layer0_outputs(4589)) and not (layer0_outputs(6503));
    layer1_outputs(10046) <= (layer0_outputs(1306)) xor (layer0_outputs(3521));
    layer1_outputs(10047) <= not((layer0_outputs(929)) or (layer0_outputs(7944)));
    layer1_outputs(10048) <= not(layer0_outputs(5572));
    layer1_outputs(10049) <= (layer0_outputs(2780)) and not (layer0_outputs(1701));
    layer1_outputs(10050) <= layer0_outputs(2140);
    layer1_outputs(10051) <= (layer0_outputs(4981)) and not (layer0_outputs(3133));
    layer1_outputs(10052) <= not(layer0_outputs(4184)) or (layer0_outputs(1859));
    layer1_outputs(10053) <= layer0_outputs(8833);
    layer1_outputs(10054) <= layer0_outputs(4208);
    layer1_outputs(10055) <= not(layer0_outputs(8288));
    layer1_outputs(10056) <= layer0_outputs(8956);
    layer1_outputs(10057) <= not((layer0_outputs(6258)) or (layer0_outputs(10182)));
    layer1_outputs(10058) <= (layer0_outputs(9472)) and not (layer0_outputs(9377));
    layer1_outputs(10059) <= not(layer0_outputs(4088));
    layer1_outputs(10060) <= not(layer0_outputs(1564));
    layer1_outputs(10061) <= not(layer0_outputs(997));
    layer1_outputs(10062) <= layer0_outputs(126);
    layer1_outputs(10063) <= not(layer0_outputs(9726));
    layer1_outputs(10064) <= layer0_outputs(3444);
    layer1_outputs(10065) <= not((layer0_outputs(8964)) or (layer0_outputs(4090)));
    layer1_outputs(10066) <= layer0_outputs(10076);
    layer1_outputs(10067) <= (layer0_outputs(6214)) and (layer0_outputs(5207));
    layer1_outputs(10068) <= not(layer0_outputs(2424));
    layer1_outputs(10069) <= (layer0_outputs(4751)) and (layer0_outputs(6989));
    layer1_outputs(10070) <= not((layer0_outputs(9471)) and (layer0_outputs(477)));
    layer1_outputs(10071) <= layer0_outputs(8233);
    layer1_outputs(10072) <= not((layer0_outputs(3560)) or (layer0_outputs(7216)));
    layer1_outputs(10073) <= not(layer0_outputs(834));
    layer1_outputs(10074) <= (layer0_outputs(4470)) and not (layer0_outputs(9456));
    layer1_outputs(10075) <= layer0_outputs(4635);
    layer1_outputs(10076) <= not((layer0_outputs(6570)) and (layer0_outputs(7676)));
    layer1_outputs(10077) <= not((layer0_outputs(3520)) and (layer0_outputs(4106)));
    layer1_outputs(10078) <= not((layer0_outputs(10054)) or (layer0_outputs(7840)));
    layer1_outputs(10079) <= not((layer0_outputs(7193)) or (layer0_outputs(10180)));
    layer1_outputs(10080) <= '0';
    layer1_outputs(10081) <= layer0_outputs(9704);
    layer1_outputs(10082) <= not(layer0_outputs(4253)) or (layer0_outputs(2171));
    layer1_outputs(10083) <= not((layer0_outputs(10223)) and (layer0_outputs(5947)));
    layer1_outputs(10084) <= not((layer0_outputs(1510)) xor (layer0_outputs(8589)));
    layer1_outputs(10085) <= '0';
    layer1_outputs(10086) <= layer0_outputs(10110);
    layer1_outputs(10087) <= layer0_outputs(775);
    layer1_outputs(10088) <= not(layer0_outputs(6096)) or (layer0_outputs(2399));
    layer1_outputs(10089) <= not(layer0_outputs(1792));
    layer1_outputs(10090) <= (layer0_outputs(5277)) and not (layer0_outputs(9950));
    layer1_outputs(10091) <= not((layer0_outputs(7354)) xor (layer0_outputs(5113)));
    layer1_outputs(10092) <= layer0_outputs(8253);
    layer1_outputs(10093) <= (layer0_outputs(2019)) and (layer0_outputs(891));
    layer1_outputs(10094) <= not(layer0_outputs(7521));
    layer1_outputs(10095) <= not(layer0_outputs(9955));
    layer1_outputs(10096) <= not(layer0_outputs(891));
    layer1_outputs(10097) <= layer0_outputs(6707);
    layer1_outputs(10098) <= (layer0_outputs(1635)) or (layer0_outputs(477));
    layer1_outputs(10099) <= (layer0_outputs(945)) or (layer0_outputs(2154));
    layer1_outputs(10100) <= not(layer0_outputs(967));
    layer1_outputs(10101) <= layer0_outputs(198);
    layer1_outputs(10102) <= not((layer0_outputs(1161)) xor (layer0_outputs(6673)));
    layer1_outputs(10103) <= not((layer0_outputs(2071)) and (layer0_outputs(7058)));
    layer1_outputs(10104) <= (layer0_outputs(6945)) or (layer0_outputs(3887));
    layer1_outputs(10105) <= layer0_outputs(6620);
    layer1_outputs(10106) <= not((layer0_outputs(9376)) xor (layer0_outputs(6826)));
    layer1_outputs(10107) <= not((layer0_outputs(6821)) and (layer0_outputs(6341)));
    layer1_outputs(10108) <= not(layer0_outputs(5861));
    layer1_outputs(10109) <= (layer0_outputs(382)) or (layer0_outputs(9967));
    layer1_outputs(10110) <= not(layer0_outputs(5667));
    layer1_outputs(10111) <= (layer0_outputs(1430)) and not (layer0_outputs(5081));
    layer1_outputs(10112) <= not((layer0_outputs(1963)) or (layer0_outputs(870)));
    layer1_outputs(10113) <= layer0_outputs(2069);
    layer1_outputs(10114) <= layer0_outputs(9287);
    layer1_outputs(10115) <= not(layer0_outputs(3446)) or (layer0_outputs(6643));
    layer1_outputs(10116) <= layer0_outputs(6823);
    layer1_outputs(10117) <= not((layer0_outputs(3485)) xor (layer0_outputs(4922)));
    layer1_outputs(10118) <= layer0_outputs(4509);
    layer1_outputs(10119) <= '1';
    layer1_outputs(10120) <= not(layer0_outputs(4392));
    layer1_outputs(10121) <= layer0_outputs(351);
    layer1_outputs(10122) <= (layer0_outputs(4012)) or (layer0_outputs(3896));
    layer1_outputs(10123) <= not(layer0_outputs(3153)) or (layer0_outputs(5955));
    layer1_outputs(10124) <= not(layer0_outputs(5306));
    layer1_outputs(10125) <= (layer0_outputs(6731)) or (layer0_outputs(2557));
    layer1_outputs(10126) <= (layer0_outputs(5766)) xor (layer0_outputs(4689));
    layer1_outputs(10127) <= not((layer0_outputs(8462)) and (layer0_outputs(1541)));
    layer1_outputs(10128) <= layer0_outputs(282);
    layer1_outputs(10129) <= (layer0_outputs(4719)) and not (layer0_outputs(4233));
    layer1_outputs(10130) <= (layer0_outputs(6763)) and not (layer0_outputs(6818));
    layer1_outputs(10131) <= (layer0_outputs(8666)) and not (layer0_outputs(255));
    layer1_outputs(10132) <= (layer0_outputs(432)) and (layer0_outputs(5239));
    layer1_outputs(10133) <= (layer0_outputs(9157)) and not (layer0_outputs(8973));
    layer1_outputs(10134) <= layer0_outputs(3497);
    layer1_outputs(10135) <= layer0_outputs(7319);
    layer1_outputs(10136) <= not(layer0_outputs(3318)) or (layer0_outputs(4816));
    layer1_outputs(10137) <= layer0_outputs(5673);
    layer1_outputs(10138) <= not(layer0_outputs(2848)) or (layer0_outputs(8460));
    layer1_outputs(10139) <= not((layer0_outputs(5447)) or (layer0_outputs(5771)));
    layer1_outputs(10140) <= layer0_outputs(4018);
    layer1_outputs(10141) <= (layer0_outputs(4968)) or (layer0_outputs(1225));
    layer1_outputs(10142) <= (layer0_outputs(954)) xor (layer0_outputs(9509));
    layer1_outputs(10143) <= not((layer0_outputs(8880)) xor (layer0_outputs(3177)));
    layer1_outputs(10144) <= (layer0_outputs(1359)) and not (layer0_outputs(502));
    layer1_outputs(10145) <= not(layer0_outputs(2708)) or (layer0_outputs(9157));
    layer1_outputs(10146) <= not((layer0_outputs(3759)) and (layer0_outputs(4828)));
    layer1_outputs(10147) <= (layer0_outputs(5951)) xor (layer0_outputs(4817));
    layer1_outputs(10148) <= layer0_outputs(4335);
    layer1_outputs(10149) <= (layer0_outputs(2820)) and not (layer0_outputs(9242));
    layer1_outputs(10150) <= not(layer0_outputs(7729));
    layer1_outputs(10151) <= layer0_outputs(1077);
    layer1_outputs(10152) <= (layer0_outputs(8530)) or (layer0_outputs(4523));
    layer1_outputs(10153) <= not(layer0_outputs(907));
    layer1_outputs(10154) <= layer0_outputs(6761);
    layer1_outputs(10155) <= layer0_outputs(1057);
    layer1_outputs(10156) <= not(layer0_outputs(4214)) or (layer0_outputs(1970));
    layer1_outputs(10157) <= layer0_outputs(2374);
    layer1_outputs(10158) <= layer0_outputs(2213);
    layer1_outputs(10159) <= (layer0_outputs(487)) or (layer0_outputs(7350));
    layer1_outputs(10160) <= (layer0_outputs(5861)) and not (layer0_outputs(538));
    layer1_outputs(10161) <= (layer0_outputs(4301)) and not (layer0_outputs(4625));
    layer1_outputs(10162) <= layer0_outputs(6091);
    layer1_outputs(10163) <= (layer0_outputs(3119)) or (layer0_outputs(2410));
    layer1_outputs(10164) <= layer0_outputs(2584);
    layer1_outputs(10165) <= layer0_outputs(2722);
    layer1_outputs(10166) <= (layer0_outputs(4306)) xor (layer0_outputs(2390));
    layer1_outputs(10167) <= not(layer0_outputs(6665)) or (layer0_outputs(6972));
    layer1_outputs(10168) <= (layer0_outputs(8073)) and (layer0_outputs(5548));
    layer1_outputs(10169) <= (layer0_outputs(7143)) xor (layer0_outputs(276));
    layer1_outputs(10170) <= not(layer0_outputs(5951));
    layer1_outputs(10171) <= layer0_outputs(4280);
    layer1_outputs(10172) <= not(layer0_outputs(679)) or (layer0_outputs(1566));
    layer1_outputs(10173) <= layer0_outputs(8927);
    layer1_outputs(10174) <= not(layer0_outputs(1436));
    layer1_outputs(10175) <= not(layer0_outputs(3458));
    layer1_outputs(10176) <= not(layer0_outputs(9925));
    layer1_outputs(10177) <= (layer0_outputs(8783)) xor (layer0_outputs(7829));
    layer1_outputs(10178) <= layer0_outputs(1475);
    layer1_outputs(10179) <= not(layer0_outputs(462)) or (layer0_outputs(4741));
    layer1_outputs(10180) <= layer0_outputs(2516);
    layer1_outputs(10181) <= '1';
    layer1_outputs(10182) <= not(layer0_outputs(1151)) or (layer0_outputs(4281));
    layer1_outputs(10183) <= (layer0_outputs(8873)) and not (layer0_outputs(2885));
    layer1_outputs(10184) <= not(layer0_outputs(330));
    layer1_outputs(10185) <= (layer0_outputs(815)) and (layer0_outputs(46));
    layer1_outputs(10186) <= not(layer0_outputs(5348));
    layer1_outputs(10187) <= not(layer0_outputs(1383));
    layer1_outputs(10188) <= layer0_outputs(1199);
    layer1_outputs(10189) <= (layer0_outputs(4112)) and (layer0_outputs(2568));
    layer1_outputs(10190) <= not(layer0_outputs(4293));
    layer1_outputs(10191) <= layer0_outputs(1410);
    layer1_outputs(10192) <= (layer0_outputs(1145)) and not (layer0_outputs(4749));
    layer1_outputs(10193) <= not((layer0_outputs(2579)) and (layer0_outputs(6008)));
    layer1_outputs(10194) <= not(layer0_outputs(1129)) or (layer0_outputs(6065));
    layer1_outputs(10195) <= not(layer0_outputs(1674));
    layer1_outputs(10196) <= layer0_outputs(1455);
    layer1_outputs(10197) <= '0';
    layer1_outputs(10198) <= (layer0_outputs(7217)) and (layer0_outputs(7540));
    layer1_outputs(10199) <= layer0_outputs(5898);
    layer1_outputs(10200) <= not(layer0_outputs(4509));
    layer1_outputs(10201) <= (layer0_outputs(131)) and not (layer0_outputs(5659));
    layer1_outputs(10202) <= not(layer0_outputs(7614));
    layer1_outputs(10203) <= not(layer0_outputs(7249));
    layer1_outputs(10204) <= (layer0_outputs(7817)) and not (layer0_outputs(71));
    layer1_outputs(10205) <= '1';
    layer1_outputs(10206) <= not((layer0_outputs(3544)) or (layer0_outputs(8107)));
    layer1_outputs(10207) <= (layer0_outputs(2245)) or (layer0_outputs(7410));
    layer1_outputs(10208) <= layer0_outputs(5953);
    layer1_outputs(10209) <= (layer0_outputs(6320)) or (layer0_outputs(2019));
    layer1_outputs(10210) <= layer0_outputs(7979);
    layer1_outputs(10211) <= (layer0_outputs(2295)) and (layer0_outputs(1011));
    layer1_outputs(10212) <= '0';
    layer1_outputs(10213) <= not((layer0_outputs(7103)) and (layer0_outputs(7894)));
    layer1_outputs(10214) <= layer0_outputs(299);
    layer1_outputs(10215) <= (layer0_outputs(4300)) and not (layer0_outputs(9141));
    layer1_outputs(10216) <= not((layer0_outputs(9667)) and (layer0_outputs(9026)));
    layer1_outputs(10217) <= not(layer0_outputs(5961)) or (layer0_outputs(1128));
    layer1_outputs(10218) <= (layer0_outputs(5498)) or (layer0_outputs(6705));
    layer1_outputs(10219) <= layer0_outputs(8099);
    layer1_outputs(10220) <= (layer0_outputs(4969)) xor (layer0_outputs(4066));
    layer1_outputs(10221) <= layer0_outputs(2806);
    layer1_outputs(10222) <= not((layer0_outputs(8502)) and (layer0_outputs(3704)));
    layer1_outputs(10223) <= (layer0_outputs(7044)) xor (layer0_outputs(3803));
    layer1_outputs(10224) <= not((layer0_outputs(3404)) or (layer0_outputs(7375)));
    layer1_outputs(10225) <= not(layer0_outputs(3515)) or (layer0_outputs(205));
    layer1_outputs(10226) <= not((layer0_outputs(4743)) and (layer0_outputs(2461)));
    layer1_outputs(10227) <= not(layer0_outputs(6516));
    layer1_outputs(10228) <= layer0_outputs(7843);
    layer1_outputs(10229) <= layer0_outputs(4437);
    layer1_outputs(10230) <= (layer0_outputs(5914)) xor (layer0_outputs(2076));
    layer1_outputs(10231) <= not(layer0_outputs(5305)) or (layer0_outputs(4725));
    layer1_outputs(10232) <= layer0_outputs(7039);
    layer1_outputs(10233) <= layer0_outputs(8375);
    layer1_outputs(10234) <= not((layer0_outputs(4302)) xor (layer0_outputs(4987)));
    layer1_outputs(10235) <= not((layer0_outputs(746)) or (layer0_outputs(3009)));
    layer1_outputs(10236) <= not((layer0_outputs(503)) and (layer0_outputs(7722)));
    layer1_outputs(10237) <= not(layer0_outputs(6641)) or (layer0_outputs(7592));
    layer1_outputs(10238) <= not(layer0_outputs(4032));
    layer1_outputs(10239) <= not((layer0_outputs(786)) and (layer0_outputs(4608)));
    layer2_outputs(0) <= layer1_outputs(4968);
    layer2_outputs(1) <= layer1_outputs(7563);
    layer2_outputs(2) <= (layer1_outputs(325)) or (layer1_outputs(3006));
    layer2_outputs(3) <= (layer1_outputs(8653)) xor (layer1_outputs(1662));
    layer2_outputs(4) <= (layer1_outputs(3358)) xor (layer1_outputs(306));
    layer2_outputs(5) <= layer1_outputs(5247);
    layer2_outputs(6) <= layer1_outputs(5722);
    layer2_outputs(7) <= (layer1_outputs(6749)) and not (layer1_outputs(8465));
    layer2_outputs(8) <= not((layer1_outputs(7352)) and (layer1_outputs(9117)));
    layer2_outputs(9) <= layer1_outputs(7263);
    layer2_outputs(10) <= not(layer1_outputs(9712));
    layer2_outputs(11) <= not(layer1_outputs(10011)) or (layer1_outputs(2061));
    layer2_outputs(12) <= layer1_outputs(6778);
    layer2_outputs(13) <= not((layer1_outputs(7471)) xor (layer1_outputs(1704)));
    layer2_outputs(14) <= not(layer1_outputs(3897)) or (layer1_outputs(7067));
    layer2_outputs(15) <= layer1_outputs(8474);
    layer2_outputs(16) <= (layer1_outputs(6479)) and (layer1_outputs(6839));
    layer2_outputs(17) <= not(layer1_outputs(5676)) or (layer1_outputs(1807));
    layer2_outputs(18) <= not(layer1_outputs(4422));
    layer2_outputs(19) <= (layer1_outputs(3910)) and not (layer1_outputs(9711));
    layer2_outputs(20) <= not(layer1_outputs(612));
    layer2_outputs(21) <= (layer1_outputs(8414)) xor (layer1_outputs(6816));
    layer2_outputs(22) <= not(layer1_outputs(5857)) or (layer1_outputs(6310));
    layer2_outputs(23) <= not(layer1_outputs(6386));
    layer2_outputs(24) <= layer1_outputs(8106);
    layer2_outputs(25) <= not(layer1_outputs(5701));
    layer2_outputs(26) <= not(layer1_outputs(2085));
    layer2_outputs(27) <= layer1_outputs(5270);
    layer2_outputs(28) <= not(layer1_outputs(5873));
    layer2_outputs(29) <= (layer1_outputs(2810)) and not (layer1_outputs(3242));
    layer2_outputs(30) <= not((layer1_outputs(1606)) or (layer1_outputs(833)));
    layer2_outputs(31) <= not((layer1_outputs(7095)) and (layer1_outputs(6140)));
    layer2_outputs(32) <= (layer1_outputs(2290)) and not (layer1_outputs(10090));
    layer2_outputs(33) <= not(layer1_outputs(2230));
    layer2_outputs(34) <= layer1_outputs(5049);
    layer2_outputs(35) <= not((layer1_outputs(3179)) or (layer1_outputs(6296)));
    layer2_outputs(36) <= (layer1_outputs(1028)) and not (layer1_outputs(6077));
    layer2_outputs(37) <= not(layer1_outputs(5654));
    layer2_outputs(38) <= layer1_outputs(3025);
    layer2_outputs(39) <= not(layer1_outputs(7565));
    layer2_outputs(40) <= not(layer1_outputs(5133)) or (layer1_outputs(9445));
    layer2_outputs(41) <= layer1_outputs(3285);
    layer2_outputs(42) <= (layer1_outputs(4125)) xor (layer1_outputs(3559));
    layer2_outputs(43) <= layer1_outputs(7671);
    layer2_outputs(44) <= layer1_outputs(8839);
    layer2_outputs(45) <= layer1_outputs(9015);
    layer2_outputs(46) <= not(layer1_outputs(5605)) or (layer1_outputs(468));
    layer2_outputs(47) <= (layer1_outputs(5790)) xor (layer1_outputs(8613));
    layer2_outputs(48) <= (layer1_outputs(9768)) and (layer1_outputs(9189));
    layer2_outputs(49) <= '1';
    layer2_outputs(50) <= layer1_outputs(3211);
    layer2_outputs(51) <= layer1_outputs(1579);
    layer2_outputs(52) <= (layer1_outputs(8471)) and not (layer1_outputs(4190));
    layer2_outputs(53) <= not(layer1_outputs(6560));
    layer2_outputs(54) <= not(layer1_outputs(9730)) or (layer1_outputs(6579));
    layer2_outputs(55) <= (layer1_outputs(5105)) xor (layer1_outputs(9510));
    layer2_outputs(56) <= (layer1_outputs(8226)) or (layer1_outputs(8755));
    layer2_outputs(57) <= layer1_outputs(906);
    layer2_outputs(58) <= not((layer1_outputs(8170)) xor (layer1_outputs(8483)));
    layer2_outputs(59) <= (layer1_outputs(4962)) and not (layer1_outputs(4470));
    layer2_outputs(60) <= layer1_outputs(3542);
    layer2_outputs(61) <= not(layer1_outputs(7972));
    layer2_outputs(62) <= not((layer1_outputs(2068)) xor (layer1_outputs(2430)));
    layer2_outputs(63) <= not(layer1_outputs(7108));
    layer2_outputs(64) <= (layer1_outputs(1599)) and (layer1_outputs(8081));
    layer2_outputs(65) <= layer1_outputs(6918);
    layer2_outputs(66) <= layer1_outputs(6917);
    layer2_outputs(67) <= layer1_outputs(477);
    layer2_outputs(68) <= (layer1_outputs(2584)) or (layer1_outputs(2084));
    layer2_outputs(69) <= (layer1_outputs(6544)) and not (layer1_outputs(3267));
    layer2_outputs(70) <= layer1_outputs(8938);
    layer2_outputs(71) <= not(layer1_outputs(3833)) or (layer1_outputs(8249));
    layer2_outputs(72) <= not(layer1_outputs(1166));
    layer2_outputs(73) <= (layer1_outputs(6221)) xor (layer1_outputs(8773));
    layer2_outputs(74) <= layer1_outputs(9532);
    layer2_outputs(75) <= not((layer1_outputs(6167)) and (layer1_outputs(1689)));
    layer2_outputs(76) <= not(layer1_outputs(9769));
    layer2_outputs(77) <= not(layer1_outputs(10000));
    layer2_outputs(78) <= layer1_outputs(5852);
    layer2_outputs(79) <= not(layer1_outputs(9367));
    layer2_outputs(80) <= (layer1_outputs(3203)) xor (layer1_outputs(1844));
    layer2_outputs(81) <= (layer1_outputs(4365)) and not (layer1_outputs(7466));
    layer2_outputs(82) <= layer1_outputs(4847);
    layer2_outputs(83) <= (layer1_outputs(6846)) and not (layer1_outputs(3729));
    layer2_outputs(84) <= layer1_outputs(9224);
    layer2_outputs(85) <= not(layer1_outputs(4139));
    layer2_outputs(86) <= layer1_outputs(3801);
    layer2_outputs(87) <= not(layer1_outputs(9646)) or (layer1_outputs(2447));
    layer2_outputs(88) <= not(layer1_outputs(6160)) or (layer1_outputs(2553));
    layer2_outputs(89) <= not((layer1_outputs(3687)) or (layer1_outputs(6952)));
    layer2_outputs(90) <= not(layer1_outputs(904)) or (layer1_outputs(2957));
    layer2_outputs(91) <= not((layer1_outputs(10182)) and (layer1_outputs(2298)));
    layer2_outputs(92) <= layer1_outputs(411);
    layer2_outputs(93) <= layer1_outputs(5833);
    layer2_outputs(94) <= not(layer1_outputs(5025));
    layer2_outputs(95) <= not((layer1_outputs(9056)) and (layer1_outputs(572)));
    layer2_outputs(96) <= (layer1_outputs(10227)) and not (layer1_outputs(6970));
    layer2_outputs(97) <= not(layer1_outputs(9818));
    layer2_outputs(98) <= layer1_outputs(4854);
    layer2_outputs(99) <= (layer1_outputs(8875)) or (layer1_outputs(5579));
    layer2_outputs(100) <= not((layer1_outputs(5086)) and (layer1_outputs(9340)));
    layer2_outputs(101) <= layer1_outputs(3514);
    layer2_outputs(102) <= (layer1_outputs(8520)) or (layer1_outputs(4790));
    layer2_outputs(103) <= not(layer1_outputs(222)) or (layer1_outputs(465));
    layer2_outputs(104) <= (layer1_outputs(9017)) and not (layer1_outputs(6235));
    layer2_outputs(105) <= layer1_outputs(3826);
    layer2_outputs(106) <= layer1_outputs(9650);
    layer2_outputs(107) <= not((layer1_outputs(6955)) xor (layer1_outputs(488)));
    layer2_outputs(108) <= not(layer1_outputs(6386));
    layer2_outputs(109) <= layer1_outputs(8618);
    layer2_outputs(110) <= not((layer1_outputs(8518)) or (layer1_outputs(10025)));
    layer2_outputs(111) <= not(layer1_outputs(1326));
    layer2_outputs(112) <= layer1_outputs(1246);
    layer2_outputs(113) <= not(layer1_outputs(5246));
    layer2_outputs(114) <= not(layer1_outputs(2767));
    layer2_outputs(115) <= not((layer1_outputs(8298)) and (layer1_outputs(10063)));
    layer2_outputs(116) <= (layer1_outputs(165)) and not (layer1_outputs(8195));
    layer2_outputs(117) <= not(layer1_outputs(7697));
    layer2_outputs(118) <= not(layer1_outputs(8319));
    layer2_outputs(119) <= '0';
    layer2_outputs(120) <= layer1_outputs(7794);
    layer2_outputs(121) <= '0';
    layer2_outputs(122) <= not(layer1_outputs(2934));
    layer2_outputs(123) <= not(layer1_outputs(602));
    layer2_outputs(124) <= layer1_outputs(6024);
    layer2_outputs(125) <= (layer1_outputs(940)) xor (layer1_outputs(1601));
    layer2_outputs(126) <= not(layer1_outputs(3703));
    layer2_outputs(127) <= (layer1_outputs(51)) and not (layer1_outputs(8797));
    layer2_outputs(128) <= not(layer1_outputs(8614)) or (layer1_outputs(9147));
    layer2_outputs(129) <= not(layer1_outputs(328));
    layer2_outputs(130) <= layer1_outputs(6770);
    layer2_outputs(131) <= not(layer1_outputs(10023)) or (layer1_outputs(2433));
    layer2_outputs(132) <= not(layer1_outputs(9919));
    layer2_outputs(133) <= not(layer1_outputs(7336)) or (layer1_outputs(2465));
    layer2_outputs(134) <= '1';
    layer2_outputs(135) <= layer1_outputs(4775);
    layer2_outputs(136) <= not(layer1_outputs(7342)) or (layer1_outputs(5471));
    layer2_outputs(137) <= not(layer1_outputs(1409));
    layer2_outputs(138) <= (layer1_outputs(9532)) or (layer1_outputs(84));
    layer2_outputs(139) <= not(layer1_outputs(2406));
    layer2_outputs(140) <= not(layer1_outputs(7556));
    layer2_outputs(141) <= (layer1_outputs(6837)) xor (layer1_outputs(9720));
    layer2_outputs(142) <= (layer1_outputs(1824)) and not (layer1_outputs(7007));
    layer2_outputs(143) <= (layer1_outputs(2472)) and not (layer1_outputs(7860));
    layer2_outputs(144) <= (layer1_outputs(9804)) xor (layer1_outputs(5769));
    layer2_outputs(145) <= layer1_outputs(9201);
    layer2_outputs(146) <= not(layer1_outputs(7494));
    layer2_outputs(147) <= '0';
    layer2_outputs(148) <= layer1_outputs(9758);
    layer2_outputs(149) <= not(layer1_outputs(9524)) or (layer1_outputs(1001));
    layer2_outputs(150) <= (layer1_outputs(5265)) xor (layer1_outputs(1842));
    layer2_outputs(151) <= layer1_outputs(231);
    layer2_outputs(152) <= (layer1_outputs(4456)) and (layer1_outputs(2964));
    layer2_outputs(153) <= not(layer1_outputs(7051));
    layer2_outputs(154) <= not(layer1_outputs(4575));
    layer2_outputs(155) <= layer1_outputs(5929);
    layer2_outputs(156) <= (layer1_outputs(8320)) xor (layer1_outputs(5384));
    layer2_outputs(157) <= not(layer1_outputs(3428));
    layer2_outputs(158) <= not(layer1_outputs(7789));
    layer2_outputs(159) <= layer1_outputs(5800);
    layer2_outputs(160) <= not(layer1_outputs(6334));
    layer2_outputs(161) <= layer1_outputs(2505);
    layer2_outputs(162) <= not(layer1_outputs(3936));
    layer2_outputs(163) <= not(layer1_outputs(8862));
    layer2_outputs(164) <= not(layer1_outputs(7075));
    layer2_outputs(165) <= not(layer1_outputs(1201));
    layer2_outputs(166) <= layer1_outputs(8289);
    layer2_outputs(167) <= not((layer1_outputs(6292)) or (layer1_outputs(2350)));
    layer2_outputs(168) <= not(layer1_outputs(1983));
    layer2_outputs(169) <= (layer1_outputs(8500)) xor (layer1_outputs(8470));
    layer2_outputs(170) <= not(layer1_outputs(4760));
    layer2_outputs(171) <= layer1_outputs(1335);
    layer2_outputs(172) <= layer1_outputs(626);
    layer2_outputs(173) <= (layer1_outputs(2510)) and not (layer1_outputs(7970));
    layer2_outputs(174) <= not(layer1_outputs(9374)) or (layer1_outputs(8604));
    layer2_outputs(175) <= not((layer1_outputs(7537)) xor (layer1_outputs(9217)));
    layer2_outputs(176) <= not(layer1_outputs(1849));
    layer2_outputs(177) <= not(layer1_outputs(4950));
    layer2_outputs(178) <= '0';
    layer2_outputs(179) <= layer1_outputs(4205);
    layer2_outputs(180) <= layer1_outputs(6205);
    layer2_outputs(181) <= not(layer1_outputs(9326));
    layer2_outputs(182) <= not(layer1_outputs(4527));
    layer2_outputs(183) <= not((layer1_outputs(9620)) xor (layer1_outputs(1167)));
    layer2_outputs(184) <= (layer1_outputs(5747)) or (layer1_outputs(2569));
    layer2_outputs(185) <= layer1_outputs(2281);
    layer2_outputs(186) <= (layer1_outputs(1717)) and not (layer1_outputs(6433));
    layer2_outputs(187) <= layer1_outputs(3739);
    layer2_outputs(188) <= layer1_outputs(3127);
    layer2_outputs(189) <= not((layer1_outputs(10009)) or (layer1_outputs(8125)));
    layer2_outputs(190) <= (layer1_outputs(9840)) or (layer1_outputs(2973));
    layer2_outputs(191) <= layer1_outputs(733);
    layer2_outputs(192) <= not(layer1_outputs(9687)) or (layer1_outputs(6454));
    layer2_outputs(193) <= layer1_outputs(8684);
    layer2_outputs(194) <= not((layer1_outputs(9564)) or (layer1_outputs(8906)));
    layer2_outputs(195) <= not(layer1_outputs(7105)) or (layer1_outputs(7001));
    layer2_outputs(196) <= layer1_outputs(5137);
    layer2_outputs(197) <= (layer1_outputs(7833)) xor (layer1_outputs(6640));
    layer2_outputs(198) <= not(layer1_outputs(9955)) or (layer1_outputs(2879));
    layer2_outputs(199) <= not(layer1_outputs(1256));
    layer2_outputs(200) <= not(layer1_outputs(2867)) or (layer1_outputs(5415));
    layer2_outputs(201) <= not(layer1_outputs(3072));
    layer2_outputs(202) <= layer1_outputs(6866);
    layer2_outputs(203) <= layer1_outputs(2514);
    layer2_outputs(204) <= layer1_outputs(10074);
    layer2_outputs(205) <= not((layer1_outputs(8465)) xor (layer1_outputs(3743)));
    layer2_outputs(206) <= not(layer1_outputs(9139)) or (layer1_outputs(1721));
    layer2_outputs(207) <= layer1_outputs(7474);
    layer2_outputs(208) <= not(layer1_outputs(2248));
    layer2_outputs(209) <= layer1_outputs(7469);
    layer2_outputs(210) <= not(layer1_outputs(6775)) or (layer1_outputs(9659));
    layer2_outputs(211) <= not((layer1_outputs(8498)) and (layer1_outputs(451)));
    layer2_outputs(212) <= not(layer1_outputs(1842));
    layer2_outputs(213) <= (layer1_outputs(4795)) and not (layer1_outputs(7224));
    layer2_outputs(214) <= layer1_outputs(10078);
    layer2_outputs(215) <= layer1_outputs(1995);
    layer2_outputs(216) <= not(layer1_outputs(6962));
    layer2_outputs(217) <= not((layer1_outputs(4447)) or (layer1_outputs(7719)));
    layer2_outputs(218) <= not(layer1_outputs(4314));
    layer2_outputs(219) <= layer1_outputs(6350);
    layer2_outputs(220) <= layer1_outputs(5569);
    layer2_outputs(221) <= not((layer1_outputs(7366)) xor (layer1_outputs(2790)));
    layer2_outputs(222) <= layer1_outputs(1586);
    layer2_outputs(223) <= not(layer1_outputs(10117));
    layer2_outputs(224) <= not((layer1_outputs(3832)) xor (layer1_outputs(10202)));
    layer2_outputs(225) <= layer1_outputs(8531);
    layer2_outputs(226) <= not(layer1_outputs(467));
    layer2_outputs(227) <= (layer1_outputs(3089)) xor (layer1_outputs(2446));
    layer2_outputs(228) <= (layer1_outputs(3171)) and not (layer1_outputs(3091));
    layer2_outputs(229) <= not((layer1_outputs(8488)) or (layer1_outputs(9029)));
    layer2_outputs(230) <= not(layer1_outputs(5313));
    layer2_outputs(231) <= layer1_outputs(4045);
    layer2_outputs(232) <= layer1_outputs(5578);
    layer2_outputs(233) <= not(layer1_outputs(6672));
    layer2_outputs(234) <= (layer1_outputs(6420)) and not (layer1_outputs(380));
    layer2_outputs(235) <= not((layer1_outputs(9773)) xor (layer1_outputs(2649)));
    layer2_outputs(236) <= '0';
    layer2_outputs(237) <= layer1_outputs(6613);
    layer2_outputs(238) <= (layer1_outputs(5319)) xor (layer1_outputs(3825));
    layer2_outputs(239) <= layer1_outputs(4607);
    layer2_outputs(240) <= layer1_outputs(5981);
    layer2_outputs(241) <= layer1_outputs(4693);
    layer2_outputs(242) <= layer1_outputs(994);
    layer2_outputs(243) <= not(layer1_outputs(2424));
    layer2_outputs(244) <= not(layer1_outputs(7819));
    layer2_outputs(245) <= (layer1_outputs(2240)) and not (layer1_outputs(3013));
    layer2_outputs(246) <= not(layer1_outputs(1796)) or (layer1_outputs(2158));
    layer2_outputs(247) <= not(layer1_outputs(5481));
    layer2_outputs(248) <= not(layer1_outputs(9468));
    layer2_outputs(249) <= not((layer1_outputs(10017)) or (layer1_outputs(1540)));
    layer2_outputs(250) <= layer1_outputs(6443);
    layer2_outputs(251) <= (layer1_outputs(6032)) and (layer1_outputs(7539));
    layer2_outputs(252) <= layer1_outputs(6711);
    layer2_outputs(253) <= (layer1_outputs(9201)) and not (layer1_outputs(4739));
    layer2_outputs(254) <= layer1_outputs(4017);
    layer2_outputs(255) <= layer1_outputs(6776);
    layer2_outputs(256) <= not(layer1_outputs(2601)) or (layer1_outputs(2009));
    layer2_outputs(257) <= not(layer1_outputs(9202));
    layer2_outputs(258) <= layer1_outputs(265);
    layer2_outputs(259) <= (layer1_outputs(2142)) and not (layer1_outputs(2073));
    layer2_outputs(260) <= not(layer1_outputs(706));
    layer2_outputs(261) <= not((layer1_outputs(1535)) or (layer1_outputs(4690)));
    layer2_outputs(262) <= layer1_outputs(2057);
    layer2_outputs(263) <= (layer1_outputs(3558)) and not (layer1_outputs(4354));
    layer2_outputs(264) <= layer1_outputs(7524);
    layer2_outputs(265) <= (layer1_outputs(5919)) or (layer1_outputs(353));
    layer2_outputs(266) <= not(layer1_outputs(417));
    layer2_outputs(267) <= layer1_outputs(1822);
    layer2_outputs(268) <= not(layer1_outputs(10049)) or (layer1_outputs(4050));
    layer2_outputs(269) <= layer1_outputs(2572);
    layer2_outputs(270) <= not(layer1_outputs(3917));
    layer2_outputs(271) <= not(layer1_outputs(9036));
    layer2_outputs(272) <= layer1_outputs(5407);
    layer2_outputs(273) <= not(layer1_outputs(8457));
    layer2_outputs(274) <= not(layer1_outputs(5492));
    layer2_outputs(275) <= (layer1_outputs(3383)) or (layer1_outputs(3855));
    layer2_outputs(276) <= layer1_outputs(5201);
    layer2_outputs(277) <= not(layer1_outputs(9050));
    layer2_outputs(278) <= not(layer1_outputs(9618));
    layer2_outputs(279) <= not(layer1_outputs(281));
    layer2_outputs(280) <= not(layer1_outputs(9631));
    layer2_outputs(281) <= (layer1_outputs(3953)) and (layer1_outputs(717));
    layer2_outputs(282) <= not((layer1_outputs(8203)) and (layer1_outputs(9475)));
    layer2_outputs(283) <= layer1_outputs(9);
    layer2_outputs(284) <= not(layer1_outputs(9961)) or (layer1_outputs(2082));
    layer2_outputs(285) <= layer1_outputs(10172);
    layer2_outputs(286) <= layer1_outputs(8192);
    layer2_outputs(287) <= layer1_outputs(5404);
    layer2_outputs(288) <= layer1_outputs(1702);
    layer2_outputs(289) <= layer1_outputs(3096);
    layer2_outputs(290) <= not(layer1_outputs(7191)) or (layer1_outputs(10055));
    layer2_outputs(291) <= (layer1_outputs(5443)) xor (layer1_outputs(3627));
    layer2_outputs(292) <= not(layer1_outputs(5264));
    layer2_outputs(293) <= (layer1_outputs(2084)) and not (layer1_outputs(8821));
    layer2_outputs(294) <= not(layer1_outputs(2938));
    layer2_outputs(295) <= not(layer1_outputs(10124));
    layer2_outputs(296) <= (layer1_outputs(5755)) xor (layer1_outputs(5339));
    layer2_outputs(297) <= layer1_outputs(1475);
    layer2_outputs(298) <= layer1_outputs(7449);
    layer2_outputs(299) <= not(layer1_outputs(9840));
    layer2_outputs(300) <= not((layer1_outputs(6106)) and (layer1_outputs(7954)));
    layer2_outputs(301) <= not(layer1_outputs(2717));
    layer2_outputs(302) <= (layer1_outputs(3410)) xor (layer1_outputs(6624));
    layer2_outputs(303) <= (layer1_outputs(1423)) and (layer1_outputs(4833));
    layer2_outputs(304) <= not((layer1_outputs(9531)) or (layer1_outputs(249)));
    layer2_outputs(305) <= not(layer1_outputs(4307));
    layer2_outputs(306) <= not(layer1_outputs(1588)) or (layer1_outputs(494));
    layer2_outputs(307) <= (layer1_outputs(9798)) and not (layer1_outputs(1921));
    layer2_outputs(308) <= (layer1_outputs(4518)) and (layer1_outputs(7520));
    layer2_outputs(309) <= not(layer1_outputs(2558)) or (layer1_outputs(2194));
    layer2_outputs(310) <= not((layer1_outputs(5054)) xor (layer1_outputs(1859)));
    layer2_outputs(311) <= layer1_outputs(3708);
    layer2_outputs(312) <= (layer1_outputs(9358)) xor (layer1_outputs(2731));
    layer2_outputs(313) <= layer1_outputs(747);
    layer2_outputs(314) <= layer1_outputs(100);
    layer2_outputs(315) <= not((layer1_outputs(7312)) and (layer1_outputs(9387)));
    layer2_outputs(316) <= (layer1_outputs(7850)) xor (layer1_outputs(1323));
    layer2_outputs(317) <= not(layer1_outputs(3514));
    layer2_outputs(318) <= not(layer1_outputs(5161));
    layer2_outputs(319) <= not((layer1_outputs(1181)) or (layer1_outputs(6064)));
    layer2_outputs(320) <= layer1_outputs(2449);
    layer2_outputs(321) <= not(layer1_outputs(5017));
    layer2_outputs(322) <= not(layer1_outputs(8970));
    layer2_outputs(323) <= layer1_outputs(3343);
    layer2_outputs(324) <= not((layer1_outputs(163)) or (layer1_outputs(120)));
    layer2_outputs(325) <= layer1_outputs(2856);
    layer2_outputs(326) <= not(layer1_outputs(425));
    layer2_outputs(327) <= not((layer1_outputs(4355)) xor (layer1_outputs(7391)));
    layer2_outputs(328) <= layer1_outputs(9872);
    layer2_outputs(329) <= not(layer1_outputs(7939));
    layer2_outputs(330) <= (layer1_outputs(6096)) and not (layer1_outputs(6028));
    layer2_outputs(331) <= layer1_outputs(9425);
    layer2_outputs(332) <= not((layer1_outputs(9442)) xor (layer1_outputs(10239)));
    layer2_outputs(333) <= layer1_outputs(5117);
    layer2_outputs(334) <= not(layer1_outputs(3301));
    layer2_outputs(335) <= layer1_outputs(654);
    layer2_outputs(336) <= (layer1_outputs(2952)) and not (layer1_outputs(3790));
    layer2_outputs(337) <= (layer1_outputs(4700)) and not (layer1_outputs(8954));
    layer2_outputs(338) <= (layer1_outputs(7819)) and not (layer1_outputs(2393));
    layer2_outputs(339) <= layer1_outputs(1974);
    layer2_outputs(340) <= layer1_outputs(315);
    layer2_outputs(341) <= (layer1_outputs(6700)) or (layer1_outputs(3651));
    layer2_outputs(342) <= (layer1_outputs(8442)) xor (layer1_outputs(8750));
    layer2_outputs(343) <= (layer1_outputs(3216)) and not (layer1_outputs(5678));
    layer2_outputs(344) <= not((layer1_outputs(1445)) xor (layer1_outputs(5649)));
    layer2_outputs(345) <= not(layer1_outputs(1674));
    layer2_outputs(346) <= not(layer1_outputs(8817)) or (layer1_outputs(5587));
    layer2_outputs(347) <= not(layer1_outputs(2365));
    layer2_outputs(348) <= not(layer1_outputs(7736));
    layer2_outputs(349) <= layer1_outputs(9458);
    layer2_outputs(350) <= not((layer1_outputs(4758)) xor (layer1_outputs(4312)));
    layer2_outputs(351) <= not((layer1_outputs(2048)) xor (layer1_outputs(9934)));
    layer2_outputs(352) <= not(layer1_outputs(1979)) or (layer1_outputs(2635));
    layer2_outputs(353) <= not(layer1_outputs(7338));
    layer2_outputs(354) <= layer1_outputs(6865);
    layer2_outputs(355) <= layer1_outputs(4732);
    layer2_outputs(356) <= layer1_outputs(9510);
    layer2_outputs(357) <= layer1_outputs(3314);
    layer2_outputs(358) <= layer1_outputs(4294);
    layer2_outputs(359) <= layer1_outputs(7245);
    layer2_outputs(360) <= not((layer1_outputs(10225)) or (layer1_outputs(8704)));
    layer2_outputs(361) <= not(layer1_outputs(327));
    layer2_outputs(362) <= not(layer1_outputs(3065)) or (layer1_outputs(10135));
    layer2_outputs(363) <= not(layer1_outputs(6849));
    layer2_outputs(364) <= (layer1_outputs(10130)) and not (layer1_outputs(2815));
    layer2_outputs(365) <= (layer1_outputs(6984)) and not (layer1_outputs(1558));
    layer2_outputs(366) <= not(layer1_outputs(6868));
    layer2_outputs(367) <= layer1_outputs(835);
    layer2_outputs(368) <= (layer1_outputs(3279)) and (layer1_outputs(7476));
    layer2_outputs(369) <= not(layer1_outputs(2644)) or (layer1_outputs(5964));
    layer2_outputs(370) <= layer1_outputs(4526);
    layer2_outputs(371) <= not(layer1_outputs(5833));
    layer2_outputs(372) <= layer1_outputs(10024);
    layer2_outputs(373) <= layer1_outputs(5725);
    layer2_outputs(374) <= layer1_outputs(1973);
    layer2_outputs(375) <= layer1_outputs(5412);
    layer2_outputs(376) <= (layer1_outputs(6357)) and (layer1_outputs(550));
    layer2_outputs(377) <= not(layer1_outputs(9548));
    layer2_outputs(378) <= not((layer1_outputs(8400)) or (layer1_outputs(9596)));
    layer2_outputs(379) <= (layer1_outputs(9084)) and not (layer1_outputs(6298));
    layer2_outputs(380) <= not(layer1_outputs(5102));
    layer2_outputs(381) <= not((layer1_outputs(1204)) or (layer1_outputs(558)));
    layer2_outputs(382) <= layer1_outputs(3958);
    layer2_outputs(383) <= layer1_outputs(73);
    layer2_outputs(384) <= layer1_outputs(1251);
    layer2_outputs(385) <= not(layer1_outputs(3935));
    layer2_outputs(386) <= not(layer1_outputs(10217)) or (layer1_outputs(1840));
    layer2_outputs(387) <= not(layer1_outputs(4642));
    layer2_outputs(388) <= (layer1_outputs(4036)) and not (layer1_outputs(8385));
    layer2_outputs(389) <= not(layer1_outputs(4930));
    layer2_outputs(390) <= not(layer1_outputs(4977));
    layer2_outputs(391) <= not((layer1_outputs(1015)) or (layer1_outputs(9166)));
    layer2_outputs(392) <= (layer1_outputs(5492)) or (layer1_outputs(8544));
    layer2_outputs(393) <= not(layer1_outputs(5747));
    layer2_outputs(394) <= not(layer1_outputs(4948));
    layer2_outputs(395) <= layer1_outputs(4484);
    layer2_outputs(396) <= layer1_outputs(625);
    layer2_outputs(397) <= not(layer1_outputs(1668));
    layer2_outputs(398) <= (layer1_outputs(4519)) or (layer1_outputs(874));
    layer2_outputs(399) <= layer1_outputs(9855);
    layer2_outputs(400) <= (layer1_outputs(1929)) xor (layer1_outputs(1104));
    layer2_outputs(401) <= (layer1_outputs(4143)) xor (layer1_outputs(4871));
    layer2_outputs(402) <= not((layer1_outputs(5513)) xor (layer1_outputs(1683)));
    layer2_outputs(403) <= (layer1_outputs(8651)) and not (layer1_outputs(1246));
    layer2_outputs(404) <= not(layer1_outputs(6291));
    layer2_outputs(405) <= layer1_outputs(5232);
    layer2_outputs(406) <= not(layer1_outputs(8141));
    layer2_outputs(407) <= layer1_outputs(4336);
    layer2_outputs(408) <= layer1_outputs(292);
    layer2_outputs(409) <= not(layer1_outputs(6574)) or (layer1_outputs(7021));
    layer2_outputs(410) <= layer1_outputs(1353);
    layer2_outputs(411) <= layer1_outputs(7585);
    layer2_outputs(412) <= not((layer1_outputs(5118)) xor (layer1_outputs(7452)));
    layer2_outputs(413) <= layer1_outputs(2835);
    layer2_outputs(414) <= not((layer1_outputs(3255)) xor (layer1_outputs(5291)));
    layer2_outputs(415) <= (layer1_outputs(214)) and not (layer1_outputs(2804));
    layer2_outputs(416) <= not(layer1_outputs(7960)) or (layer1_outputs(1391));
    layer2_outputs(417) <= not(layer1_outputs(9068));
    layer2_outputs(418) <= layer1_outputs(2716);
    layer2_outputs(419) <= (layer1_outputs(6491)) xor (layer1_outputs(1159));
    layer2_outputs(420) <= not((layer1_outputs(4102)) or (layer1_outputs(6904)));
    layer2_outputs(421) <= not((layer1_outputs(9770)) or (layer1_outputs(1997)));
    layer2_outputs(422) <= not((layer1_outputs(790)) or (layer1_outputs(2218)));
    layer2_outputs(423) <= layer1_outputs(2822);
    layer2_outputs(424) <= not(layer1_outputs(3485));
    layer2_outputs(425) <= '1';
    layer2_outputs(426) <= layer1_outputs(9031);
    layer2_outputs(427) <= not(layer1_outputs(5437));
    layer2_outputs(428) <= not(layer1_outputs(1300));
    layer2_outputs(429) <= layer1_outputs(2755);
    layer2_outputs(430) <= not(layer1_outputs(9288)) or (layer1_outputs(7991));
    layer2_outputs(431) <= not(layer1_outputs(4358));
    layer2_outputs(432) <= not(layer1_outputs(4303));
    layer2_outputs(433) <= not(layer1_outputs(582));
    layer2_outputs(434) <= not(layer1_outputs(6903)) or (layer1_outputs(10228));
    layer2_outputs(435) <= layer1_outputs(2266);
    layer2_outputs(436) <= layer1_outputs(1032);
    layer2_outputs(437) <= not(layer1_outputs(6872));
    layer2_outputs(438) <= layer1_outputs(7329);
    layer2_outputs(439) <= not(layer1_outputs(6328));
    layer2_outputs(440) <= not(layer1_outputs(1933));
    layer2_outputs(441) <= (layer1_outputs(2055)) xor (layer1_outputs(721));
    layer2_outputs(442) <= not(layer1_outputs(6356));
    layer2_outputs(443) <= (layer1_outputs(4696)) or (layer1_outputs(4778));
    layer2_outputs(444) <= not(layer1_outputs(9678));
    layer2_outputs(445) <= (layer1_outputs(1105)) and not (layer1_outputs(360));
    layer2_outputs(446) <= (layer1_outputs(9217)) and not (layer1_outputs(1434));
    layer2_outputs(447) <= layer1_outputs(344);
    layer2_outputs(448) <= not((layer1_outputs(4582)) xor (layer1_outputs(1808)));
    layer2_outputs(449) <= layer1_outputs(378);
    layer2_outputs(450) <= not(layer1_outputs(3557));
    layer2_outputs(451) <= (layer1_outputs(4813)) xor (layer1_outputs(6397));
    layer2_outputs(452) <= layer1_outputs(6566);
    layer2_outputs(453) <= (layer1_outputs(7977)) or (layer1_outputs(4971));
    layer2_outputs(454) <= layer1_outputs(8036);
    layer2_outputs(455) <= (layer1_outputs(571)) or (layer1_outputs(164));
    layer2_outputs(456) <= not((layer1_outputs(7838)) xor (layer1_outputs(4601)));
    layer2_outputs(457) <= layer1_outputs(2307);
    layer2_outputs(458) <= not(layer1_outputs(10200));
    layer2_outputs(459) <= (layer1_outputs(3120)) and not (layer1_outputs(9998));
    layer2_outputs(460) <= not(layer1_outputs(6591));
    layer2_outputs(461) <= layer1_outputs(9059);
    layer2_outputs(462) <= not((layer1_outputs(6265)) xor (layer1_outputs(2705)));
    layer2_outputs(463) <= not(layer1_outputs(7608));
    layer2_outputs(464) <= layer1_outputs(2609);
    layer2_outputs(465) <= layer1_outputs(147);
    layer2_outputs(466) <= not(layer1_outputs(4181));
    layer2_outputs(467) <= not((layer1_outputs(9379)) or (layer1_outputs(5430)));
    layer2_outputs(468) <= not((layer1_outputs(9343)) xor (layer1_outputs(3098)));
    layer2_outputs(469) <= not(layer1_outputs(3721));
    layer2_outputs(470) <= not((layer1_outputs(3181)) xor (layer1_outputs(5561)));
    layer2_outputs(471) <= not(layer1_outputs(6660));
    layer2_outputs(472) <= (layer1_outputs(556)) xor (layer1_outputs(3018));
    layer2_outputs(473) <= not(layer1_outputs(8569));
    layer2_outputs(474) <= layer1_outputs(7109);
    layer2_outputs(475) <= (layer1_outputs(422)) xor (layer1_outputs(3880));
    layer2_outputs(476) <= (layer1_outputs(4629)) xor (layer1_outputs(1035));
    layer2_outputs(477) <= not(layer1_outputs(7776));
    layer2_outputs(478) <= not((layer1_outputs(1452)) or (layer1_outputs(10058)));
    layer2_outputs(479) <= layer1_outputs(9753);
    layer2_outputs(480) <= layer1_outputs(8426);
    layer2_outputs(481) <= layer1_outputs(4221);
    layer2_outputs(482) <= not(layer1_outputs(7233));
    layer2_outputs(483) <= layer1_outputs(1330);
    layer2_outputs(484) <= not(layer1_outputs(1431)) or (layer1_outputs(1099));
    layer2_outputs(485) <= not((layer1_outputs(285)) and (layer1_outputs(7460)));
    layer2_outputs(486) <= not(layer1_outputs(6704));
    layer2_outputs(487) <= not(layer1_outputs(7853));
    layer2_outputs(488) <= not(layer1_outputs(9467));
    layer2_outputs(489) <= not((layer1_outputs(9563)) or (layer1_outputs(2959)));
    layer2_outputs(490) <= not(layer1_outputs(954));
    layer2_outputs(491) <= not(layer1_outputs(934));
    layer2_outputs(492) <= (layer1_outputs(3341)) or (layer1_outputs(885));
    layer2_outputs(493) <= not(layer1_outputs(4767));
    layer2_outputs(494) <= not(layer1_outputs(4725));
    layer2_outputs(495) <= (layer1_outputs(6398)) or (layer1_outputs(5501));
    layer2_outputs(496) <= layer1_outputs(7249);
    layer2_outputs(497) <= layer1_outputs(7220);
    layer2_outputs(498) <= not(layer1_outputs(8029)) or (layer1_outputs(9252));
    layer2_outputs(499) <= not(layer1_outputs(969)) or (layer1_outputs(5736));
    layer2_outputs(500) <= (layer1_outputs(9449)) xor (layer1_outputs(6298));
    layer2_outputs(501) <= not((layer1_outputs(3312)) and (layer1_outputs(779)));
    layer2_outputs(502) <= not(layer1_outputs(7032));
    layer2_outputs(503) <= (layer1_outputs(3636)) and not (layer1_outputs(6300));
    layer2_outputs(504) <= layer1_outputs(8263);
    layer2_outputs(505) <= not(layer1_outputs(419));
    layer2_outputs(506) <= layer1_outputs(5748);
    layer2_outputs(507) <= (layer1_outputs(6252)) or (layer1_outputs(551));
    layer2_outputs(508) <= layer1_outputs(9039);
    layer2_outputs(509) <= not((layer1_outputs(447)) or (layer1_outputs(3618)));
    layer2_outputs(510) <= not(layer1_outputs(3378)) or (layer1_outputs(2318));
    layer2_outputs(511) <= not(layer1_outputs(3798)) or (layer1_outputs(8050));
    layer2_outputs(512) <= not(layer1_outputs(1913));
    layer2_outputs(513) <= not(layer1_outputs(9799));
    layer2_outputs(514) <= not((layer1_outputs(5862)) xor (layer1_outputs(8527)));
    layer2_outputs(515) <= not((layer1_outputs(9070)) or (layer1_outputs(9951)));
    layer2_outputs(516) <= layer1_outputs(2323);
    layer2_outputs(517) <= (layer1_outputs(3907)) and not (layer1_outputs(7398));
    layer2_outputs(518) <= not(layer1_outputs(4488));
    layer2_outputs(519) <= layer1_outputs(371);
    layer2_outputs(520) <= layer1_outputs(5963);
    layer2_outputs(521) <= (layer1_outputs(7401)) xor (layer1_outputs(3616));
    layer2_outputs(522) <= not(layer1_outputs(9909)) or (layer1_outputs(4289));
    layer2_outputs(523) <= not(layer1_outputs(7063));
    layer2_outputs(524) <= layer1_outputs(3219);
    layer2_outputs(525) <= not(layer1_outputs(4746));
    layer2_outputs(526) <= '0';
    layer2_outputs(527) <= layer1_outputs(1458);
    layer2_outputs(528) <= (layer1_outputs(52)) and (layer1_outputs(9014));
    layer2_outputs(529) <= layer1_outputs(7966);
    layer2_outputs(530) <= (layer1_outputs(6085)) and not (layer1_outputs(5804));
    layer2_outputs(531) <= layer1_outputs(7887);
    layer2_outputs(532) <= layer1_outputs(6766);
    layer2_outputs(533) <= layer1_outputs(6005);
    layer2_outputs(534) <= not(layer1_outputs(6684)) or (layer1_outputs(1554));
    layer2_outputs(535) <= not(layer1_outputs(5537)) or (layer1_outputs(6902));
    layer2_outputs(536) <= layer1_outputs(1944);
    layer2_outputs(537) <= (layer1_outputs(3085)) xor (layer1_outputs(7865));
    layer2_outputs(538) <= layer1_outputs(7655);
    layer2_outputs(539) <= not(layer1_outputs(9891));
    layer2_outputs(540) <= layer1_outputs(5420);
    layer2_outputs(541) <= not(layer1_outputs(6994));
    layer2_outputs(542) <= not(layer1_outputs(587));
    layer2_outputs(543) <= layer1_outputs(46);
    layer2_outputs(544) <= not(layer1_outputs(1107));
    layer2_outputs(545) <= (layer1_outputs(103)) xor (layer1_outputs(6975));
    layer2_outputs(546) <= layer1_outputs(5409);
    layer2_outputs(547) <= not(layer1_outputs(5286));
    layer2_outputs(548) <= (layer1_outputs(6369)) and (layer1_outputs(6272));
    layer2_outputs(549) <= (layer1_outputs(4120)) and not (layer1_outputs(1659));
    layer2_outputs(550) <= (layer1_outputs(2003)) xor (layer1_outputs(3550));
    layer2_outputs(551) <= (layer1_outputs(7790)) xor (layer1_outputs(5284));
    layer2_outputs(552) <= not(layer1_outputs(5233));
    layer2_outputs(553) <= layer1_outputs(9400);
    layer2_outputs(554) <= not((layer1_outputs(2931)) xor (layer1_outputs(50)));
    layer2_outputs(555) <= not((layer1_outputs(10104)) or (layer1_outputs(7399)));
    layer2_outputs(556) <= (layer1_outputs(1517)) and not (layer1_outputs(9319));
    layer2_outputs(557) <= not(layer1_outputs(9657));
    layer2_outputs(558) <= (layer1_outputs(2596)) and not (layer1_outputs(6862));
    layer2_outputs(559) <= (layer1_outputs(3416)) or (layer1_outputs(3982));
    layer2_outputs(560) <= layer1_outputs(4689);
    layer2_outputs(561) <= not((layer1_outputs(664)) xor (layer1_outputs(2955)));
    layer2_outputs(562) <= not(layer1_outputs(9009)) or (layer1_outputs(8800));
    layer2_outputs(563) <= layer1_outputs(1190);
    layer2_outputs(564) <= layer1_outputs(8538);
    layer2_outputs(565) <= not(layer1_outputs(6326)) or (layer1_outputs(801));
    layer2_outputs(566) <= layer1_outputs(5478);
    layer2_outputs(567) <= layer1_outputs(8256);
    layer2_outputs(568) <= layer1_outputs(6351);
    layer2_outputs(569) <= not(layer1_outputs(811)) or (layer1_outputs(7803));
    layer2_outputs(570) <= not(layer1_outputs(8719)) or (layer1_outputs(6300));
    layer2_outputs(571) <= not((layer1_outputs(6073)) xor (layer1_outputs(3984)));
    layer2_outputs(572) <= not(layer1_outputs(203));
    layer2_outputs(573) <= (layer1_outputs(2862)) and not (layer1_outputs(6129));
    layer2_outputs(574) <= not(layer1_outputs(3951)) or (layer1_outputs(6229));
    layer2_outputs(575) <= not(layer1_outputs(145)) or (layer1_outputs(3315));
    layer2_outputs(576) <= layer1_outputs(5684);
    layer2_outputs(577) <= not(layer1_outputs(2138)) or (layer1_outputs(5039));
    layer2_outputs(578) <= '1';
    layer2_outputs(579) <= not(layer1_outputs(4292));
    layer2_outputs(580) <= not(layer1_outputs(3746));
    layer2_outputs(581) <= (layer1_outputs(9081)) or (layer1_outputs(7115));
    layer2_outputs(582) <= not((layer1_outputs(5181)) and (layer1_outputs(3792)));
    layer2_outputs(583) <= (layer1_outputs(3614)) and not (layer1_outputs(10081));
    layer2_outputs(584) <= layer1_outputs(4428);
    layer2_outputs(585) <= not(layer1_outputs(862)) or (layer1_outputs(2927));
    layer2_outputs(586) <= layer1_outputs(3912);
    layer2_outputs(587) <= layer1_outputs(6492);
    layer2_outputs(588) <= '1';
    layer2_outputs(589) <= not((layer1_outputs(3045)) or (layer1_outputs(5811)));
    layer2_outputs(590) <= not((layer1_outputs(4867)) and (layer1_outputs(1590)));
    layer2_outputs(591) <= not((layer1_outputs(6537)) xor (layer1_outputs(3804)));
    layer2_outputs(592) <= (layer1_outputs(8894)) and not (layer1_outputs(6814));
    layer2_outputs(593) <= (layer1_outputs(4919)) xor (layer1_outputs(639));
    layer2_outputs(594) <= not(layer1_outputs(6468));
    layer2_outputs(595) <= not((layer1_outputs(9239)) and (layer1_outputs(3861)));
    layer2_outputs(596) <= '0';
    layer2_outputs(597) <= layer1_outputs(6199);
    layer2_outputs(598) <= not(layer1_outputs(2911)) or (layer1_outputs(3966));
    layer2_outputs(599) <= not(layer1_outputs(2795)) or (layer1_outputs(620));
    layer2_outputs(600) <= layer1_outputs(3766);
    layer2_outputs(601) <= layer1_outputs(7613);
    layer2_outputs(602) <= (layer1_outputs(172)) and not (layer1_outputs(1262));
    layer2_outputs(603) <= not((layer1_outputs(3281)) xor (layer1_outputs(6581)));
    layer2_outputs(604) <= not(layer1_outputs(7931));
    layer2_outputs(605) <= not(layer1_outputs(9499));
    layer2_outputs(606) <= not(layer1_outputs(7484)) or (layer1_outputs(5539));
    layer2_outputs(607) <= not(layer1_outputs(6980));
    layer2_outputs(608) <= not(layer1_outputs(7524));
    layer2_outputs(609) <= (layer1_outputs(7090)) or (layer1_outputs(9572));
    layer2_outputs(610) <= not((layer1_outputs(6351)) or (layer1_outputs(3840)));
    layer2_outputs(611) <= not(layer1_outputs(5854));
    layer2_outputs(612) <= (layer1_outputs(5872)) and not (layer1_outputs(9109));
    layer2_outputs(613) <= not(layer1_outputs(4862));
    layer2_outputs(614) <= not(layer1_outputs(1841));
    layer2_outputs(615) <= not(layer1_outputs(4135)) or (layer1_outputs(5763));
    layer2_outputs(616) <= layer1_outputs(8156);
    layer2_outputs(617) <= (layer1_outputs(4098)) or (layer1_outputs(3892));
    layer2_outputs(618) <= not(layer1_outputs(2447));
    layer2_outputs(619) <= layer1_outputs(1405);
    layer2_outputs(620) <= not(layer1_outputs(5091)) or (layer1_outputs(580));
    layer2_outputs(621) <= not(layer1_outputs(8706));
    layer2_outputs(622) <= not(layer1_outputs(4199));
    layer2_outputs(623) <= not(layer1_outputs(9795));
    layer2_outputs(624) <= (layer1_outputs(4948)) xor (layer1_outputs(8276));
    layer2_outputs(625) <= not(layer1_outputs(1754)) or (layer1_outputs(1587));
    layer2_outputs(626) <= not((layer1_outputs(7527)) and (layer1_outputs(4163)));
    layer2_outputs(627) <= (layer1_outputs(2485)) and (layer1_outputs(4902));
    layer2_outputs(628) <= not(layer1_outputs(6609));
    layer2_outputs(629) <= (layer1_outputs(9621)) xor (layer1_outputs(8783));
    layer2_outputs(630) <= not(layer1_outputs(6347));
    layer2_outputs(631) <= layer1_outputs(6254);
    layer2_outputs(632) <= layer1_outputs(9309);
    layer2_outputs(633) <= (layer1_outputs(3166)) or (layer1_outputs(5598));
    layer2_outputs(634) <= layer1_outputs(6213);
    layer2_outputs(635) <= (layer1_outputs(7341)) and (layer1_outputs(6983));
    layer2_outputs(636) <= not(layer1_outputs(7778)) or (layer1_outputs(5954));
    layer2_outputs(637) <= layer1_outputs(3820);
    layer2_outputs(638) <= not((layer1_outputs(980)) or (layer1_outputs(465)));
    layer2_outputs(639) <= layer1_outputs(3232);
    layer2_outputs(640) <= (layer1_outputs(7570)) or (layer1_outputs(1711));
    layer2_outputs(641) <= not(layer1_outputs(2743)) or (layer1_outputs(7465));
    layer2_outputs(642) <= not(layer1_outputs(2479)) or (layer1_outputs(734));
    layer2_outputs(643) <= layer1_outputs(4006);
    layer2_outputs(644) <= (layer1_outputs(5558)) and not (layer1_outputs(10155));
    layer2_outputs(645) <= not(layer1_outputs(7455));
    layer2_outputs(646) <= layer1_outputs(6497);
    layer2_outputs(647) <= layer1_outputs(6624);
    layer2_outputs(648) <= (layer1_outputs(7705)) and not (layer1_outputs(4301));
    layer2_outputs(649) <= not((layer1_outputs(10176)) xor (layer1_outputs(7922)));
    layer2_outputs(650) <= not((layer1_outputs(6089)) or (layer1_outputs(6859)));
    layer2_outputs(651) <= not(layer1_outputs(5868));
    layer2_outputs(652) <= (layer1_outputs(3413)) or (layer1_outputs(3750));
    layer2_outputs(653) <= layer1_outputs(1969);
    layer2_outputs(654) <= not(layer1_outputs(5279));
    layer2_outputs(655) <= not((layer1_outputs(5425)) or (layer1_outputs(7282)));
    layer2_outputs(656) <= (layer1_outputs(196)) and not (layer1_outputs(2410));
    layer2_outputs(657) <= not(layer1_outputs(1114));
    layer2_outputs(658) <= layer1_outputs(7198);
    layer2_outputs(659) <= not((layer1_outputs(4031)) xor (layer1_outputs(4156)));
    layer2_outputs(660) <= layer1_outputs(1405);
    layer2_outputs(661) <= (layer1_outputs(6822)) and not (layer1_outputs(2606));
    layer2_outputs(662) <= not(layer1_outputs(3716));
    layer2_outputs(663) <= not(layer1_outputs(6877));
    layer2_outputs(664) <= (layer1_outputs(8587)) and (layer1_outputs(5398));
    layer2_outputs(665) <= (layer1_outputs(4654)) xor (layer1_outputs(9098));
    layer2_outputs(666) <= not(layer1_outputs(6650));
    layer2_outputs(667) <= not(layer1_outputs(2275));
    layer2_outputs(668) <= not(layer1_outputs(4622)) or (layer1_outputs(8169));
    layer2_outputs(669) <= layer1_outputs(5129);
    layer2_outputs(670) <= (layer1_outputs(28)) xor (layer1_outputs(5644));
    layer2_outputs(671) <= layer1_outputs(3570);
    layer2_outputs(672) <= layer1_outputs(5082);
    layer2_outputs(673) <= not((layer1_outputs(7748)) and (layer1_outputs(405)));
    layer2_outputs(674) <= not(layer1_outputs(3375)) or (layer1_outputs(2157));
    layer2_outputs(675) <= layer1_outputs(9592);
    layer2_outputs(676) <= layer1_outputs(6706);
    layer2_outputs(677) <= not((layer1_outputs(8449)) and (layer1_outputs(4198)));
    layer2_outputs(678) <= layer1_outputs(5429);
    layer2_outputs(679) <= '1';
    layer2_outputs(680) <= (layer1_outputs(872)) and not (layer1_outputs(3484));
    layer2_outputs(681) <= layer1_outputs(322);
    layer2_outputs(682) <= not((layer1_outputs(8415)) and (layer1_outputs(3258)));
    layer2_outputs(683) <= not((layer1_outputs(1888)) and (layer1_outputs(431)));
    layer2_outputs(684) <= not(layer1_outputs(2843));
    layer2_outputs(685) <= not((layer1_outputs(514)) xor (layer1_outputs(4878)));
    layer2_outputs(686) <= layer1_outputs(1418);
    layer2_outputs(687) <= layer1_outputs(6928);
    layer2_outputs(688) <= not(layer1_outputs(8608));
    layer2_outputs(689) <= '0';
    layer2_outputs(690) <= not(layer1_outputs(5733));
    layer2_outputs(691) <= (layer1_outputs(9753)) and not (layer1_outputs(1313));
    layer2_outputs(692) <= (layer1_outputs(3963)) and (layer1_outputs(5520));
    layer2_outputs(693) <= not(layer1_outputs(4367));
    layer2_outputs(694) <= layer1_outputs(7387);
    layer2_outputs(695) <= not((layer1_outputs(3)) or (layer1_outputs(2479)));
    layer2_outputs(696) <= (layer1_outputs(8753)) and not (layer1_outputs(2219));
    layer2_outputs(697) <= not(layer1_outputs(5614));
    layer2_outputs(698) <= not(layer1_outputs(2206));
    layer2_outputs(699) <= not((layer1_outputs(7156)) xor (layer1_outputs(2899)));
    layer2_outputs(700) <= (layer1_outputs(4314)) or (layer1_outputs(390));
    layer2_outputs(701) <= layer1_outputs(3186);
    layer2_outputs(702) <= not(layer1_outputs(2090)) or (layer1_outputs(7034));
    layer2_outputs(703) <= not(layer1_outputs(2829)) or (layer1_outputs(299));
    layer2_outputs(704) <= not(layer1_outputs(7339));
    layer2_outputs(705) <= not(layer1_outputs(8022));
    layer2_outputs(706) <= not(layer1_outputs(5040));
    layer2_outputs(707) <= (layer1_outputs(5476)) and not (layer1_outputs(6434));
    layer2_outputs(708) <= not(layer1_outputs(1597));
    layer2_outputs(709) <= not(layer1_outputs(4040));
    layer2_outputs(710) <= not(layer1_outputs(10077)) or (layer1_outputs(795));
    layer2_outputs(711) <= (layer1_outputs(4865)) xor (layer1_outputs(7653));
    layer2_outputs(712) <= layer1_outputs(4761);
    layer2_outputs(713) <= (layer1_outputs(5583)) and not (layer1_outputs(9253));
    layer2_outputs(714) <= layer1_outputs(1410);
    layer2_outputs(715) <= not(layer1_outputs(1898));
    layer2_outputs(716) <= layer1_outputs(781);
    layer2_outputs(717) <= not((layer1_outputs(3617)) xor (layer1_outputs(8914)));
    layer2_outputs(718) <= not(layer1_outputs(7108)) or (layer1_outputs(7304));
    layer2_outputs(719) <= not(layer1_outputs(2403)) or (layer1_outputs(6851));
    layer2_outputs(720) <= layer1_outputs(6848);
    layer2_outputs(721) <= (layer1_outputs(7237)) xor (layer1_outputs(2441));
    layer2_outputs(722) <= not(layer1_outputs(4383));
    layer2_outputs(723) <= not(layer1_outputs(8315));
    layer2_outputs(724) <= (layer1_outputs(2292)) and not (layer1_outputs(1866));
    layer2_outputs(725) <= not((layer1_outputs(3932)) xor (layer1_outputs(5577)));
    layer2_outputs(726) <= (layer1_outputs(1587)) xor (layer1_outputs(3993));
    layer2_outputs(727) <= not(layer1_outputs(5801)) or (layer1_outputs(4677));
    layer2_outputs(728) <= not(layer1_outputs(9460));
    layer2_outputs(729) <= not((layer1_outputs(4474)) xor (layer1_outputs(1611)));
    layer2_outputs(730) <= not(layer1_outputs(5347));
    layer2_outputs(731) <= not(layer1_outputs(4516));
    layer2_outputs(732) <= not(layer1_outputs(3841));
    layer2_outputs(733) <= not(layer1_outputs(930));
    layer2_outputs(734) <= not(layer1_outputs(2687)) or (layer1_outputs(5172));
    layer2_outputs(735) <= layer1_outputs(5408);
    layer2_outputs(736) <= layer1_outputs(5668);
    layer2_outputs(737) <= (layer1_outputs(2614)) and not (layer1_outputs(3964));
    layer2_outputs(738) <= not(layer1_outputs(6783));
    layer2_outputs(739) <= not(layer1_outputs(9526));
    layer2_outputs(740) <= not((layer1_outputs(9503)) or (layer1_outputs(8637)));
    layer2_outputs(741) <= layer1_outputs(7589);
    layer2_outputs(742) <= (layer1_outputs(3148)) xor (layer1_outputs(6576));
    layer2_outputs(743) <= layer1_outputs(4715);
    layer2_outputs(744) <= not(layer1_outputs(7810));
    layer2_outputs(745) <= not(layer1_outputs(279));
    layer2_outputs(746) <= not(layer1_outputs(3819));
    layer2_outputs(747) <= not(layer1_outputs(5716));
    layer2_outputs(748) <= (layer1_outputs(8265)) xor (layer1_outputs(7292));
    layer2_outputs(749) <= layer1_outputs(3920);
    layer2_outputs(750) <= layer1_outputs(1970);
    layer2_outputs(751) <= not((layer1_outputs(5701)) xor (layer1_outputs(6604)));
    layer2_outputs(752) <= not(layer1_outputs(4193));
    layer2_outputs(753) <= (layer1_outputs(731)) or (layer1_outputs(8535));
    layer2_outputs(754) <= layer1_outputs(1719);
    layer2_outputs(755) <= not(layer1_outputs(3344));
    layer2_outputs(756) <= layer1_outputs(6515);
    layer2_outputs(757) <= (layer1_outputs(7784)) xor (layer1_outputs(9580));
    layer2_outputs(758) <= not(layer1_outputs(9813));
    layer2_outputs(759) <= not(layer1_outputs(3709));
    layer2_outputs(760) <= not((layer1_outputs(8586)) or (layer1_outputs(4117)));
    layer2_outputs(761) <= not(layer1_outputs(5073));
    layer2_outputs(762) <= not((layer1_outputs(473)) or (layer1_outputs(369)));
    layer2_outputs(763) <= not(layer1_outputs(6628)) or (layer1_outputs(8135));
    layer2_outputs(764) <= not(layer1_outputs(2566)) or (layer1_outputs(1195));
    layer2_outputs(765) <= not(layer1_outputs(5609)) or (layer1_outputs(8417));
    layer2_outputs(766) <= not(layer1_outputs(1796));
    layer2_outputs(767) <= not((layer1_outputs(4561)) and (layer1_outputs(2506)));
    layer2_outputs(768) <= '0';
    layer2_outputs(769) <= not(layer1_outputs(2942));
    layer2_outputs(770) <= not((layer1_outputs(5779)) or (layer1_outputs(4312)));
    layer2_outputs(771) <= (layer1_outputs(2286)) xor (layer1_outputs(4736));
    layer2_outputs(772) <= not((layer1_outputs(3023)) xor (layer1_outputs(7723)));
    layer2_outputs(773) <= layer1_outputs(6010);
    layer2_outputs(774) <= (layer1_outputs(10181)) and not (layer1_outputs(6275));
    layer2_outputs(775) <= layer1_outputs(3229);
    layer2_outputs(776) <= layer1_outputs(2662);
    layer2_outputs(777) <= not((layer1_outputs(9624)) and (layer1_outputs(9236)));
    layer2_outputs(778) <= not((layer1_outputs(3287)) xor (layer1_outputs(453)));
    layer2_outputs(779) <= (layer1_outputs(1918)) xor (layer1_outputs(8087));
    layer2_outputs(780) <= not(layer1_outputs(5646));
    layer2_outputs(781) <= layer1_outputs(2679);
    layer2_outputs(782) <= (layer1_outputs(1595)) xor (layer1_outputs(8791));
    layer2_outputs(783) <= not((layer1_outputs(3679)) or (layer1_outputs(8013)));
    layer2_outputs(784) <= (layer1_outputs(6639)) xor (layer1_outputs(5159));
    layer2_outputs(785) <= layer1_outputs(1927);
    layer2_outputs(786) <= layer1_outputs(4399);
    layer2_outputs(787) <= not((layer1_outputs(7882)) xor (layer1_outputs(7704)));
    layer2_outputs(788) <= not(layer1_outputs(971));
    layer2_outputs(789) <= layer1_outputs(5767);
    layer2_outputs(790) <= layer1_outputs(5469);
    layer2_outputs(791) <= not((layer1_outputs(7017)) or (layer1_outputs(657)));
    layer2_outputs(792) <= not(layer1_outputs(2769));
    layer2_outputs(793) <= not(layer1_outputs(7790)) or (layer1_outputs(3943));
    layer2_outputs(794) <= (layer1_outputs(119)) or (layer1_outputs(911));
    layer2_outputs(795) <= not(layer1_outputs(5688)) or (layer1_outputs(7353));
    layer2_outputs(796) <= not(layer1_outputs(4044));
    layer2_outputs(797) <= not(layer1_outputs(8128));
    layer2_outputs(798) <= (layer1_outputs(7590)) or (layer1_outputs(5799));
    layer2_outputs(799) <= not(layer1_outputs(3758)) or (layer1_outputs(5914));
    layer2_outputs(800) <= (layer1_outputs(4200)) xor (layer1_outputs(6774));
    layer2_outputs(801) <= not(layer1_outputs(8982));
    layer2_outputs(802) <= not(layer1_outputs(4625));
    layer2_outputs(803) <= not(layer1_outputs(5916));
    layer2_outputs(804) <= not((layer1_outputs(585)) xor (layer1_outputs(804)));
    layer2_outputs(805) <= layer1_outputs(9447);
    layer2_outputs(806) <= not(layer1_outputs(159));
    layer2_outputs(807) <= not(layer1_outputs(3250)) or (layer1_outputs(7884));
    layer2_outputs(808) <= layer1_outputs(6585);
    layer2_outputs(809) <= not(layer1_outputs(1394));
    layer2_outputs(810) <= layer1_outputs(6025);
    layer2_outputs(811) <= not(layer1_outputs(584)) or (layer1_outputs(2912));
    layer2_outputs(812) <= layer1_outputs(4534);
    layer2_outputs(813) <= not(layer1_outputs(832)) or (layer1_outputs(9748));
    layer2_outputs(814) <= (layer1_outputs(7989)) xor (layer1_outputs(176));
    layer2_outputs(815) <= (layer1_outputs(7553)) or (layer1_outputs(8009));
    layer2_outputs(816) <= (layer1_outputs(5883)) and (layer1_outputs(3800));
    layer2_outputs(817) <= not(layer1_outputs(1339));
    layer2_outputs(818) <= layer1_outputs(10021);
    layer2_outputs(819) <= not(layer1_outputs(5845));
    layer2_outputs(820) <= layer1_outputs(9537);
    layer2_outputs(821) <= not(layer1_outputs(984));
    layer2_outputs(822) <= not((layer1_outputs(803)) or (layer1_outputs(9666)));
    layer2_outputs(823) <= not(layer1_outputs(3024));
    layer2_outputs(824) <= not(layer1_outputs(4008));
    layer2_outputs(825) <= not(layer1_outputs(16));
    layer2_outputs(826) <= (layer1_outputs(2490)) and not (layer1_outputs(1433));
    layer2_outputs(827) <= not(layer1_outputs(9168));
    layer2_outputs(828) <= not(layer1_outputs(3096)) or (layer1_outputs(4425));
    layer2_outputs(829) <= layer1_outputs(3095);
    layer2_outputs(830) <= (layer1_outputs(5800)) or (layer1_outputs(2522));
    layer2_outputs(831) <= (layer1_outputs(4008)) xor (layer1_outputs(347));
    layer2_outputs(832) <= not((layer1_outputs(7212)) and (layer1_outputs(2952)));
    layer2_outputs(833) <= not(layer1_outputs(8346));
    layer2_outputs(834) <= layer1_outputs(9930);
    layer2_outputs(835) <= layer1_outputs(8087);
    layer2_outputs(836) <= not(layer1_outputs(3134)) or (layer1_outputs(6738));
    layer2_outputs(837) <= '1';
    layer2_outputs(838) <= (layer1_outputs(2476)) and (layer1_outputs(5853));
    layer2_outputs(839) <= not(layer1_outputs(6585));
    layer2_outputs(840) <= (layer1_outputs(5398)) and not (layer1_outputs(5219));
    layer2_outputs(841) <= not((layer1_outputs(6780)) and (layer1_outputs(9063)));
    layer2_outputs(842) <= layer1_outputs(9128);
    layer2_outputs(843) <= layer1_outputs(5427);
    layer2_outputs(844) <= not(layer1_outputs(4480));
    layer2_outputs(845) <= layer1_outputs(9330);
    layer2_outputs(846) <= (layer1_outputs(3027)) and not (layer1_outputs(4278));
    layer2_outputs(847) <= not(layer1_outputs(4821));
    layer2_outputs(848) <= layer1_outputs(613);
    layer2_outputs(849) <= not(layer1_outputs(5366));
    layer2_outputs(850) <= not((layer1_outputs(2080)) xor (layer1_outputs(1724)));
    layer2_outputs(851) <= not(layer1_outputs(513));
    layer2_outputs(852) <= not(layer1_outputs(9359));
    layer2_outputs(853) <= layer1_outputs(2502);
    layer2_outputs(854) <= not(layer1_outputs(9838));
    layer2_outputs(855) <= not(layer1_outputs(10143));
    layer2_outputs(856) <= layer1_outputs(10206);
    layer2_outputs(857) <= not(layer1_outputs(1840));
    layer2_outputs(858) <= not(layer1_outputs(1681));
    layer2_outputs(859) <= (layer1_outputs(2703)) xor (layer1_outputs(5946));
    layer2_outputs(860) <= not(layer1_outputs(321)) or (layer1_outputs(8208));
    layer2_outputs(861) <= layer1_outputs(2806);
    layer2_outputs(862) <= not(layer1_outputs(554));
    layer2_outputs(863) <= layer1_outputs(9727);
    layer2_outputs(864) <= layer1_outputs(8910);
    layer2_outputs(865) <= (layer1_outputs(5439)) xor (layer1_outputs(8051));
    layer2_outputs(866) <= layer1_outputs(7017);
    layer2_outputs(867) <= not(layer1_outputs(3254));
    layer2_outputs(868) <= not(layer1_outputs(7288));
    layer2_outputs(869) <= '1';
    layer2_outputs(870) <= layer1_outputs(629);
    layer2_outputs(871) <= layer1_outputs(5222);
    layer2_outputs(872) <= (layer1_outputs(3288)) and not (layer1_outputs(9716));
    layer2_outputs(873) <= layer1_outputs(7905);
    layer2_outputs(874) <= not(layer1_outputs(1361));
    layer2_outputs(875) <= not((layer1_outputs(313)) and (layer1_outputs(6559)));
    layer2_outputs(876) <= (layer1_outputs(4719)) xor (layer1_outputs(8973));
    layer2_outputs(877) <= layer1_outputs(948);
    layer2_outputs(878) <= layer1_outputs(8622);
    layer2_outputs(879) <= layer1_outputs(7458);
    layer2_outputs(880) <= not(layer1_outputs(8919)) or (layer1_outputs(199));
    layer2_outputs(881) <= not(layer1_outputs(10083));
    layer2_outputs(882) <= not(layer1_outputs(3414));
    layer2_outputs(883) <= not(layer1_outputs(1342));
    layer2_outputs(884) <= (layer1_outputs(3041)) and not (layer1_outputs(2308));
    layer2_outputs(885) <= not((layer1_outputs(4619)) and (layer1_outputs(8359)));
    layer2_outputs(886) <= layer1_outputs(10230);
    layer2_outputs(887) <= (layer1_outputs(7319)) and not (layer1_outputs(8333));
    layer2_outputs(888) <= not(layer1_outputs(4516)) or (layer1_outputs(1293));
    layer2_outputs(889) <= (layer1_outputs(8493)) and not (layer1_outputs(1127));
    layer2_outputs(890) <= not((layer1_outputs(7480)) or (layer1_outputs(6093)));
    layer2_outputs(891) <= layer1_outputs(3951);
    layer2_outputs(892) <= layer1_outputs(6996);
    layer2_outputs(893) <= (layer1_outputs(1497)) xor (layer1_outputs(3321));
    layer2_outputs(894) <= layer1_outputs(5380);
    layer2_outputs(895) <= not((layer1_outputs(988)) or (layer1_outputs(6400)));
    layer2_outputs(896) <= not(layer1_outputs(2204));
    layer2_outputs(897) <= not(layer1_outputs(2480));
    layer2_outputs(898) <= not((layer1_outputs(6031)) xor (layer1_outputs(1452)));
    layer2_outputs(899) <= (layer1_outputs(673)) xor (layer1_outputs(9155));
    layer2_outputs(900) <= layer1_outputs(7205);
    layer2_outputs(901) <= not(layer1_outputs(9954));
    layer2_outputs(902) <= not(layer1_outputs(10052));
    layer2_outputs(903) <= (layer1_outputs(3409)) xor (layer1_outputs(2944));
    layer2_outputs(904) <= not(layer1_outputs(7685));
    layer2_outputs(905) <= not(layer1_outputs(3111)) or (layer1_outputs(2849));
    layer2_outputs(906) <= not(layer1_outputs(3586));
    layer2_outputs(907) <= not(layer1_outputs(1958));
    layer2_outputs(908) <= '0';
    layer2_outputs(909) <= not((layer1_outputs(74)) xor (layer1_outputs(6291)));
    layer2_outputs(910) <= layer1_outputs(3477);
    layer2_outputs(911) <= not(layer1_outputs(8794));
    layer2_outputs(912) <= not(layer1_outputs(1727)) or (layer1_outputs(9311));
    layer2_outputs(913) <= layer1_outputs(1732);
    layer2_outputs(914) <= (layer1_outputs(2928)) or (layer1_outputs(7151));
    layer2_outputs(915) <= layer1_outputs(9254);
    layer2_outputs(916) <= not((layer1_outputs(8858)) xor (layer1_outputs(6529)));
    layer2_outputs(917) <= not(layer1_outputs(8770)) or (layer1_outputs(5974));
    layer2_outputs(918) <= layer1_outputs(3797);
    layer2_outputs(919) <= not(layer1_outputs(573));
    layer2_outputs(920) <= not((layer1_outputs(4459)) xor (layer1_outputs(5160)));
    layer2_outputs(921) <= not(layer1_outputs(741));
    layer2_outputs(922) <= not(layer1_outputs(2106)) or (layer1_outputs(5539));
    layer2_outputs(923) <= (layer1_outputs(6662)) xor (layer1_outputs(6715));
    layer2_outputs(924) <= not(layer1_outputs(1755)) or (layer1_outputs(9490));
    layer2_outputs(925) <= not((layer1_outputs(9726)) xor (layer1_outputs(1232)));
    layer2_outputs(926) <= not(layer1_outputs(1569)) or (layer1_outputs(6644));
    layer2_outputs(927) <= not(layer1_outputs(4888)) or (layer1_outputs(9420));
    layer2_outputs(928) <= (layer1_outputs(3879)) or (layer1_outputs(9774));
    layer2_outputs(929) <= not((layer1_outputs(7336)) xor (layer1_outputs(9153)));
    layer2_outputs(930) <= (layer1_outputs(1955)) and not (layer1_outputs(3328));
    layer2_outputs(931) <= not(layer1_outputs(1346));
    layer2_outputs(932) <= not((layer1_outputs(6023)) and (layer1_outputs(6338)));
    layer2_outputs(933) <= layer1_outputs(1512);
    layer2_outputs(934) <= not((layer1_outputs(3657)) and (layer1_outputs(8607)));
    layer2_outputs(935) <= not(layer1_outputs(6809));
    layer2_outputs(936) <= layer1_outputs(6589);
    layer2_outputs(937) <= layer1_outputs(7110);
    layer2_outputs(938) <= not(layer1_outputs(2555));
    layer2_outputs(939) <= (layer1_outputs(6368)) and not (layer1_outputs(8122));
    layer2_outputs(940) <= not(layer1_outputs(5740)) or (layer1_outputs(9378));
    layer2_outputs(941) <= not(layer1_outputs(5419)) or (layer1_outputs(8221));
    layer2_outputs(942) <= not((layer1_outputs(1225)) xor (layer1_outputs(6020)));
    layer2_outputs(943) <= layer1_outputs(1561);
    layer2_outputs(944) <= (layer1_outputs(8768)) and (layer1_outputs(3560));
    layer2_outputs(945) <= not((layer1_outputs(5446)) xor (layer1_outputs(2551)));
    layer2_outputs(946) <= not((layer1_outputs(7661)) and (layer1_outputs(2356)));
    layer2_outputs(947) <= (layer1_outputs(1954)) xor (layer1_outputs(2206));
    layer2_outputs(948) <= layer1_outputs(3105);
    layer2_outputs(949) <= not(layer1_outputs(6564)) or (layer1_outputs(9210));
    layer2_outputs(950) <= (layer1_outputs(6141)) and not (layer1_outputs(9905));
    layer2_outputs(951) <= not(layer1_outputs(7125));
    layer2_outputs(952) <= not(layer1_outputs(9810)) or (layer1_outputs(5180));
    layer2_outputs(953) <= not(layer1_outputs(1820));
    layer2_outputs(954) <= not(layer1_outputs(2703));
    layer2_outputs(955) <= not(layer1_outputs(8010)) or (layer1_outputs(2182));
    layer2_outputs(956) <= not(layer1_outputs(6895));
    layer2_outputs(957) <= not((layer1_outputs(9856)) xor (layer1_outputs(69)));
    layer2_outputs(958) <= not(layer1_outputs(8579));
    layer2_outputs(959) <= layer1_outputs(2718);
    layer2_outputs(960) <= (layer1_outputs(4655)) and not (layer1_outputs(965));
    layer2_outputs(961) <= layer1_outputs(10084);
    layer2_outputs(962) <= (layer1_outputs(4223)) xor (layer1_outputs(3818));
    layer2_outputs(963) <= (layer1_outputs(10156)) and (layer1_outputs(1572));
    layer2_outputs(964) <= layer1_outputs(5617);
    layer2_outputs(965) <= (layer1_outputs(8737)) and not (layer1_outputs(7402));
    layer2_outputs(966) <= layer1_outputs(9694);
    layer2_outputs(967) <= layer1_outputs(5204);
    layer2_outputs(968) <= (layer1_outputs(9873)) and (layer1_outputs(7213));
    layer2_outputs(969) <= not((layer1_outputs(551)) or (layer1_outputs(7732)));
    layer2_outputs(970) <= layer1_outputs(10218);
    layer2_outputs(971) <= not(layer1_outputs(2956));
    layer2_outputs(972) <= (layer1_outputs(4268)) and not (layer1_outputs(2532));
    layer2_outputs(973) <= layer1_outputs(7876);
    layer2_outputs(974) <= not(layer1_outputs(7729)) or (layer1_outputs(7226));
    layer2_outputs(975) <= not((layer1_outputs(9971)) xor (layer1_outputs(7564)));
    layer2_outputs(976) <= layer1_outputs(6022);
    layer2_outputs(977) <= not(layer1_outputs(9611));
    layer2_outputs(978) <= not(layer1_outputs(8616)) or (layer1_outputs(7849));
    layer2_outputs(979) <= (layer1_outputs(54)) xor (layer1_outputs(9302));
    layer2_outputs(980) <= (layer1_outputs(6262)) and not (layer1_outputs(1001));
    layer2_outputs(981) <= (layer1_outputs(1610)) and (layer1_outputs(1446));
    layer2_outputs(982) <= not(layer1_outputs(9451));
    layer2_outputs(983) <= (layer1_outputs(9600)) and not (layer1_outputs(5361));
    layer2_outputs(984) <= not(layer1_outputs(10084)) or (layer1_outputs(1632));
    layer2_outputs(985) <= not(layer1_outputs(8245)) or (layer1_outputs(6795));
    layer2_outputs(986) <= layer1_outputs(2078);
    layer2_outputs(987) <= not((layer1_outputs(1230)) xor (layer1_outputs(9135)));
    layer2_outputs(988) <= not(layer1_outputs(6390));
    layer2_outputs(989) <= not(layer1_outputs(7020)) or (layer1_outputs(3155));
    layer2_outputs(990) <= '1';
    layer2_outputs(991) <= layer1_outputs(1526);
    layer2_outputs(992) <= not(layer1_outputs(4119));
    layer2_outputs(993) <= not(layer1_outputs(8173)) or (layer1_outputs(5143));
    layer2_outputs(994) <= not(layer1_outputs(6773));
    layer2_outputs(995) <= not(layer1_outputs(8575));
    layer2_outputs(996) <= (layer1_outputs(3192)) and not (layer1_outputs(4178));
    layer2_outputs(997) <= not((layer1_outputs(2516)) and (layer1_outputs(8509)));
    layer2_outputs(998) <= layer1_outputs(720);
    layer2_outputs(999) <= layer1_outputs(3140);
    layer2_outputs(1000) <= '0';
    layer2_outputs(1001) <= not((layer1_outputs(8248)) or (layer1_outputs(7305)));
    layer2_outputs(1002) <= (layer1_outputs(3320)) and (layer1_outputs(6266));
    layer2_outputs(1003) <= not((layer1_outputs(8708)) and (layer1_outputs(4800)));
    layer2_outputs(1004) <= (layer1_outputs(4443)) xor (layer1_outputs(3624));
    layer2_outputs(1005) <= not(layer1_outputs(7213)) or (layer1_outputs(8891));
    layer2_outputs(1006) <= (layer1_outputs(2550)) xor (layer1_outputs(4606));
    layer2_outputs(1007) <= layer1_outputs(6966);
    layer2_outputs(1008) <= not(layer1_outputs(2273)) or (layer1_outputs(2020));
    layer2_outputs(1009) <= not(layer1_outputs(8588)) or (layer1_outputs(5214));
    layer2_outputs(1010) <= not(layer1_outputs(790));
    layer2_outputs(1011) <= layer1_outputs(5340);
    layer2_outputs(1012) <= not(layer1_outputs(8867));
    layer2_outputs(1013) <= not(layer1_outputs(6444));
    layer2_outputs(1014) <= not((layer1_outputs(4607)) or (layer1_outputs(2245)));
    layer2_outputs(1015) <= not((layer1_outputs(5681)) or (layer1_outputs(5127)));
    layer2_outputs(1016) <= (layer1_outputs(3506)) and not (layer1_outputs(4376));
    layer2_outputs(1017) <= (layer1_outputs(6604)) xor (layer1_outputs(2000));
    layer2_outputs(1018) <= '1';
    layer2_outputs(1019) <= layer1_outputs(9116);
    layer2_outputs(1020) <= not(layer1_outputs(6773)) or (layer1_outputs(7301));
    layer2_outputs(1021) <= layer1_outputs(202);
    layer2_outputs(1022) <= not(layer1_outputs(8485)) or (layer1_outputs(6471));
    layer2_outputs(1023) <= layer1_outputs(9922);
    layer2_outputs(1024) <= layer1_outputs(3973);
    layer2_outputs(1025) <= layer1_outputs(8944);
    layer2_outputs(1026) <= layer1_outputs(9606);
    layer2_outputs(1027) <= not(layer1_outputs(9997)) or (layer1_outputs(5295));
    layer2_outputs(1028) <= (layer1_outputs(6330)) or (layer1_outputs(1758));
    layer2_outputs(1029) <= not(layer1_outputs(38));
    layer2_outputs(1030) <= layer1_outputs(931);
    layer2_outputs(1031) <= layer1_outputs(6326);
    layer2_outputs(1032) <= not(layer1_outputs(4652));
    layer2_outputs(1033) <= (layer1_outputs(8838)) and not (layer1_outputs(8898));
    layer2_outputs(1034) <= layer1_outputs(5925);
    layer2_outputs(1035) <= not(layer1_outputs(7390));
    layer2_outputs(1036) <= not(layer1_outputs(2053));
    layer2_outputs(1037) <= not(layer1_outputs(9077));
    layer2_outputs(1038) <= layer1_outputs(2568);
    layer2_outputs(1039) <= (layer1_outputs(4258)) or (layer1_outputs(1068));
    layer2_outputs(1040) <= not((layer1_outputs(9301)) xor (layer1_outputs(10114)));
    layer2_outputs(1041) <= not(layer1_outputs(8041));
    layer2_outputs(1042) <= layer1_outputs(9976);
    layer2_outputs(1043) <= not((layer1_outputs(6880)) and (layer1_outputs(1897)));
    layer2_outputs(1044) <= layer1_outputs(301);
    layer2_outputs(1045) <= layer1_outputs(8951);
    layer2_outputs(1046) <= not((layer1_outputs(7152)) or (layer1_outputs(7937)));
    layer2_outputs(1047) <= not(layer1_outputs(3303)) or (layer1_outputs(3972));
    layer2_outputs(1048) <= layer1_outputs(2493);
    layer2_outputs(1049) <= not(layer1_outputs(3031)) or (layer1_outputs(686));
    layer2_outputs(1050) <= not((layer1_outputs(5884)) and (layer1_outputs(6848)));
    layer2_outputs(1051) <= layer1_outputs(9024);
    layer2_outputs(1052) <= not(layer1_outputs(7080));
    layer2_outputs(1053) <= layer1_outputs(7761);
    layer2_outputs(1054) <= not(layer1_outputs(2908)) or (layer1_outputs(4562));
    layer2_outputs(1055) <= not((layer1_outputs(5548)) and (layer1_outputs(5868)));
    layer2_outputs(1056) <= (layer1_outputs(5586)) and (layer1_outputs(8281));
    layer2_outputs(1057) <= (layer1_outputs(9037)) xor (layer1_outputs(10008));
    layer2_outputs(1058) <= (layer1_outputs(4832)) and not (layer1_outputs(3226));
    layer2_outputs(1059) <= layer1_outputs(5131);
    layer2_outputs(1060) <= not(layer1_outputs(2074));
    layer2_outputs(1061) <= not(layer1_outputs(4030));
    layer2_outputs(1062) <= not((layer1_outputs(6099)) xor (layer1_outputs(4768)));
    layer2_outputs(1063) <= not(layer1_outputs(6514));
    layer2_outputs(1064) <= (layer1_outputs(1941)) and not (layer1_outputs(9702));
    layer2_outputs(1065) <= layer1_outputs(1264);
    layer2_outputs(1066) <= not(layer1_outputs(7952));
    layer2_outputs(1067) <= not(layer1_outputs(2026));
    layer2_outputs(1068) <= not(layer1_outputs(376));
    layer2_outputs(1069) <= (layer1_outputs(1479)) and not (layer1_outputs(4809));
    layer2_outputs(1070) <= (layer1_outputs(3286)) xor (layer1_outputs(8234));
    layer2_outputs(1071) <= not(layer1_outputs(5052));
    layer2_outputs(1072) <= (layer1_outputs(2890)) and not (layer1_outputs(1257));
    layer2_outputs(1073) <= layer1_outputs(4057);
    layer2_outputs(1074) <= not(layer1_outputs(3475));
    layer2_outputs(1075) <= (layer1_outputs(4896)) and not (layer1_outputs(1857));
    layer2_outputs(1076) <= not(layer1_outputs(2177));
    layer2_outputs(1077) <= (layer1_outputs(8479)) and not (layer1_outputs(9914));
    layer2_outputs(1078) <= not((layer1_outputs(2546)) and (layer1_outputs(8695)));
    layer2_outputs(1079) <= not(layer1_outputs(10145)) or (layer1_outputs(4886));
    layer2_outputs(1080) <= '0';
    layer2_outputs(1081) <= not(layer1_outputs(363));
    layer2_outputs(1082) <= '0';
    layer2_outputs(1083) <= (layer1_outputs(282)) or (layer1_outputs(4568));
    layer2_outputs(1084) <= not(layer1_outputs(2021));
    layer2_outputs(1085) <= not((layer1_outputs(2877)) and (layer1_outputs(2999)));
    layer2_outputs(1086) <= layer1_outputs(6993);
    layer2_outputs(1087) <= not((layer1_outputs(6006)) or (layer1_outputs(2672)));
    layer2_outputs(1088) <= not((layer1_outputs(3519)) and (layer1_outputs(2965)));
    layer2_outputs(1089) <= layer1_outputs(10086);
    layer2_outputs(1090) <= layer1_outputs(2034);
    layer2_outputs(1091) <= not((layer1_outputs(6361)) or (layer1_outputs(2201)));
    layer2_outputs(1092) <= not((layer1_outputs(7628)) and (layer1_outputs(9465)));
    layer2_outputs(1093) <= not((layer1_outputs(10080)) xor (layer1_outputs(6427)));
    layer2_outputs(1094) <= layer1_outputs(9851);
    layer2_outputs(1095) <= layer1_outputs(7264);
    layer2_outputs(1096) <= not(layer1_outputs(1961));
    layer2_outputs(1097) <= layer1_outputs(9141);
    layer2_outputs(1098) <= not(layer1_outputs(8775));
    layer2_outputs(1099) <= not((layer1_outputs(3625)) xor (layer1_outputs(4038)));
    layer2_outputs(1100) <= not(layer1_outputs(2306));
    layer2_outputs(1101) <= layer1_outputs(3526);
    layer2_outputs(1102) <= layer1_outputs(5642);
    layer2_outputs(1103) <= (layer1_outputs(10158)) and not (layer1_outputs(9363));
    layer2_outputs(1104) <= (layer1_outputs(4260)) or (layer1_outputs(10100));
    layer2_outputs(1105) <= not((layer1_outputs(4753)) or (layer1_outputs(8545)));
    layer2_outputs(1106) <= not(layer1_outputs(9095));
    layer2_outputs(1107) <= not(layer1_outputs(5838));
    layer2_outputs(1108) <= not(layer1_outputs(9158));
    layer2_outputs(1109) <= layer1_outputs(6830);
    layer2_outputs(1110) <= (layer1_outputs(6581)) and (layer1_outputs(6488));
    layer2_outputs(1111) <= layer1_outputs(7625);
    layer2_outputs(1112) <= not((layer1_outputs(229)) xor (layer1_outputs(4254)));
    layer2_outputs(1113) <= not((layer1_outputs(2968)) or (layer1_outputs(3859)));
    layer2_outputs(1114) <= (layer1_outputs(5468)) and not (layer1_outputs(2315));
    layer2_outputs(1115) <= not(layer1_outputs(9154));
    layer2_outputs(1116) <= layer1_outputs(8716);
    layer2_outputs(1117) <= layer1_outputs(6413);
    layer2_outputs(1118) <= layer1_outputs(57);
    layer2_outputs(1119) <= layer1_outputs(2443);
    layer2_outputs(1120) <= not(layer1_outputs(1573)) or (layer1_outputs(8352));
    layer2_outputs(1121) <= not(layer1_outputs(7363));
    layer2_outputs(1122) <= (layer1_outputs(4150)) and not (layer1_outputs(102));
    layer2_outputs(1123) <= not((layer1_outputs(7011)) xor (layer1_outputs(7713)));
    layer2_outputs(1124) <= layer1_outputs(3966);
    layer2_outputs(1125) <= not(layer1_outputs(457));
    layer2_outputs(1126) <= layer1_outputs(10234);
    layer2_outputs(1127) <= layer1_outputs(4654);
    layer2_outputs(1128) <= not(layer1_outputs(2007));
    layer2_outputs(1129) <= not(layer1_outputs(7889)) or (layer1_outputs(8309));
    layer2_outputs(1130) <= not(layer1_outputs(1777)) or (layer1_outputs(7355));
    layer2_outputs(1131) <= layer1_outputs(9207);
    layer2_outputs(1132) <= not(layer1_outputs(1765));
    layer2_outputs(1133) <= (layer1_outputs(1053)) and not (layer1_outputs(7295));
    layer2_outputs(1134) <= layer1_outputs(1696);
    layer2_outputs(1135) <= layer1_outputs(3034);
    layer2_outputs(1136) <= layer1_outputs(8730);
    layer2_outputs(1137) <= not((layer1_outputs(989)) xor (layer1_outputs(8371)));
    layer2_outputs(1138) <= layer1_outputs(8030);
    layer2_outputs(1139) <= (layer1_outputs(3669)) or (layer1_outputs(1056));
    layer2_outputs(1140) <= not((layer1_outputs(9182)) or (layer1_outputs(9046)));
    layer2_outputs(1141) <= not(layer1_outputs(8924));
    layer2_outputs(1142) <= not((layer1_outputs(8538)) xor (layer1_outputs(458)));
    layer2_outputs(1143) <= layer1_outputs(4286);
    layer2_outputs(1144) <= layer1_outputs(6938);
    layer2_outputs(1145) <= not(layer1_outputs(6675)) or (layer1_outputs(9769));
    layer2_outputs(1146) <= not(layer1_outputs(6736));
    layer2_outputs(1147) <= not(layer1_outputs(1037));
    layer2_outputs(1148) <= (layer1_outputs(6813)) xor (layer1_outputs(8667));
    layer2_outputs(1149) <= not(layer1_outputs(5092)) or (layer1_outputs(512));
    layer2_outputs(1150) <= not(layer1_outputs(1799));
    layer2_outputs(1151) <= layer1_outputs(5878);
    layer2_outputs(1152) <= layer1_outputs(1783);
    layer2_outputs(1153) <= (layer1_outputs(4563)) and (layer1_outputs(5772));
    layer2_outputs(1154) <= layer1_outputs(2610);
    layer2_outputs(1155) <= (layer1_outputs(2295)) or (layer1_outputs(7221));
    layer2_outputs(1156) <= not(layer1_outputs(6804));
    layer2_outputs(1157) <= layer1_outputs(3083);
    layer2_outputs(1158) <= (layer1_outputs(832)) and (layer1_outputs(410));
    layer2_outputs(1159) <= not(layer1_outputs(9913)) or (layer1_outputs(2656));
    layer2_outputs(1160) <= (layer1_outputs(7027)) or (layer1_outputs(844));
    layer2_outputs(1161) <= layer1_outputs(8550);
    layer2_outputs(1162) <= layer1_outputs(4619);
    layer2_outputs(1163) <= not(layer1_outputs(3694)) or (layer1_outputs(5382));
    layer2_outputs(1164) <= not(layer1_outputs(9622)) or (layer1_outputs(9483));
    layer2_outputs(1165) <= not(layer1_outputs(9697));
    layer2_outputs(1166) <= layer1_outputs(2163);
    layer2_outputs(1167) <= not(layer1_outputs(5192)) or (layer1_outputs(9812));
    layer2_outputs(1168) <= not(layer1_outputs(7219));
    layer2_outputs(1169) <= layer1_outputs(3208);
    layer2_outputs(1170) <= layer1_outputs(5785);
    layer2_outputs(1171) <= layer1_outputs(7954);
    layer2_outputs(1172) <= not(layer1_outputs(659)) or (layer1_outputs(3736));
    layer2_outputs(1173) <= (layer1_outputs(3040)) xor (layer1_outputs(3498));
    layer2_outputs(1174) <= not(layer1_outputs(6954));
    layer2_outputs(1175) <= layer1_outputs(2378);
    layer2_outputs(1176) <= '0';
    layer2_outputs(1177) <= (layer1_outputs(258)) and not (layer1_outputs(8617));
    layer2_outputs(1178) <= (layer1_outputs(1274)) xor (layer1_outputs(3213));
    layer2_outputs(1179) <= layer1_outputs(917);
    layer2_outputs(1180) <= not((layer1_outputs(7811)) xor (layer1_outputs(5491)));
    layer2_outputs(1181) <= not((layer1_outputs(5786)) or (layer1_outputs(10237)));
    layer2_outputs(1182) <= not(layer1_outputs(658));
    layer2_outputs(1183) <= '1';
    layer2_outputs(1184) <= layer1_outputs(6896);
    layer2_outputs(1185) <= not(layer1_outputs(4554));
    layer2_outputs(1186) <= not(layer1_outputs(8758));
    layer2_outputs(1187) <= not(layer1_outputs(6486));
    layer2_outputs(1188) <= not(layer1_outputs(10002));
    layer2_outputs(1189) <= not(layer1_outputs(9133));
    layer2_outputs(1190) <= (layer1_outputs(887)) and not (layer1_outputs(9080));
    layer2_outputs(1191) <= not(layer1_outputs(6021));
    layer2_outputs(1192) <= not(layer1_outputs(5160));
    layer2_outputs(1193) <= not(layer1_outputs(3592));
    layer2_outputs(1194) <= layer1_outputs(8975);
    layer2_outputs(1195) <= (layer1_outputs(7751)) and not (layer1_outputs(4946));
    layer2_outputs(1196) <= not(layer1_outputs(7873));
    layer2_outputs(1197) <= not((layer1_outputs(487)) or (layer1_outputs(7816)));
    layer2_outputs(1198) <= (layer1_outputs(5475)) or (layer1_outputs(7029));
    layer2_outputs(1199) <= layer1_outputs(4503);
    layer2_outputs(1200) <= not(layer1_outputs(5938));
    layer2_outputs(1201) <= not((layer1_outputs(9156)) or (layer1_outputs(9135)));
    layer2_outputs(1202) <= layer1_outputs(946);
    layer2_outputs(1203) <= (layer1_outputs(3696)) and not (layer1_outputs(1728));
    layer2_outputs(1204) <= (layer1_outputs(803)) or (layer1_outputs(7256));
    layer2_outputs(1205) <= not((layer1_outputs(5095)) or (layer1_outputs(1474)));
    layer2_outputs(1206) <= (layer1_outputs(232)) and not (layer1_outputs(8405));
    layer2_outputs(1207) <= layer1_outputs(2398);
    layer2_outputs(1208) <= (layer1_outputs(5629)) or (layer1_outputs(8174));
    layer2_outputs(1209) <= layer1_outputs(8859);
    layer2_outputs(1210) <= not(layer1_outputs(7151));
    layer2_outputs(1211) <= layer1_outputs(7868);
    layer2_outputs(1212) <= layer1_outputs(10018);
    layer2_outputs(1213) <= layer1_outputs(544);
    layer2_outputs(1214) <= (layer1_outputs(2451)) and not (layer1_outputs(3178));
    layer2_outputs(1215) <= not(layer1_outputs(4015));
    layer2_outputs(1216) <= layer1_outputs(8244);
    layer2_outputs(1217) <= layer1_outputs(5760);
    layer2_outputs(1218) <= not(layer1_outputs(4706)) or (layer1_outputs(880));
    layer2_outputs(1219) <= layer1_outputs(5212);
    layer2_outputs(1220) <= (layer1_outputs(3940)) and (layer1_outputs(4257));
    layer2_outputs(1221) <= not(layer1_outputs(7425)) or (layer1_outputs(6478));
    layer2_outputs(1222) <= not(layer1_outputs(6172));
    layer2_outputs(1223) <= not(layer1_outputs(9265)) or (layer1_outputs(3691));
    layer2_outputs(1224) <= layer1_outputs(1471);
    layer2_outputs(1225) <= layer1_outputs(2100);
    layer2_outputs(1226) <= (layer1_outputs(7911)) xor (layer1_outputs(2056));
    layer2_outputs(1227) <= (layer1_outputs(6352)) or (layer1_outputs(7673));
    layer2_outputs(1228) <= (layer1_outputs(6728)) and not (layer1_outputs(5104));
    layer2_outputs(1229) <= not(layer1_outputs(8676)) or (layer1_outputs(5861));
    layer2_outputs(1230) <= not(layer1_outputs(9399));
    layer2_outputs(1231) <= not(layer1_outputs(6718));
    layer2_outputs(1232) <= (layer1_outputs(3620)) and (layer1_outputs(2791));
    layer2_outputs(1233) <= layer1_outputs(10220);
    layer2_outputs(1234) <= (layer1_outputs(6043)) and (layer1_outputs(8210));
    layer2_outputs(1235) <= not((layer1_outputs(10001)) xor (layer1_outputs(5107)));
    layer2_outputs(1236) <= layer1_outputs(848);
    layer2_outputs(1237) <= (layer1_outputs(514)) and (layer1_outputs(6850));
    layer2_outputs(1238) <= layer1_outputs(7714);
    layer2_outputs(1239) <= layer1_outputs(10104);
    layer2_outputs(1240) <= not(layer1_outputs(2299));
    layer2_outputs(1241) <= not(layer1_outputs(6706)) or (layer1_outputs(2604));
    layer2_outputs(1242) <= not(layer1_outputs(5293)) or (layer1_outputs(1386));
    layer2_outputs(1243) <= not((layer1_outputs(7553)) or (layer1_outputs(5396)));
    layer2_outputs(1244) <= not((layer1_outputs(9392)) and (layer1_outputs(495)));
    layer2_outputs(1245) <= (layer1_outputs(6098)) and (layer1_outputs(1524));
    layer2_outputs(1246) <= layer1_outputs(2261);
    layer2_outputs(1247) <= layer1_outputs(5428);
    layer2_outputs(1248) <= layer1_outputs(695);
    layer2_outputs(1249) <= (layer1_outputs(9120)) and (layer1_outputs(1034));
    layer2_outputs(1250) <= (layer1_outputs(2713)) or (layer1_outputs(3443));
    layer2_outputs(1251) <= layer1_outputs(1640);
    layer2_outputs(1252) <= layer1_outputs(7407);
    layer2_outputs(1253) <= not(layer1_outputs(3436)) or (layer1_outputs(5140));
    layer2_outputs(1254) <= layer1_outputs(6682);
    layer2_outputs(1255) <= not(layer1_outputs(3385)) or (layer1_outputs(5088));
    layer2_outputs(1256) <= (layer1_outputs(7384)) and not (layer1_outputs(2472));
    layer2_outputs(1257) <= not(layer1_outputs(9911)) or (layer1_outputs(4581));
    layer2_outputs(1258) <= not(layer1_outputs(9576));
    layer2_outputs(1259) <= not(layer1_outputs(2221));
    layer2_outputs(1260) <= not(layer1_outputs(2232));
    layer2_outputs(1261) <= (layer1_outputs(8496)) or (layer1_outputs(5250));
    layer2_outputs(1262) <= (layer1_outputs(8294)) and not (layer1_outputs(7473));
    layer2_outputs(1263) <= layer1_outputs(6135);
    layer2_outputs(1264) <= layer1_outputs(8629);
    layer2_outputs(1265) <= (layer1_outputs(1317)) and (layer1_outputs(8180));
    layer2_outputs(1266) <= not((layer1_outputs(9141)) and (layer1_outputs(4179)));
    layer2_outputs(1267) <= not(layer1_outputs(6429)) or (layer1_outputs(8573));
    layer2_outputs(1268) <= not(layer1_outputs(4282)) or (layer1_outputs(3340));
    layer2_outputs(1269) <= (layer1_outputs(5753)) xor (layer1_outputs(3399));
    layer2_outputs(1270) <= not(layer1_outputs(6052));
    layer2_outputs(1271) <= layer1_outputs(4025);
    layer2_outputs(1272) <= not(layer1_outputs(6341));
    layer2_outputs(1273) <= not((layer1_outputs(9758)) and (layer1_outputs(4486)));
    layer2_outputs(1274) <= layer1_outputs(7078);
    layer2_outputs(1275) <= (layer1_outputs(8309)) and not (layer1_outputs(3530));
    layer2_outputs(1276) <= not((layer1_outputs(9709)) xor (layer1_outputs(1419)));
    layer2_outputs(1277) <= layer1_outputs(7756);
    layer2_outputs(1278) <= not((layer1_outputs(2883)) xor (layer1_outputs(6484)));
    layer2_outputs(1279) <= (layer1_outputs(5034)) or (layer1_outputs(3722));
    layer2_outputs(1280) <= layer1_outputs(9907);
    layer2_outputs(1281) <= not(layer1_outputs(9691));
    layer2_outputs(1282) <= (layer1_outputs(4497)) and (layer1_outputs(745));
    layer2_outputs(1283) <= (layer1_outputs(1291)) and not (layer1_outputs(8635));
    layer2_outputs(1284) <= (layer1_outputs(6083)) and (layer1_outputs(5958));
    layer2_outputs(1285) <= layer1_outputs(9892);
    layer2_outputs(1286) <= not(layer1_outputs(4391));
    layer2_outputs(1287) <= (layer1_outputs(4844)) xor (layer1_outputs(2343));
    layer2_outputs(1288) <= layer1_outputs(9);
    layer2_outputs(1289) <= layer1_outputs(4005);
    layer2_outputs(1290) <= not((layer1_outputs(6081)) and (layer1_outputs(5346)));
    layer2_outputs(1291) <= not((layer1_outputs(7132)) xor (layer1_outputs(5179)));
    layer2_outputs(1292) <= layer1_outputs(1666);
    layer2_outputs(1293) <= not(layer1_outputs(978)) or (layer1_outputs(4489));
    layer2_outputs(1294) <= not(layer1_outputs(5489));
    layer2_outputs(1295) <= not(layer1_outputs(4949));
    layer2_outputs(1296) <= not(layer1_outputs(6850));
    layer2_outputs(1297) <= (layer1_outputs(6281)) xor (layer1_outputs(5774));
    layer2_outputs(1298) <= (layer1_outputs(7902)) and not (layer1_outputs(5846));
    layer2_outputs(1299) <= not((layer1_outputs(9209)) and (layer1_outputs(1536)));
    layer2_outputs(1300) <= layer1_outputs(3829);
    layer2_outputs(1301) <= (layer1_outputs(3907)) or (layer1_outputs(1529));
    layer2_outputs(1302) <= not((layer1_outputs(5611)) xor (layer1_outputs(4236)));
    layer2_outputs(1303) <= not(layer1_outputs(2898));
    layer2_outputs(1304) <= not((layer1_outputs(10192)) and (layer1_outputs(8437)));
    layer2_outputs(1305) <= not((layer1_outputs(6762)) or (layer1_outputs(8510)));
    layer2_outputs(1306) <= not((layer1_outputs(2096)) or (layer1_outputs(848)));
    layer2_outputs(1307) <= not(layer1_outputs(1734));
    layer2_outputs(1308) <= not(layer1_outputs(8178)) or (layer1_outputs(7225));
    layer2_outputs(1309) <= layer1_outputs(1394);
    layer2_outputs(1310) <= layer1_outputs(605);
    layer2_outputs(1311) <= layer1_outputs(8740);
    layer2_outputs(1312) <= layer1_outputs(6263);
    layer2_outputs(1313) <= layer1_outputs(9808);
    layer2_outputs(1314) <= layer1_outputs(6883);
    layer2_outputs(1315) <= layer1_outputs(7886);
    layer2_outputs(1316) <= not(layer1_outputs(4837));
    layer2_outputs(1317) <= (layer1_outputs(4444)) or (layer1_outputs(6696));
    layer2_outputs(1318) <= (layer1_outputs(4079)) xor (layer1_outputs(21));
    layer2_outputs(1319) <= not(layer1_outputs(2695)) or (layer1_outputs(6959));
    layer2_outputs(1320) <= not((layer1_outputs(4742)) or (layer1_outputs(463)));
    layer2_outputs(1321) <= layer1_outputs(8918);
    layer2_outputs(1322) <= (layer1_outputs(7271)) xor (layer1_outputs(7571));
    layer2_outputs(1323) <= (layer1_outputs(1652)) xor (layer1_outputs(6106));
    layer2_outputs(1324) <= layer1_outputs(1036);
    layer2_outputs(1325) <= layer1_outputs(3930);
    layer2_outputs(1326) <= not(layer1_outputs(1279));
    layer2_outputs(1327) <= (layer1_outputs(8540)) xor (layer1_outputs(7573));
    layer2_outputs(1328) <= (layer1_outputs(148)) and not (layer1_outputs(9935));
    layer2_outputs(1329) <= not(layer1_outputs(6009));
    layer2_outputs(1330) <= layer1_outputs(4237);
    layer2_outputs(1331) <= (layer1_outputs(5488)) xor (layer1_outputs(3019));
    layer2_outputs(1332) <= '1';
    layer2_outputs(1333) <= not((layer1_outputs(2841)) xor (layer1_outputs(7397)));
    layer2_outputs(1334) <= (layer1_outputs(3714)) and (layer1_outputs(4846));
    layer2_outputs(1335) <= layer1_outputs(2650);
    layer2_outputs(1336) <= not(layer1_outputs(3314));
    layer2_outputs(1337) <= (layer1_outputs(5905)) xor (layer1_outputs(7458));
    layer2_outputs(1338) <= (layer1_outputs(9744)) or (layer1_outputs(490));
    layer2_outputs(1339) <= layer1_outputs(5806);
    layer2_outputs(1340) <= not((layer1_outputs(6515)) xor (layer1_outputs(6133)));
    layer2_outputs(1341) <= not(layer1_outputs(3193));
    layer2_outputs(1342) <= not(layer1_outputs(8728)) or (layer1_outputs(4993));
    layer2_outputs(1343) <= not((layer1_outputs(9183)) xor (layer1_outputs(7618)));
    layer2_outputs(1344) <= (layer1_outputs(559)) and (layer1_outputs(368));
    layer2_outputs(1345) <= not(layer1_outputs(3076)) or (layer1_outputs(9278));
    layer2_outputs(1346) <= not(layer1_outputs(5781)) or (layer1_outputs(7347));
    layer2_outputs(1347) <= (layer1_outputs(6464)) and not (layer1_outputs(1142));
    layer2_outputs(1348) <= not(layer1_outputs(4492));
    layer2_outputs(1349) <= layer1_outputs(1097);
    layer2_outputs(1350) <= not(layer1_outputs(4050));
    layer2_outputs(1351) <= layer1_outputs(4819);
    layer2_outputs(1352) <= not(layer1_outputs(6117));
    layer2_outputs(1353) <= not(layer1_outputs(856));
    layer2_outputs(1354) <= not((layer1_outputs(8149)) or (layer1_outputs(4828)));
    layer2_outputs(1355) <= not(layer1_outputs(2526));
    layer2_outputs(1356) <= not(layer1_outputs(10168));
    layer2_outputs(1357) <= not(layer1_outputs(4403)) or (layer1_outputs(5954));
    layer2_outputs(1358) <= (layer1_outputs(7810)) or (layer1_outputs(7522));
    layer2_outputs(1359) <= layer1_outputs(8883);
    layer2_outputs(1360) <= (layer1_outputs(7833)) xor (layer1_outputs(310));
    layer2_outputs(1361) <= not(layer1_outputs(7768));
    layer2_outputs(1362) <= (layer1_outputs(4022)) and not (layer1_outputs(1843));
    layer2_outputs(1363) <= not(layer1_outputs(9745));
    layer2_outputs(1364) <= not(layer1_outputs(378));
    layer2_outputs(1365) <= not(layer1_outputs(8280)) or (layer1_outputs(3908));
    layer2_outputs(1366) <= layer1_outputs(1017);
    layer2_outputs(1367) <= layer1_outputs(9087);
    layer2_outputs(1368) <= not(layer1_outputs(1910));
    layer2_outputs(1369) <= layer1_outputs(2875);
    layer2_outputs(1370) <= (layer1_outputs(1732)) or (layer1_outputs(8951));
    layer2_outputs(1371) <= not((layer1_outputs(4947)) xor (layer1_outputs(211)));
    layer2_outputs(1372) <= not(layer1_outputs(4842));
    layer2_outputs(1373) <= layer1_outputs(2624);
    layer2_outputs(1374) <= not(layer1_outputs(4885));
    layer2_outputs(1375) <= layer1_outputs(8278);
    layer2_outputs(1376) <= layer1_outputs(716);
    layer2_outputs(1377) <= layer1_outputs(710);
    layer2_outputs(1378) <= layer1_outputs(6749);
    layer2_outputs(1379) <= not((layer1_outputs(9296)) and (layer1_outputs(4941)));
    layer2_outputs(1380) <= not((layer1_outputs(8161)) and (layer1_outputs(3697)));
    layer2_outputs(1381) <= not((layer1_outputs(9939)) or (layer1_outputs(9761)));
    layer2_outputs(1382) <= not((layer1_outputs(1294)) xor (layer1_outputs(5734)));
    layer2_outputs(1383) <= (layer1_outputs(8222)) xor (layer1_outputs(9984));
    layer2_outputs(1384) <= not(layer1_outputs(2057));
    layer2_outputs(1385) <= not(layer1_outputs(4194));
    layer2_outputs(1386) <= (layer1_outputs(5407)) or (layer1_outputs(6248));
    layer2_outputs(1387) <= not((layer1_outputs(4090)) or (layer1_outputs(2370)));
    layer2_outputs(1388) <= not(layer1_outputs(3566));
    layer2_outputs(1389) <= not(layer1_outputs(7538));
    layer2_outputs(1390) <= (layer1_outputs(8736)) and not (layer1_outputs(3337));
    layer2_outputs(1391) <= not(layer1_outputs(7376));
    layer2_outputs(1392) <= not(layer1_outputs(79));
    layer2_outputs(1393) <= (layer1_outputs(1150)) and not (layer1_outputs(8889));
    layer2_outputs(1394) <= not((layer1_outputs(5718)) xor (layer1_outputs(5077)));
    layer2_outputs(1395) <= layer1_outputs(3449);
    layer2_outputs(1396) <= not(layer1_outputs(6916)) or (layer1_outputs(9349));
    layer2_outputs(1397) <= not(layer1_outputs(3690));
    layer2_outputs(1398) <= layer1_outputs(4145);
    layer2_outputs(1399) <= layer1_outputs(6249);
    layer2_outputs(1400) <= layer1_outputs(9820);
    layer2_outputs(1401) <= not(layer1_outputs(3494));
    layer2_outputs(1402) <= (layer1_outputs(8788)) and not (layer1_outputs(2990));
    layer2_outputs(1403) <= layer1_outputs(2008);
    layer2_outputs(1404) <= not(layer1_outputs(9816)) or (layer1_outputs(35));
    layer2_outputs(1405) <= not(layer1_outputs(2738));
    layer2_outputs(1406) <= not(layer1_outputs(3890));
    layer2_outputs(1407) <= not((layer1_outputs(9373)) or (layer1_outputs(1382)));
    layer2_outputs(1408) <= (layer1_outputs(9688)) or (layer1_outputs(5157));
    layer2_outputs(1409) <= layer1_outputs(6785);
    layer2_outputs(1410) <= not(layer1_outputs(8224));
    layer2_outputs(1411) <= not((layer1_outputs(111)) or (layer1_outputs(9796)));
    layer2_outputs(1412) <= not(layer1_outputs(1509)) or (layer1_outputs(1193));
    layer2_outputs(1413) <= not(layer1_outputs(1816));
    layer2_outputs(1414) <= not(layer1_outputs(1979));
    layer2_outputs(1415) <= not(layer1_outputs(2623)) or (layer1_outputs(3499));
    layer2_outputs(1416) <= not(layer1_outputs(2774)) or (layer1_outputs(3187));
    layer2_outputs(1417) <= not(layer1_outputs(834)) or (layer1_outputs(5933));
    layer2_outputs(1418) <= (layer1_outputs(5659)) and not (layer1_outputs(7818));
    layer2_outputs(1419) <= not(layer1_outputs(4869)) or (layer1_outputs(8792));
    layer2_outputs(1420) <= not(layer1_outputs(171));
    layer2_outputs(1421) <= layer1_outputs(8560);
    layer2_outputs(1422) <= layer1_outputs(8832);
    layer2_outputs(1423) <= layer1_outputs(821);
    layer2_outputs(1424) <= not((layer1_outputs(802)) and (layer1_outputs(1221)));
    layer2_outputs(1425) <= (layer1_outputs(7792)) and (layer1_outputs(3784));
    layer2_outputs(1426) <= layer1_outputs(7389);
    layer2_outputs(1427) <= (layer1_outputs(3866)) and not (layer1_outputs(6058));
    layer2_outputs(1428) <= layer1_outputs(1676);
    layer2_outputs(1429) <= layer1_outputs(1776);
    layer2_outputs(1430) <= not(layer1_outputs(6550));
    layer2_outputs(1431) <= not(layer1_outputs(9191));
    layer2_outputs(1432) <= layer1_outputs(2170);
    layer2_outputs(1433) <= layer1_outputs(6090);
    layer2_outputs(1434) <= not(layer1_outputs(5858));
    layer2_outputs(1435) <= layer1_outputs(3611);
    layer2_outputs(1436) <= layer1_outputs(1970);
    layer2_outputs(1437) <= not((layer1_outputs(6612)) xor (layer1_outputs(389)));
    layer2_outputs(1438) <= not((layer1_outputs(5095)) xor (layer1_outputs(8966)));
    layer2_outputs(1439) <= (layer1_outputs(1314)) xor (layer1_outputs(5582));
    layer2_outputs(1440) <= layer1_outputs(7040);
    layer2_outputs(1441) <= layer1_outputs(5751);
    layer2_outputs(1442) <= not(layer1_outputs(5113));
    layer2_outputs(1443) <= (layer1_outputs(3676)) and not (layer1_outputs(5999));
    layer2_outputs(1444) <= layer1_outputs(3554);
    layer2_outputs(1445) <= layer1_outputs(3067);
    layer2_outputs(1446) <= not((layer1_outputs(9939)) xor (layer1_outputs(2963)));
    layer2_outputs(1447) <= (layer1_outputs(8055)) or (layer1_outputs(555));
    layer2_outputs(1448) <= layer1_outputs(2172);
    layer2_outputs(1449) <= not(layer1_outputs(4412)) or (layer1_outputs(3521));
    layer2_outputs(1450) <= not(layer1_outputs(1385));
    layer2_outputs(1451) <= not(layer1_outputs(661));
    layer2_outputs(1452) <= not(layer1_outputs(9391)) or (layer1_outputs(8242));
    layer2_outputs(1453) <= not(layer1_outputs(8595)) or (layer1_outputs(2169));
    layer2_outputs(1454) <= not(layer1_outputs(6843)) or (layer1_outputs(4524));
    layer2_outputs(1455) <= (layer1_outputs(2833)) and not (layer1_outputs(9723));
    layer2_outputs(1456) <= not(layer1_outputs(6820)) or (layer1_outputs(7420));
    layer2_outputs(1457) <= not((layer1_outputs(4729)) and (layer1_outputs(2282)));
    layer2_outputs(1458) <= not(layer1_outputs(2842));
    layer2_outputs(1459) <= layer1_outputs(9963);
    layer2_outputs(1460) <= not(layer1_outputs(10205)) or (layer1_outputs(1152));
    layer2_outputs(1461) <= not(layer1_outputs(7184));
    layer2_outputs(1462) <= layer1_outputs(7815);
    layer2_outputs(1463) <= not(layer1_outputs(6128)) or (layer1_outputs(7675));
    layer2_outputs(1464) <= (layer1_outputs(7077)) and not (layer1_outputs(7117));
    layer2_outputs(1465) <= layer1_outputs(2511);
    layer2_outputs(1466) <= not(layer1_outputs(8177));
    layer2_outputs(1467) <= layer1_outputs(2181);
    layer2_outputs(1468) <= not(layer1_outputs(3369));
    layer2_outputs(1469) <= layer1_outputs(776);
    layer2_outputs(1470) <= layer1_outputs(3768);
    layer2_outputs(1471) <= (layer1_outputs(456)) and (layer1_outputs(4331));
    layer2_outputs(1472) <= (layer1_outputs(6335)) or (layer1_outputs(8370));
    layer2_outputs(1473) <= not(layer1_outputs(3229)) or (layer1_outputs(2448));
    layer2_outputs(1474) <= layer1_outputs(8505);
    layer2_outputs(1475) <= layer1_outputs(5176);
    layer2_outputs(1476) <= (layer1_outputs(5634)) and not (layer1_outputs(4290));
    layer2_outputs(1477) <= not(layer1_outputs(2544));
    layer2_outputs(1478) <= not(layer1_outputs(363));
    layer2_outputs(1479) <= not(layer1_outputs(8473));
    layer2_outputs(1480) <= (layer1_outputs(914)) and not (layer1_outputs(6573));
    layer2_outputs(1481) <= layer1_outputs(246);
    layer2_outputs(1482) <= layer1_outputs(9518);
    layer2_outputs(1483) <= layer1_outputs(4586);
    layer2_outputs(1484) <= not((layer1_outputs(8692)) and (layer1_outputs(8163)));
    layer2_outputs(1485) <= (layer1_outputs(4718)) and (layer1_outputs(9282));
    layer2_outputs(1486) <= (layer1_outputs(8475)) xor (layer1_outputs(3536));
    layer2_outputs(1487) <= (layer1_outputs(2871)) and not (layer1_outputs(2147));
    layer2_outputs(1488) <= (layer1_outputs(878)) xor (layer1_outputs(7285));
    layer2_outputs(1489) <= not((layer1_outputs(3427)) or (layer1_outputs(4598)));
    layer2_outputs(1490) <= not((layer1_outputs(6778)) xor (layer1_outputs(7073)));
    layer2_outputs(1491) <= layer1_outputs(8112);
    layer2_outputs(1492) <= (layer1_outputs(1779)) or (layer1_outputs(5627));
    layer2_outputs(1493) <= not(layer1_outputs(7220));
    layer2_outputs(1494) <= not((layer1_outputs(6065)) xor (layer1_outputs(5523)));
    layer2_outputs(1495) <= layer1_outputs(1037);
    layer2_outputs(1496) <= not(layer1_outputs(5298));
    layer2_outputs(1497) <= (layer1_outputs(7245)) and not (layer1_outputs(3495));
    layer2_outputs(1498) <= (layer1_outputs(2554)) or (layer1_outputs(6155));
    layer2_outputs(1499) <= layer1_outputs(6727);
    layer2_outputs(1500) <= (layer1_outputs(6127)) or (layer1_outputs(6470));
    layer2_outputs(1501) <= not(layer1_outputs(5058)) or (layer1_outputs(2184));
    layer2_outputs(1502) <= (layer1_outputs(5399)) xor (layer1_outputs(6950));
    layer2_outputs(1503) <= layer1_outputs(5370);
    layer2_outputs(1504) <= not(layer1_outputs(2940));
    layer2_outputs(1505) <= (layer1_outputs(5032)) xor (layer1_outputs(6978));
    layer2_outputs(1506) <= not((layer1_outputs(7760)) or (layer1_outputs(8649)));
    layer2_outputs(1507) <= not(layer1_outputs(8948)) or (layer1_outputs(1980));
    layer2_outputs(1508) <= (layer1_outputs(2534)) or (layer1_outputs(161));
    layer2_outputs(1509) <= layer1_outputs(7107);
    layer2_outputs(1510) <= not(layer1_outputs(9346));
    layer2_outputs(1511) <= (layer1_outputs(2991)) xor (layer1_outputs(1812));
    layer2_outputs(1512) <= not(layer1_outputs(3786));
    layer2_outputs(1513) <= not(layer1_outputs(4877));
    layer2_outputs(1514) <= (layer1_outputs(6175)) and (layer1_outputs(7619));
    layer2_outputs(1515) <= layer1_outputs(9630);
    layer2_outputs(1516) <= layer1_outputs(5957);
    layer2_outputs(1517) <= not((layer1_outputs(2847)) xor (layer1_outputs(4733)));
    layer2_outputs(1518) <= not(layer1_outputs(1910));
    layer2_outputs(1519) <= not(layer1_outputs(5450));
    layer2_outputs(1520) <= (layer1_outputs(1367)) and (layer1_outputs(1745));
    layer2_outputs(1521) <= not(layer1_outputs(831));
    layer2_outputs(1522) <= layer1_outputs(2074);
    layer2_outputs(1523) <= layer1_outputs(7887);
    layer2_outputs(1524) <= (layer1_outputs(6276)) and not (layer1_outputs(4346));
    layer2_outputs(1525) <= not(layer1_outputs(3077));
    layer2_outputs(1526) <= not(layer1_outputs(7499));
    layer2_outputs(1527) <= not(layer1_outputs(1623)) or (layer1_outputs(1234));
    layer2_outputs(1528) <= (layer1_outputs(5603)) xor (layer1_outputs(302));
    layer2_outputs(1529) <= not(layer1_outputs(1568));
    layer2_outputs(1530) <= not(layer1_outputs(8300)) or (layer1_outputs(3602));
    layer2_outputs(1531) <= '0';
    layer2_outputs(1532) <= layer1_outputs(2588);
    layer2_outputs(1533) <= not(layer1_outputs(5732));
    layer2_outputs(1534) <= not(layer1_outputs(2975)) or (layer1_outputs(5353));
    layer2_outputs(1535) <= (layer1_outputs(4137)) or (layer1_outputs(65));
    layer2_outputs(1536) <= layer1_outputs(5240);
    layer2_outputs(1537) <= not(layer1_outputs(943));
    layer2_outputs(1538) <= (layer1_outputs(2029)) xor (layer1_outputs(7636));
    layer2_outputs(1539) <= not(layer1_outputs(3554));
    layer2_outputs(1540) <= (layer1_outputs(8228)) and (layer1_outputs(5983));
    layer2_outputs(1541) <= layer1_outputs(7688);
    layer2_outputs(1542) <= layer1_outputs(8169);
    layer2_outputs(1543) <= not(layer1_outputs(4818));
    layer2_outputs(1544) <= (layer1_outputs(737)) and not (layer1_outputs(1096));
    layer2_outputs(1545) <= not(layer1_outputs(3015));
    layer2_outputs(1546) <= layer1_outputs(5059);
    layer2_outputs(1547) <= not(layer1_outputs(2539));
    layer2_outputs(1548) <= not((layer1_outputs(1095)) xor (layer1_outputs(4594)));
    layer2_outputs(1549) <= (layer1_outputs(1985)) and not (layer1_outputs(7558));
    layer2_outputs(1550) <= not((layer1_outputs(9899)) xor (layer1_outputs(1617)));
    layer2_outputs(1551) <= layer1_outputs(10102);
    layer2_outputs(1552) <= (layer1_outputs(9895)) xor (layer1_outputs(3453));
    layer2_outputs(1553) <= (layer1_outputs(8603)) and (layer1_outputs(936));
    layer2_outputs(1554) <= not((layer1_outputs(6686)) and (layer1_outputs(6473)));
    layer2_outputs(1555) <= not(layer1_outputs(9036));
    layer2_outputs(1556) <= not((layer1_outputs(6331)) and (layer1_outputs(7154)));
    layer2_outputs(1557) <= not(layer1_outputs(4366)) or (layer1_outputs(3913));
    layer2_outputs(1558) <= (layer1_outputs(8563)) xor (layer1_outputs(7844));
    layer2_outputs(1559) <= (layer1_outputs(1135)) xor (layer1_outputs(9778));
    layer2_outputs(1560) <= '0';
    layer2_outputs(1561) <= (layer1_outputs(6244)) xor (layer1_outputs(3283));
    layer2_outputs(1562) <= layer1_outputs(6763);
    layer2_outputs(1563) <= not(layer1_outputs(7681));
    layer2_outputs(1564) <= not((layer1_outputs(6135)) xor (layer1_outputs(9227)));
    layer2_outputs(1565) <= not(layer1_outputs(9942));
    layer2_outputs(1566) <= not(layer1_outputs(2383));
    layer2_outputs(1567) <= not(layer1_outputs(1352));
    layer2_outputs(1568) <= layer1_outputs(108);
    layer2_outputs(1569) <= not(layer1_outputs(10002));
    layer2_outputs(1570) <= (layer1_outputs(4105)) and not (layer1_outputs(1905));
    layer2_outputs(1571) <= layer1_outputs(4367);
    layer2_outputs(1572) <= layer1_outputs(5112);
    layer2_outputs(1573) <= (layer1_outputs(9637)) and not (layer1_outputs(8024));
    layer2_outputs(1574) <= not(layer1_outputs(6682));
    layer2_outputs(1575) <= '0';
    layer2_outputs(1576) <= '0';
    layer2_outputs(1577) <= layer1_outputs(6694);
    layer2_outputs(1578) <= not((layer1_outputs(2647)) and (layer1_outputs(8183)));
    layer2_outputs(1579) <= (layer1_outputs(3423)) and not (layer1_outputs(6997));
    layer2_outputs(1580) <= not((layer1_outputs(3172)) or (layer1_outputs(5968)));
    layer2_outputs(1581) <= not(layer1_outputs(5441));
    layer2_outputs(1582) <= not(layer1_outputs(8477));
    layer2_outputs(1583) <= not(layer1_outputs(4315));
    layer2_outputs(1584) <= not(layer1_outputs(8616));
    layer2_outputs(1585) <= (layer1_outputs(5423)) and (layer1_outputs(6237));
    layer2_outputs(1586) <= not(layer1_outputs(8405)) or (layer1_outputs(593));
    layer2_outputs(1587) <= not(layer1_outputs(5004));
    layer2_outputs(1588) <= (layer1_outputs(8690)) and (layer1_outputs(7698));
    layer2_outputs(1589) <= not(layer1_outputs(425));
    layer2_outputs(1590) <= not((layer1_outputs(1199)) and (layer1_outputs(293)));
    layer2_outputs(1591) <= (layer1_outputs(5496)) and not (layer1_outputs(1459));
    layer2_outputs(1592) <= layer1_outputs(2504);
    layer2_outputs(1593) <= layer1_outputs(953);
    layer2_outputs(1594) <= layer1_outputs(522);
    layer2_outputs(1595) <= not(layer1_outputs(3107));
    layer2_outputs(1596) <= (layer1_outputs(219)) or (layer1_outputs(8435));
    layer2_outputs(1597) <= layer1_outputs(9977);
    layer2_outputs(1598) <= '0';
    layer2_outputs(1599) <= not((layer1_outputs(3782)) or (layer1_outputs(2752)));
    layer2_outputs(1600) <= not(layer1_outputs(1669)) or (layer1_outputs(2616));
    layer2_outputs(1601) <= not(layer1_outputs(7016));
    layer2_outputs(1602) <= not(layer1_outputs(4208));
    layer2_outputs(1603) <= not(layer1_outputs(686));
    layer2_outputs(1604) <= (layer1_outputs(5351)) or (layer1_outputs(8914));
    layer2_outputs(1605) <= layer1_outputs(9127);
    layer2_outputs(1606) <= (layer1_outputs(9669)) and not (layer1_outputs(3402));
    layer2_outputs(1607) <= (layer1_outputs(9670)) xor (layer1_outputs(6003));
    layer2_outputs(1608) <= not((layer1_outputs(4670)) xor (layer1_outputs(1907)));
    layer2_outputs(1609) <= (layer1_outputs(4153)) or (layer1_outputs(8217));
    layer2_outputs(1610) <= not(layer1_outputs(1258)) or (layer1_outputs(9497));
    layer2_outputs(1611) <= not((layer1_outputs(3278)) or (layer1_outputs(2414)));
    layer2_outputs(1612) <= layer1_outputs(2523);
    layer2_outputs(1613) <= layer1_outputs(4600);
    layer2_outputs(1614) <= layer1_outputs(866);
    layer2_outputs(1615) <= not(layer1_outputs(9182));
    layer2_outputs(1616) <= not(layer1_outputs(4984)) or (layer1_outputs(2419));
    layer2_outputs(1617) <= layer1_outputs(5632);
    layer2_outputs(1618) <= not((layer1_outputs(943)) or (layer1_outputs(10207)));
    layer2_outputs(1619) <= not(layer1_outputs(8630));
    layer2_outputs(1620) <= not(layer1_outputs(3425));
    layer2_outputs(1621) <= layer1_outputs(10154);
    layer2_outputs(1622) <= not(layer1_outputs(5727));
    layer2_outputs(1623) <= layer1_outputs(173);
    layer2_outputs(1624) <= (layer1_outputs(1577)) xor (layer1_outputs(7025));
    layer2_outputs(1625) <= not(layer1_outputs(8791));
    layer2_outputs(1626) <= layer1_outputs(516);
    layer2_outputs(1627) <= not(layer1_outputs(8858));
    layer2_outputs(1628) <= (layer1_outputs(4583)) xor (layer1_outputs(3777));
    layer2_outputs(1629) <= layer1_outputs(5305);
    layer2_outputs(1630) <= not(layer1_outputs(1894)) or (layer1_outputs(4811));
    layer2_outputs(1631) <= not(layer1_outputs(2739));
    layer2_outputs(1632) <= not(layer1_outputs(7351)) or (layer1_outputs(912));
    layer2_outputs(1633) <= not((layer1_outputs(4959)) or (layer1_outputs(1154)));
    layer2_outputs(1634) <= layer1_outputs(6680);
    layer2_outputs(1635) <= not((layer1_outputs(3183)) xor (layer1_outputs(3979)));
    layer2_outputs(1636) <= not((layer1_outputs(7081)) xor (layer1_outputs(9328)));
    layer2_outputs(1637) <= '1';
    layer2_outputs(1638) <= not(layer1_outputs(3029));
    layer2_outputs(1639) <= layer1_outputs(8210);
    layer2_outputs(1640) <= not((layer1_outputs(7498)) and (layer1_outputs(4396)));
    layer2_outputs(1641) <= layer1_outputs(1527);
    layer2_outputs(1642) <= layer1_outputs(6736);
    layer2_outputs(1643) <= layer1_outputs(7969);
    layer2_outputs(1644) <= layer1_outputs(8758);
    layer2_outputs(1645) <= layer1_outputs(6058);
    layer2_outputs(1646) <= layer1_outputs(9130);
    layer2_outputs(1647) <= not(layer1_outputs(2782));
    layer2_outputs(1648) <= layer1_outputs(274);
    layer2_outputs(1649) <= not(layer1_outputs(9674));
    layer2_outputs(1650) <= not(layer1_outputs(9399));
    layer2_outputs(1651) <= layer1_outputs(5908);
    layer2_outputs(1652) <= layer1_outputs(9248);
    layer2_outputs(1653) <= not(layer1_outputs(207));
    layer2_outputs(1654) <= (layer1_outputs(1967)) xor (layer1_outputs(1592));
    layer2_outputs(1655) <= not((layer1_outputs(1993)) xor (layer1_outputs(9846)));
    layer2_outputs(1656) <= not(layer1_outputs(922));
    layer2_outputs(1657) <= layer1_outputs(7082);
    layer2_outputs(1658) <= layer1_outputs(2041);
    layer2_outputs(1659) <= layer1_outputs(5507);
    layer2_outputs(1660) <= layer1_outputs(9318);
    layer2_outputs(1661) <= not(layer1_outputs(2375));
    layer2_outputs(1662) <= not(layer1_outputs(6123));
    layer2_outputs(1663) <= not(layer1_outputs(6486)) or (layer1_outputs(1233));
    layer2_outputs(1664) <= not(layer1_outputs(2788));
    layer2_outputs(1665) <= (layer1_outputs(4741)) and not (layer1_outputs(2742));
    layer2_outputs(1666) <= layer1_outputs(10072);
    layer2_outputs(1667) <= layer1_outputs(1111);
    layer2_outputs(1668) <= not(layer1_outputs(9204));
    layer2_outputs(1669) <= layer1_outputs(4684);
    layer2_outputs(1670) <= not(layer1_outputs(946));
    layer2_outputs(1671) <= not((layer1_outputs(1360)) and (layer1_outputs(8890)));
    layer2_outputs(1672) <= layer1_outputs(7315);
    layer2_outputs(1673) <= not(layer1_outputs(8214)) or (layer1_outputs(2495));
    layer2_outputs(1674) <= layer1_outputs(9963);
    layer2_outputs(1675) <= (layer1_outputs(8112)) and (layer1_outputs(3253));
    layer2_outputs(1676) <= not(layer1_outputs(1660)) or (layer1_outputs(8803));
    layer2_outputs(1677) <= layer1_outputs(2187);
    layer2_outputs(1678) <= (layer1_outputs(9777)) and (layer1_outputs(5459));
    layer2_outputs(1679) <= not(layer1_outputs(9366)) or (layer1_outputs(144));
    layer2_outputs(1680) <= (layer1_outputs(4542)) xor (layer1_outputs(7188));
    layer2_outputs(1681) <= not(layer1_outputs(8208));
    layer2_outputs(1682) <= (layer1_outputs(8252)) and (layer1_outputs(8996));
    layer2_outputs(1683) <= not((layer1_outputs(6645)) xor (layer1_outputs(3474)));
    layer2_outputs(1684) <= not(layer1_outputs(9798)) or (layer1_outputs(8189));
    layer2_outputs(1685) <= not(layer1_outputs(5352));
    layer2_outputs(1686) <= not((layer1_outputs(1747)) xor (layer1_outputs(2023)));
    layer2_outputs(1687) <= not(layer1_outputs(8232));
    layer2_outputs(1688) <= (layer1_outputs(5809)) and not (layer1_outputs(4400));
    layer2_outputs(1689) <= not(layer1_outputs(1661));
    layer2_outputs(1690) <= layer1_outputs(4299);
    layer2_outputs(1691) <= not((layer1_outputs(3194)) xor (layer1_outputs(2618)));
    layer2_outputs(1692) <= not((layer1_outputs(9282)) xor (layer1_outputs(4678)));
    layer2_outputs(1693) <= not(layer1_outputs(5062));
    layer2_outputs(1694) <= (layer1_outputs(9034)) and not (layer1_outputs(3296));
    layer2_outputs(1695) <= (layer1_outputs(3265)) and not (layer1_outputs(8342));
    layer2_outputs(1696) <= not((layer1_outputs(8431)) or (layer1_outputs(7324)));
    layer2_outputs(1697) <= not(layer1_outputs(2087));
    layer2_outputs(1698) <= not(layer1_outputs(5890));
    layer2_outputs(1699) <= (layer1_outputs(5341)) and (layer1_outputs(3981));
    layer2_outputs(1700) <= not(layer1_outputs(3878));
    layer2_outputs(1701) <= not(layer1_outputs(730)) or (layer1_outputs(6760));
    layer2_outputs(1702) <= layer1_outputs(9331);
    layer2_outputs(1703) <= layer1_outputs(8773);
    layer2_outputs(1704) <= not(layer1_outputs(1831));
    layer2_outputs(1705) <= layer1_outputs(9542);
    layer2_outputs(1706) <= not((layer1_outputs(1027)) xor (layer1_outputs(8003)));
    layer2_outputs(1707) <= not((layer1_outputs(6126)) xor (layer1_outputs(4318)));
    layer2_outputs(1708) <= not(layer1_outputs(142));
    layer2_outputs(1709) <= (layer1_outputs(3218)) and not (layer1_outputs(6917));
    layer2_outputs(1710) <= (layer1_outputs(9933)) and not (layer1_outputs(4019));
    layer2_outputs(1711) <= (layer1_outputs(7641)) and (layer1_outputs(8590));
    layer2_outputs(1712) <= (layer1_outputs(6879)) and not (layer1_outputs(2432));
    layer2_outputs(1713) <= (layer1_outputs(3047)) and not (layer1_outputs(1556));
    layer2_outputs(1714) <= layer1_outputs(4463);
    layer2_outputs(1715) <= layer1_outputs(4231);
    layer2_outputs(1716) <= not(layer1_outputs(7826));
    layer2_outputs(1717) <= not(layer1_outputs(7696));
    layer2_outputs(1718) <= not(layer1_outputs(3720));
    layer2_outputs(1719) <= (layer1_outputs(2992)) or (layer1_outputs(5452));
    layer2_outputs(1720) <= not((layer1_outputs(10152)) or (layer1_outputs(1018)));
    layer2_outputs(1721) <= not((layer1_outputs(5648)) xor (layer1_outputs(7568)));
    layer2_outputs(1722) <= not((layer1_outputs(2652)) or (layer1_outputs(7461)));
    layer2_outputs(1723) <= not(layer1_outputs(6002));
    layer2_outputs(1724) <= layer1_outputs(6324);
    layer2_outputs(1725) <= layer1_outputs(1005);
    layer2_outputs(1726) <= (layer1_outputs(2017)) and (layer1_outputs(7966));
    layer2_outputs(1727) <= not(layer1_outputs(1824));
    layer2_outputs(1728) <= (layer1_outputs(9421)) and not (layer1_outputs(1814));
    layer2_outputs(1729) <= not((layer1_outputs(6983)) xor (layer1_outputs(1711)));
    layer2_outputs(1730) <= layer1_outputs(1184);
    layer2_outputs(1731) <= not(layer1_outputs(1556)) or (layer1_outputs(3553));
    layer2_outputs(1732) <= layer1_outputs(334);
    layer2_outputs(1733) <= not(layer1_outputs(84));
    layer2_outputs(1734) <= (layer1_outputs(4794)) or (layer1_outputs(5231));
    layer2_outputs(1735) <= (layer1_outputs(1173)) and (layer1_outputs(7364));
    layer2_outputs(1736) <= not(layer1_outputs(224)) or (layer1_outputs(2399));
    layer2_outputs(1737) <= not(layer1_outputs(738));
    layer2_outputs(1738) <= not(layer1_outputs(7832)) or (layer1_outputs(1420));
    layer2_outputs(1739) <= not(layer1_outputs(3984)) or (layer1_outputs(9395));
    layer2_outputs(1740) <= layer1_outputs(5871);
    layer2_outputs(1741) <= (layer1_outputs(2354)) or (layer1_outputs(5301));
    layer2_outputs(1742) <= not(layer1_outputs(6816));
    layer2_outputs(1743) <= not(layer1_outputs(605));
    layer2_outputs(1744) <= layer1_outputs(6264);
    layer2_outputs(1745) <= not(layer1_outputs(393));
    layer2_outputs(1746) <= not(layer1_outputs(1312)) or (layer1_outputs(9428));
    layer2_outputs(1747) <= (layer1_outputs(841)) or (layer1_outputs(7801));
    layer2_outputs(1748) <= not((layer1_outputs(5369)) or (layer1_outputs(5880)));
    layer2_outputs(1749) <= layer1_outputs(4325);
    layer2_outputs(1750) <= (layer1_outputs(7793)) or (layer1_outputs(5261));
    layer2_outputs(1751) <= not(layer1_outputs(10115));
    layer2_outputs(1752) <= layer1_outputs(1647);
    layer2_outputs(1753) <= '0';
    layer2_outputs(1754) <= not(layer1_outputs(5937)) or (layer1_outputs(201));
    layer2_outputs(1755) <= (layer1_outputs(9978)) or (layer1_outputs(4801));
    layer2_outputs(1756) <= not(layer1_outputs(9519));
    layer2_outputs(1757) <= not(layer1_outputs(5288));
    layer2_outputs(1758) <= layer1_outputs(3056);
    layer2_outputs(1759) <= (layer1_outputs(9581)) or (layer1_outputs(4305));
    layer2_outputs(1760) <= (layer1_outputs(3846)) and (layer1_outputs(631));
    layer2_outputs(1761) <= not(layer1_outputs(8287));
    layer2_outputs(1762) <= not(layer1_outputs(366));
    layer2_outputs(1763) <= not(layer1_outputs(8375));
    layer2_outputs(1764) <= not(layer1_outputs(2246)) or (layer1_outputs(6156));
    layer2_outputs(1765) <= layer1_outputs(1483);
    layer2_outputs(1766) <= not(layer1_outputs(6520));
    layer2_outputs(1767) <= not(layer1_outputs(6874));
    layer2_outputs(1768) <= layer1_outputs(5544);
    layer2_outputs(1769) <= (layer1_outputs(10175)) xor (layer1_outputs(6950));
    layer2_outputs(1770) <= (layer1_outputs(7111)) and (layer1_outputs(4598));
    layer2_outputs(1771) <= not(layer1_outputs(1180));
    layer2_outputs(1772) <= not(layer1_outputs(7935));
    layer2_outputs(1773) <= not(layer1_outputs(9879));
    layer2_outputs(1774) <= layer1_outputs(4040);
    layer2_outputs(1775) <= (layer1_outputs(5670)) and not (layer1_outputs(637));
    layer2_outputs(1776) <= not((layer1_outputs(3802)) xor (layer1_outputs(442)));
    layer2_outputs(1777) <= not((layer1_outputs(5795)) and (layer1_outputs(3106)));
    layer2_outputs(1778) <= not(layer1_outputs(651));
    layer2_outputs(1779) <= not(layer1_outputs(4681)) or (layer1_outputs(9061));
    layer2_outputs(1780) <= not(layer1_outputs(7250));
    layer2_outputs(1781) <= not(layer1_outputs(9491));
    layer2_outputs(1782) <= layer1_outputs(6001);
    layer2_outputs(1783) <= not(layer1_outputs(3291));
    layer2_outputs(1784) <= (layer1_outputs(4334)) and (layer1_outputs(1428));
    layer2_outputs(1785) <= not(layer1_outputs(9443));
    layer2_outputs(1786) <= layer1_outputs(6349);
    layer2_outputs(1787) <= (layer1_outputs(2254)) and not (layer1_outputs(5416));
    layer2_outputs(1788) <= not((layer1_outputs(3292)) xor (layer1_outputs(6696)));
    layer2_outputs(1789) <= not(layer1_outputs(4742));
    layer2_outputs(1790) <= layer1_outputs(155);
    layer2_outputs(1791) <= (layer1_outputs(4266)) and (layer1_outputs(7805));
    layer2_outputs(1792) <= (layer1_outputs(1522)) and not (layer1_outputs(8009));
    layer2_outputs(1793) <= layer1_outputs(8952);
    layer2_outputs(1794) <= layer1_outputs(7059);
    layer2_outputs(1795) <= (layer1_outputs(8156)) and (layer1_outputs(7294));
    layer2_outputs(1796) <= (layer1_outputs(9219)) and not (layer1_outputs(8246));
    layer2_outputs(1797) <= layer1_outputs(3804);
    layer2_outputs(1798) <= layer1_outputs(8678);
    layer2_outputs(1799) <= layer1_outputs(2836);
    layer2_outputs(1800) <= (layer1_outputs(8744)) and (layer1_outputs(4343));
    layer2_outputs(1801) <= layer1_outputs(4270);
    layer2_outputs(1802) <= not(layer1_outputs(7344));
    layer2_outputs(1803) <= layer1_outputs(897);
    layer2_outputs(1804) <= layer1_outputs(813);
    layer2_outputs(1805) <= layer1_outputs(1029);
    layer2_outputs(1806) <= (layer1_outputs(4549)) xor (layer1_outputs(7505));
    layer2_outputs(1807) <= not((layer1_outputs(10208)) xor (layer1_outputs(3947)));
    layer2_outputs(1808) <= not(layer1_outputs(1947));
    layer2_outputs(1809) <= (layer1_outputs(6739)) and (layer1_outputs(7298));
    layer2_outputs(1810) <= (layer1_outputs(3072)) and not (layer1_outputs(2855));
    layer2_outputs(1811) <= not((layer1_outputs(2001)) and (layer1_outputs(3435)));
    layer2_outputs(1812) <= (layer1_outputs(2387)) and (layer1_outputs(7014));
    layer2_outputs(1813) <= layer1_outputs(630);
    layer2_outputs(1814) <= not(layer1_outputs(9828));
    layer2_outputs(1815) <= layer1_outputs(5464);
    layer2_outputs(1816) <= layer1_outputs(4979);
    layer2_outputs(1817) <= layer1_outputs(5257);
    layer2_outputs(1818) <= '0';
    layer2_outputs(1819) <= not(layer1_outputs(4020));
    layer2_outputs(1820) <= layer1_outputs(91);
    layer2_outputs(1821) <= layer1_outputs(4603);
    layer2_outputs(1822) <= layer1_outputs(9641);
    layer2_outputs(1823) <= (layer1_outputs(3745)) and not (layer1_outputs(5664));
    layer2_outputs(1824) <= not((layer1_outputs(9772)) or (layer1_outputs(740)));
    layer2_outputs(1825) <= layer1_outputs(1285);
    layer2_outputs(1826) <= layer1_outputs(6337);
    layer2_outputs(1827) <= (layer1_outputs(6576)) xor (layer1_outputs(10044));
    layer2_outputs(1828) <= not((layer1_outputs(10009)) or (layer1_outputs(2513)));
    layer2_outputs(1829) <= not(layer1_outputs(588));
    layer2_outputs(1830) <= (layer1_outputs(2196)) and not (layer1_outputs(5410));
    layer2_outputs(1831) <= not(layer1_outputs(2695)) or (layer1_outputs(1827));
    layer2_outputs(1832) <= layer1_outputs(4583);
    layer2_outputs(1833) <= (layer1_outputs(8430)) and not (layer1_outputs(6453));
    layer2_outputs(1834) <= layer1_outputs(8492);
    layer2_outputs(1835) <= not(layer1_outputs(1132));
    layer2_outputs(1836) <= not((layer1_outputs(5710)) or (layer1_outputs(4651)));
    layer2_outputs(1837) <= (layer1_outputs(6115)) and not (layer1_outputs(142));
    layer2_outputs(1838) <= (layer1_outputs(4574)) and not (layer1_outputs(5299));
    layer2_outputs(1839) <= not(layer1_outputs(1427)) or (layer1_outputs(2208));
    layer2_outputs(1840) <= layer1_outputs(3866);
    layer2_outputs(1841) <= (layer1_outputs(9791)) and (layer1_outputs(4769));
    layer2_outputs(1842) <= not((layer1_outputs(4157)) or (layer1_outputs(10144)));
    layer2_outputs(1843) <= not(layer1_outputs(167));
    layer2_outputs(1844) <= not(layer1_outputs(1650));
    layer2_outputs(1845) <= (layer1_outputs(4167)) and not (layer1_outputs(1839));
    layer2_outputs(1846) <= (layer1_outputs(386)) or (layer1_outputs(6034));
    layer2_outputs(1847) <= not(layer1_outputs(4877));
    layer2_outputs(1848) <= not(layer1_outputs(4369));
    layer2_outputs(1849) <= (layer1_outputs(9097)) xor (layer1_outputs(10140));
    layer2_outputs(1850) <= layer1_outputs(8424);
    layer2_outputs(1851) <= not(layer1_outputs(2987));
    layer2_outputs(1852) <= (layer1_outputs(9083)) and not (layer1_outputs(9922));
    layer2_outputs(1853) <= not((layer1_outputs(1594)) xor (layer1_outputs(5924)));
    layer2_outputs(1854) <= not(layer1_outputs(4730));
    layer2_outputs(1855) <= not(layer1_outputs(6962));
    layer2_outputs(1856) <= not(layer1_outputs(7607));
    layer2_outputs(1857) <= not((layer1_outputs(10229)) xor (layer1_outputs(580)));
    layer2_outputs(1858) <= (layer1_outputs(6203)) and not (layer1_outputs(6980));
    layer2_outputs(1859) <= (layer1_outputs(714)) xor (layer1_outputs(4061));
    layer2_outputs(1860) <= layer1_outputs(6136);
    layer2_outputs(1861) <= (layer1_outputs(6139)) or (layer1_outputs(8588));
    layer2_outputs(1862) <= '1';
    layer2_outputs(1863) <= layer1_outputs(5979);
    layer2_outputs(1864) <= (layer1_outputs(597)) and (layer1_outputs(3082));
    layer2_outputs(1865) <= (layer1_outputs(6321)) and not (layer1_outputs(7808));
    layer2_outputs(1866) <= not(layer1_outputs(2309)) or (layer1_outputs(8497));
    layer2_outputs(1867) <= layer1_outputs(4538);
    layer2_outputs(1868) <= not(layer1_outputs(5542));
    layer2_outputs(1869) <= (layer1_outputs(5322)) xor (layer1_outputs(9763));
    layer2_outputs(1870) <= (layer1_outputs(1372)) and not (layer1_outputs(9121));
    layer2_outputs(1871) <= layer1_outputs(10001);
    layer2_outputs(1872) <= layer1_outputs(158);
    layer2_outputs(1873) <= layer1_outputs(63);
    layer2_outputs(1874) <= layer1_outputs(1024);
    layer2_outputs(1875) <= not(layer1_outputs(4658));
    layer2_outputs(1876) <= (layer1_outputs(3305)) or (layer1_outputs(6322));
    layer2_outputs(1877) <= (layer1_outputs(5025)) and not (layer1_outputs(7395));
    layer2_outputs(1878) <= (layer1_outputs(4464)) or (layer1_outputs(4759));
    layer2_outputs(1879) <= layer1_outputs(3958);
    layer2_outputs(1880) <= (layer1_outputs(1484)) xor (layer1_outputs(9413));
    layer2_outputs(1881) <= layer1_outputs(10121);
    layer2_outputs(1882) <= not(layer1_outputs(3587));
    layer2_outputs(1883) <= (layer1_outputs(3959)) and (layer1_outputs(9026));
    layer2_outputs(1884) <= not((layer1_outputs(4787)) xor (layer1_outputs(3473)));
    layer2_outputs(1885) <= layer1_outputs(2201);
    layer2_outputs(1886) <= not((layer1_outputs(4414)) and (layer1_outputs(975)));
    layer2_outputs(1887) <= not(layer1_outputs(2962));
    layer2_outputs(1888) <= not((layer1_outputs(8336)) xor (layer1_outputs(5550)));
    layer2_outputs(1889) <= (layer1_outputs(9160)) and not (layer1_outputs(6233));
    layer2_outputs(1890) <= not((layer1_outputs(4969)) xor (layer1_outputs(6675)));
    layer2_outputs(1891) <= not((layer1_outputs(6105)) or (layer1_outputs(8171)));
    layer2_outputs(1892) <= (layer1_outputs(5115)) and not (layer1_outputs(1333));
    layer2_outputs(1893) <= (layer1_outputs(4373)) xor (layer1_outputs(6413));
    layer2_outputs(1894) <= not(layer1_outputs(6084)) or (layer1_outputs(8689));
    layer2_outputs(1895) <= layer1_outputs(962);
    layer2_outputs(1896) <= (layer1_outputs(6258)) xor (layer1_outputs(9887));
    layer2_outputs(1897) <= (layer1_outputs(3133)) and not (layer1_outputs(7549));
    layer2_outputs(1898) <= not(layer1_outputs(441));
    layer2_outputs(1899) <= layer1_outputs(7021);
    layer2_outputs(1900) <= layer1_outputs(9560);
    layer2_outputs(1901) <= (layer1_outputs(4827)) and not (layer1_outputs(2314));
    layer2_outputs(1902) <= not(layer1_outputs(6290));
    layer2_outputs(1903) <= not((layer1_outputs(6598)) and (layer1_outputs(4169)));
    layer2_outputs(1904) <= layer1_outputs(5393);
    layer2_outputs(1905) <= layer1_outputs(10142);
    layer2_outputs(1906) <= (layer1_outputs(8967)) xor (layer1_outputs(507));
    layer2_outputs(1907) <= not(layer1_outputs(10173));
    layer2_outputs(1908) <= not(layer1_outputs(10165));
    layer2_outputs(1909) <= layer1_outputs(4783);
    layer2_outputs(1910) <= (layer1_outputs(4393)) and (layer1_outputs(4478));
    layer2_outputs(1911) <= layer1_outputs(9754);
    layer2_outputs(1912) <= not((layer1_outputs(7472)) xor (layer1_outputs(7301)));
    layer2_outputs(1913) <= not((layer1_outputs(345)) or (layer1_outputs(4467)));
    layer2_outputs(1914) <= (layer1_outputs(10109)) and not (layer1_outputs(4182));
    layer2_outputs(1915) <= layer1_outputs(750);
    layer2_outputs(1916) <= not((layer1_outputs(3285)) xor (layer1_outputs(7765)));
    layer2_outputs(1917) <= layer1_outputs(9459);
    layer2_outputs(1918) <= layer1_outputs(6288);
    layer2_outputs(1919) <= not((layer1_outputs(1653)) and (layer1_outputs(6195)));
    layer2_outputs(1920) <= (layer1_outputs(618)) and not (layer1_outputs(2464));
    layer2_outputs(1921) <= layer1_outputs(9601);
    layer2_outputs(1922) <= not(layer1_outputs(2250));
    layer2_outputs(1923) <= not(layer1_outputs(10051));
    layer2_outputs(1924) <= not(layer1_outputs(9965)) or (layer1_outputs(536));
    layer2_outputs(1925) <= not((layer1_outputs(7157)) xor (layer1_outputs(6283)));
    layer2_outputs(1926) <= layer1_outputs(4884);
    layer2_outputs(1927) <= not(layer1_outputs(5859));
    layer2_outputs(1928) <= (layer1_outputs(5636)) and (layer1_outputs(2745));
    layer2_outputs(1929) <= layer1_outputs(3549);
    layer2_outputs(1930) <= not(layer1_outputs(8347));
    layer2_outputs(1931) <= not(layer1_outputs(6634));
    layer2_outputs(1932) <= (layer1_outputs(2347)) and not (layer1_outputs(1946));
    layer2_outputs(1933) <= not(layer1_outputs(662));
    layer2_outputs(1934) <= (layer1_outputs(8692)) xor (layer1_outputs(7186));
    layer2_outputs(1935) <= (layer1_outputs(9074)) or (layer1_outputs(1811));
    layer2_outputs(1936) <= not((layer1_outputs(2978)) and (layer1_outputs(9847)));
    layer2_outputs(1937) <= not(layer1_outputs(8946));
    layer2_outputs(1938) <= (layer1_outputs(311)) and (layer1_outputs(624));
    layer2_outputs(1939) <= (layer1_outputs(9723)) xor (layer1_outputs(8323));
    layer2_outputs(1940) <= (layer1_outputs(886)) and not (layer1_outputs(5652));
    layer2_outputs(1941) <= layer1_outputs(1961);
    layer2_outputs(1942) <= not(layer1_outputs(8742)) or (layer1_outputs(1641));
    layer2_outputs(1943) <= layer1_outputs(3778);
    layer2_outputs(1944) <= (layer1_outputs(4640)) or (layer1_outputs(2933));
    layer2_outputs(1945) <= layer1_outputs(6220);
    layer2_outputs(1946) <= not(layer1_outputs(3452)) or (layer1_outputs(466));
    layer2_outputs(1947) <= not(layer1_outputs(226));
    layer2_outputs(1948) <= not(layer1_outputs(9422));
    layer2_outputs(1949) <= layer1_outputs(3917);
    layer2_outputs(1950) <= not(layer1_outputs(2375)) or (layer1_outputs(8834));
    layer2_outputs(1951) <= not((layer1_outputs(2445)) xor (layer1_outputs(4285)));
    layer2_outputs(1952) <= not(layer1_outputs(952));
    layer2_outputs(1953) <= (layer1_outputs(777)) and not (layer1_outputs(3349));
    layer2_outputs(1954) <= not((layer1_outputs(9004)) or (layer1_outputs(5417)));
    layer2_outputs(1955) <= not((layer1_outputs(7015)) or (layer1_outputs(7908)));
    layer2_outputs(1956) <= not(layer1_outputs(2061));
    layer2_outputs(1957) <= layer1_outputs(9933);
    layer2_outputs(1958) <= not(layer1_outputs(2385)) or (layer1_outputs(793));
    layer2_outputs(1959) <= (layer1_outputs(7857)) xor (layer1_outputs(4370));
    layer2_outputs(1960) <= not((layer1_outputs(4553)) or (layer1_outputs(3251)));
    layer2_outputs(1961) <= (layer1_outputs(9130)) or (layer1_outputs(5277));
    layer2_outputs(1962) <= layer1_outputs(1807);
    layer2_outputs(1963) <= not(layer1_outputs(2143));
    layer2_outputs(1964) <= layer1_outputs(6788);
    layer2_outputs(1965) <= (layer1_outputs(3362)) xor (layer1_outputs(2905));
    layer2_outputs(1966) <= layer1_outputs(209);
    layer2_outputs(1967) <= not(layer1_outputs(9461)) or (layer1_outputs(4989));
    layer2_outputs(1968) <= not(layer1_outputs(9604));
    layer2_outputs(1969) <= (layer1_outputs(2750)) and not (layer1_outputs(2609));
    layer2_outputs(1970) <= layer1_outputs(4324);
    layer2_outputs(1971) <= not(layer1_outputs(3080));
    layer2_outputs(1972) <= not((layer1_outputs(1163)) or (layer1_outputs(3547)));
    layer2_outputs(1973) <= layer1_outputs(2885);
    layer2_outputs(1974) <= not(layer1_outputs(8624));
    layer2_outputs(1975) <= not(layer1_outputs(131));
    layer2_outputs(1976) <= (layer1_outputs(1224)) and not (layer1_outputs(8668));
    layer2_outputs(1977) <= not(layer1_outputs(5221));
    layer2_outputs(1978) <= (layer1_outputs(5251)) or (layer1_outputs(3776));
    layer2_outputs(1979) <= not(layer1_outputs(6947)) or (layer1_outputs(8809));
    layer2_outputs(1980) <= (layer1_outputs(4743)) and (layer1_outputs(2506));
    layer2_outputs(1981) <= layer1_outputs(8218);
    layer2_outputs(1982) <= not(layer1_outputs(8874)) or (layer1_outputs(5017));
    layer2_outputs(1983) <= not(layer1_outputs(6569));
    layer2_outputs(1984) <= (layer1_outputs(7327)) and not (layer1_outputs(9185));
    layer2_outputs(1985) <= not(layer1_outputs(8842)) or (layer1_outputs(8429));
    layer2_outputs(1986) <= layer1_outputs(9889);
    layer2_outputs(1987) <= not((layer1_outputs(6823)) or (layer1_outputs(4779)));
    layer2_outputs(1988) <= not(layer1_outputs(5080));
    layer2_outputs(1989) <= layer1_outputs(3787);
    layer2_outputs(1990) <= not((layer1_outputs(3876)) and (layer1_outputs(3498)));
    layer2_outputs(1991) <= not(layer1_outputs(6138));
    layer2_outputs(1992) <= (layer1_outputs(1296)) and not (layer1_outputs(4311));
    layer2_outputs(1993) <= layer1_outputs(4175);
    layer2_outputs(1994) <= layer1_outputs(501);
    layer2_outputs(1995) <= not((layer1_outputs(240)) and (layer1_outputs(4763)));
    layer2_outputs(1996) <= not(layer1_outputs(1139));
    layer2_outputs(1997) <= not(layer1_outputs(5592));
    layer2_outputs(1998) <= layer1_outputs(2872);
    layer2_outputs(1999) <= (layer1_outputs(3578)) and not (layer1_outputs(3513));
    layer2_outputs(2000) <= layer1_outputs(5764);
    layer2_outputs(2001) <= (layer1_outputs(4465)) or (layer1_outputs(4));
    layer2_outputs(2002) <= layer1_outputs(2581);
    layer2_outputs(2003) <= not(layer1_outputs(7962));
    layer2_outputs(2004) <= not(layer1_outputs(3507));
    layer2_outputs(2005) <= not(layer1_outputs(562));
    layer2_outputs(2006) <= not(layer1_outputs(8042));
    layer2_outputs(2007) <= (layer1_outputs(2423)) xor (layer1_outputs(744));
    layer2_outputs(2008) <= not((layer1_outputs(3029)) or (layer1_outputs(9471)));
    layer2_outputs(2009) <= (layer1_outputs(3217)) and not (layer1_outputs(7143));
    layer2_outputs(2010) <= layer1_outputs(7753);
    layer2_outputs(2011) <= (layer1_outputs(3205)) and (layer1_outputs(7186));
    layer2_outputs(2012) <= (layer1_outputs(7924)) and not (layer1_outputs(7325));
    layer2_outputs(2013) <= layer1_outputs(2516);
    layer2_outputs(2014) <= not((layer1_outputs(7897)) or (layer1_outputs(4243)));
    layer2_outputs(2015) <= not((layer1_outputs(2793)) and (layer1_outputs(3357)));
    layer2_outputs(2016) <= layer1_outputs(10063);
    layer2_outputs(2017) <= not(layer1_outputs(8695));
    layer2_outputs(2018) <= not((layer1_outputs(2957)) xor (layer1_outputs(8307)));
    layer2_outputs(2019) <= layer1_outputs(7563);
    layer2_outputs(2020) <= layer1_outputs(3414);
    layer2_outputs(2021) <= not(layer1_outputs(9599));
    layer2_outputs(2022) <= not(layer1_outputs(9093));
    layer2_outputs(2023) <= layer1_outputs(10004);
    layer2_outputs(2024) <= (layer1_outputs(3009)) xor (layer1_outputs(247));
    layer2_outputs(2025) <= not(layer1_outputs(3677));
    layer2_outputs(2026) <= not(layer1_outputs(2874)) or (layer1_outputs(3980));
    layer2_outputs(2027) <= not(layer1_outputs(5109));
    layer2_outputs(2028) <= not(layer1_outputs(8443));
    layer2_outputs(2029) <= layer1_outputs(3654);
    layer2_outputs(2030) <= not(layer1_outputs(5365));
    layer2_outputs(2031) <= layer1_outputs(4070);
    layer2_outputs(2032) <= not((layer1_outputs(2502)) xor (layer1_outputs(5955)));
    layer2_outputs(2033) <= (layer1_outputs(6799)) and not (layer1_outputs(7701));
    layer2_outputs(2034) <= layer1_outputs(7402);
    layer2_outputs(2035) <= not(layer1_outputs(5831));
    layer2_outputs(2036) <= not((layer1_outputs(972)) xor (layer1_outputs(628)));
    layer2_outputs(2037) <= layer1_outputs(10072);
    layer2_outputs(2038) <= layer1_outputs(6942);
    layer2_outputs(2039) <= not(layer1_outputs(892)) or (layer1_outputs(2586));
    layer2_outputs(2040) <= not(layer1_outputs(2124));
    layer2_outputs(2041) <= (layer1_outputs(4057)) and not (layer1_outputs(8339));
    layer2_outputs(2042) <= layer1_outputs(2845);
    layer2_outputs(2043) <= not((layer1_outputs(4502)) and (layer1_outputs(3690)));
    layer2_outputs(2044) <= (layer1_outputs(2977)) and (layer1_outputs(8968));
    layer2_outputs(2045) <= layer1_outputs(8930);
    layer2_outputs(2046) <= (layer1_outputs(1056)) and (layer1_outputs(1817));
    layer2_outputs(2047) <= not((layer1_outputs(6190)) and (layer1_outputs(7771)));
    layer2_outputs(2048) <= (layer1_outputs(9511)) and not (layer1_outputs(2391));
    layer2_outputs(2049) <= layer1_outputs(1620);
    layer2_outputs(2050) <= not(layer1_outputs(9032));
    layer2_outputs(2051) <= '1';
    layer2_outputs(2052) <= not(layer1_outputs(8544));
    layer2_outputs(2053) <= (layer1_outputs(3365)) and (layer1_outputs(7974));
    layer2_outputs(2054) <= layer1_outputs(1871);
    layer2_outputs(2055) <= layer1_outputs(2309);
    layer2_outputs(2056) <= not(layer1_outputs(5992)) or (layer1_outputs(2973));
    layer2_outputs(2057) <= (layer1_outputs(5307)) or (layer1_outputs(4695));
    layer2_outputs(2058) <= not(layer1_outputs(9576)) or (layer1_outputs(3927));
    layer2_outputs(2059) <= (layer1_outputs(5520)) xor (layer1_outputs(495));
    layer2_outputs(2060) <= not(layer1_outputs(6270));
    layer2_outputs(2061) <= (layer1_outputs(2854)) and not (layer1_outputs(452));
    layer2_outputs(2062) <= layer1_outputs(3381);
    layer2_outputs(2063) <= layer1_outputs(5127);
    layer2_outputs(2064) <= not(layer1_outputs(1823));
    layer2_outputs(2065) <= not(layer1_outputs(5764));
    layer2_outputs(2066) <= not((layer1_outputs(629)) and (layer1_outputs(3648)));
    layer2_outputs(2067) <= not(layer1_outputs(9348));
    layer2_outputs(2068) <= layer1_outputs(9515);
    layer2_outputs(2069) <= not(layer1_outputs(3430));
    layer2_outputs(2070) <= (layer1_outputs(2953)) or (layer1_outputs(2401));
    layer2_outputs(2071) <= (layer1_outputs(4171)) and not (layer1_outputs(6941));
    layer2_outputs(2072) <= (layer1_outputs(8160)) or (layer1_outputs(3018));
    layer2_outputs(2073) <= layer1_outputs(5308);
    layer2_outputs(2074) <= not(layer1_outputs(4487)) or (layer1_outputs(1400));
    layer2_outputs(2075) <= not(layer1_outputs(1516));
    layer2_outputs(2076) <= not((layer1_outputs(7316)) xor (layer1_outputs(5702)));
    layer2_outputs(2077) <= not((layer1_outputs(5478)) and (layer1_outputs(4781)));
    layer2_outputs(2078) <= not((layer1_outputs(1976)) and (layer1_outputs(7265)));
    layer2_outputs(2079) <= (layer1_outputs(6730)) or (layer1_outputs(7923));
    layer2_outputs(2080) <= layer1_outputs(4902);
    layer2_outputs(2081) <= layer1_outputs(9346);
    layer2_outputs(2082) <= not((layer1_outputs(8358)) xor (layer1_outputs(1306)));
    layer2_outputs(2083) <= not(layer1_outputs(9350));
    layer2_outputs(2084) <= layer1_outputs(7929);
    layer2_outputs(2085) <= layer1_outputs(7536);
    layer2_outputs(2086) <= (layer1_outputs(4202)) and not (layer1_outputs(5700));
    layer2_outputs(2087) <= (layer1_outputs(7208)) and not (layer1_outputs(4293));
    layer2_outputs(2088) <= layer1_outputs(295);
    layer2_outputs(2089) <= layer1_outputs(4353);
    layer2_outputs(2090) <= not((layer1_outputs(2253)) and (layer1_outputs(6230)));
    layer2_outputs(2091) <= not((layer1_outputs(9844)) and (layer1_outputs(5758)));
    layer2_outputs(2092) <= not(layer1_outputs(3384)) or (layer1_outputs(2664));
    layer2_outputs(2093) <= layer1_outputs(821);
    layer2_outputs(2094) <= not(layer1_outputs(540));
    layer2_outputs(2095) <= not(layer1_outputs(3040));
    layer2_outputs(2096) <= layer1_outputs(3233);
    layer2_outputs(2097) <= layer1_outputs(3051);
    layer2_outputs(2098) <= not((layer1_outputs(8257)) or (layer1_outputs(8966)));
    layer2_outputs(2099) <= layer1_outputs(2392);
    layer2_outputs(2100) <= layer1_outputs(175);
    layer2_outputs(2101) <= (layer1_outputs(5444)) and not (layer1_outputs(4795));
    layer2_outputs(2102) <= not(layer1_outputs(2013));
    layer2_outputs(2103) <= not(layer1_outputs(3129));
    layer2_outputs(2104) <= not(layer1_outputs(10128));
    layer2_outputs(2105) <= (layer1_outputs(1347)) and not (layer1_outputs(3160));
    layer2_outputs(2106) <= (layer1_outputs(6672)) xor (layer1_outputs(1716));
    layer2_outputs(2107) <= layer1_outputs(5992);
    layer2_outputs(2108) <= layer1_outputs(643);
    layer2_outputs(2109) <= (layer1_outputs(6658)) and (layer1_outputs(5303));
    layer2_outputs(2110) <= not(layer1_outputs(3581));
    layer2_outputs(2111) <= layer1_outputs(9344);
    layer2_outputs(2112) <= layer1_outputs(9194);
    layer2_outputs(2113) <= not((layer1_outputs(2052)) and (layer1_outputs(6532)));
    layer2_outputs(2114) <= not(layer1_outputs(10105)) or (layer1_outputs(3558));
    layer2_outputs(2115) <= not(layer1_outputs(3831));
    layer2_outputs(2116) <= not(layer1_outputs(7127));
    layer2_outputs(2117) <= layer1_outputs(6046);
    layer2_outputs(2118) <= (layer1_outputs(9670)) and (layer1_outputs(9229));
    layer2_outputs(2119) <= layer1_outputs(6483);
    layer2_outputs(2120) <= not((layer1_outputs(9367)) xor (layer1_outputs(4979)));
    layer2_outputs(2121) <= (layer1_outputs(2958)) and not (layer1_outputs(6584));
    layer2_outputs(2122) <= not(layer1_outputs(5262));
    layer2_outputs(2123) <= not((layer1_outputs(2327)) xor (layer1_outputs(6808)));
    layer2_outputs(2124) <= not((layer1_outputs(1303)) and (layer1_outputs(5960)));
    layer2_outputs(2125) <= layer1_outputs(8512);
    layer2_outputs(2126) <= (layer1_outputs(9690)) and (layer1_outputs(8039));
    layer2_outputs(2127) <= not((layer1_outputs(2766)) and (layer1_outputs(4188)));
    layer2_outputs(2128) <= not((layer1_outputs(1256)) or (layer1_outputs(8782)));
    layer2_outputs(2129) <= not(layer1_outputs(8980));
    layer2_outputs(2130) <= not(layer1_outputs(5033));
    layer2_outputs(2131) <= layer1_outputs(1278);
    layer2_outputs(2132) <= not(layer1_outputs(2646));
    layer2_outputs(2133) <= (layer1_outputs(6595)) and (layer1_outputs(9949));
    layer2_outputs(2134) <= not((layer1_outputs(5089)) xor (layer1_outputs(20)));
    layer2_outputs(2135) <= not(layer1_outputs(4563)) or (layer1_outputs(2671));
    layer2_outputs(2136) <= not(layer1_outputs(239));
    layer2_outputs(2137) <= not(layer1_outputs(10028));
    layer2_outputs(2138) <= layer1_outputs(3391);
    layer2_outputs(2139) <= not(layer1_outputs(5979)) or (layer1_outputs(553));
    layer2_outputs(2140) <= layer1_outputs(7975);
    layer2_outputs(2141) <= not(layer1_outputs(538));
    layer2_outputs(2142) <= not(layer1_outputs(437));
    layer2_outputs(2143) <= not(layer1_outputs(6463)) or (layer1_outputs(7261));
    layer2_outputs(2144) <= not(layer1_outputs(7742)) or (layer1_outputs(9044));
    layer2_outputs(2145) <= not((layer1_outputs(4963)) and (layer1_outputs(8144)));
    layer2_outputs(2146) <= not(layer1_outputs(7411));
    layer2_outputs(2147) <= (layer1_outputs(5143)) xor (layer1_outputs(8397));
    layer2_outputs(2148) <= not((layer1_outputs(3888)) xor (layer1_outputs(6577)));
    layer2_outputs(2149) <= (layer1_outputs(132)) and not (layer1_outputs(6108));
    layer2_outputs(2150) <= not(layer1_outputs(2762));
    layer2_outputs(2151) <= not(layer1_outputs(1643));
    layer2_outputs(2152) <= layer1_outputs(10089);
    layer2_outputs(2153) <= layer1_outputs(7657);
    layer2_outputs(2154) <= not(layer1_outputs(1486));
    layer2_outputs(2155) <= layer1_outputs(307);
    layer2_outputs(2156) <= layer1_outputs(4498);
    layer2_outputs(2157) <= not(layer1_outputs(5309));
    layer2_outputs(2158) <= layer1_outputs(1852);
    layer2_outputs(2159) <= layer1_outputs(3361);
    layer2_outputs(2160) <= layer1_outputs(6553);
    layer2_outputs(2161) <= not(layer1_outputs(9394)) or (layer1_outputs(3382));
    layer2_outputs(2162) <= not(layer1_outputs(8571));
    layer2_outputs(2163) <= not(layer1_outputs(7896));
    layer2_outputs(2164) <= layer1_outputs(8897);
    layer2_outputs(2165) <= (layer1_outputs(6766)) or (layer1_outputs(1538));
    layer2_outputs(2166) <= layer1_outputs(1624);
    layer2_outputs(2167) <= layer1_outputs(1258);
    layer2_outputs(2168) <= (layer1_outputs(5342)) xor (layer1_outputs(4762));
    layer2_outputs(2169) <= layer1_outputs(7014);
    layer2_outputs(2170) <= layer1_outputs(2284);
    layer2_outputs(2171) <= not((layer1_outputs(5663)) and (layer1_outputs(2429)));
    layer2_outputs(2172) <= layer1_outputs(4178);
    layer2_outputs(2173) <= layer1_outputs(4064);
    layer2_outputs(2174) <= (layer1_outputs(94)) or (layer1_outputs(9666));
    layer2_outputs(2175) <= '1';
    layer2_outputs(2176) <= layer1_outputs(9233);
    layer2_outputs(2177) <= not(layer1_outputs(9397));
    layer2_outputs(2178) <= layer1_outputs(1043);
    layer2_outputs(2179) <= (layer1_outputs(4509)) or (layer1_outputs(4639));
    layer2_outputs(2180) <= (layer1_outputs(48)) and not (layer1_outputs(5616));
    layer2_outputs(2181) <= (layer1_outputs(8191)) and not (layer1_outputs(6040));
    layer2_outputs(2182) <= not((layer1_outputs(8623)) xor (layer1_outputs(7064)));
    layer2_outputs(2183) <= layer1_outputs(3260);
    layer2_outputs(2184) <= layer1_outputs(9658);
    layer2_outputs(2185) <= not(layer1_outputs(7284));
    layer2_outputs(2186) <= not((layer1_outputs(7713)) xor (layer1_outputs(3500)));
    layer2_outputs(2187) <= layer1_outputs(1754);
    layer2_outputs(2188) <= layer1_outputs(3461);
    layer2_outputs(2189) <= not(layer1_outputs(2875));
    layer2_outputs(2190) <= not(layer1_outputs(8944));
    layer2_outputs(2191) <= not(layer1_outputs(6228));
    layer2_outputs(2192) <= not((layer1_outputs(252)) and (layer1_outputs(4983)));
    layer2_outputs(2193) <= (layer1_outputs(1833)) and not (layer1_outputs(10203));
    layer2_outputs(2194) <= not(layer1_outputs(1116)) or (layer1_outputs(7135));
    layer2_outputs(2195) <= (layer1_outputs(5720)) or (layer1_outputs(9674));
    layer2_outputs(2196) <= layer1_outputs(921);
    layer2_outputs(2197) <= not((layer1_outputs(7269)) or (layer1_outputs(5074)));
    layer2_outputs(2198) <= layer1_outputs(98);
    layer2_outputs(2199) <= not(layer1_outputs(5893));
    layer2_outputs(2200) <= not(layer1_outputs(2317)) or (layer1_outputs(6885));
    layer2_outputs(2201) <= not((layer1_outputs(43)) and (layer1_outputs(6887)));
    layer2_outputs(2202) <= not(layer1_outputs(10010));
    layer2_outputs(2203) <= not(layer1_outputs(1225)) or (layer1_outputs(10004));
    layer2_outputs(2204) <= layer1_outputs(1447);
    layer2_outputs(2205) <= not(layer1_outputs(2409));
    layer2_outputs(2206) <= layer1_outputs(2348);
    layer2_outputs(2207) <= not(layer1_outputs(1980));
    layer2_outputs(2208) <= (layer1_outputs(3735)) xor (layer1_outputs(7698));
    layer2_outputs(2209) <= not(layer1_outputs(2038)) or (layer1_outputs(9756));
    layer2_outputs(2210) <= not((layer1_outputs(4591)) and (layer1_outputs(2810)));
    layer2_outputs(2211) <= not((layer1_outputs(4196)) and (layer1_outputs(1542)));
    layer2_outputs(2212) <= layer1_outputs(8728);
    layer2_outputs(2213) <= not(layer1_outputs(2205)) or (layer1_outputs(728));
    layer2_outputs(2214) <= not((layer1_outputs(5726)) xor (layer1_outputs(9613)));
    layer2_outputs(2215) <= (layer1_outputs(9881)) and (layer1_outputs(6433));
    layer2_outputs(2216) <= (layer1_outputs(3647)) xor (layer1_outputs(9314));
    layer2_outputs(2217) <= (layer1_outputs(7211)) and not (layer1_outputs(6829));
    layer2_outputs(2218) <= not(layer1_outputs(5590));
    layer2_outputs(2219) <= not(layer1_outputs(1318));
    layer2_outputs(2220) <= not((layer1_outputs(9183)) and (layer1_outputs(4631)));
    layer2_outputs(2221) <= layer1_outputs(23);
    layer2_outputs(2222) <= not((layer1_outputs(910)) or (layer1_outputs(9628)));
    layer2_outputs(2223) <= layer1_outputs(7871);
    layer2_outputs(2224) <= layer1_outputs(704);
    layer2_outputs(2225) <= not(layer1_outputs(6771));
    layer2_outputs(2226) <= layer1_outputs(7318);
    layer2_outputs(2227) <= layer1_outputs(9965);
    layer2_outputs(2228) <= layer1_outputs(1477);
    layer2_outputs(2229) <= not(layer1_outputs(2865));
    layer2_outputs(2230) <= layer1_outputs(8277);
    layer2_outputs(2231) <= layer1_outputs(1259);
    layer2_outputs(2232) <= not((layer1_outputs(5121)) or (layer1_outputs(5933)));
    layer2_outputs(2233) <= layer1_outputs(2853);
    layer2_outputs(2234) <= not((layer1_outputs(817)) xor (layer1_outputs(4666)));
    layer2_outputs(2235) <= layer1_outputs(9162);
    layer2_outputs(2236) <= not(layer1_outputs(544));
    layer2_outputs(2237) <= layer1_outputs(7271);
    layer2_outputs(2238) <= not(layer1_outputs(9522)) or (layer1_outputs(2136));
    layer2_outputs(2239) <= layer1_outputs(10159);
    layer2_outputs(2240) <= layer1_outputs(4520);
    layer2_outputs(2241) <= not(layer1_outputs(2937));
    layer2_outputs(2242) <= not(layer1_outputs(3499));
    layer2_outputs(2243) <= not(layer1_outputs(6462));
    layer2_outputs(2244) <= (layer1_outputs(4772)) xor (layer1_outputs(9289));
    layer2_outputs(2245) <= not((layer1_outputs(471)) and (layer1_outputs(4095)));
    layer2_outputs(2246) <= not(layer1_outputs(964)) or (layer1_outputs(846));
    layer2_outputs(2247) <= layer1_outputs(3881);
    layer2_outputs(2248) <= '0';
    layer2_outputs(2249) <= not(layer1_outputs(8702));
    layer2_outputs(2250) <= layer1_outputs(10040);
    layer2_outputs(2251) <= not(layer1_outputs(2452)) or (layer1_outputs(959));
    layer2_outputs(2252) <= not(layer1_outputs(9851));
    layer2_outputs(2253) <= not(layer1_outputs(1860));
    layer2_outputs(2254) <= not(layer1_outputs(8514));
    layer2_outputs(2255) <= not(layer1_outputs(3649));
    layer2_outputs(2256) <= (layer1_outputs(10192)) or (layer1_outputs(8374));
    layer2_outputs(2257) <= (layer1_outputs(6158)) xor (layer1_outputs(9521));
    layer2_outputs(2258) <= (layer1_outputs(4889)) and (layer1_outputs(8671));
    layer2_outputs(2259) <= not(layer1_outputs(5454)) or (layer1_outputs(4919));
    layer2_outputs(2260) <= not((layer1_outputs(665)) or (layer1_outputs(3238)));
    layer2_outputs(2261) <= not(layer1_outputs(6758));
    layer2_outputs(2262) <= not(layer1_outputs(7632));
    layer2_outputs(2263) <= layer1_outputs(7950);
    layer2_outputs(2264) <= layer1_outputs(7866);
    layer2_outputs(2265) <= not((layer1_outputs(5165)) and (layer1_outputs(5907)));
    layer2_outputs(2266) <= not(layer1_outputs(3445));
    layer2_outputs(2267) <= (layer1_outputs(4229)) and not (layer1_outputs(6525));
    layer2_outputs(2268) <= (layer1_outputs(4060)) and (layer1_outputs(5929));
    layer2_outputs(2269) <= not(layer1_outputs(9397));
    layer2_outputs(2270) <= not(layer1_outputs(6613));
    layer2_outputs(2271) <= (layer1_outputs(3748)) xor (layer1_outputs(5165));
    layer2_outputs(2272) <= layer1_outputs(10176);
    layer2_outputs(2273) <= not(layer1_outputs(691));
    layer2_outputs(2274) <= not(layer1_outputs(6181));
    layer2_outputs(2275) <= not(layer1_outputs(3100));
    layer2_outputs(2276) <= layer1_outputs(7435);
    layer2_outputs(2277) <= layer1_outputs(1217);
    layer2_outputs(2278) <= layer1_outputs(5211);
    layer2_outputs(2279) <= not(layer1_outputs(5411)) or (layer1_outputs(6293));
    layer2_outputs(2280) <= not(layer1_outputs(9517));
    layer2_outputs(2281) <= layer1_outputs(682);
    layer2_outputs(2282) <= not((layer1_outputs(3948)) xor (layer1_outputs(6598)));
    layer2_outputs(2283) <= layer1_outputs(4408);
    layer2_outputs(2284) <= not(layer1_outputs(10096));
    layer2_outputs(2285) <= not(layer1_outputs(9677));
    layer2_outputs(2286) <= (layer1_outputs(10)) and (layer1_outputs(9486));
    layer2_outputs(2287) <= not((layer1_outputs(7430)) xor (layer1_outputs(2893)));
    layer2_outputs(2288) <= not(layer1_outputs(8864));
    layer2_outputs(2289) <= layer1_outputs(8900);
    layer2_outputs(2290) <= layer1_outputs(8273);
    layer2_outputs(2291) <= layer1_outputs(2930);
    layer2_outputs(2292) <= layer1_outputs(9127);
    layer2_outputs(2293) <= layer1_outputs(5786);
    layer2_outputs(2294) <= layer1_outputs(3655);
    layer2_outputs(2295) <= not(layer1_outputs(796));
    layer2_outputs(2296) <= '0';
    layer2_outputs(2297) <= '1';
    layer2_outputs(2298) <= not(layer1_outputs(7957));
    layer2_outputs(2299) <= not(layer1_outputs(3297));
    layer2_outputs(2300) <= layer1_outputs(2293);
    layer2_outputs(2301) <= (layer1_outputs(2871)) xor (layer1_outputs(6809));
    layer2_outputs(2302) <= layer1_outputs(1850);
    layer2_outputs(2303) <= (layer1_outputs(4985)) and not (layer1_outputs(9633));
    layer2_outputs(2304) <= layer1_outputs(1514);
    layer2_outputs(2305) <= not(layer1_outputs(2981));
    layer2_outputs(2306) <= '1';
    layer2_outputs(2307) <= layer1_outputs(6636);
    layer2_outputs(2308) <= (layer1_outputs(305)) and not (layer1_outputs(2548));
    layer2_outputs(2309) <= (layer1_outputs(10125)) and not (layer1_outputs(8661));
    layer2_outputs(2310) <= layer1_outputs(1537);
    layer2_outputs(2311) <= layer1_outputs(9703);
    layer2_outputs(2312) <= (layer1_outputs(6712)) xor (layer1_outputs(5738));
    layer2_outputs(2313) <= (layer1_outputs(3144)) and not (layer1_outputs(7932));
    layer2_outputs(2314) <= layer1_outputs(3567);
    layer2_outputs(2315) <= '0';
    layer2_outputs(2316) <= layer1_outputs(9883);
    layer2_outputs(2317) <= not((layer1_outputs(2277)) xor (layer1_outputs(4226)));
    layer2_outputs(2318) <= not((layer1_outputs(8294)) xor (layer1_outputs(831)));
    layer2_outputs(2319) <= not(layer1_outputs(2329));
    layer2_outputs(2320) <= not((layer1_outputs(6882)) and (layer1_outputs(8683)));
    layer2_outputs(2321) <= not(layer1_outputs(4609));
    layer2_outputs(2322) <= not(layer1_outputs(3433)) or (layer1_outputs(4935));
    layer2_outputs(2323) <= not((layer1_outputs(9380)) or (layer1_outputs(3293)));
    layer2_outputs(2324) <= layer1_outputs(7091);
    layer2_outputs(2325) <= layer1_outputs(8132);
    layer2_outputs(2326) <= layer1_outputs(1089);
    layer2_outputs(2327) <= (layer1_outputs(1859)) and not (layer1_outputs(563));
    layer2_outputs(2328) <= layer1_outputs(2357);
    layer2_outputs(2329) <= layer1_outputs(7547);
    layer2_outputs(2330) <= not(layer1_outputs(7638));
    layer2_outputs(2331) <= layer1_outputs(6294);
    layer2_outputs(2332) <= layer1_outputs(2279);
    layer2_outputs(2333) <= not(layer1_outputs(3496));
    layer2_outputs(2334) <= not(layer1_outputs(3942)) or (layer1_outputs(3975));
    layer2_outputs(2335) <= (layer1_outputs(9331)) and (layer1_outputs(7949));
    layer2_outputs(2336) <= not(layer1_outputs(6241));
    layer2_outputs(2337) <= not(layer1_outputs(9967));
    layer2_outputs(2338) <= not(layer1_outputs(9834));
    layer2_outputs(2339) <= not((layer1_outputs(5514)) xor (layer1_outputs(5114)));
    layer2_outputs(2340) <= (layer1_outputs(3574)) and (layer1_outputs(4661));
    layer2_outputs(2341) <= '0';
    layer2_outputs(2342) <= (layer1_outputs(9737)) or (layer1_outputs(6385));
    layer2_outputs(2343) <= not(layer1_outputs(1631));
    layer2_outputs(2344) <= layer1_outputs(3961);
    layer2_outputs(2345) <= (layer1_outputs(7535)) and not (layer1_outputs(7870));
    layer2_outputs(2346) <= (layer1_outputs(5554)) xor (layer1_outputs(961));
    layer2_outputs(2347) <= (layer1_outputs(5595)) or (layer1_outputs(3267));
    layer2_outputs(2348) <= layer1_outputs(6447);
    layer2_outputs(2349) <= not(layer1_outputs(10078)) or (layer1_outputs(2800));
    layer2_outputs(2350) <= not(layer1_outputs(2286)) or (layer1_outputs(10047));
    layer2_outputs(2351) <= not(layer1_outputs(7114));
    layer2_outputs(2352) <= (layer1_outputs(7542)) xor (layer1_outputs(1501));
    layer2_outputs(2353) <= not((layer1_outputs(10111)) or (layer1_outputs(2130)));
    layer2_outputs(2354) <= layer1_outputs(4072);
    layer2_outputs(2355) <= '1';
    layer2_outputs(2356) <= not(layer1_outputs(5782));
    layer2_outputs(2357) <= not(layer1_outputs(5618));
    layer2_outputs(2358) <= not((layer1_outputs(996)) or (layer1_outputs(8724)));
    layer2_outputs(2359) <= not(layer1_outputs(1247));
    layer2_outputs(2360) <= not(layer1_outputs(6719)) or (layer1_outputs(1206));
    layer2_outputs(2361) <= not(layer1_outputs(5050));
    layer2_outputs(2362) <= layer1_outputs(3568);
    layer2_outputs(2363) <= (layer1_outputs(9995)) and not (layer1_outputs(3551));
    layer2_outputs(2364) <= not(layer1_outputs(5962));
    layer2_outputs(2365) <= '1';
    layer2_outputs(2366) <= layer1_outputs(1695);
    layer2_outputs(2367) <= layer1_outputs(5439);
    layer2_outputs(2368) <= not(layer1_outputs(1277)) or (layer1_outputs(2950));
    layer2_outputs(2369) <= layer1_outputs(5097);
    layer2_outputs(2370) <= layer1_outputs(5003);
    layer2_outputs(2371) <= not(layer1_outputs(5177));
    layer2_outputs(2372) <= layer1_outputs(6998);
    layer2_outputs(2373) <= not(layer1_outputs(2818));
    layer2_outputs(2374) <= not(layer1_outputs(1355)) or (layer1_outputs(6890));
    layer2_outputs(2375) <= not(layer1_outputs(6231));
    layer2_outputs(2376) <= not((layer1_outputs(3855)) xor (layer1_outputs(4806)));
    layer2_outputs(2377) <= not(layer1_outputs(1429));
    layer2_outputs(2378) <= (layer1_outputs(8540)) xor (layer1_outputs(5827));
    layer2_outputs(2379) <= layer1_outputs(4643);
    layer2_outputs(2380) <= not((layer1_outputs(6092)) and (layer1_outputs(6698)));
    layer2_outputs(2381) <= (layer1_outputs(8283)) or (layer1_outputs(6425));
    layer2_outputs(2382) <= (layer1_outputs(7387)) and not (layer1_outputs(4189));
    layer2_outputs(2383) <= layer1_outputs(8668);
    layer2_outputs(2384) <= not((layer1_outputs(3637)) xor (layer1_outputs(9093)));
    layer2_outputs(2385) <= not((layer1_outputs(6930)) xor (layer1_outputs(7975)));
    layer2_outputs(2386) <= not((layer1_outputs(2544)) or (layer1_outputs(6689)));
    layer2_outputs(2387) <= not(layer1_outputs(4530));
    layer2_outputs(2388) <= layer1_outputs(8866);
    layer2_outputs(2389) <= (layer1_outputs(1459)) and (layer1_outputs(8916));
    layer2_outputs(2390) <= layer1_outputs(2306);
    layer2_outputs(2391) <= not((layer1_outputs(2265)) or (layer1_outputs(8328)));
    layer2_outputs(2392) <= not((layer1_outputs(598)) and (layer1_outputs(840)));
    layer2_outputs(2393) <= not(layer1_outputs(7114)) or (layer1_outputs(3371));
    layer2_outputs(2394) <= (layer1_outputs(2546)) xor (layer1_outputs(2414));
    layer2_outputs(2395) <= not(layer1_outputs(1853));
    layer2_outputs(2396) <= '1';
    layer2_outputs(2397) <= not((layer1_outputs(4368)) xor (layer1_outputs(9750)));
    layer2_outputs(2398) <= layer1_outputs(4891);
    layer2_outputs(2399) <= not(layer1_outputs(7860));
    layer2_outputs(2400) <= not(layer1_outputs(270));
    layer2_outputs(2401) <= not(layer1_outputs(1301));
    layer2_outputs(2402) <= not(layer1_outputs(5365));
    layer2_outputs(2403) <= layer1_outputs(6396);
    layer2_outputs(2404) <= layer1_outputs(2765);
    layer2_outputs(2405) <= layer1_outputs(5486);
    layer2_outputs(2406) <= not(layer1_outputs(8403));
    layer2_outputs(2407) <= not((layer1_outputs(8025)) or (layer1_outputs(6425)));
    layer2_outputs(2408) <= not(layer1_outputs(809)) or (layer1_outputs(2935));
    layer2_outputs(2409) <= (layer1_outputs(6963)) xor (layer1_outputs(8589));
    layer2_outputs(2410) <= layer1_outputs(905);
    layer2_outputs(2411) <= (layer1_outputs(4938)) xor (layer1_outputs(2251));
    layer2_outputs(2412) <= layer1_outputs(7593);
    layer2_outputs(2413) <= not(layer1_outputs(3893)) or (layer1_outputs(8971));
    layer2_outputs(2414) <= (layer1_outputs(4831)) xor (layer1_outputs(7260));
    layer2_outputs(2415) <= (layer1_outputs(1471)) xor (layer1_outputs(3700));
    layer2_outputs(2416) <= not(layer1_outputs(7280));
    layer2_outputs(2417) <= not(layer1_outputs(8259));
    layer2_outputs(2418) <= not(layer1_outputs(1463)) or (layer1_outputs(475));
    layer2_outputs(2419) <= not(layer1_outputs(7979));
    layer2_outputs(2420) <= layer1_outputs(324);
    layer2_outputs(2421) <= not((layer1_outputs(920)) and (layer1_outputs(9410)));
    layer2_outputs(2422) <= not(layer1_outputs(641)) or (layer1_outputs(2847));
    layer2_outputs(2423) <= not(layer1_outputs(10232));
    layer2_outputs(2424) <= layer1_outputs(5899);
    layer2_outputs(2425) <= layer1_outputs(445);
    layer2_outputs(2426) <= layer1_outputs(2970);
    layer2_outputs(2427) <= (layer1_outputs(9574)) xor (layer1_outputs(7231));
    layer2_outputs(2428) <= not(layer1_outputs(8059));
    layer2_outputs(2429) <= not(layer1_outputs(4377)) or (layer1_outputs(5087));
    layer2_outputs(2430) <= layer1_outputs(10141);
    layer2_outputs(2431) <= not(layer1_outputs(5581)) or (layer1_outputs(6423));
    layer2_outputs(2432) <= not(layer1_outputs(8803));
    layer2_outputs(2433) <= (layer1_outputs(6363)) or (layer1_outputs(1773));
    layer2_outputs(2434) <= not(layer1_outputs(5674));
    layer2_outputs(2435) <= layer1_outputs(2658);
    layer2_outputs(2436) <= not(layer1_outputs(4545)) or (layer1_outputs(3061));
    layer2_outputs(2437) <= layer1_outputs(6004);
    layer2_outputs(2438) <= not(layer1_outputs(290));
    layer2_outputs(2439) <= layer1_outputs(6723);
    layer2_outputs(2440) <= layer1_outputs(8388);
    layer2_outputs(2441) <= not(layer1_outputs(489));
    layer2_outputs(2442) <= (layer1_outputs(6059)) or (layer1_outputs(2852));
    layer2_outputs(2443) <= layer1_outputs(3585);
    layer2_outputs(2444) <= layer1_outputs(3668);
    layer2_outputs(2445) <= not((layer1_outputs(7600)) xor (layer1_outputs(8063)));
    layer2_outputs(2446) <= (layer1_outputs(9173)) and not (layer1_outputs(814));
    layer2_outputs(2447) <= not((layer1_outputs(5869)) and (layer1_outputs(3275)));
    layer2_outputs(2448) <= not(layer1_outputs(367));
    layer2_outputs(2449) <= layer1_outputs(217);
    layer2_outputs(2450) <= layer1_outputs(2752);
    layer2_outputs(2451) <= not(layer1_outputs(7085));
    layer2_outputs(2452) <= layer1_outputs(5847);
    layer2_outputs(2453) <= not((layer1_outputs(6535)) xor (layer1_outputs(364)));
    layer2_outputs(2454) <= layer1_outputs(6678);
    layer2_outputs(2455) <= not(layer1_outputs(7883)) or (layer1_outputs(2664));
    layer2_outputs(2456) <= layer1_outputs(1525);
    layer2_outputs(2457) <= not(layer1_outputs(5171));
    layer2_outputs(2458) <= layer1_outputs(1345);
    layer2_outputs(2459) <= not(layer1_outputs(8645));
    layer2_outputs(2460) <= not(layer1_outputs(7895));
    layer2_outputs(2461) <= not(layer1_outputs(1276));
    layer2_outputs(2462) <= (layer1_outputs(4942)) xor (layer1_outputs(3404));
    layer2_outputs(2463) <= layer1_outputs(3132);
    layer2_outputs(2464) <= not((layer1_outputs(1045)) xor (layer1_outputs(5233)));
    layer2_outputs(2465) <= (layer1_outputs(9901)) and not (layer1_outputs(10160));
    layer2_outputs(2466) <= layer1_outputs(671);
    layer2_outputs(2467) <= not(layer1_outputs(9161));
    layer2_outputs(2468) <= not(layer1_outputs(5074)) or (layer1_outputs(8445));
    layer2_outputs(2469) <= layer1_outputs(1309);
    layer2_outputs(2470) <= layer1_outputs(6746);
    layer2_outputs(2471) <= not(layer1_outputs(1158));
    layer2_outputs(2472) <= (layer1_outputs(7506)) xor (layer1_outputs(3619));
    layer2_outputs(2473) <= not((layer1_outputs(5819)) and (layer1_outputs(6482)));
    layer2_outputs(2474) <= '0';
    layer2_outputs(2475) <= not((layer1_outputs(8467)) xor (layer1_outputs(9555)));
    layer2_outputs(2476) <= not(layer1_outputs(630));
    layer2_outputs(2477) <= not(layer1_outputs(3480));
    layer2_outputs(2478) <= not(layer1_outputs(5144)) or (layer1_outputs(5297));
    layer2_outputs(2479) <= layer1_outputs(2066);
    layer2_outputs(2480) <= layer1_outputs(7762);
    layer2_outputs(2481) <= (layer1_outputs(4811)) and (layer1_outputs(2859));
    layer2_outputs(2482) <= layer1_outputs(2262);
    layer2_outputs(2483) <= layer1_outputs(2797);
    layer2_outputs(2484) <= (layer1_outputs(8012)) and (layer1_outputs(6527));
    layer2_outputs(2485) <= layer1_outputs(7891);
    layer2_outputs(2486) <= (layer1_outputs(42)) and not (layer1_outputs(10127));
    layer2_outputs(2487) <= layer1_outputs(2572);
    layer2_outputs(2488) <= layer1_outputs(6475);
    layer2_outputs(2489) <= not(layer1_outputs(8543));
    layer2_outputs(2490) <= not(layer1_outputs(3802));
    layer2_outputs(2491) <= layer1_outputs(4427);
    layer2_outputs(2492) <= layer1_outputs(153);
    layer2_outputs(2493) <= not(layer1_outputs(9509));
    layer2_outputs(2494) <= (layer1_outputs(8972)) and not (layer1_outputs(6921));
    layer2_outputs(2495) <= not(layer1_outputs(342));
    layer2_outputs(2496) <= not((layer1_outputs(7813)) and (layer1_outputs(8978)));
    layer2_outputs(2497) <= not(layer1_outputs(4591));
    layer2_outputs(2498) <= not((layer1_outputs(6941)) and (layer1_outputs(3744)));
    layer2_outputs(2499) <= (layer1_outputs(1021)) and (layer1_outputs(7046));
    layer2_outputs(2500) <= not(layer1_outputs(6807));
    layer2_outputs(2501) <= (layer1_outputs(9848)) and not (layer1_outputs(223));
    layer2_outputs(2502) <= layer1_outputs(7588);
    layer2_outputs(2503) <= not(layer1_outputs(8212)) or (layer1_outputs(9108));
    layer2_outputs(2504) <= not(layer1_outputs(1598));
    layer2_outputs(2505) <= not(layer1_outputs(9053));
    layer2_outputs(2506) <= not((layer1_outputs(1427)) and (layer1_outputs(4495)));
    layer2_outputs(2507) <= not(layer1_outputs(7502));
    layer2_outputs(2508) <= not((layer1_outputs(7559)) or (layer1_outputs(4248)));
    layer2_outputs(2509) <= (layer1_outputs(7501)) xor (layer1_outputs(5940));
    layer2_outputs(2510) <= not(layer1_outputs(330)) or (layer1_outputs(7008));
    layer2_outputs(2511) <= (layer1_outputs(9035)) and not (layer1_outputs(6977));
    layer2_outputs(2512) <= layer1_outputs(8652);
    layer2_outputs(2513) <= layer1_outputs(9776);
    layer2_outputs(2514) <= not(layer1_outputs(3025)) or (layer1_outputs(10235));
    layer2_outputs(2515) <= not(layer1_outputs(4799));
    layer2_outputs(2516) <= layer1_outputs(7303);
    layer2_outputs(2517) <= layer1_outputs(9947);
    layer2_outputs(2518) <= not(layer1_outputs(8515));
    layer2_outputs(2519) <= not(layer1_outputs(2654));
    layer2_outputs(2520) <= not((layer1_outputs(884)) and (layer1_outputs(12)));
    layer2_outputs(2521) <= not(layer1_outputs(322));
    layer2_outputs(2522) <= layer1_outputs(9629);
    layer2_outputs(2523) <= layer1_outputs(6797);
    layer2_outputs(2524) <= (layer1_outputs(7206)) and not (layer1_outputs(5013));
    layer2_outputs(2525) <= layer1_outputs(3788);
    layer2_outputs(2526) <= (layer1_outputs(7193)) and not (layer1_outputs(9469));
    layer2_outputs(2527) <= not(layer1_outputs(5579));
    layer2_outputs(2528) <= layer1_outputs(7750);
    layer2_outputs(2529) <= (layer1_outputs(9464)) and not (layer1_outputs(8928));
    layer2_outputs(2530) <= (layer1_outputs(6472)) and (layer1_outputs(5716));
    layer2_outputs(2531) <= (layer1_outputs(6678)) and not (layer1_outputs(1845));
    layer2_outputs(2532) <= (layer1_outputs(2215)) xor (layer1_outputs(10007));
    layer2_outputs(2533) <= not(layer1_outputs(7705)) or (layer1_outputs(582));
    layer2_outputs(2534) <= layer1_outputs(10048);
    layer2_outputs(2535) <= not(layer1_outputs(7496)) or (layer1_outputs(2768));
    layer2_outputs(2536) <= not(layer1_outputs(698));
    layer2_outputs(2537) <= not(layer1_outputs(8379)) or (layer1_outputs(3432));
    layer2_outputs(2538) <= not(layer1_outputs(5991));
    layer2_outputs(2539) <= not((layer1_outputs(5081)) and (layer1_outputs(2432)));
    layer2_outputs(2540) <= not(layer1_outputs(4059));
    layer2_outputs(2541) <= (layer1_outputs(4693)) and (layer1_outputs(9407));
    layer2_outputs(2542) <= (layer1_outputs(2096)) and not (layer1_outputs(8462));
    layer2_outputs(2543) <= layer1_outputs(2159);
    layer2_outputs(2544) <= '1';
    layer2_outputs(2545) <= (layer1_outputs(7889)) or (layer1_outputs(5093));
    layer2_outputs(2546) <= (layer1_outputs(4733)) or (layer1_outputs(4429));
    layer2_outputs(2547) <= (layer1_outputs(3038)) and not (layer1_outputs(4801));
    layer2_outputs(2548) <= (layer1_outputs(537)) xor (layer1_outputs(5643));
    layer2_outputs(2549) <= not(layer1_outputs(8435));
    layer2_outputs(2550) <= layer1_outputs(6439);
    layer2_outputs(2551) <= layer1_outputs(614);
    layer2_outputs(2552) <= layer1_outputs(1544);
    layer2_outputs(2553) <= not((layer1_outputs(7663)) or (layer1_outputs(9837)));
    layer2_outputs(2554) <= not(layer1_outputs(1371));
    layer2_outputs(2555) <= layer1_outputs(6253);
    layer2_outputs(2556) <= not(layer1_outputs(2520));
    layer2_outputs(2557) <= layer1_outputs(3117);
    layer2_outputs(2558) <= (layer1_outputs(10185)) or (layer1_outputs(1784));
    layer2_outputs(2559) <= layer1_outputs(4987);
    layer2_outputs(2560) <= layer1_outputs(8255);
    layer2_outputs(2561) <= (layer1_outputs(5855)) or (layer1_outputs(6554));
    layer2_outputs(2562) <= layer1_outputs(6049);
    layer2_outputs(2563) <= (layer1_outputs(2431)) or (layer1_outputs(6993));
    layer2_outputs(2564) <= layer1_outputs(7415);
    layer2_outputs(2565) <= not((layer1_outputs(7308)) or (layer1_outputs(8316)));
    layer2_outputs(2566) <= not((layer1_outputs(1578)) xor (layer1_outputs(2589)));
    layer2_outputs(2567) <= not(layer1_outputs(5789));
    layer2_outputs(2568) <= not((layer1_outputs(9588)) or (layer1_outputs(6873)));
    layer2_outputs(2569) <= (layer1_outputs(10015)) and (layer1_outputs(8278));
    layer2_outputs(2570) <= layer1_outputs(5138);
    layer2_outputs(2571) <= layer1_outputs(3962);
    layer2_outputs(2572) <= (layer1_outputs(5395)) and not (layer1_outputs(9775));
    layer2_outputs(2573) <= not(layer1_outputs(1115)) or (layer1_outputs(3042));
    layer2_outputs(2574) <= not(layer1_outputs(8367));
    layer2_outputs(2575) <= layer1_outputs(4590);
    layer2_outputs(2576) <= not(layer1_outputs(6339));
    layer2_outputs(2577) <= layer1_outputs(1461);
    layer2_outputs(2578) <= layer1_outputs(2788);
    layer2_outputs(2579) <= '0';
    layer2_outputs(2580) <= layer1_outputs(6343);
    layer2_outputs(2581) <= not((layer1_outputs(1769)) and (layer1_outputs(7546)));
    layer2_outputs(2582) <= (layer1_outputs(4246)) and not (layer1_outputs(3052));
    layer2_outputs(2583) <= not(layer1_outputs(5384));
    layer2_outputs(2584) <= '0';
    layer2_outputs(2585) <= layer1_outputs(4372);
    layer2_outputs(2586) <= (layer1_outputs(5543)) and not (layer1_outputs(4372));
    layer2_outputs(2587) <= not(layer1_outputs(3075)) or (layer1_outputs(3682));
    layer2_outputs(2588) <= not(layer1_outputs(6151)) or (layer1_outputs(7109));
    layer2_outputs(2589) <= (layer1_outputs(6414)) and not (layer1_outputs(7433));
    layer2_outputs(2590) <= not(layer1_outputs(779));
    layer2_outputs(2591) <= layer1_outputs(4274);
    layer2_outputs(2592) <= layer1_outputs(9137);
    layer2_outputs(2593) <= not(layer1_outputs(1482));
    layer2_outputs(2594) <= not(layer1_outputs(3462));
    layer2_outputs(2595) <= not((layer1_outputs(2351)) or (layer1_outputs(3856)));
    layer2_outputs(2596) <= not(layer1_outputs(3884));
    layer2_outputs(2597) <= layer1_outputs(5765);
    layer2_outputs(2598) <= not(layer1_outputs(3048));
    layer2_outputs(2599) <= (layer1_outputs(7653)) and (layer1_outputs(162));
    layer2_outputs(2600) <= (layer1_outputs(99)) and not (layer1_outputs(7251));
    layer2_outputs(2601) <= layer1_outputs(8448);
    layer2_outputs(2602) <= not((layer1_outputs(5842)) or (layer1_outputs(2562)));
    layer2_outputs(2603) <= not(layer1_outputs(2357));
    layer2_outputs(2604) <= (layer1_outputs(7817)) and (layer1_outputs(10209));
    layer2_outputs(2605) <= not(layer1_outputs(9462));
    layer2_outputs(2606) <= layer1_outputs(2757);
    layer2_outputs(2607) <= (layer1_outputs(1780)) and not (layer1_outputs(7690));
    layer2_outputs(2608) <= not(layer1_outputs(5495));
    layer2_outputs(2609) <= not((layer1_outputs(4360)) and (layer1_outputs(212)));
    layer2_outputs(2610) <= not(layer1_outputs(2373));
    layer2_outputs(2611) <= layer1_outputs(1359);
    layer2_outputs(2612) <= not(layer1_outputs(1952));
    layer2_outputs(2613) <= layer1_outputs(3128);
    layer2_outputs(2614) <= (layer1_outputs(5770)) or (layer1_outputs(609));
    layer2_outputs(2615) <= (layer1_outputs(3622)) and (layer1_outputs(9113));
    layer2_outputs(2616) <= layer1_outputs(6511);
    layer2_outputs(2617) <= not(layer1_outputs(4398));
    layer2_outputs(2618) <= (layer1_outputs(7990)) and not (layer1_outputs(1895));
    layer2_outputs(2619) <= layer1_outputs(245);
    layer2_outputs(2620) <= layer1_outputs(6320);
    layer2_outputs(2621) <= (layer1_outputs(481)) or (layer1_outputs(5245));
    layer2_outputs(2622) <= not(layer1_outputs(9680));
    layer2_outputs(2623) <= layer1_outputs(6608);
    layer2_outputs(2624) <= layer1_outputs(6426);
    layer2_outputs(2625) <= not((layer1_outputs(7408)) xor (layer1_outputs(1978)));
    layer2_outputs(2626) <= layer1_outputs(2112);
    layer2_outputs(2627) <= (layer1_outputs(1900)) and (layer1_outputs(8393));
    layer2_outputs(2628) <= layer1_outputs(4529);
    layer2_outputs(2629) <= (layer1_outputs(3223)) and not (layer1_outputs(71));
    layer2_outputs(2630) <= not((layer1_outputs(822)) or (layer1_outputs(2784)));
    layer2_outputs(2631) <= layer1_outputs(121);
    layer2_outputs(2632) <= not(layer1_outputs(8099));
    layer2_outputs(2633) <= not(layer1_outputs(9022));
    layer2_outputs(2634) <= (layer1_outputs(2399)) or (layer1_outputs(7453));
    layer2_outputs(2635) <= not(layer1_outputs(7129));
    layer2_outputs(2636) <= not(layer1_outputs(8314));
    layer2_outputs(2637) <= layer1_outputs(8436);
    layer2_outputs(2638) <= layer1_outputs(8220);
    layer2_outputs(2639) <= layer1_outputs(4592);
    layer2_outputs(2640) <= not(layer1_outputs(2300));
    layer2_outputs(2641) <= not(layer1_outputs(4993));
    layer2_outputs(2642) <= not(layer1_outputs(4151));
    layer2_outputs(2643) <= not((layer1_outputs(2340)) and (layer1_outputs(1369)));
    layer2_outputs(2644) <= not((layer1_outputs(3542)) xor (layer1_outputs(6754)));
    layer2_outputs(2645) <= not(layer1_outputs(8394));
    layer2_outputs(2646) <= not(layer1_outputs(5805));
    layer2_outputs(2647) <= not((layer1_outputs(3419)) or (layer1_outputs(5146)));
    layer2_outputs(2648) <= not(layer1_outputs(1089));
    layer2_outputs(2649) <= not(layer1_outputs(4415));
    layer2_outputs(2650) <= (layer1_outputs(6583)) and not (layer1_outputs(8398));
    layer2_outputs(2651) <= not((layer1_outputs(8048)) or (layer1_outputs(3540)));
    layer2_outputs(2652) <= not(layer1_outputs(9918));
    layer2_outputs(2653) <= not(layer1_outputs(5424));
    layer2_outputs(2654) <= not(layer1_outputs(9904));
    layer2_outputs(2655) <= (layer1_outputs(1321)) or (layer1_outputs(5091));
    layer2_outputs(2656) <= layer1_outputs(1272);
    layer2_outputs(2657) <= not(layer1_outputs(2727)) or (layer1_outputs(8108));
    layer2_outputs(2658) <= layer1_outputs(7542);
    layer2_outputs(2659) <= not(layer1_outputs(5855));
    layer2_outputs(2660) <= (layer1_outputs(6733)) xor (layer1_outputs(4222));
    layer2_outputs(2661) <= layer1_outputs(9239);
    layer2_outputs(2662) <= not(layer1_outputs(5293));
    layer2_outputs(2663) <= layer1_outputs(6508);
    layer2_outputs(2664) <= (layer1_outputs(3640)) and (layer1_outputs(3073));
    layer2_outputs(2665) <= not(layer1_outputs(6064));
    layer2_outputs(2666) <= not(layer1_outputs(824));
    layer2_outputs(2667) <= not(layer1_outputs(9176));
    layer2_outputs(2668) <= not(layer1_outputs(1183)) or (layer1_outputs(6033));
    layer2_outputs(2669) <= not((layer1_outputs(4620)) or (layer1_outputs(1032)));
    layer2_outputs(2670) <= layer1_outputs(5741);
    layer2_outputs(2671) <= layer1_outputs(7687);
    layer2_outputs(2672) <= not(layer1_outputs(5167)) or (layer1_outputs(3601));
    layer2_outputs(2673) <= (layer1_outputs(1249)) and not (layer1_outputs(7489));
    layer2_outputs(2674) <= (layer1_outputs(8482)) or (layer1_outputs(5052));
    layer2_outputs(2675) <= not(layer1_outputs(8934));
    layer2_outputs(2676) <= not(layer1_outputs(5835));
    layer2_outputs(2677) <= layer1_outputs(4141);
    layer2_outputs(2678) <= not(layer1_outputs(5996));
    layer2_outputs(2679) <= layer1_outputs(8681);
    layer2_outputs(2680) <= (layer1_outputs(9263)) xor (layer1_outputs(5807));
    layer2_outputs(2681) <= layer1_outputs(3177);
    layer2_outputs(2682) <= not(layer1_outputs(1141)) or (layer1_outputs(10147));
    layer2_outputs(2683) <= (layer1_outputs(1491)) and not (layer1_outputs(3650));
    layer2_outputs(2684) <= not((layer1_outputs(9869)) xor (layer1_outputs(1636)));
    layer2_outputs(2685) <= not(layer1_outputs(1487));
    layer2_outputs(2686) <= not((layer1_outputs(7226)) and (layer1_outputs(3323)));
    layer2_outputs(2687) <= (layer1_outputs(8907)) and (layer1_outputs(8321));
    layer2_outputs(2688) <= not(layer1_outputs(3310));
    layer2_outputs(2689) <= not(layer1_outputs(9158));
    layer2_outputs(2690) <= layer1_outputs(9326);
    layer2_outputs(2691) <= not(layer1_outputs(4190));
    layer2_outputs(2692) <= (layer1_outputs(6039)) or (layer1_outputs(3678));
    layer2_outputs(2693) <= '0';
    layer2_outputs(2694) <= not((layer1_outputs(6556)) and (layer1_outputs(5597)));
    layer2_outputs(2695) <= not(layer1_outputs(9357));
    layer2_outputs(2696) <= not(layer1_outputs(9405));
    layer2_outputs(2697) <= layer1_outputs(4798);
    layer2_outputs(2698) <= (layer1_outputs(7787)) and not (layer1_outputs(7063));
    layer2_outputs(2699) <= layer1_outputs(2636);
    layer2_outputs(2700) <= not((layer1_outputs(3115)) and (layer1_outputs(8361)));
    layer2_outputs(2701) <= layer1_outputs(2467);
    layer2_outputs(2702) <= layer1_outputs(990);
    layer2_outputs(2703) <= not((layer1_outputs(1654)) and (layer1_outputs(3717)));
    layer2_outputs(2704) <= (layer1_outputs(6280)) or (layer1_outputs(8905));
    layer2_outputs(2705) <= (layer1_outputs(1080)) or (layer1_outputs(7421));
    layer2_outputs(2706) <= (layer1_outputs(929)) and not (layer1_outputs(9981));
    layer2_outputs(2707) <= layer1_outputs(3057);
    layer2_outputs(2708) <= not(layer1_outputs(6665)) or (layer1_outputs(190));
    layer2_outputs(2709) <= not(layer1_outputs(6147)) or (layer1_outputs(4595));
    layer2_outputs(2710) <= not(layer1_outputs(9784));
    layer2_outputs(2711) <= not(layer1_outputs(5188)) or (layer1_outputs(303));
    layer2_outputs(2712) <= not(layer1_outputs(1454));
    layer2_outputs(2713) <= (layer1_outputs(7886)) xor (layer1_outputs(4378));
    layer2_outputs(2714) <= not((layer1_outputs(8217)) xor (layer1_outputs(4879)));
    layer2_outputs(2715) <= layer1_outputs(8188);
    layer2_outputs(2716) <= (layer1_outputs(9923)) and not (layer1_outputs(2460));
    layer2_outputs(2717) <= not(layer1_outputs(3662));
    layer2_outputs(2718) <= not(layer1_outputs(3895));
    layer2_outputs(2719) <= not((layer1_outputs(8014)) or (layer1_outputs(8426)));
    layer2_outputs(2720) <= not(layer1_outputs(5966)) or (layer1_outputs(2443));
    layer2_outputs(2721) <= layer1_outputs(676);
    layer2_outputs(2722) <= not(layer1_outputs(870));
    layer2_outputs(2723) <= not((layer1_outputs(3767)) xor (layer1_outputs(7018)));
    layer2_outputs(2724) <= (layer1_outputs(4018)) or (layer1_outputs(3968));
    layer2_outputs(2725) <= not(layer1_outputs(5374));
    layer2_outputs(2726) <= not(layer1_outputs(9859));
    layer2_outputs(2727) <= layer1_outputs(6311);
    layer2_outputs(2728) <= not(layer1_outputs(6449)) or (layer1_outputs(2197));
    layer2_outputs(2729) <= layer1_outputs(4906);
    layer2_outputs(2730) <= not(layer1_outputs(4302)) or (layer1_outputs(10076));
    layer2_outputs(2731) <= (layer1_outputs(8049)) or (layer1_outputs(5695));
    layer2_outputs(2732) <= layer1_outputs(5057);
    layer2_outputs(2733) <= not((layer1_outputs(7900)) or (layer1_outputs(2474)));
    layer2_outputs(2734) <= not(layer1_outputs(1727)) or (layer1_outputs(9299));
    layer2_outputs(2735) <= (layer1_outputs(9105)) and (layer1_outputs(6387));
    layer2_outputs(2736) <= not(layer1_outputs(7359));
    layer2_outputs(2737) <= (layer1_outputs(3308)) and not (layer1_outputs(9340));
    layer2_outputs(2738) <= '0';
    layer2_outputs(2739) <= layer1_outputs(5654);
    layer2_outputs(2740) <= not((layer1_outputs(2133)) and (layer1_outputs(9396)));
    layer2_outputs(2741) <= (layer1_outputs(4016)) or (layer1_outputs(5135));
    layer2_outputs(2742) <= not(layer1_outputs(8506)) or (layer1_outputs(8068));
    layer2_outputs(2743) <= (layer1_outputs(4144)) and (layer1_outputs(5397));
    layer2_outputs(2744) <= not((layer1_outputs(7816)) or (layer1_outputs(9384)));
    layer2_outputs(2745) <= layer1_outputs(4389);
    layer2_outputs(2746) <= not((layer1_outputs(8395)) or (layer1_outputs(6395)));
    layer2_outputs(2747) <= layer1_outputs(4126);
    layer2_outputs(2748) <= not((layer1_outputs(10168)) xor (layer1_outputs(9570)));
    layer2_outputs(2749) <= layer1_outputs(1295);
    layer2_outputs(2750) <= (layer1_outputs(6382)) and not (layer1_outputs(4211));
    layer2_outputs(2751) <= (layer1_outputs(2247)) xor (layer1_outputs(1206));
    layer2_outputs(2752) <= not((layer1_outputs(8978)) xor (layer1_outputs(7560)));
    layer2_outputs(2753) <= (layer1_outputs(9440)) and (layer1_outputs(9602));
    layer2_outputs(2754) <= not(layer1_outputs(6641)) or (layer1_outputs(7087));
    layer2_outputs(2755) <= (layer1_outputs(4632)) and (layer1_outputs(7658));
    layer2_outputs(2756) <= layer1_outputs(3288);
    layer2_outputs(2757) <= not(layer1_outputs(7958));
    layer2_outputs(2758) <= layer1_outputs(10031);
    layer2_outputs(2759) <= (layer1_outputs(478)) or (layer1_outputs(780));
    layer2_outputs(2760) <= layer1_outputs(5047);
    layer2_outputs(2761) <= not(layer1_outputs(6878));
    layer2_outputs(2762) <= layer1_outputs(7634);
    layer2_outputs(2763) <= (layer1_outputs(9801)) and not (layer1_outputs(8574));
    layer2_outputs(2764) <= not(layer1_outputs(9682));
    layer2_outputs(2765) <= not(layer1_outputs(496)) or (layer1_outputs(7817));
    layer2_outputs(2766) <= (layer1_outputs(2291)) and (layer1_outputs(5713));
    layer2_outputs(2767) <= layer1_outputs(1629);
    layer2_outputs(2768) <= not(layer1_outputs(1646));
    layer2_outputs(2769) <= (layer1_outputs(9263)) and (layer1_outputs(2408));
    layer2_outputs(2770) <= (layer1_outputs(6260)) xor (layer1_outputs(4240));
    layer2_outputs(2771) <= layer1_outputs(3967);
    layer2_outputs(2772) <= layer1_outputs(1880);
    layer2_outputs(2773) <= not((layer1_outputs(8748)) xor (layer1_outputs(4327)));
    layer2_outputs(2774) <= not(layer1_outputs(7765));
    layer2_outputs(2775) <= not(layer1_outputs(9396));
    layer2_outputs(2776) <= not(layer1_outputs(4387));
    layer2_outputs(2777) <= not(layer1_outputs(2597)) or (layer1_outputs(248));
    layer2_outputs(2778) <= (layer1_outputs(3269)) or (layer1_outputs(8984));
    layer2_outputs(2779) <= not((layer1_outputs(5667)) or (layer1_outputs(3272)));
    layer2_outputs(2780) <= not(layer1_outputs(3568)) or (layer1_outputs(3046));
    layer2_outputs(2781) <= (layer1_outputs(3978)) or (layer1_outputs(6165));
    layer2_outputs(2782) <= not((layer1_outputs(1338)) and (layer1_outputs(5780)));
    layer2_outputs(2783) <= not(layer1_outputs(9639));
    layer2_outputs(2784) <= not(layer1_outputs(596));
    layer2_outputs(2785) <= layer1_outputs(196);
    layer2_outputs(2786) <= (layer1_outputs(3132)) xor (layer1_outputs(3594));
    layer2_outputs(2787) <= (layer1_outputs(2740)) and not (layer1_outputs(8509));
    layer2_outputs(2788) <= layer1_outputs(5794);
    layer2_outputs(2789) <= layer1_outputs(4713);
    layer2_outputs(2790) <= (layer1_outputs(642)) or (layer1_outputs(1207));
    layer2_outputs(2791) <= (layer1_outputs(3531)) xor (layer1_outputs(2860));
    layer2_outputs(2792) <= not(layer1_outputs(143));
    layer2_outputs(2793) <= layer1_outputs(8384);
    layer2_outputs(2794) <= not(layer1_outputs(5721));
    layer2_outputs(2795) <= not(layer1_outputs(7596));
    layer2_outputs(2796) <= not((layer1_outputs(2982)) xor (layer1_outputs(124)));
    layer2_outputs(2797) <= layer1_outputs(4246);
    layer2_outputs(2798) <= not(layer1_outputs(1778)) or (layer1_outputs(1971));
    layer2_outputs(2799) <= layer1_outputs(8372);
    layer2_outputs(2800) <= (layer1_outputs(1943)) and not (layer1_outputs(61));
    layer2_outputs(2801) <= not(layer1_outputs(8286));
    layer2_outputs(2802) <= (layer1_outputs(9899)) xor (layer1_outputs(3084));
    layer2_outputs(2803) <= not(layer1_outputs(9175));
    layer2_outputs(2804) <= not(layer1_outputs(3571)) or (layer1_outputs(2503));
    layer2_outputs(2805) <= not(layer1_outputs(1991)) or (layer1_outputs(3891));
    layer2_outputs(2806) <= (layer1_outputs(1671)) and (layer1_outputs(5624));
    layer2_outputs(2807) <= layer1_outputs(4440);
    layer2_outputs(2808) <= not(layer1_outputs(3150));
    layer2_outputs(2809) <= not(layer1_outputs(7692));
    layer2_outputs(2810) <= (layer1_outputs(999)) xor (layer1_outputs(8909));
    layer2_outputs(2811) <= not(layer1_outputs(4609));
    layer2_outputs(2812) <= not(layer1_outputs(2217)) or (layer1_outputs(4323));
    layer2_outputs(2813) <= (layer1_outputs(1582)) and (layer1_outputs(2152));
    layer2_outputs(2814) <= not((layer1_outputs(1115)) xor (layer1_outputs(6648)));
    layer2_outputs(2815) <= not(layer1_outputs(7444));
    layer2_outputs(2816) <= layer1_outputs(10204);
    layer2_outputs(2817) <= layer1_outputs(3478);
    layer2_outputs(2818) <= not(layer1_outputs(2932));
    layer2_outputs(2819) <= layer1_outputs(5155);
    layer2_outputs(2820) <= not(layer1_outputs(962));
    layer2_outputs(2821) <= not((layer1_outputs(2175)) or (layer1_outputs(5324)));
    layer2_outputs(2822) <= (layer1_outputs(5697)) and not (layer1_outputs(7217));
    layer2_outputs(2823) <= layer1_outputs(9208);
    layer2_outputs(2824) <= layer1_outputs(1252);
    layer2_outputs(2825) <= not((layer1_outputs(3330)) or (layer1_outputs(1794)));
    layer2_outputs(2826) <= (layer1_outputs(239)) and not (layer1_outputs(6516));
    layer2_outputs(2827) <= layer1_outputs(3103);
    layer2_outputs(2828) <= layer1_outputs(10177);
    layer2_outputs(2829) <= (layer1_outputs(8799)) xor (layer1_outputs(2719));
    layer2_outputs(2830) <= layer1_outputs(6268);
    layer2_outputs(2831) <= not(layer1_outputs(2237));
    layer2_outputs(2832) <= not(layer1_outputs(28));
    layer2_outputs(2833) <= (layer1_outputs(3901)) xor (layer1_outputs(693));
    layer2_outputs(2834) <= not(layer1_outputs(5358));
    layer2_outputs(2835) <= not(layer1_outputs(9759));
    layer2_outputs(2836) <= not(layer1_outputs(6418));
    layer2_outputs(2837) <= not(layer1_outputs(7405));
    layer2_outputs(2838) <= layer1_outputs(6752);
    layer2_outputs(2839) <= layer1_outputs(6052);
    layer2_outputs(2840) <= (layer1_outputs(750)) and (layer1_outputs(1491));
    layer2_outputs(2841) <= not(layer1_outputs(7545));
    layer2_outputs(2842) <= '1';
    layer2_outputs(2843) <= not(layer1_outputs(3068));
    layer2_outputs(2844) <= (layer1_outputs(7943)) xor (layer1_outputs(5871));
    layer2_outputs(2845) <= layer1_outputs(6514);
    layer2_outputs(2846) <= not(layer1_outputs(7666));
    layer2_outputs(2847) <= not((layer1_outputs(8576)) or (layer1_outputs(6173)));
    layer2_outputs(2848) <= layer1_outputs(6070);
    layer2_outputs(2849) <= layer1_outputs(3487);
    layer2_outputs(2850) <= not((layer1_outputs(6910)) or (layer1_outputs(3429)));
    layer2_outputs(2851) <= not((layer1_outputs(2120)) and (layer1_outputs(4680)));
    layer2_outputs(2852) <= layer1_outputs(9700);
    layer2_outputs(2853) <= not(layer1_outputs(5752));
    layer2_outputs(2854) <= layer1_outputs(1302);
    layer2_outputs(2855) <= not(layer1_outputs(8802));
    layer2_outputs(2856) <= layer1_outputs(8764);
    layer2_outputs(2857) <= layer1_outputs(9081);
    layer2_outputs(2858) <= not(layer1_outputs(7126));
    layer2_outputs(2859) <= layer1_outputs(575);
    layer2_outputs(2860) <= not(layer1_outputs(8061));
    layer2_outputs(2861) <= not(layer1_outputs(1369));
    layer2_outputs(2862) <= (layer1_outputs(3041)) and not (layer1_outputs(7645));
    layer2_outputs(2863) <= (layer1_outputs(5457)) xor (layer1_outputs(1008));
    layer2_outputs(2864) <= layer1_outputs(8350);
    layer2_outputs(2865) <= not((layer1_outputs(4810)) or (layer1_outputs(4004)));
    layer2_outputs(2866) <= not((layer1_outputs(6866)) and (layer1_outputs(6620)));
    layer2_outputs(2867) <= layer1_outputs(4649);
    layer2_outputs(2868) <= not(layer1_outputs(9896));
    layer2_outputs(2869) <= (layer1_outputs(4173)) and not (layer1_outputs(5110));
    layer2_outputs(2870) <= not(layer1_outputs(22));
    layer2_outputs(2871) <= not((layer1_outputs(5698)) and (layer1_outputs(392)));
    layer2_outputs(2872) <= not((layer1_outputs(388)) xor (layer1_outputs(6906)));
    layer2_outputs(2873) <= not(layer1_outputs(7566));
    layer2_outputs(2874) <= layer1_outputs(8814);
    layer2_outputs(2875) <= not(layer1_outputs(9659));
    layer2_outputs(2876) <= (layer1_outputs(4519)) xor (layer1_outputs(5971));
    layer2_outputs(2877) <= (layer1_outputs(4396)) xor (layer1_outputs(6952));
    layer2_outputs(2878) <= layer1_outputs(6198);
    layer2_outputs(2879) <= layer1_outputs(5161);
    layer2_outputs(2880) <= not(layer1_outputs(52));
    layer2_outputs(2881) <= not(layer1_outputs(1468)) or (layer1_outputs(4195));
    layer2_outputs(2882) <= layer1_outputs(4751);
    layer2_outputs(2883) <= not(layer1_outputs(7464));
    layer2_outputs(2884) <= not((layer1_outputs(1948)) and (layer1_outputs(9411)));
    layer2_outputs(2885) <= not(layer1_outputs(9111));
    layer2_outputs(2886) <= not(layer1_outputs(100)) or (layer1_outputs(1214));
    layer2_outputs(2887) <= not(layer1_outputs(403));
    layer2_outputs(2888) <= not(layer1_outputs(3126)) or (layer1_outputs(7583));
    layer2_outputs(2889) <= not(layer1_outputs(1765)) or (layer1_outputs(9188));
    layer2_outputs(2890) <= '1';
    layer2_outputs(2891) <= layer1_outputs(5552);
    layer2_outputs(2892) <= not(layer1_outputs(2288)) or (layer1_outputs(4482));
    layer2_outputs(2893) <= layer1_outputs(3334);
    layer2_outputs(2894) <= not(layer1_outputs(7814));
    layer2_outputs(2895) <= not(layer1_outputs(5824));
    layer2_outputs(2896) <= not(layer1_outputs(717));
    layer2_outputs(2897) <= layer1_outputs(4261);
    layer2_outputs(2898) <= not(layer1_outputs(7572)) or (layer1_outputs(5619));
    layer2_outputs(2899) <= '0';
    layer2_outputs(2900) <= layer1_outputs(1589);
    layer2_outputs(2901) <= layer1_outputs(2036);
    layer2_outputs(2902) <= not(layer1_outputs(979));
    layer2_outputs(2903) <= (layer1_outputs(8396)) and not (layer1_outputs(873));
    layer2_outputs(2904) <= not(layer1_outputs(6646));
    layer2_outputs(2905) <= not(layer1_outputs(4412));
    layer2_outputs(2906) <= (layer1_outputs(2673)) and (layer1_outputs(1411));
    layer2_outputs(2907) <= not((layer1_outputs(2324)) xor (layer1_outputs(3603)));
    layer2_outputs(2908) <= layer1_outputs(647);
    layer2_outputs(2909) <= layer1_outputs(6030);
    layer2_outputs(2910) <= not((layer1_outputs(9180)) or (layer1_outputs(2576)));
    layer2_outputs(2911) <= layer1_outputs(4191);
    layer2_outputs(2912) <= not((layer1_outputs(4930)) xor (layer1_outputs(2200)));
    layer2_outputs(2913) <= not((layer1_outputs(1708)) or (layer1_outputs(5903)));
    layer2_outputs(2914) <= layer1_outputs(3081);
    layer2_outputs(2915) <= layer1_outputs(7328);
    layer2_outputs(2916) <= (layer1_outputs(9655)) and not (layer1_outputs(5895));
    layer2_outputs(2917) <= (layer1_outputs(2510)) xor (layer1_outputs(1686));
    layer2_outputs(2918) <= '1';
    layer2_outputs(2919) <= not(layer1_outputs(305));
    layer2_outputs(2920) <= not(layer1_outputs(8645)) or (layer1_outputs(7295));
    layer2_outputs(2921) <= not((layer1_outputs(8499)) xor (layer1_outputs(157)));
    layer2_outputs(2922) <= not(layer1_outputs(977));
    layer2_outputs(2923) <= not(layer1_outputs(3974)) or (layer1_outputs(8756));
    layer2_outputs(2924) <= layer1_outputs(1563);
    layer2_outputs(2925) <= not((layer1_outputs(6787)) xor (layer1_outputs(2154)));
    layer2_outputs(2926) <= not((layer1_outputs(2450)) or (layer1_outputs(7770)));
    layer2_outputs(2927) <= layer1_outputs(6472);
    layer2_outputs(2928) <= layer1_outputs(1336);
    layer2_outputs(2929) <= layer1_outputs(3244);
    layer2_outputs(2930) <= (layer1_outputs(9948)) and not (layer1_outputs(6010));
    layer2_outputs(2931) <= not(layer1_outputs(3918));
    layer2_outputs(2932) <= not(layer1_outputs(1879));
    layer2_outputs(2933) <= (layer1_outputs(7208)) xor (layer1_outputs(6639));
    layer2_outputs(2934) <= not(layer1_outputs(5780)) or (layer1_outputs(7462));
    layer2_outputs(2935) <= '1';
    layer2_outputs(2936) <= not(layer1_outputs(2092));
    layer2_outputs(2937) <= layer1_outputs(7699);
    layer2_outputs(2938) <= layer1_outputs(8699);
    layer2_outputs(2939) <= layer1_outputs(9649);
    layer2_outputs(2940) <= not(layer1_outputs(1212));
    layer2_outputs(2941) <= layer1_outputs(4924);
    layer2_outputs(2942) <= (layer1_outputs(2351)) xor (layer1_outputs(7096));
    layer2_outputs(2943) <= (layer1_outputs(8001)) xor (layer1_outputs(7188));
    layer2_outputs(2944) <= layer1_outputs(7811);
    layer2_outputs(2945) <= layer1_outputs(221);
    layer2_outputs(2946) <= (layer1_outputs(8552)) xor (layer1_outputs(8084));
    layer2_outputs(2947) <= not((layer1_outputs(146)) or (layer1_outputs(6225)));
    layer2_outputs(2948) <= layer1_outputs(6487);
    layer2_outputs(2949) <= not(layer1_outputs(64)) or (layer1_outputs(6927));
    layer2_outputs(2950) <= layer1_outputs(3059);
    layer2_outputs(2951) <= layer1_outputs(9843);
    layer2_outputs(2952) <= not(layer1_outputs(7674));
    layer2_outputs(2953) <= not(layer1_outputs(7059));
    layer2_outputs(2954) <= (layer1_outputs(443)) xor (layer1_outputs(8661));
    layer2_outputs(2955) <= layer1_outputs(9863);
    layer2_outputs(2956) <= not(layer1_outputs(4865));
    layer2_outputs(2957) <= not((layer1_outputs(2817)) xor (layer1_outputs(3789)));
    layer2_outputs(2958) <= layer1_outputs(6665);
    layer2_outputs(2959) <= layer1_outputs(688);
    layer2_outputs(2960) <= not((layer1_outputs(9852)) xor (layer1_outputs(591)));
    layer2_outputs(2961) <= layer1_outputs(7523);
    layer2_outputs(2962) <= layer1_outputs(701);
    layer2_outputs(2963) <= (layer1_outputs(4508)) and not (layer1_outputs(1909));
    layer2_outputs(2964) <= not((layer1_outputs(7761)) xor (layer1_outputs(1891)));
    layer2_outputs(2965) <= not((layer1_outputs(6324)) and (layer1_outputs(9002)));
    layer2_outputs(2966) <= layer1_outputs(7055);
    layer2_outputs(2967) <= not(layer1_outputs(2736));
    layer2_outputs(2968) <= layer1_outputs(6747);
    layer2_outputs(2969) <= not(layer1_outputs(7825));
    layer2_outputs(2970) <= layer1_outputs(7133);
    layer2_outputs(2971) <= not((layer1_outputs(999)) xor (layer1_outputs(7475)));
    layer2_outputs(2972) <= not(layer1_outputs(154)) or (layer1_outputs(2668));
    layer2_outputs(2973) <= layer1_outputs(711);
    layer2_outputs(2974) <= (layer1_outputs(554)) and (layer1_outputs(3441));
    layer2_outputs(2975) <= layer1_outputs(7340);
    layer2_outputs(2976) <= layer1_outputs(4298);
    layer2_outputs(2977) <= not((layer1_outputs(6632)) xor (layer1_outputs(7516)));
    layer2_outputs(2978) <= layer1_outputs(10043);
    layer2_outputs(2979) <= not(layer1_outputs(9414));
    layer2_outputs(2980) <= layer1_outputs(5977);
    layer2_outputs(2981) <= layer1_outputs(9942);
    layer2_outputs(2982) <= layer1_outputs(9275);
    layer2_outputs(2983) <= layer1_outputs(792);
    layer2_outputs(2984) <= (layer1_outputs(7739)) and not (layer1_outputs(752));
    layer2_outputs(2985) <= layer1_outputs(8903);
    layer2_outputs(2986) <= layer1_outputs(374);
    layer2_outputs(2987) <= layer1_outputs(9683);
    layer2_outputs(2988) <= layer1_outputs(1475);
    layer2_outputs(2989) <= not(layer1_outputs(681));
    layer2_outputs(2990) <= not(layer1_outputs(4893));
    layer2_outputs(2991) <= not(layer1_outputs(397));
    layer2_outputs(2992) <= layer1_outputs(1583);
    layer2_outputs(2993) <= (layer1_outputs(10186)) xor (layer1_outputs(2247));
    layer2_outputs(2994) <= not(layer1_outputs(6666));
    layer2_outputs(2995) <= layer1_outputs(3103);
    layer2_outputs(2996) <= layer1_outputs(3113);
    layer2_outputs(2997) <= not((layer1_outputs(9983)) and (layer1_outputs(7722)));
    layer2_outputs(2998) <= not(layer1_outputs(6513));
    layer2_outputs(2999) <= not(layer1_outputs(5462));
    layer2_outputs(3000) <= (layer1_outputs(1726)) xor (layer1_outputs(7511));
    layer2_outputs(3001) <= not(layer1_outputs(3386));
    layer2_outputs(3002) <= not(layer1_outputs(4341)) or (layer1_outputs(5321));
    layer2_outputs(3003) <= layer1_outputs(3590);
    layer2_outputs(3004) <= layer1_outputs(4566);
    layer2_outputs(3005) <= not((layer1_outputs(6173)) or (layer1_outputs(9762)));
    layer2_outputs(3006) <= not(layer1_outputs(8828));
    layer2_outputs(3007) <= layer1_outputs(4636);
    layer2_outputs(3008) <= not(layer1_outputs(8602));
    layer2_outputs(3009) <= (layer1_outputs(9893)) xor (layer1_outputs(5547));
    layer2_outputs(3010) <= (layer1_outputs(3793)) and (layer1_outputs(6949));
    layer2_outputs(3011) <= not(layer1_outputs(7076)) or (layer1_outputs(1370));
    layer2_outputs(3012) <= (layer1_outputs(937)) or (layer1_outputs(6960));
    layer2_outputs(3013) <= layer1_outputs(9427);
    layer2_outputs(3014) <= not(layer1_outputs(3533));
    layer2_outputs(3015) <= not(layer1_outputs(3282));
    layer2_outputs(3016) <= not(layer1_outputs(9577));
    layer2_outputs(3017) <= not(layer1_outputs(2680));
    layer2_outputs(3018) <= layer1_outputs(4141);
    layer2_outputs(3019) <= layer1_outputs(687);
    layer2_outputs(3020) <= '1';
    layer2_outputs(3021) <= (layer1_outputs(3552)) and not (layer1_outputs(2025));
    layer2_outputs(3022) <= (layer1_outputs(1070)) xor (layer1_outputs(10153));
    layer2_outputs(3023) <= not((layer1_outputs(8312)) or (layer1_outputs(4860)));
    layer2_outputs(3024) <= not(layer1_outputs(1649));
    layer2_outputs(3025) <= layer1_outputs(3123);
    layer2_outputs(3026) <= layer1_outputs(5337);
    layer2_outputs(3027) <= not((layer1_outputs(549)) or (layer1_outputs(3133)));
    layer2_outputs(3028) <= not(layer1_outputs(1534));
    layer2_outputs(3029) <= layer1_outputs(7266);
    layer2_outputs(3030) <= layer1_outputs(260);
    layer2_outputs(3031) <= layer1_outputs(3473);
    layer2_outputs(3032) <= layer1_outputs(5288);
    layer2_outputs(3033) <= not((layer1_outputs(3635)) or (layer1_outputs(10133)));
    layer2_outputs(3034) <= (layer1_outputs(3964)) and not (layer1_outputs(1942));
    layer2_outputs(3035) <= not((layer1_outputs(2935)) xor (layer1_outputs(3405)));
    layer2_outputs(3036) <= layer1_outputs(6839);
    layer2_outputs(3037) <= layer1_outputs(2614);
    layer2_outputs(3038) <= (layer1_outputs(2915)) and not (layer1_outputs(2313));
    layer2_outputs(3039) <= not(layer1_outputs(1105));
    layer2_outputs(3040) <= not(layer1_outputs(8146));
    layer2_outputs(3041) <= not((layer1_outputs(6812)) xor (layer1_outputs(2725)));
    layer2_outputs(3042) <= layer1_outputs(2235);
    layer2_outputs(3043) <= not(layer1_outputs(7519)) or (layer1_outputs(3668));
    layer2_outputs(3044) <= not(layer1_outputs(3271));
    layer2_outputs(3045) <= not(layer1_outputs(3182));
    layer2_outputs(3046) <= (layer1_outputs(7473)) and (layer1_outputs(8725));
    layer2_outputs(3047) <= not((layer1_outputs(7443)) and (layer1_outputs(5997)));
    layer2_outputs(3048) <= layer1_outputs(3886);
    layer2_outputs(3049) <= not(layer1_outputs(7127));
    layer2_outputs(3050) <= (layer1_outputs(2930)) xor (layer1_outputs(3931));
    layer2_outputs(3051) <= layer1_outputs(6540);
    layer2_outputs(3052) <= not(layer1_outputs(1615));
    layer2_outputs(3053) <= (layer1_outputs(7672)) and not (layer1_outputs(3973));
    layer2_outputs(3054) <= not(layer1_outputs(5154));
    layer2_outputs(3055) <= not((layer1_outputs(6380)) xor (layer1_outputs(75)));
    layer2_outputs(3056) <= not(layer1_outputs(6793)) or (layer1_outputs(9636));
    layer2_outputs(3057) <= (layer1_outputs(3887)) xor (layer1_outputs(3342));
    layer2_outputs(3058) <= (layer1_outputs(49)) and not (layer1_outputs(4413));
    layer2_outputs(3059) <= (layer1_outputs(4340)) and (layer1_outputs(4673));
    layer2_outputs(3060) <= layer1_outputs(4296);
    layer2_outputs(3061) <= not(layer1_outputs(6494));
    layer2_outputs(3062) <= (layer1_outputs(3220)) or (layer1_outputs(7768));
    layer2_outputs(3063) <= (layer1_outputs(5620)) xor (layer1_outputs(2948));
    layer2_outputs(3064) <= (layer1_outputs(8832)) and (layer1_outputs(8943));
    layer2_outputs(3065) <= not(layer1_outputs(4529)) or (layer1_outputs(8483));
    layer2_outputs(3066) <= layer1_outputs(8077);
    layer2_outputs(3067) <= layer1_outputs(3661);
    layer2_outputs(3068) <= not(layer1_outputs(3035));
    layer2_outputs(3069) <= (layer1_outputs(8466)) and not (layer1_outputs(7674));
    layer2_outputs(3070) <= not((layer1_outputs(10090)) and (layer1_outputs(8609)));
    layer2_outputs(3071) <= not((layer1_outputs(9498)) or (layer1_outputs(4892)));
    layer2_outputs(3072) <= layer1_outputs(5166);
    layer2_outputs(3073) <= (layer1_outputs(4920)) and not (layer1_outputs(6379));
    layer2_outputs(3074) <= (layer1_outputs(1585)) or (layer1_outputs(7299));
    layer2_outputs(3075) <= not((layer1_outputs(3825)) xor (layer1_outputs(1207)));
    layer2_outputs(3076) <= not((layer1_outputs(4224)) and (layer1_outputs(2007)));
    layer2_outputs(3077) <= not(layer1_outputs(3854));
    layer2_outputs(3078) <= not(layer1_outputs(7682));
    layer2_outputs(3079) <= not((layer1_outputs(4025)) xor (layer1_outputs(7782)));
    layer2_outputs(3080) <= not(layer1_outputs(1641));
    layer2_outputs(3081) <= (layer1_outputs(1846)) xor (layer1_outputs(6476));
    layer2_outputs(3082) <= not((layer1_outputs(1602)) and (layer1_outputs(8192)));
    layer2_outputs(3083) <= not((layer1_outputs(9478)) and (layer1_outputs(3128)));
    layer2_outputs(3084) <= (layer1_outputs(5848)) and (layer1_outputs(7041));
    layer2_outputs(3085) <= layer1_outputs(2589);
    layer2_outputs(3086) <= (layer1_outputs(4447)) and not (layer1_outputs(1751));
    layer2_outputs(3087) <= not((layer1_outputs(3938)) and (layer1_outputs(417)));
    layer2_outputs(3088) <= not(layer1_outputs(6559)) or (layer1_outputs(9678));
    layer2_outputs(3089) <= not(layer1_outputs(696));
    layer2_outputs(3090) <= layer1_outputs(6402);
    layer2_outputs(3091) <= not(layer1_outputs(2988));
    layer2_outputs(3092) <= layer1_outputs(6045);
    layer2_outputs(3093) <= not((layer1_outputs(9732)) and (layer1_outputs(5461)));
    layer2_outputs(3094) <= layer1_outputs(9001);
    layer2_outputs(3095) <= layer1_outputs(9728);
    layer2_outputs(3096) <= not((layer1_outputs(1514)) xor (layer1_outputs(7291)));
    layer2_outputs(3097) <= not(layer1_outputs(304));
    layer2_outputs(3098) <= not((layer1_outputs(10006)) and (layer1_outputs(9272)));
    layer2_outputs(3099) <= not(layer1_outputs(690)) or (layer1_outputs(7738));
    layer2_outputs(3100) <= (layer1_outputs(2511)) and (layer1_outputs(7587));
    layer2_outputs(3101) <= not((layer1_outputs(660)) and (layer1_outputs(6392)));
    layer2_outputs(3102) <= (layer1_outputs(4863)) and (layer1_outputs(9747));
    layer2_outputs(3103) <= not(layer1_outputs(1440));
    layer2_outputs(3104) <= (layer1_outputs(3362)) and not (layer1_outputs(6145));
    layer2_outputs(3105) <= not(layer1_outputs(287)) or (layer1_outputs(4404));
    layer2_outputs(3106) <= (layer1_outputs(5391)) and not (layer1_outputs(7923));
    layer2_outputs(3107) <= not((layer1_outputs(2756)) or (layer1_outputs(8350)));
    layer2_outputs(3108) <= (layer1_outputs(3947)) and not (layer1_outputs(5219));
    layer2_outputs(3109) <= layer1_outputs(6367);
    layer2_outputs(3110) <= not((layer1_outputs(1420)) xor (layer1_outputs(8416)));
    layer2_outputs(3111) <= not(layer1_outputs(5907));
    layer2_outputs(3112) <= not(layer1_outputs(2557));
    layer2_outputs(3113) <= not(layer1_outputs(2830)) or (layer1_outputs(15));
    layer2_outputs(3114) <= layer1_outputs(2653);
    layer2_outputs(3115) <= not(layer1_outputs(8094));
    layer2_outputs(3116) <= not(layer1_outputs(4335));
    layer2_outputs(3117) <= (layer1_outputs(1517)) and not (layer1_outputs(2677));
    layer2_outputs(3118) <= '0';
    layer2_outputs(3119) <= not(layer1_outputs(7055)) or (layer1_outputs(9434));
    layer2_outputs(3120) <= not(layer1_outputs(9443));
    layer2_outputs(3121) <= '0';
    layer2_outputs(3122) <= not(layer1_outputs(2580)) or (layer1_outputs(8759));
    layer2_outputs(3123) <= (layer1_outputs(76)) and (layer1_outputs(6860));
    layer2_outputs(3124) <= layer1_outputs(3872);
    layer2_outputs(3125) <= not((layer1_outputs(1208)) or (layer1_outputs(369)));
    layer2_outputs(3126) <= not((layer1_outputs(8338)) and (layer1_outputs(2831)));
    layer2_outputs(3127) <= not(layer1_outputs(7315));
    layer2_outputs(3128) <= (layer1_outputs(8229)) and not (layer1_outputs(3423));
    layer2_outputs(3129) <= not(layer1_outputs(5408));
    layer2_outputs(3130) <= (layer1_outputs(7665)) xor (layer1_outputs(9198));
    layer2_outputs(3131) <= not((layer1_outputs(2933)) xor (layer1_outputs(895)));
    layer2_outputs(3132) <= not(layer1_outputs(3835));
    layer2_outputs(3133) <= layer1_outputs(6532);
    layer2_outputs(3134) <= not(layer1_outputs(9694));
    layer2_outputs(3135) <= layer1_outputs(1734);
    layer2_outputs(3136) <= layer1_outputs(4258);
    layer2_outputs(3137) <= (layer1_outputs(7987)) and (layer1_outputs(7565));
    layer2_outputs(3138) <= not(layer1_outputs(6061));
    layer2_outputs(3139) <= not(layer1_outputs(8629)) or (layer1_outputs(6564));
    layer2_outputs(3140) <= (layer1_outputs(9849)) and (layer1_outputs(4623));
    layer2_outputs(3141) <= (layer1_outputs(8444)) and not (layer1_outputs(6097));
    layer2_outputs(3142) <= layer1_outputs(3490);
    layer2_outputs(3143) <= not(layer1_outputs(1492));
    layer2_outputs(3144) <= (layer1_outputs(8079)) or (layer1_outputs(5584));
    layer2_outputs(3145) <= not(layer1_outputs(7540));
    layer2_outputs(3146) <= layer1_outputs(6113);
    layer2_outputs(3147) <= layer1_outputs(2258);
    layer2_outputs(3148) <= (layer1_outputs(4482)) or (layer1_outputs(534));
    layer2_outputs(3149) <= not((layer1_outputs(1832)) and (layer1_outputs(7116)));
    layer2_outputs(3150) <= not(layer1_outputs(1879)) or (layer1_outputs(1851));
    layer2_outputs(3151) <= (layer1_outputs(2439)) and not (layer1_outputs(4547));
    layer2_outputs(3152) <= layer1_outputs(830);
    layer2_outputs(3153) <= (layer1_outputs(5887)) xor (layer1_outputs(7622));
    layer2_outputs(3154) <= layer1_outputs(2028);
    layer2_outputs(3155) <= not(layer1_outputs(8065));
    layer2_outputs(3156) <= not((layer1_outputs(1312)) or (layer1_outputs(2568)));
    layer2_outputs(3157) <= (layer1_outputs(4618)) and not (layer1_outputs(4496));
    layer2_outputs(3158) <= (layer1_outputs(5375)) and not (layer1_outputs(8640));
    layer2_outputs(3159) <= (layer1_outputs(4559)) and not (layer1_outputs(7404));
    layer2_outputs(3160) <= not(layer1_outputs(6519));
    layer2_outputs(3161) <= not(layer1_outputs(7772));
    layer2_outputs(3162) <= (layer1_outputs(3925)) and (layer1_outputs(3614));
    layer2_outputs(3163) <= (layer1_outputs(7714)) or (layer1_outputs(352));
    layer2_outputs(3164) <= not(layer1_outputs(4341)) or (layer1_outputs(215));
    layer2_outputs(3165) <= layer1_outputs(852);
    layer2_outputs(3166) <= layer1_outputs(8404);
    layer2_outputs(3167) <= layer1_outputs(6546);
    layer2_outputs(3168) <= (layer1_outputs(7058)) xor (layer1_outputs(825));
    layer2_outputs(3169) <= not(layer1_outputs(220));
    layer2_outputs(3170) <= (layer1_outputs(7607)) xor (layer1_outputs(1870));
    layer2_outputs(3171) <= not(layer1_outputs(3001));
    layer2_outputs(3172) <= layer1_outputs(2553);
    layer2_outputs(3173) <= not(layer1_outputs(8878));
    layer2_outputs(3174) <= not(layer1_outputs(741));
    layer2_outputs(3175) <= not(layer1_outputs(10108));
    layer2_outputs(3176) <= layer1_outputs(4104);
    layer2_outputs(3177) <= layer1_outputs(8434);
    layer2_outputs(3178) <= not(layer1_outputs(3634));
    layer2_outputs(3179) <= (layer1_outputs(3728)) or (layer1_outputs(7982));
    layer2_outputs(3180) <= not(layer1_outputs(7960));
    layer2_outputs(3181) <= not(layer1_outputs(4434));
    layer2_outputs(3182) <= layer1_outputs(7602);
    layer2_outputs(3183) <= not(layer1_outputs(1984));
    layer2_outputs(3184) <= not(layer1_outputs(4552));
    layer2_outputs(3185) <= not(layer1_outputs(6609));
    layer2_outputs(3186) <= (layer1_outputs(4860)) xor (layer1_outputs(1193));
    layer2_outputs(3187) <= layer1_outputs(4452);
    layer2_outputs(3188) <= not(layer1_outputs(6518));
    layer2_outputs(3189) <= layer1_outputs(4392);
    layer2_outputs(3190) <= not(layer1_outputs(4601));
    layer2_outputs(3191) <= not(layer1_outputs(8611));
    layer2_outputs(3192) <= not((layer1_outputs(4076)) xor (layer1_outputs(1672)));
    layer2_outputs(3193) <= (layer1_outputs(3953)) and not (layer1_outputs(1963));
    layer2_outputs(3194) <= (layer1_outputs(8040)) and (layer1_outputs(9225));
    layer2_outputs(3195) <= layer1_outputs(1597);
    layer2_outputs(3196) <= not(layer1_outputs(5414));
    layer2_outputs(3197) <= (layer1_outputs(8282)) and not (layer1_outputs(8525));
    layer2_outputs(3198) <= not(layer1_outputs(6838));
    layer2_outputs(3199) <= layer1_outputs(1301);
    layer2_outputs(3200) <= layer1_outputs(8175);
    layer2_outputs(3201) <= layer1_outputs(8908);
    layer2_outputs(3202) <= not(layer1_outputs(3065));
    layer2_outputs(3203) <= (layer1_outputs(9905)) or (layer1_outputs(6416));
    layer2_outputs(3204) <= layer1_outputs(8909);
    layer2_outputs(3205) <= not(layer1_outputs(3864));
    layer2_outputs(3206) <= (layer1_outputs(4306)) and (layer1_outputs(5844));
    layer2_outputs(3207) <= (layer1_outputs(8076)) and not (layer1_outputs(6942));
    layer2_outputs(3208) <= layer1_outputs(2852);
    layer2_outputs(3209) <= not(layer1_outputs(4045)) or (layer1_outputs(1320));
    layer2_outputs(3210) <= layer1_outputs(3946);
    layer2_outputs(3211) <= (layer1_outputs(2236)) and not (layer1_outputs(5473));
    layer2_outputs(3212) <= not(layer1_outputs(2945));
    layer2_outputs(3213) <= layer1_outputs(2953);
    layer2_outputs(3214) <= layer1_outputs(7733);
    layer2_outputs(3215) <= not((layer1_outputs(7946)) and (layer1_outputs(3325)));
    layer2_outputs(3216) <= not(layer1_outputs(5065));
    layer2_outputs(3217) <= not(layer1_outputs(4111));
    layer2_outputs(3218) <= (layer1_outputs(7636)) and (layer1_outputs(5400));
    layer2_outputs(3219) <= layer1_outputs(2170);
    layer2_outputs(3220) <= '1';
    layer2_outputs(3221) <= not(layer1_outputs(8191));
    layer2_outputs(3222) <= not(layer1_outputs(8840)) or (layer1_outputs(1739));
    layer2_outputs(3223) <= not(layer1_outputs(7272));
    layer2_outputs(3224) <= layer1_outputs(179);
    layer2_outputs(3225) <= (layer1_outputs(675)) and (layer1_outputs(2581));
    layer2_outputs(3226) <= not(layer1_outputs(358));
    layer2_outputs(3227) <= not(layer1_outputs(2746));
    layer2_outputs(3228) <= (layer1_outputs(6694)) and (layer1_outputs(1507));
    layer2_outputs(3229) <= layer1_outputs(2263);
    layer2_outputs(3230) <= (layer1_outputs(4595)) and (layer1_outputs(7830));
    layer2_outputs(3231) <= layer1_outputs(10098);
    layer2_outputs(3232) <= not(layer1_outputs(3360));
    layer2_outputs(3233) <= not(layer1_outputs(423)) or (layer1_outputs(1519));
    layer2_outputs(3234) <= not(layer1_outputs(1499));
    layer2_outputs(3235) <= not(layer1_outputs(6934));
    layer2_outputs(3236) <= (layer1_outputs(3389)) and not (layer1_outputs(1179));
    layer2_outputs(3237) <= layer1_outputs(2807);
    layer2_outputs(3238) <= not(layer1_outputs(4653)) or (layer1_outputs(5996));
    layer2_outputs(3239) <= layer1_outputs(8079);
    layer2_outputs(3240) <= not(layer1_outputs(2806));
    layer2_outputs(3241) <= not(layer1_outputs(5941));
    layer2_outputs(3242) <= not(layer1_outputs(2186)) or (layer1_outputs(2704));
    layer2_outputs(3243) <= layer1_outputs(4900);
    layer2_outputs(3244) <= layer1_outputs(3325);
    layer2_outputs(3245) <= not(layer1_outputs(4869));
    layer2_outputs(3246) <= not(layer1_outputs(9313));
    layer2_outputs(3247) <= layer1_outputs(4251);
    layer2_outputs(3248) <= not(layer1_outputs(3544)) or (layer1_outputs(188));
    layer2_outputs(3249) <= layer1_outputs(3767);
    layer2_outputs(3250) <= not(layer1_outputs(4637));
    layer2_outputs(3251) <= (layer1_outputs(8269)) and not (layer1_outputs(9167));
    layer2_outputs(3252) <= (layer1_outputs(2906)) xor (layer1_outputs(1996));
    layer2_outputs(3253) <= not(layer1_outputs(9083));
    layer2_outputs(3254) <= (layer1_outputs(1531)) xor (layer1_outputs(7606));
    layer2_outputs(3255) <= layer1_outputs(8114);
    layer2_outputs(3256) <= (layer1_outputs(2512)) and (layer1_outputs(3428));
    layer2_outputs(3257) <= '0';
    layer2_outputs(3258) <= not((layer1_outputs(10132)) and (layer1_outputs(9616)));
    layer2_outputs(3259) <= not(layer1_outputs(4782));
    layer2_outputs(3260) <= (layer1_outputs(3122)) and (layer1_outputs(508));
    layer2_outputs(3261) <= not(layer1_outputs(6430));
    layer2_outputs(3262) <= layer1_outputs(4974);
    layer2_outputs(3263) <= not(layer1_outputs(39)) or (layer1_outputs(6937));
    layer2_outputs(3264) <= not(layer1_outputs(4790));
    layer2_outputs(3265) <= (layer1_outputs(3627)) and not (layer1_outputs(804));
    layer2_outputs(3266) <= layer1_outputs(4641);
    layer2_outputs(3267) <= not(layer1_outputs(4884));
    layer2_outputs(3268) <= layer1_outputs(6596);
    layer2_outputs(3269) <= layer1_outputs(4281);
    layer2_outputs(3270) <= not(layer1_outputs(3910));
    layer2_outputs(3271) <= layer1_outputs(6630);
    layer2_outputs(3272) <= not(layer1_outputs(2470));
    layer2_outputs(3273) <= not(layer1_outputs(3440));
    layer2_outputs(3274) <= not(layer1_outputs(6289));
    layer2_outputs(3275) <= (layer1_outputs(4250)) and not (layer1_outputs(4641));
    layer2_outputs(3276) <= not(layer1_outputs(7110));
    layer2_outputs(3277) <= layer1_outputs(8900);
    layer2_outputs(3278) <= not(layer1_outputs(3537));
    layer2_outputs(3279) <= not(layer1_outputs(119));
    layer2_outputs(3280) <= layer1_outputs(3169);
    layer2_outputs(3281) <= (layer1_outputs(4138)) and not (layer1_outputs(4923));
    layer2_outputs(3282) <= not(layer1_outputs(7263));
    layer2_outputs(3283) <= not((layer1_outputs(3998)) or (layer1_outputs(10069)));
    layer2_outputs(3284) <= not((layer1_outputs(2006)) or (layer1_outputs(2487)));
    layer2_outputs(3285) <= (layer1_outputs(6899)) xor (layer1_outputs(8921));
    layer2_outputs(3286) <= not(layer1_outputs(4446));
    layer2_outputs(3287) <= (layer1_outputs(6297)) xor (layer1_outputs(7968));
    layer2_outputs(3288) <= layer1_outputs(9287);
    layer2_outputs(3289) <= not(layer1_outputs(730));
    layer2_outputs(3290) <= layer1_outputs(19);
    layer2_outputs(3291) <= layer1_outputs(3468);
    layer2_outputs(3292) <= not(layer1_outputs(528));
    layer2_outputs(3293) <= not(layer1_outputs(7867));
    layer2_outputs(3294) <= (layer1_outputs(8615)) and (layer1_outputs(8455));
    layer2_outputs(3295) <= not(layer1_outputs(7648)) or (layer1_outputs(5756));
    layer2_outputs(3296) <= not((layer1_outputs(984)) or (layer1_outputs(4385)));
    layer2_outputs(3297) <= layer1_outputs(3146);
    layer2_outputs(3298) <= not(layer1_outputs(4804));
    layer2_outputs(3299) <= (layer1_outputs(5972)) and (layer1_outputs(7436));
    layer2_outputs(3300) <= layer1_outputs(3206);
    layer2_outputs(3301) <= not(layer1_outputs(2135));
    layer2_outputs(3302) <= (layer1_outputs(172)) xor (layer1_outputs(10171));
    layer2_outputs(3303) <= '0';
    layer2_outputs(3304) <= '1';
    layer2_outputs(3305) <= layer1_outputs(1721);
    layer2_outputs(3306) <= layer1_outputs(2481);
    layer2_outputs(3307) <= not((layer1_outputs(7103)) and (layer1_outputs(6806)));
    layer2_outputs(3308) <= not(layer1_outputs(1639));
    layer2_outputs(3309) <= layer1_outputs(4669);
    layer2_outputs(3310) <= (layer1_outputs(2909)) xor (layer1_outputs(9067));
    layer2_outputs(3311) <= not((layer1_outputs(3844)) xor (layer1_outputs(429)));
    layer2_outputs(3312) <= not((layer1_outputs(9809)) xor (layer1_outputs(6448)));
    layer2_outputs(3313) <= layer1_outputs(8790);
    layer2_outputs(3314) <= not(layer1_outputs(7423));
    layer2_outputs(3315) <= not((layer1_outputs(719)) and (layer1_outputs(7132)));
    layer2_outputs(3316) <= not((layer1_outputs(715)) or (layer1_outputs(7822)));
    layer2_outputs(3317) <= '1';
    layer2_outputs(3318) <= not(layer1_outputs(7757)) or (layer1_outputs(2519));
    layer2_outputs(3319) <= not(layer1_outputs(5557));
    layer2_outputs(3320) <= not((layer1_outputs(8777)) xor (layer1_outputs(1020)));
    layer2_outputs(3321) <= (layer1_outputs(1955)) and not (layer1_outputs(3019));
    layer2_outputs(3322) <= (layer1_outputs(8681)) and (layer1_outputs(1396));
    layer2_outputs(3323) <= not(layer1_outputs(1971));
    layer2_outputs(3324) <= layer1_outputs(1334);
    layer2_outputs(3325) <= layer1_outputs(3896);
    layer2_outputs(3326) <= not(layer1_outputs(2657));
    layer2_outputs(3327) <= layer1_outputs(5187);
    layer2_outputs(3328) <= not(layer1_outputs(6849)) or (layer1_outputs(2346));
    layer2_outputs(3329) <= not(layer1_outputs(3162));
    layer2_outputs(3330) <= not((layer1_outputs(9264)) and (layer1_outputs(1122)));
    layer2_outputs(3331) <= (layer1_outputs(3762)) and (layer1_outputs(9254));
    layer2_outputs(3332) <= not(layer1_outputs(3942));
    layer2_outputs(3333) <= not(layer1_outputs(3606));
    layer2_outputs(3334) <= not(layer1_outputs(99)) or (layer1_outputs(3480));
    layer2_outputs(3335) <= layer1_outputs(5540);
    layer2_outputs(3336) <= layer1_outputs(2558);
    layer2_outputs(3337) <= not(layer1_outputs(7551)) or (layer1_outputs(1568));
    layer2_outputs(3338) <= not(layer1_outputs(1918));
    layer2_outputs(3339) <= not((layer1_outputs(2983)) xor (layer1_outputs(5530)));
    layer2_outputs(3340) <= not(layer1_outputs(2951)) or (layer1_outputs(3042));
    layer2_outputs(3341) <= not(layer1_outputs(8369));
    layer2_outputs(3342) <= layer1_outputs(5297);
    layer2_outputs(3343) <= (layer1_outputs(5496)) and (layer1_outputs(1951));
    layer2_outputs(3344) <= layer1_outputs(1368);
    layer2_outputs(3345) <= not(layer1_outputs(4748));
    layer2_outputs(3346) <= not(layer1_outputs(637));
    layer2_outputs(3347) <= not(layer1_outputs(9353));
    layer2_outputs(3348) <= layer1_outputs(4349);
    layer2_outputs(3349) <= '1';
    layer2_outputs(3350) <= not(layer1_outputs(8772));
    layer2_outputs(3351) <= (layer1_outputs(5433)) and not (layer1_outputs(5613));
    layer2_outputs(3352) <= not(layer1_outputs(5152));
    layer2_outputs(3353) <= (layer1_outputs(2010)) and (layer1_outputs(3169));
    layer2_outputs(3354) <= not(layer1_outputs(8186));
    layer2_outputs(3355) <= layer1_outputs(4822);
    layer2_outputs(3356) <= (layer1_outputs(4081)) or (layer1_outputs(692));
    layer2_outputs(3357) <= layer1_outputs(4769);
    layer2_outputs(3358) <= not(layer1_outputs(293));
    layer2_outputs(3359) <= not(layer1_outputs(1323));
    layer2_outputs(3360) <= (layer1_outputs(2435)) and not (layer1_outputs(7340));
    layer2_outputs(3361) <= layer1_outputs(9560);
    layer2_outputs(3362) <= layer1_outputs(724);
    layer2_outputs(3363) <= layer1_outputs(8161);
    layer2_outputs(3364) <= not(layer1_outputs(1374)) or (layer1_outputs(2046));
    layer2_outputs(3365) <= (layer1_outputs(2653)) xor (layer1_outputs(5294));
    layer2_outputs(3366) <= not(layer1_outputs(4451));
    layer2_outputs(3367) <= layer1_outputs(7656);
    layer2_outputs(3368) <= not((layer1_outputs(10088)) or (layer1_outputs(2110)));
    layer2_outputs(3369) <= (layer1_outputs(9781)) and not (layer1_outputs(349));
    layer2_outputs(3370) <= not(layer1_outputs(2678));
    layer2_outputs(3371) <= not(layer1_outputs(2947)) or (layer1_outputs(8905));
    layer2_outputs(3372) <= (layer1_outputs(9355)) and not (layer1_outputs(9341));
    layer2_outputs(3373) <= (layer1_outputs(8331)) and not (layer1_outputs(134));
    layer2_outputs(3374) <= layer1_outputs(9089);
    layer2_outputs(3375) <= not(layer1_outputs(1449));
    layer2_outputs(3376) <= not(layer1_outputs(5559));
    layer2_outputs(3377) <= not((layer1_outputs(4291)) xor (layer1_outputs(4537)));
    layer2_outputs(3378) <= not((layer1_outputs(1739)) or (layer1_outputs(3027)));
    layer2_outputs(3379) <= layer1_outputs(5474);
    layer2_outputs(3380) <= (layer1_outputs(7879)) and (layer1_outputs(1351));
    layer2_outputs(3381) <= not(layer1_outputs(1061));
    layer2_outputs(3382) <= (layer1_outputs(2129)) and not (layer1_outputs(3666));
    layer2_outputs(3383) <= not((layer1_outputs(4615)) xor (layer1_outputs(10156)));
    layer2_outputs(3384) <= not((layer1_outputs(1997)) xor (layer1_outputs(9333)));
    layer2_outputs(3385) <= (layer1_outputs(3712)) and not (layer1_outputs(8127));
    layer2_outputs(3386) <= layer1_outputs(95);
    layer2_outputs(3387) <= not(layer1_outputs(2134)) or (layer1_outputs(851));
    layer2_outputs(3388) <= layer1_outputs(7526);
    layer2_outputs(3389) <= not((layer1_outputs(1580)) or (layer1_outputs(2477)));
    layer2_outputs(3390) <= layer1_outputs(3516);
    layer2_outputs(3391) <= (layer1_outputs(7717)) xor (layer1_outputs(4324));
    layer2_outputs(3392) <= layer1_outputs(7677);
    layer2_outputs(3393) <= layer1_outputs(9586);
    layer2_outputs(3394) <= layer1_outputs(7159);
    layer2_outputs(3395) <= layer1_outputs(9660);
    layer2_outputs(3396) <= layer1_outputs(5608);
    layer2_outputs(3397) <= not((layer1_outputs(5621)) xor (layer1_outputs(3723)));
    layer2_outputs(3398) <= layer1_outputs(4823);
    layer2_outputs(3399) <= layer1_outputs(9632);
    layer2_outputs(3400) <= not(layer1_outputs(6316));
    layer2_outputs(3401) <= not(layer1_outputs(1368));
    layer2_outputs(3402) <= layer1_outputs(8598);
    layer2_outputs(3403) <= not((layer1_outputs(1288)) xor (layer1_outputs(6553)));
    layer2_outputs(3404) <= (layer1_outputs(673)) xor (layer1_outputs(3805));
    layer2_outputs(3405) <= not((layer1_outputs(6183)) or (layer1_outputs(5156)));
    layer2_outputs(3406) <= not(layer1_outputs(859)) or (layer1_outputs(1819));
    layer2_outputs(3407) <= not(layer1_outputs(296));
    layer2_outputs(3408) <= layer1_outputs(3837);
    layer2_outputs(3409) <= layer1_outputs(5367);
    layer2_outputs(3410) <= not(layer1_outputs(5171));
    layer2_outputs(3411) <= layer1_outputs(422);
    layer2_outputs(3412) <= not((layer1_outputs(6863)) xor (layer1_outputs(4796)));
    layer2_outputs(3413) <= not(layer1_outputs(10095));
    layer2_outputs(3414) <= not(layer1_outputs(9071));
    layer2_outputs(3415) <= layer1_outputs(3366);
    layer2_outputs(3416) <= not(layer1_outputs(5276));
    layer2_outputs(3417) <= not(layer1_outputs(6366));
    layer2_outputs(3418) <= not(layer1_outputs(9729));
    layer2_outputs(3419) <= layer1_outputs(4379);
    layer2_outputs(3420) <= (layer1_outputs(545)) xor (layer1_outputs(7307));
    layer2_outputs(3421) <= (layer1_outputs(3005)) or (layer1_outputs(10065));
    layer2_outputs(3422) <= (layer1_outputs(2152)) and not (layer1_outputs(4102));
    layer2_outputs(3423) <= not(layer1_outputs(406));
    layer2_outputs(3424) <= (layer1_outputs(7877)) and not (layer1_outputs(9072));
    layer2_outputs(3425) <= layer1_outputs(3332);
    layer2_outputs(3426) <= not(layer1_outputs(6390));
    layer2_outputs(3427) <= not(layer1_outputs(6557));
    layer2_outputs(3428) <= not(layer1_outputs(10020));
    layer2_outputs(3429) <= not(layer1_outputs(6281));
    layer2_outputs(3430) <= '0';
    layer2_outputs(3431) <= (layer1_outputs(5315)) or (layer1_outputs(282));
    layer2_outputs(3432) <= not(layer1_outputs(8932)) or (layer1_outputs(5347));
    layer2_outputs(3433) <= not((layer1_outputs(1685)) xor (layer1_outputs(564)));
    layer2_outputs(3434) <= (layer1_outputs(6178)) and (layer1_outputs(7113));
    layer2_outputs(3435) <= not((layer1_outputs(7874)) and (layer1_outputs(1865)));
    layer2_outputs(3436) <= layer1_outputs(7169);
    layer2_outputs(3437) <= layer1_outputs(7529);
    layer2_outputs(3438) <= not((layer1_outputs(3316)) xor (layer1_outputs(1538)));
    layer2_outputs(3439) <= layer1_outputs(4417);
    layer2_outputs(3440) <= not(layer1_outputs(8240));
    layer2_outputs(3441) <= layer1_outputs(4623);
    layer2_outputs(3442) <= (layer1_outputs(8945)) xor (layer1_outputs(7610));
    layer2_outputs(3443) <= (layer1_outputs(6779)) xor (layer1_outputs(3832));
    layer2_outputs(3444) <= not(layer1_outputs(9569)) or (layer1_outputs(314));
    layer2_outputs(3445) <= (layer1_outputs(900)) or (layer1_outputs(763));
    layer2_outputs(3446) <= not(layer1_outputs(3905));
    layer2_outputs(3447) <= layer1_outputs(8397);
    layer2_outputs(3448) <= not((layer1_outputs(9002)) xor (layer1_outputs(5267)));
    layer2_outputs(3449) <= not((layer1_outputs(2525)) xor (layer1_outputs(5732)));
    layer2_outputs(3450) <= layer1_outputs(3821);
    layer2_outputs(3451) <= (layer1_outputs(8742)) and not (layer1_outputs(9764));
    layer2_outputs(3452) <= layer1_outputs(7530);
    layer2_outputs(3453) <= not((layer1_outputs(4473)) xor (layer1_outputs(940)));
    layer2_outputs(3454) <= (layer1_outputs(519)) and not (layer1_outputs(1341));
    layer2_outputs(3455) <= (layer1_outputs(5773)) or (layer1_outputs(6206));
    layer2_outputs(3456) <= not(layer1_outputs(2638));
    layer2_outputs(3457) <= layer1_outputs(6995);
    layer2_outputs(3458) <= layer1_outputs(1856);
    layer2_outputs(3459) <= (layer1_outputs(6861)) or (layer1_outputs(1015));
    layer2_outputs(3460) <= not(layer1_outputs(9969));
    layer2_outputs(3461) <= not(layer1_outputs(3270)) or (layer1_outputs(1636));
    layer2_outputs(3462) <= (layer1_outputs(1485)) and (layer1_outputs(9853));
    layer2_outputs(3463) <= layer1_outputs(6540);
    layer2_outputs(3464) <= not(layer1_outputs(8358)) or (layer1_outputs(2418));
    layer2_outputs(3465) <= layer1_outputs(9741);
    layer2_outputs(3466) <= not(layer1_outputs(3266)) or (layer1_outputs(762));
    layer2_outputs(3467) <= not((layer1_outputs(6951)) and (layer1_outputs(2371)));
    layer2_outputs(3468) <= not((layer1_outputs(2252)) xor (layer1_outputs(5646)));
    layer2_outputs(3469) <= layer1_outputs(4413);
    layer2_outputs(3470) <= not(layer1_outputs(6724)) or (layer1_outputs(4723));
    layer2_outputs(3471) <= not(layer1_outputs(5210));
    layer2_outputs(3472) <= not(layer1_outputs(2485));
    layer2_outputs(3473) <= (layer1_outputs(7309)) and not (layer1_outputs(8533));
    layer2_outputs(3474) <= not(layer1_outputs(2584));
    layer2_outputs(3475) <= not(layer1_outputs(2427));
    layer2_outputs(3476) <= layer1_outputs(9354);
    layer2_outputs(3477) <= layer1_outputs(6914);
    layer2_outputs(3478) <= layer1_outputs(4503);
    layer2_outputs(3479) <= not(layer1_outputs(6570));
    layer2_outputs(3480) <= layer1_outputs(1692);
    layer2_outputs(3481) <= (layer1_outputs(538)) and not (layer1_outputs(5657));
    layer2_outputs(3482) <= not(layer1_outputs(5918));
    layer2_outputs(3483) <= not(layer1_outputs(4681));
    layer2_outputs(3484) <= not(layer1_outputs(8286));
    layer2_outputs(3485) <= layer1_outputs(3834);
    layer2_outputs(3486) <= not(layer1_outputs(3109));
    layer2_outputs(3487) <= (layer1_outputs(5730)) and not (layer1_outputs(7376));
    layer2_outputs(3488) <= not(layer1_outputs(433)) or (layer1_outputs(4259));
    layer2_outputs(3489) <= (layer1_outputs(6501)) or (layer1_outputs(3116));
    layer2_outputs(3490) <= layer1_outputs(9696);
    layer2_outputs(3491) <= not(layer1_outputs(4435));
    layer2_outputs(3492) <= (layer1_outputs(6446)) xor (layer1_outputs(2395));
    layer2_outputs(3493) <= layer1_outputs(1282);
    layer2_outputs(3494) <= (layer1_outputs(5951)) and not (layer1_outputs(1088));
    layer2_outputs(3495) <= not(layer1_outputs(3153));
    layer2_outputs(3496) <= layer1_outputs(7030);
    layer2_outputs(3497) <= not((layer1_outputs(524)) and (layer1_outputs(9566)));
    layer2_outputs(3498) <= '0';
    layer2_outputs(3499) <= not(layer1_outputs(6695)) or (layer1_outputs(714));
    layer2_outputs(3500) <= not((layer1_outputs(945)) xor (layer1_outputs(2089)));
    layer2_outputs(3501) <= layer1_outputs(1883);
    layer2_outputs(3502) <= layer1_outputs(298);
    layer2_outputs(3503) <= (layer1_outputs(3848)) and not (layer1_outputs(6373));
    layer2_outputs(3504) <= '1';
    layer2_outputs(3505) <= not((layer1_outputs(5445)) and (layer1_outputs(4395)));
    layer2_outputs(3506) <= layer1_outputs(2778);
    layer2_outputs(3507) <= not(layer1_outputs(5456)) or (layer1_outputs(6084));
    layer2_outputs(3508) <= not((layer1_outputs(8583)) and (layer1_outputs(7380)));
    layer2_outputs(3509) <= not((layer1_outputs(242)) and (layer1_outputs(4074)));
    layer2_outputs(3510) <= layer1_outputs(760);
    layer2_outputs(3511) <= not((layer1_outputs(416)) or (layer1_outputs(2449)));
    layer2_outputs(3512) <= layer1_outputs(1712);
    layer2_outputs(3513) <= not(layer1_outputs(7957));
    layer2_outputs(3514) <= (layer1_outputs(17)) and (layer1_outputs(5731));
    layer2_outputs(3515) <= layer1_outputs(2369);
    layer2_outputs(3516) <= not(layer1_outputs(7712));
    layer2_outputs(3517) <= '1';
    layer2_outputs(3518) <= not(layer1_outputs(3858)) or (layer1_outputs(10026));
    layer2_outputs(3519) <= (layer1_outputs(2185)) and not (layer1_outputs(5708));
    layer2_outputs(3520) <= layer1_outputs(6633);
    layer2_outputs(3521) <= layer1_outputs(1797);
    layer2_outputs(3522) <= (layer1_outputs(10216)) and not (layer1_outputs(8807));
    layer2_outputs(3523) <= not((layer1_outputs(7357)) xor (layer1_outputs(1135)));
    layer2_outputs(3524) <= not((layer1_outputs(9536)) xor (layer1_outputs(5892)));
    layer2_outputs(3525) <= layer1_outputs(4183);
    layer2_outputs(3526) <= layer1_outputs(3760);
    layer2_outputs(3527) <= not(layer1_outputs(9057));
    layer2_outputs(3528) <= layer1_outputs(6764);
    layer2_outputs(3529) <= not(layer1_outputs(3765));
    layer2_outputs(3530) <= not(layer1_outputs(6510)) or (layer1_outputs(6476));
    layer2_outputs(3531) <= not(layer1_outputs(10213));
    layer2_outputs(3532) <= (layer1_outputs(6643)) xor (layer1_outputs(8998));
    layer2_outputs(3533) <= layer1_outputs(8440);
    layer2_outputs(3534) <= not((layer1_outputs(3843)) xor (layer1_outputs(1048)));
    layer2_outputs(3535) <= layer1_outputs(4231);
    layer2_outputs(3536) <= (layer1_outputs(8702)) and (layer1_outputs(9413));
    layer2_outputs(3537) <= not(layer1_outputs(4954));
    layer2_outputs(3538) <= not(layer1_outputs(6396));
    layer2_outputs(3539) <= not(layer1_outputs(4866));
    layer2_outputs(3540) <= layer1_outputs(4753);
    layer2_outputs(3541) <= not(layer1_outputs(4488));
    layer2_outputs(3542) <= (layer1_outputs(9063)) and not (layer1_outputs(7225));
    layer2_outputs(3543) <= not((layer1_outputs(5746)) and (layer1_outputs(4085)));
    layer2_outputs(3544) <= (layer1_outputs(2436)) and not (layer1_outputs(113));
    layer2_outputs(3545) <= (layer1_outputs(3059)) or (layer1_outputs(8754));
    layer2_outputs(3546) <= layer1_outputs(3711);
    layer2_outputs(3547) <= layer1_outputs(5947);
    layer2_outputs(3548) <= not(layer1_outputs(2387)) or (layer1_outputs(5137));
    layer2_outputs(3549) <= not(layer1_outputs(6269));
    layer2_outputs(3550) <= not((layer1_outputs(5466)) and (layer1_outputs(4955)));
    layer2_outputs(3551) <= (layer1_outputs(4402)) or (layer1_outputs(2475));
    layer2_outputs(3552) <= (layer1_outputs(7083)) or (layer1_outputs(8143));
    layer2_outputs(3553) <= not(layer1_outputs(4386));
    layer2_outputs(3554) <= '0';
    layer2_outputs(3555) <= layer1_outputs(3523);
    layer2_outputs(3556) <= (layer1_outputs(3842)) and not (layer1_outputs(4904));
    layer2_outputs(3557) <= (layer1_outputs(4798)) or (layer1_outputs(5396));
    layer2_outputs(3558) <= (layer1_outputs(3094)) xor (layer1_outputs(8075));
    layer2_outputs(3559) <= not((layer1_outputs(7100)) xor (layer1_outputs(5830)));
    layer2_outputs(3560) <= not((layer1_outputs(3604)) and (layer1_outputs(4505)));
    layer2_outputs(3561) <= (layer1_outputs(4153)) and not (layer1_outputs(8865));
    layer2_outputs(3562) <= (layer1_outputs(0)) and not (layer1_outputs(5447));
    layer2_outputs(3563) <= not(layer1_outputs(6214)) or (layer1_outputs(4886));
    layer2_outputs(3564) <= not((layer1_outputs(3941)) or (layer1_outputs(60)));
    layer2_outputs(3565) <= not(layer1_outputs(9428));
    layer2_outputs(3566) <= not(layer1_outputs(1795)) or (layer1_outputs(1606));
    layer2_outputs(3567) <= layer1_outputs(2382);
    layer2_outputs(3568) <= (layer1_outputs(3012)) and not (layer1_outputs(2054));
    layer2_outputs(3569) <= layer1_outputs(4368);
    layer2_outputs(3570) <= not((layer1_outputs(6707)) or (layer1_outputs(5215)));
    layer2_outputs(3571) <= layer1_outputs(5842);
    layer2_outputs(3572) <= '0';
    layer2_outputs(3573) <= not(layer1_outputs(4674));
    layer2_outputs(3574) <= layer1_outputs(7539);
    layer2_outputs(3575) <= (layer1_outputs(6898)) xor (layer1_outputs(9415));
    layer2_outputs(3576) <= not((layer1_outputs(8043)) or (layer1_outputs(2726)));
    layer2_outputs(3577) <= not(layer1_outputs(3733));
    layer2_outputs(3578) <= not(layer1_outputs(5234));
    layer2_outputs(3579) <= not(layer1_outputs(1925)) or (layer1_outputs(2460));
    layer2_outputs(3580) <= layer1_outputs(2028);
    layer2_outputs(3581) <= layer1_outputs(6999);
    layer2_outputs(3582) <= (layer1_outputs(6137)) xor (layer1_outputs(4887));
    layer2_outputs(3583) <= not(layer1_outputs(1176)) or (layer1_outputs(4206));
    layer2_outputs(3584) <= (layer1_outputs(5316)) and (layer1_outputs(6528));
    layer2_outputs(3585) <= not(layer1_outputs(3518));
    layer2_outputs(3586) <= not(layer1_outputs(6168));
    layer2_outputs(3587) <= not(layer1_outputs(574));
    layer2_outputs(3588) <= layer1_outputs(8383);
    layer2_outputs(3589) <= not(layer1_outputs(8100));
    layer2_outputs(3590) <= not(layer1_outputs(6313));
    layer2_outputs(3591) <= (layer1_outputs(8310)) xor (layer1_outputs(5915));
    layer2_outputs(3592) <= (layer1_outputs(5234)) xor (layer1_outputs(10157));
    layer2_outputs(3593) <= not(layer1_outputs(10082));
    layer2_outputs(3594) <= layer1_outputs(6791);
    layer2_outputs(3595) <= not(layer1_outputs(8584));
    layer2_outputs(3596) <= not((layer1_outputs(8241)) or (layer1_outputs(7024)));
    layer2_outputs(3597) <= layer1_outputs(1657);
    layer2_outputs(3598) <= layer1_outputs(1670);
    layer2_outputs(3599) <= (layer1_outputs(3564)) and not (layer1_outputs(4075));
    layer2_outputs(3600) <= layer1_outputs(2682);
    layer2_outputs(3601) <= not((layer1_outputs(5169)) xor (layer1_outputs(7236)));
    layer2_outputs(3602) <= not((layer1_outputs(6209)) and (layer1_outputs(8602)));
    layer2_outputs(3603) <= layer1_outputs(1226);
    layer2_outputs(3604) <= not(layer1_outputs(3189));
    layer2_outputs(3605) <= not(layer1_outputs(1412));
    layer2_outputs(3606) <= layer1_outputs(7776);
    layer2_outputs(3607) <= not(layer1_outputs(3363));
    layer2_outputs(3608) <= not(layer1_outputs(7797));
    layer2_outputs(3609) <= not(layer1_outputs(3561)) or (layer1_outputs(1730));
    layer2_outputs(3610) <= (layer1_outputs(1827)) and (layer1_outputs(2444));
    layer2_outputs(3611) <= layer1_outputs(9146);
    layer2_outputs(3612) <= layer1_outputs(9136);
    layer2_outputs(3613) <= not((layer1_outputs(6531)) and (layer1_outputs(892)));
    layer2_outputs(3614) <= layer1_outputs(228);
    layer2_outputs(3615) <= not(layer1_outputs(7244));
    layer2_outputs(3616) <= layer1_outputs(9256);
    layer2_outputs(3617) <= layer1_outputs(4555);
    layer2_outputs(3618) <= not(layer1_outputs(6086));
    layer2_outputs(3619) <= layer1_outputs(7731);
    layer2_outputs(3620) <= not((layer1_outputs(474)) xor (layer1_outputs(1091)));
    layer2_outputs(3621) <= not(layer1_outputs(1421));
    layer2_outputs(3622) <= (layer1_outputs(190)) xor (layer1_outputs(7560));
    layer2_outputs(3623) <= layer1_outputs(9786);
    layer2_outputs(3624) <= not(layer1_outputs(4551));
    layer2_outputs(3625) <= (layer1_outputs(4698)) and not (layer1_outputs(3882));
    layer2_outputs(3626) <= not((layer1_outputs(3511)) or (layer1_outputs(788)));
    layer2_outputs(3627) <= layer1_outputs(241);
    layer2_outputs(3628) <= layer1_outputs(671);
    layer2_outputs(3629) <= (layer1_outputs(10068)) and (layer1_outputs(9248));
    layer2_outputs(3630) <= layer1_outputs(10204);
    layer2_outputs(3631) <= layer1_outputs(7382);
    layer2_outputs(3632) <= layer1_outputs(5225);
    layer2_outputs(3633) <= not(layer1_outputs(6976));
    layer2_outputs(3634) <= not(layer1_outputs(2858));
    layer2_outputs(3635) <= (layer1_outputs(7999)) or (layer1_outputs(5183));
    layer2_outputs(3636) <= not((layer1_outputs(9938)) xor (layer1_outputs(3791)));
    layer2_outputs(3637) <= (layer1_outputs(3164)) and (layer1_outputs(854));
    layer2_outputs(3638) <= layer1_outputs(3437);
    layer2_outputs(3639) <= layer1_outputs(3200);
    layer2_outputs(3640) <= layer1_outputs(806);
    layer2_outputs(3641) <= layer1_outputs(3182);
    layer2_outputs(3642) <= (layer1_outputs(2494)) xor (layer1_outputs(4485));
    layer2_outputs(3643) <= not(layer1_outputs(5386));
    layer2_outputs(3644) <= not(layer1_outputs(2552));
    layer2_outputs(3645) <= not(layer1_outputs(5423)) or (layer1_outputs(1118));
    layer2_outputs(3646) <= not(layer1_outputs(6016));
    layer2_outputs(3647) <= not((layer1_outputs(7230)) and (layer1_outputs(7900)));
    layer2_outputs(3648) <= layer1_outputs(276);
    layer2_outputs(3649) <= not(layer1_outputs(5097));
    layer2_outputs(3650) <= not(layer1_outputs(9327)) or (layer1_outputs(8368));
    layer2_outputs(3651) <= layer1_outputs(6069);
    layer2_outputs(3652) <= not(layer1_outputs(8083));
    layer2_outputs(3653) <= not(layer1_outputs(193)) or (layer1_outputs(2144));
    layer2_outputs(3654) <= layer1_outputs(4757);
    layer2_outputs(3655) <= not(layer1_outputs(2350));
    layer2_outputs(3656) <= not(layer1_outputs(6789));
    layer2_outputs(3657) <= not(layer1_outputs(6834));
    layer2_outputs(3658) <= layer1_outputs(7485);
    layer2_outputs(3659) <= layer1_outputs(4565);
    layer2_outputs(3660) <= layer1_outputs(9685);
    layer2_outputs(3661) <= layer1_outputs(3915);
    layer2_outputs(3662) <= not(layer1_outputs(8152));
    layer2_outputs(3663) <= layer1_outputs(4247);
    layer2_outputs(3664) <= layer1_outputs(705);
    layer2_outputs(3665) <= (layer1_outputs(9134)) xor (layer1_outputs(7379));
    layer2_outputs(3666) <= layer1_outputs(6842);
    layer2_outputs(3667) <= not(layer1_outputs(7574));
    layer2_outputs(3668) <= (layer1_outputs(391)) xor (layer1_outputs(1571));
    layer2_outputs(3669) <= (layer1_outputs(5468)) and (layer1_outputs(3469));
    layer2_outputs(3670) <= not(layer1_outputs(5961));
    layer2_outputs(3671) <= (layer1_outputs(1289)) and (layer1_outputs(947));
    layer2_outputs(3672) <= (layer1_outputs(2149)) or (layer1_outputs(6732));
    layer2_outputs(3673) <= (layer1_outputs(7802)) or (layer1_outputs(6679));
    layer2_outputs(3674) <= layer1_outputs(30);
    layer2_outputs(3675) <= layer1_outputs(8480);
    layer2_outputs(3676) <= (layer1_outputs(10017)) and not (layer1_outputs(6910));
    layer2_outputs(3677) <= layer1_outputs(3078);
    layer2_outputs(3678) <= not(layer1_outputs(3139));
    layer2_outputs(3679) <= (layer1_outputs(10099)) and not (layer1_outputs(2421));
    layer2_outputs(3680) <= layer1_outputs(2478);
    layer2_outputs(3681) <= not(layer1_outputs(4351)) or (layer1_outputs(8075));
    layer2_outputs(3682) <= not(layer1_outputs(7492));
    layer2_outputs(3683) <= layer1_outputs(5541);
    layer2_outputs(3684) <= layer1_outputs(7311);
    layer2_outputs(3685) <= not(layer1_outputs(10129));
    layer2_outputs(3686) <= not((layer1_outputs(3329)) xor (layer1_outputs(9826)));
    layer2_outputs(3687) <= not(layer1_outputs(7062));
    layer2_outputs(3688) <= not(layer1_outputs(6670));
    layer2_outputs(3689) <= (layer1_outputs(8064)) xor (layer1_outputs(2577));
    layer2_outputs(3690) <= layer1_outputs(5073);
    layer2_outputs(3691) <= not((layer1_outputs(5500)) and (layer1_outputs(7523)));
    layer2_outputs(3692) <= not((layer1_outputs(7492)) or (layer1_outputs(7081)));
    layer2_outputs(3693) <= not(layer1_outputs(9915));
    layer2_outputs(3694) <= not((layer1_outputs(8297)) or (layer1_outputs(9892)));
    layer2_outputs(3695) <= layer1_outputs(9388);
    layer2_outputs(3696) <= layer1_outputs(6320);
    layer2_outputs(3697) <= (layer1_outputs(7527)) and not (layer1_outputs(5523));
    layer2_outputs(3698) <= layer1_outputs(9949);
    layer2_outputs(3699) <= (layer1_outputs(2271)) xor (layer1_outputs(4994));
    layer2_outputs(3700) <= not(layer1_outputs(3364)) or (layer1_outputs(5455));
    layer2_outputs(3701) <= not(layer1_outputs(9710));
    layer2_outputs(3702) <= (layer1_outputs(3711)) xor (layer1_outputs(2287));
    layer2_outputs(3703) <= not((layer1_outputs(9314)) or (layer1_outputs(3653)));
    layer2_outputs(3704) <= not(layer1_outputs(9864)) or (layer1_outputs(5420));
    layer2_outputs(3705) <= (layer1_outputs(1963)) or (layer1_outputs(7642));
    layer2_outputs(3706) <= layer1_outputs(6719);
    layer2_outputs(3707) <= not((layer1_outputs(6722)) and (layer1_outputs(6266)));
    layer2_outputs(3708) <= (layer1_outputs(8363)) xor (layer1_outputs(2531));
    layer2_outputs(3709) <= not(layer1_outputs(6994));
    layer2_outputs(3710) <= layer1_outputs(929);
    layer2_outputs(3711) <= layer1_outputs(4507);
    layer2_outputs(3712) <= layer1_outputs(1379);
    layer2_outputs(3713) <= not(layer1_outputs(600)) or (layer1_outputs(5941));
    layer2_outputs(3714) <= layer1_outputs(421);
    layer2_outputs(3715) <= (layer1_outputs(9704)) and (layer1_outputs(5619));
    layer2_outputs(3716) <= not(layer1_outputs(9111)) or (layer1_outputs(7079));
    layer2_outputs(3717) <= layer1_outputs(4469);
    layer2_outputs(3718) <= layer1_outputs(384);
    layer2_outputs(3719) <= not(layer1_outputs(9281));
    layer2_outputs(3720) <= not(layer1_outputs(9916));
    layer2_outputs(3721) <= not(layer1_outputs(4342));
    layer2_outputs(3722) <= (layer1_outputs(4817)) and not (layer1_outputs(1302));
    layer2_outputs(3723) <= layer1_outputs(3456);
    layer2_outputs(3724) <= not(layer1_outputs(7875));
    layer2_outputs(3725) <= layer1_outputs(7448);
    layer2_outputs(3726) <= (layer1_outputs(1447)) xor (layer1_outputs(3280));
    layer2_outputs(3727) <= (layer1_outputs(6080)) and not (layer1_outputs(6714));
    layer2_outputs(3728) <= not(layer1_outputs(8738));
    layer2_outputs(3729) <= not((layer1_outputs(2002)) xor (layer1_outputs(849)));
    layer2_outputs(3730) <= (layer1_outputs(7988)) or (layer1_outputs(3780));
    layer2_outputs(3731) <= not(layer1_outputs(9818));
    layer2_outputs(3732) <= layer1_outputs(5098);
    layer2_outputs(3733) <= (layer1_outputs(6216)) and not (layer1_outputs(5353));
    layer2_outputs(3734) <= (layer1_outputs(7037)) xor (layer1_outputs(7266));
    layer2_outputs(3735) <= not(layer1_outputs(1007));
    layer2_outputs(3736) <= not(layer1_outputs(9398)) or (layer1_outputs(2616));
    layer2_outputs(3737) <= not(layer1_outputs(3053));
    layer2_outputs(3738) <= layer1_outputs(3112);
    layer2_outputs(3739) <= (layer1_outputs(3684)) xor (layer1_outputs(6222));
    layer2_outputs(3740) <= layer1_outputs(5986);
    layer2_outputs(3741) <= (layer1_outputs(9841)) and (layer1_outputs(521));
    layer2_outputs(3742) <= not(layer1_outputs(8625));
    layer2_outputs(3743) <= (layer1_outputs(2707)) and not (layer1_outputs(2998));
    layer2_outputs(3744) <= not(layer1_outputs(8459));
    layer2_outputs(3745) <= (layer1_outputs(4391)) or (layer1_outputs(4917));
    layer2_outputs(3746) <= not((layer1_outputs(6272)) or (layer1_outputs(9088)));
    layer2_outputs(3747) <= not((layer1_outputs(2939)) xor (layer1_outputs(5490)));
    layer2_outputs(3748) <= not(layer1_outputs(9226));
    layer2_outputs(3749) <= not((layer1_outputs(6363)) and (layer1_outputs(10038)));
    layer2_outputs(3750) <= not(layer1_outputs(7800));
    layer2_outputs(3751) <= layer1_outputs(3924);
    layer2_outputs(3752) <= not(layer1_outputs(6955));
    layer2_outputs(3753) <= not(layer1_outputs(1593));
    layer2_outputs(3754) <= (layer1_outputs(5506)) or (layer1_outputs(7410));
    layer2_outputs(3755) <= not(layer1_outputs(1990));
    layer2_outputs(3756) <= not(layer1_outputs(2361));
    layer2_outputs(3757) <= not(layer1_outputs(2535));
    layer2_outputs(3758) <= not(layer1_outputs(9010));
    layer2_outputs(3759) <= (layer1_outputs(6932)) xor (layer1_outputs(8814));
    layer2_outputs(3760) <= layer1_outputs(1867);
    layer2_outputs(3761) <= (layer1_outputs(1112)) xor (layer1_outputs(2670));
    layer2_outputs(3762) <= not((layer1_outputs(2728)) and (layer1_outputs(1782)));
    layer2_outputs(3763) <= layer1_outputs(8072);
    layer2_outputs(3764) <= layer1_outputs(922);
    layer2_outputs(3765) <= layer1_outputs(9654);
    layer2_outputs(3766) <= not(layer1_outputs(2256)) or (layer1_outputs(4326));
    layer2_outputs(3767) <= not(layer1_outputs(205));
    layer2_outputs(3768) <= not((layer1_outputs(9337)) and (layer1_outputs(2128)));
    layer2_outputs(3769) <= (layer1_outputs(4374)) and not (layer1_outputs(4142));
    layer2_outputs(3770) <= not(layer1_outputs(1815));
    layer2_outputs(3771) <= not(layer1_outputs(6101));
    layer2_outputs(3772) <= not(layer1_outputs(7893));
    layer2_outputs(3773) <= (layer1_outputs(4576)) and (layer1_outputs(1130));
    layer2_outputs(3774) <= (layer1_outputs(3626)) and (layer1_outputs(3632));
    layer2_outputs(3775) <= (layer1_outputs(10081)) and not (layer1_outputs(761));
    layer2_outputs(3776) <= not(layer1_outputs(5271));
    layer2_outputs(3777) <= layer1_outputs(5816);
    layer2_outputs(3778) <= not(layer1_outputs(160));
    layer2_outputs(3779) <= (layer1_outputs(7888)) and not (layer1_outputs(9502));
    layer2_outputs(3780) <= not(layer1_outputs(5248));
    layer2_outputs(3781) <= not(layer1_outputs(2918));
    layer2_outputs(3782) <= layer1_outputs(3658);
    layer2_outputs(3783) <= not((layer1_outputs(6547)) xor (layer1_outputs(3809)));
    layer2_outputs(3784) <= '1';
    layer2_outputs(3785) <= layer1_outputs(1287);
    layer2_outputs(3786) <= (layer1_outputs(3010)) xor (layer1_outputs(4994));
    layer2_outputs(3787) <= (layer1_outputs(131)) xor (layer1_outputs(7709));
    layer2_outputs(3788) <= not(layer1_outputs(1843));
    layer2_outputs(3789) <= layer1_outputs(3839);
    layer2_outputs(3790) <= (layer1_outputs(2295)) xor (layer1_outputs(8741));
    layer2_outputs(3791) <= layer1_outputs(7411);
    layer2_outputs(3792) <= (layer1_outputs(5374)) and not (layer1_outputs(1252));
    layer2_outputs(3793) <= (layer1_outputs(2597)) and (layer1_outputs(1584));
    layer2_outputs(3794) <= (layer1_outputs(1170)) and not (layer1_outputs(1169));
    layer2_outputs(3795) <= not(layer1_outputs(5508)) or (layer1_outputs(3176));
    layer2_outputs(3796) <= not((layer1_outputs(2989)) or (layer1_outputs(850)));
    layer2_outputs(3797) <= (layer1_outputs(1838)) and not (layer1_outputs(8566));
    layer2_outputs(3798) <= not(layer1_outputs(7888));
    layer2_outputs(3799) <= layer1_outputs(4922);
    layer2_outputs(3800) <= not(layer1_outputs(152));
    layer2_outputs(3801) <= layer1_outputs(10030);
    layer2_outputs(3802) <= not(layer1_outputs(385)) or (layer1_outputs(5913));
    layer2_outputs(3803) <= (layer1_outputs(3201)) and not (layer1_outputs(7899));
    layer2_outputs(3804) <= not((layer1_outputs(4024)) and (layer1_outputs(8089)));
    layer2_outputs(3805) <= (layer1_outputs(2274)) xor (layer1_outputs(6842));
    layer2_outputs(3806) <= (layer1_outputs(3195)) xor (layer1_outputs(150));
    layer2_outputs(3807) <= not((layer1_outputs(6781)) xor (layer1_outputs(7139)));
    layer2_outputs(3808) <= layer1_outputs(2071);
    layer2_outputs(3809) <= (layer1_outputs(1686)) xor (layer1_outputs(5401));
    layer2_outputs(3810) <= layer1_outputs(10188);
    layer2_outputs(3811) <= not(layer1_outputs(186));
    layer2_outputs(3812) <= (layer1_outputs(8712)) and not (layer1_outputs(3530));
    layer2_outputs(3813) <= not(layer1_outputs(4855));
    layer2_outputs(3814) <= (layer1_outputs(8853)) xor (layer1_outputs(3660));
    layer2_outputs(3815) <= not((layer1_outputs(3189)) and (layer1_outputs(7619)));
    layer2_outputs(3816) <= (layer1_outputs(9908)) and not (layer1_outputs(6191));
    layer2_outputs(3817) <= layer1_outputs(1215);
    layer2_outputs(3818) <= layer1_outputs(8311);
    layer2_outputs(3819) <= (layer1_outputs(8845)) and not (layer1_outputs(7601));
    layer2_outputs(3820) <= not(layer1_outputs(9173));
    layer2_outputs(3821) <= layer1_outputs(1684);
    layer2_outputs(3822) <= not(layer1_outputs(64));
    layer2_outputs(3823) <= not((layer1_outputs(3465)) xor (layer1_outputs(2592)));
    layer2_outputs(3824) <= (layer1_outputs(5479)) xor (layer1_outputs(8089));
    layer2_outputs(3825) <= not((layer1_outputs(4773)) and (layer1_outputs(7834)));
    layer2_outputs(3826) <= not(layer1_outputs(3742));
    layer2_outputs(3827) <= (layer1_outputs(9244)) or (layer1_outputs(9689));
    layer2_outputs(3828) <= layer1_outputs(6301);
    layer2_outputs(3829) <= (layer1_outputs(480)) and (layer1_outputs(10097));
    layer2_outputs(3830) <= (layer1_outputs(3979)) and not (layer1_outputs(2000));
    layer2_outputs(3831) <= layer1_outputs(1059);
    layer2_outputs(3832) <= layer1_outputs(617);
    layer2_outputs(3833) <= layer1_outputs(2577);
    layer2_outputs(3834) <= layer1_outputs(2005);
    layer2_outputs(3835) <= not((layer1_outputs(9704)) and (layer1_outputs(2665)));
    layer2_outputs(3836) <= not(layer1_outputs(5798));
    layer2_outputs(3837) <= not((layer1_outputs(3571)) or (layer1_outputs(5934)));
    layer2_outputs(3838) <= not(layer1_outputs(2730));
    layer2_outputs(3839) <= not(layer1_outputs(314));
    layer2_outputs(3840) <= not((layer1_outputs(6801)) or (layer1_outputs(1255)));
    layer2_outputs(3841) <= not(layer1_outputs(7158));
    layer2_outputs(3842) <= not(layer1_outputs(6555));
    layer2_outputs(3843) <= not(layer1_outputs(8998));
    layer2_outputs(3844) <= not(layer1_outputs(324));
    layer2_outputs(3845) <= not(layer1_outputs(4064)) or (layer1_outputs(7645));
    layer2_outputs(3846) <= not((layer1_outputs(4377)) or (layer1_outputs(1552)));
    layer2_outputs(3847) <= (layer1_outputs(9209)) xor (layer1_outputs(2367));
    layer2_outputs(3848) <= not((layer1_outputs(8184)) xor (layer1_outputs(4679)));
    layer2_outputs(3849) <= not(layer1_outputs(9152)) or (layer1_outputs(7522));
    layer2_outputs(3850) <= layer1_outputs(6785);
    layer2_outputs(3851) <= layer1_outputs(2655);
    layer2_outputs(3852) <= not(layer1_outputs(2311)) or (layer1_outputs(9950));
    layer2_outputs(3853) <= (layer1_outputs(5988)) and (layer1_outputs(7062));
    layer2_outputs(3854) <= not(layer1_outputs(3221));
    layer2_outputs(3855) <= not(layer1_outputs(8580)) or (layer1_outputs(8630));
    layer2_outputs(3856) <= (layer1_outputs(4923)) and not (layer1_outputs(8662));
    layer2_outputs(3857) <= (layer1_outputs(3376)) and not (layer1_outputs(6048));
    layer2_outputs(3858) <= layer1_outputs(4187);
    layer2_outputs(3859) <= not(layer1_outputs(2949));
    layer2_outputs(3860) <= (layer1_outputs(1778)) xor (layer1_outputs(3740));
    layer2_outputs(3861) <= layer1_outputs(9092);
    layer2_outputs(3862) <= layer1_outputs(2602);
    layer2_outputs(3863) <= not(layer1_outputs(2868));
    layer2_outputs(3864) <= not(layer1_outputs(5373));
    layer2_outputs(3865) <= (layer1_outputs(8687)) and not (layer1_outputs(9449));
    layer2_outputs(3866) <= not((layer1_outputs(5253)) xor (layer1_outputs(43)));
    layer2_outputs(3867) <= layer1_outputs(3290);
    layer2_outputs(3868) <= layer1_outputs(2156);
    layer2_outputs(3869) <= (layer1_outputs(2366)) xor (layer1_outputs(9474));
    layer2_outputs(3870) <= not(layer1_outputs(5605));
    layer2_outputs(3871) <= (layer1_outputs(5235)) and not (layer1_outputs(1088));
    layer2_outputs(3872) <= (layer1_outputs(6869)) or (layer1_outputs(3874));
    layer2_outputs(3873) <= not(layer1_outputs(434)) or (layer1_outputs(9279));
    layer2_outputs(3874) <= (layer1_outputs(4378)) and not (layer1_outputs(6992));
    layer2_outputs(3875) <= layer1_outputs(5131);
    layer2_outputs(3876) <= layer1_outputs(560);
    layer2_outputs(3877) <= layer1_outputs(5743);
    layer2_outputs(3878) <= (layer1_outputs(517)) or (layer1_outputs(4155));
    layer2_outputs(3879) <= not(layer1_outputs(194));
    layer2_outputs(3880) <= not(layer1_outputs(10087));
    layer2_outputs(3881) <= layer1_outputs(10190);
    layer2_outputs(3882) <= not(layer1_outputs(7515));
    layer2_outputs(3883) <= not((layer1_outputs(7918)) or (layer1_outputs(2515)));
    layer2_outputs(3884) <= (layer1_outputs(890)) and not (layer1_outputs(1476));
    layer2_outputs(3885) <= not(layer1_outputs(1108)) or (layer1_outputs(5902));
    layer2_outputs(3886) <= (layer1_outputs(3119)) and not (layer1_outputs(7561));
    layer2_outputs(3887) <= (layer1_outputs(2469)) and (layer1_outputs(9816));
    layer2_outputs(3888) <= not((layer1_outputs(8297)) or (layer1_outputs(6693)));
    layer2_outputs(3889) <= layer1_outputs(439);
    layer2_outputs(3890) <= not(layer1_outputs(718));
    layer2_outputs(3891) <= not(layer1_outputs(1093));
    layer2_outputs(3892) <= not(layer1_outputs(1656));
    layer2_outputs(3893) <= not((layer1_outputs(5442)) or (layer1_outputs(3088)));
    layer2_outputs(3894) <= not(layer1_outputs(5946)) or (layer1_outputs(9324));
    layer2_outputs(3895) <= layer1_outputs(7367);
    layer2_outputs(3896) <= (layer1_outputs(1419)) and (layer1_outputs(8841));
    layer2_outputs(3897) <= not(layer1_outputs(5338)) or (layer1_outputs(7049));
    layer2_outputs(3898) <= not(layer1_outputs(5090)) or (layer1_outputs(7031));
    layer2_outputs(3899) <= layer1_outputs(5486);
    layer2_outputs(3900) <= not(layer1_outputs(5226)) or (layer1_outputs(9943));
    layer2_outputs(3901) <= not(layer1_outputs(2337));
    layer2_outputs(3902) <= not(layer1_outputs(8216));
    layer2_outputs(3903) <= (layer1_outputs(866)) and not (layer1_outputs(9959));
    layer2_outputs(3904) <= not(layer1_outputs(6999));
    layer2_outputs(3905) <= layer1_outputs(5702);
    layer2_outputs(3906) <= (layer1_outputs(8796)) and (layer1_outputs(2821));
    layer2_outputs(3907) <= layer1_outputs(7510);
    layer2_outputs(3908) <= (layer1_outputs(4385)) or (layer1_outputs(7002));
    layer2_outputs(3909) <= '0';
    layer2_outputs(3910) <= layer1_outputs(1148);
    layer2_outputs(3911) <= not(layer1_outputs(6170));
    layer2_outputs(3912) <= (layer1_outputs(7584)) and not (layer1_outputs(8433));
    layer2_outputs(3913) <= layer1_outputs(7890);
    layer2_outputs(3914) <= not((layer1_outputs(2663)) and (layer1_outputs(317)));
    layer2_outputs(3915) <= layer1_outputs(3184);
    layer2_outputs(3916) <= not((layer1_outputs(4646)) and (layer1_outputs(1307)));
    layer2_outputs(3917) <= not(layer1_outputs(7258)) or (layer1_outputs(1337));
    layer2_outputs(3918) <= layer1_outputs(791);
    layer2_outputs(3919) <= layer1_outputs(9936);
    layer2_outputs(3920) <= layer1_outputs(1223);
    layer2_outputs(3921) <= not(layer1_outputs(8568));
    layer2_outputs(3922) <= '1';
    layer2_outputs(3923) <= layer1_outputs(2676);
    layer2_outputs(3924) <= layer1_outputs(2700);
    layer2_outputs(3925) <= not((layer1_outputs(8964)) and (layer1_outputs(167)));
    layer2_outputs(3926) <= not(layer1_outputs(7028)) or (layer1_outputs(4408));
    layer2_outputs(3927) <= not(layer1_outputs(6669));
    layer2_outputs(3928) <= (layer1_outputs(7836)) and not (layer1_outputs(4245));
    layer2_outputs(3929) <= (layer1_outputs(41)) and not (layer1_outputs(7685));
    layer2_outputs(3930) <= not(layer1_outputs(2389));
    layer2_outputs(3931) <= not(layer1_outputs(6488));
    layer2_outputs(3932) <= (layer1_outputs(785)) and (layer1_outputs(5063));
    layer2_outputs(3933) <= layer1_outputs(3185);
    layer2_outputs(3934) <= layer1_outputs(2288);
    layer2_outputs(3935) <= (layer1_outputs(5538)) or (layer1_outputs(7785));
    layer2_outputs(3936) <= (layer1_outputs(625)) and not (layer1_outputs(1930));
    layer2_outputs(3937) <= not(layer1_outputs(3695)) or (layer1_outputs(1086));
    layer2_outputs(3938) <= not(layer1_outputs(9996));
    layer2_outputs(3939) <= layer1_outputs(3311);
    layer2_outputs(3940) <= layer1_outputs(3424);
    layer2_outputs(3941) <= not(layer1_outputs(6617));
    layer2_outputs(3942) <= not(layer1_outputs(1804));
    layer2_outputs(3943) <= not(layer1_outputs(9648));
    layer2_outputs(3944) <= not((layer1_outputs(9612)) xor (layer1_outputs(5244)));
    layer2_outputs(3945) <= (layer1_outputs(8806)) xor (layer1_outputs(2227));
    layer2_outputs(3946) <= not((layer1_outputs(2426)) and (layer1_outputs(3380)));
    layer2_outputs(3947) <= layer1_outputs(8301);
    layer2_outputs(3948) <= (layer1_outputs(1340)) xor (layer1_outputs(7835));
    layer2_outputs(3949) <= not(layer1_outputs(8749));
    layer2_outputs(3950) <= not(layer1_outputs(4165));
    layer2_outputs(3951) <= not(layer1_outputs(3148));
    layer2_outputs(3952) <= layer1_outputs(7938);
    layer2_outputs(3953) <= not((layer1_outputs(2660)) or (layer1_outputs(7915)));
    layer2_outputs(3954) <= not(layer1_outputs(616));
    layer2_outputs(3955) <= not(layer1_outputs(9062));
    layer2_outputs(3956) <= (layer1_outputs(4728)) and not (layer1_outputs(10045));
    layer2_outputs(3957) <= not(layer1_outputs(6295)) or (layer1_outputs(3852));
    layer2_outputs(3958) <= not((layer1_outputs(2560)) and (layer1_outputs(6911)));
    layer2_outputs(3959) <= layer1_outputs(9888);
    layer2_outputs(3960) <= not(layer1_outputs(360)) or (layer1_outputs(1835));
    layer2_outputs(3961) <= not((layer1_outputs(4780)) and (layer1_outputs(6227)));
    layer2_outputs(3962) <= not((layer1_outputs(5114)) xor (layer1_outputs(6841)));
    layer2_outputs(3963) <= layer1_outputs(2413);
    layer2_outputs(3964) <= not(layer1_outputs(2842));
    layer2_outputs(3965) <= layer1_outputs(7332);
    layer2_outputs(3966) <= '0';
    layer2_outputs(3967) <= not(layer1_outputs(9072));
    layer2_outputs(3968) <= not(layer1_outputs(6033));
    layer2_outputs(3969) <= layer1_outputs(5292);
    layer2_outputs(3970) <= not(layer1_outputs(3768)) or (layer1_outputs(412));
    layer2_outputs(3971) <= not(layer1_outputs(9550));
    layer2_outputs(3972) <= not(layer1_outputs(7669));
    layer2_outputs(3973) <= (layer1_outputs(6551)) and not (layer1_outputs(5829));
    layer2_outputs(3974) <= not(layer1_outputs(5631));
    layer2_outputs(3975) <= not(layer1_outputs(525));
    layer2_outputs(3976) <= layer1_outputs(9161);
    layer2_outputs(3977) <= not(layer1_outputs(2960));
    layer2_outputs(3978) <= not(layer1_outputs(3655));
    layer2_outputs(3979) <= (layer1_outputs(976)) xor (layer1_outputs(8412));
    layer2_outputs(3980) <= layer1_outputs(2180);
    layer2_outputs(3981) <= not(layer1_outputs(10123));
    layer2_outputs(3982) <= layer1_outputs(8890);
    layer2_outputs(3983) <= layer1_outputs(9763);
    layer2_outputs(3984) <= not((layer1_outputs(7464)) and (layer1_outputs(5715)));
    layer2_outputs(3985) <= not(layer1_outputs(6424));
    layer2_outputs(3986) <= not(layer1_outputs(6536));
    layer2_outputs(3987) <= layer1_outputs(4497);
    layer2_outputs(3988) <= not(layer1_outputs(10027));
    layer2_outputs(3989) <= not((layer1_outputs(2749)) or (layer1_outputs(2483)));
    layer2_outputs(3990) <= not(layer1_outputs(4810)) or (layer1_outputs(1041));
    layer2_outputs(3991) <= (layer1_outputs(7341)) and not (layer1_outputs(54));
    layer2_outputs(3992) <= layer1_outputs(1124);
    layer2_outputs(3993) <= not((layer1_outputs(1395)) and (layer1_outputs(3501)));
    layer2_outputs(3994) <= not((layer1_outputs(2951)) and (layer1_outputs(3730)));
    layer2_outputs(3995) <= not((layer1_outputs(2783)) or (layer1_outputs(5686)));
    layer2_outputs(3996) <= not((layer1_outputs(9343)) xor (layer1_outputs(1975)));
    layer2_outputs(3997) <= (layer1_outputs(4464)) or (layer1_outputs(2051));
    layer2_outputs(3998) <= not(layer1_outputs(2954));
    layer2_outputs(3999) <= layer1_outputs(6969);
    layer2_outputs(4000) <= layer1_outputs(656);
    layer2_outputs(4001) <= not(layer1_outputs(5414));
    layer2_outputs(4002) <= not(layer1_outputs(10008));
    layer2_outputs(4003) <= (layer1_outputs(9707)) xor (layer1_outputs(1044));
    layer2_outputs(4004) <= not(layer1_outputs(7678));
    layer2_outputs(4005) <= (layer1_outputs(2263)) xor (layer1_outputs(68));
    layer2_outputs(4006) <= not(layer1_outputs(3736));
    layer2_outputs(4007) <= layer1_outputs(5498);
    layer2_outputs(4008) <= (layer1_outputs(10075)) xor (layer1_outputs(89));
    layer2_outputs(4009) <= not((layer1_outputs(1218)) or (layer1_outputs(4433)));
    layer2_outputs(4010) <= not(layer1_outputs(8270)) or (layer1_outputs(134));
    layer2_outputs(4011) <= not(layer1_outputs(5064)) or (layer1_outputs(9110));
    layer2_outputs(4012) <= not(layer1_outputs(1462));
    layer2_outputs(4013) <= not(layer1_outputs(8197));
    layer2_outputs(4014) <= not((layer1_outputs(3801)) and (layer1_outputs(1763)));
    layer2_outputs(4015) <= not(layer1_outputs(8060));
    layer2_outputs(4016) <= not((layer1_outputs(461)) xor (layer1_outputs(3163)));
    layer2_outputs(4017) <= not(layer1_outputs(930));
    layer2_outputs(4018) <= not(layer1_outputs(1147));
    layer2_outputs(4019) <= layer1_outputs(2271);
    layer2_outputs(4020) <= not(layer1_outputs(9040));
    layer2_outputs(4021) <= (layer1_outputs(5737)) and not (layer1_outputs(4491));
    layer2_outputs(4022) <= '1';
    layer2_outputs(4023) <= layer1_outputs(1059);
    layer2_outputs(4024) <= not((layer1_outputs(599)) and (layer1_outputs(7804)));
    layer2_outputs(4025) <= layer1_outputs(1425);
    layer2_outputs(4026) <= not(layer1_outputs(3944));
    layer2_outputs(4027) <= not((layer1_outputs(6021)) xor (layer1_outputs(8005)));
    layer2_outputs(4028) <= (layer1_outputs(6204)) xor (layer1_outputs(1786));
    layer2_outputs(4029) <= not(layer1_outputs(9103));
    layer2_outputs(4030) <= (layer1_outputs(6821)) xor (layer1_outputs(8016));
    layer2_outputs(4031) <= layer1_outputs(5375);
    layer2_outputs(4032) <= not(layer1_outputs(6282)) or (layer1_outputs(9754));
    layer2_outputs(4033) <= (layer1_outputs(5875)) or (layer1_outputs(653));
    layer2_outputs(4034) <= (layer1_outputs(8767)) and (layer1_outputs(645));
    layer2_outputs(4035) <= (layer1_outputs(6625)) and (layer1_outputs(2290));
    layer2_outputs(4036) <= layer1_outputs(3125);
    layer2_outputs(4037) <= layer1_outputs(6322);
    layer2_outputs(4038) <= layer1_outputs(1912);
    layer2_outputs(4039) <= (layer1_outputs(1954)) or (layer1_outputs(8667));
    layer2_outputs(4040) <= not((layer1_outputs(6202)) or (layer1_outputs(1554)));
    layer2_outputs(4041) <= (layer1_outputs(1406)) xor (layer1_outputs(2995));
    layer2_outputs(4042) <= (layer1_outputs(7071)) and not (layer1_outputs(8881));
    layer2_outputs(4043) <= not(layer1_outputs(5660));
    layer2_outputs(4044) <= not(layer1_outputs(2657)) or (layer1_outputs(4770));
    layer2_outputs(4045) <= not(layer1_outputs(6299));
    layer2_outputs(4046) <= not((layer1_outputs(5406)) or (layer1_outputs(793)));
    layer2_outputs(4047) <= layer1_outputs(5362);
    layer2_outputs(4048) <= not((layer1_outputs(5170)) xor (layer1_outputs(1924)));
    layer2_outputs(4049) <= not(layer1_outputs(6565));
    layer2_outputs(4050) <= not((layer1_outputs(7566)) and (layer1_outputs(3644)));
    layer2_outputs(4051) <= layer1_outputs(2055);
    layer2_outputs(4052) <= layer1_outputs(9197);
    layer2_outputs(4053) <= not((layer1_outputs(4986)) and (layer1_outputs(9836)));
    layer2_outputs(4054) <= not((layer1_outputs(541)) or (layer1_outputs(4471)));
    layer2_outputs(4055) <= (layer1_outputs(634)) and not (layer1_outputs(5174));
    layer2_outputs(4056) <= not(layer1_outputs(2416));
    layer2_outputs(4057) <= not(layer1_outputs(8539));
    layer2_outputs(4058) <= layer1_outputs(7436);
    layer2_outputs(4059) <= (layer1_outputs(7375)) or (layer1_outputs(2808));
    layer2_outputs(4060) <= layer1_outputs(5534);
    layer2_outputs(4061) <= layer1_outputs(539);
    layer2_outputs(4062) <= not(layer1_outputs(2386));
    layer2_outputs(4063) <= not(layer1_outputs(3123));
    layer2_outputs(4064) <= layer1_outputs(4468);
    layer2_outputs(4065) <= not((layer1_outputs(7781)) xor (layer1_outputs(3873)));
    layer2_outputs(4066) <= not(layer1_outputs(5638));
    layer2_outputs(4067) <= layer1_outputs(5237);
    layer2_outputs(4068) <= not(layer1_outputs(1640));
    layer2_outputs(4069) <= not(layer1_outputs(546));
    layer2_outputs(4070) <= (layer1_outputs(1438)) and not (layer1_outputs(2060));
    layer2_outputs(4071) <= (layer1_outputs(649)) and (layer1_outputs(5177));
    layer2_outputs(4072) <= not(layer1_outputs(6520));
    layer2_outputs(4073) <= layer1_outputs(3294);
    layer2_outputs(4074) <= layer1_outputs(3925);
    layer2_outputs(4075) <= not(layer1_outputs(6580));
    layer2_outputs(4076) <= layer1_outputs(5542);
    layer2_outputs(4077) <= (layer1_outputs(6070)) and not (layer1_outputs(2162));
    layer2_outputs(4078) <= (layer1_outputs(8983)) and (layer1_outputs(8029));
    layer2_outputs(4079) <= layer1_outputs(9815);
    layer2_outputs(4080) <= (layer1_outputs(3014)) and (layer1_outputs(2311));
    layer2_outputs(4081) <= not(layer1_outputs(6620));
    layer2_outputs(4082) <= layer1_outputs(4695);
    layer2_outputs(4083) <= not(layer1_outputs(4909));
    layer2_outputs(4084) <= not(layer1_outputs(6599));
    layer2_outputs(4085) <= not((layer1_outputs(81)) xor (layer1_outputs(6075)));
    layer2_outputs(4086) <= layer1_outputs(692);
    layer2_outputs(4087) <= not(layer1_outputs(10112)) or (layer1_outputs(4845));
    layer2_outputs(4088) <= not((layer1_outputs(483)) or (layer1_outputs(10233)));
    layer2_outputs(4089) <= not(layer1_outputs(6209));
    layer2_outputs(4090) <= (layer1_outputs(1768)) and not (layer1_outputs(8367));
    layer2_outputs(4091) <= layer1_outputs(2330);
    layer2_outputs(4092) <= not(layer1_outputs(2018));
    layer2_outputs(4093) <= (layer1_outputs(4912)) and not (layer1_outputs(833));
    layer2_outputs(4094) <= not(layer1_outputs(10193));
    layer2_outputs(4095) <= not(layer1_outputs(2593));
    layer2_outputs(4096) <= (layer1_outputs(8836)) xor (layer1_outputs(7253));
    layer2_outputs(4097) <= not((layer1_outputs(7002)) xor (layer1_outputs(333)));
    layer2_outputs(4098) <= not(layer1_outputs(2312));
    layer2_outputs(4099) <= layer1_outputs(5376);
    layer2_outputs(4100) <= layer1_outputs(6649);
    layer2_outputs(4101) <= layer1_outputs(3623);
    layer2_outputs(4102) <= not((layer1_outputs(8365)) or (layer1_outputs(9902)));
    layer2_outputs(4103) <= layer1_outputs(7896);
    layer2_outputs(4104) <= not(layer1_outputs(1324)) or (layer1_outputs(9232));
    layer2_outputs(4105) <= (layer1_outputs(8887)) and not (layer1_outputs(3689));
    layer2_outputs(4106) <= (layer1_outputs(2802)) and not (layer1_outputs(3412));
    layer2_outputs(4107) <= not(layer1_outputs(635));
    layer2_outputs(4108) <= (layer1_outputs(3865)) and (layer1_outputs(9235));
    layer2_outputs(4109) <= layer1_outputs(1725);
    layer2_outputs(4110) <= layer1_outputs(9869);
    layer2_outputs(4111) <= not(layer1_outputs(609)) or (layer1_outputs(5223));
    layer2_outputs(4112) <= not(layer1_outputs(1131)) or (layer1_outputs(7061));
    layer2_outputs(4113) <= '0';
    layer2_outputs(4114) <= layer1_outputs(2593);
    layer2_outputs(4115) <= not(layer1_outputs(8584));
    layer2_outputs(4116) <= layer1_outputs(1077);
    layer2_outputs(4117) <= not(layer1_outputs(955));
    layer2_outputs(4118) <= (layer1_outputs(2394)) xor (layer1_outputs(819));
    layer2_outputs(4119) <= not(layer1_outputs(2721)) or (layer1_outputs(7349));
    layer2_outputs(4120) <= layer1_outputs(5371);
    layer2_outputs(4121) <= layer1_outputs(7561);
    layer2_outputs(4122) <= not(layer1_outputs(9684)) or (layer1_outputs(4821));
    layer2_outputs(4123) <= not((layer1_outputs(2853)) or (layer1_outputs(9076)));
    layer2_outputs(4124) <= not(layer1_outputs(5563)) or (layer1_outputs(5596));
    layer2_outputs(4125) <= (layer1_outputs(6406)) or (layer1_outputs(1858));
    layer2_outputs(4126) <= (layer1_outputs(616)) xor (layer1_outputs(3240));
    layer2_outputs(4127) <= (layer1_outputs(783)) and not (layer1_outputs(9561));
    layer2_outputs(4128) <= layer1_outputs(8073);
    layer2_outputs(4129) <= not(layer1_outputs(9200));
    layer2_outputs(4130) <= (layer1_outputs(3675)) and (layer1_outputs(1348));
    layer2_outputs(4131) <= not(layer1_outputs(7841));
    layer2_outputs(4132) <= not(layer1_outputs(1888)) or (layer1_outputs(2713));
    layer2_outputs(4133) <= layer1_outputs(3204);
    layer2_outputs(4134) <= not(layer1_outputs(8419));
    layer2_outputs(4135) <= layer1_outputs(5098);
    layer2_outputs(4136) <= not((layer1_outputs(8145)) xor (layer1_outputs(9956)));
    layer2_outputs(4137) <= not((layer1_outputs(8833)) or (layer1_outputs(3757)));
    layer2_outputs(4138) <= not(layer1_outputs(3184));
    layer2_outputs(4139) <= layer1_outputs(344);
    layer2_outputs(4140) <= (layer1_outputs(5418)) and not (layer1_outputs(7372));
    layer2_outputs(4141) <= (layer1_outputs(3836)) and not (layer1_outputs(9321));
    layer2_outputs(4142) <= not(layer1_outputs(2535));
    layer2_outputs(4143) <= not((layer1_outputs(3600)) and (layer1_outputs(2943)));
    layer2_outputs(4144) <= layer1_outputs(784);
    layer2_outputs(4145) <= layer1_outputs(1874);
    layer2_outputs(4146) <= layer1_outputs(3815);
    layer2_outputs(4147) <= not(layer1_outputs(2922));
    layer2_outputs(4148) <= layer1_outputs(9006);
    layer2_outputs(4149) <= not(layer1_outputs(180));
    layer2_outputs(4150) <= not((layer1_outputs(3894)) or (layer1_outputs(7517)));
    layer2_outputs(4151) <= layer1_outputs(464);
    layer2_outputs(4152) <= (layer1_outputs(8372)) or (layer1_outputs(876));
    layer2_outputs(4153) <= layer1_outputs(1162);
    layer2_outputs(4154) <= layer1_outputs(2894);
    layer2_outputs(4155) <= layer1_outputs(6722);
    layer2_outputs(4156) <= (layer1_outputs(1152)) and not (layer1_outputs(1407));
    layer2_outputs(4157) <= not((layer1_outputs(2665)) xor (layer1_outputs(1306)));
    layer2_outputs(4158) <= not(layer1_outputs(2239)) or (layer1_outputs(9936));
    layer2_outputs(4159) <= (layer1_outputs(1069)) and (layer1_outputs(1870));
    layer2_outputs(4160) <= not(layer1_outputs(9205));
    layer2_outputs(4161) <= not(layer1_outputs(2340)) or (layer1_outputs(6358));
    layer2_outputs(4162) <= not(layer1_outputs(370)) or (layer1_outputs(1153));
    layer2_outputs(4163) <= layer1_outputs(6168);
    layer2_outputs(4164) <= layer1_outputs(1087);
    layer2_outputs(4165) <= (layer1_outputs(5993)) and (layer1_outputs(9429));
    layer2_outputs(4166) <= layer1_outputs(1376);
    layer2_outputs(4167) <= (layer1_outputs(7754)) and (layer1_outputs(10047));
    layer2_outputs(4168) <= (layer1_outputs(4593)) and (layer1_outputs(6881));
    layer2_outputs(4169) <= not((layer1_outputs(4409)) and (layer1_outputs(648)));
    layer2_outputs(4170) <= not((layer1_outputs(10154)) or (layer1_outputs(2571)));
    layer2_outputs(4171) <= not(layer1_outputs(674));
    layer2_outputs(4172) <= layer1_outputs(3904);
    layer2_outputs(4173) <= layer1_outputs(4608);
    layer2_outputs(4174) <= (layer1_outputs(9728)) or (layer1_outputs(5156));
    layer2_outputs(4175) <= not(layer1_outputs(1848));
    layer2_outputs(4176) <= layer1_outputs(7806);
    layer2_outputs(4177) <= (layer1_outputs(5602)) and not (layer1_outputs(8799));
    layer2_outputs(4178) <= layer1_outputs(1021);
    layer2_outputs(4179) <= not(layer1_outputs(7921));
    layer2_outputs(4180) <= not(layer1_outputs(2803));
    layer2_outputs(4181) <= layer1_outputs(1982);
    layer2_outputs(4182) <= (layer1_outputs(641)) or (layer1_outputs(5852));
    layer2_outputs(4183) <= not(layer1_outputs(1209));
    layer2_outputs(4184) <= (layer1_outputs(4726)) and (layer1_outputs(8516));
    layer2_outputs(4185) <= (layer1_outputs(5415)) and not (layer1_outputs(4773));
    layer2_outputs(4186) <= not((layer1_outputs(7041)) xor (layer1_outputs(8854)));
    layer2_outputs(4187) <= (layer1_outputs(9932)) xor (layer1_outputs(6572));
    layer2_outputs(4188) <= not(layer1_outputs(3849));
    layer2_outputs(4189) <= not(layer1_outputs(2326));
    layer2_outputs(4190) <= layer1_outputs(7551);
    layer2_outputs(4191) <= not(layer1_outputs(4134)) or (layer1_outputs(2213));
    layer2_outputs(4192) <= not((layer1_outputs(8570)) xor (layer1_outputs(642)));
    layer2_outputs(4193) <= not(layer1_outputs(3007));
    layer2_outputs(4194) <= (layer1_outputs(4295)) or (layer1_outputs(4874));
    layer2_outputs(4195) <= layer1_outputs(6932);
    layer2_outputs(4196) <= not((layer1_outputs(3406)) and (layer1_outputs(8414)));
    layer2_outputs(4197) <= not((layer1_outputs(942)) or (layer1_outputs(4467)));
    layer2_outputs(4198) <= not(layer1_outputs(2500));
    layer2_outputs(4199) <= not((layer1_outputs(1057)) xor (layer1_outputs(957)));
    layer2_outputs(4200) <= not(layer1_outputs(8307));
    layer2_outputs(4201) <= not((layer1_outputs(9423)) and (layer1_outputs(6171)));
    layer2_outputs(4202) <= not(layer1_outputs(5644));
    layer2_outputs(4203) <= not((layer1_outputs(9085)) xor (layer1_outputs(743)));
    layer2_outputs(4204) <= (layer1_outputs(5802)) and not (layer1_outputs(3724));
    layer2_outputs(4205) <= (layer1_outputs(9077)) and not (layer1_outputs(8654));
    layer2_outputs(4206) <= layer1_outputs(6419);
    layer2_outputs(4207) <= not((layer1_outputs(4204)) or (layer1_outputs(5516)));
    layer2_outputs(4208) <= (layer1_outputs(7634)) and (layer1_outputs(8527));
    layer2_outputs(4209) <= not(layer1_outputs(2771));
    layer2_outputs(4210) <= layer1_outputs(6302);
    layer2_outputs(4211) <= '0';
    layer2_outputs(4212) <= not(layer1_outputs(8253));
    layer2_outputs(4213) <= layer1_outputs(4911);
    layer2_outputs(4214) <= not(layer1_outputs(9206));
    layer2_outputs(4215) <= (layer1_outputs(7868)) and not (layer1_outputs(3680));
    layer2_outputs(4216) <= not(layer1_outputs(2547));
    layer2_outputs(4217) <= not(layer1_outputs(8022));
    layer2_outputs(4218) <= (layer1_outputs(6676)) xor (layer1_outputs(1310));
    layer2_outputs(4219) <= layer1_outputs(6522);
    layer2_outputs(4220) <= layer1_outputs(8002);
    layer2_outputs(4221) <= not(layer1_outputs(6459));
    layer2_outputs(4222) <= (layer1_outputs(277)) or (layer1_outputs(8989));
    layer2_outputs(4223) <= not(layer1_outputs(9571)) or (layer1_outputs(9473));
    layer2_outputs(4224) <= not(layer1_outputs(1476));
    layer2_outputs(4225) <= layer1_outputs(8003);
    layer2_outputs(4226) <= layer1_outputs(5010);
    layer2_outputs(4227) <= not(layer1_outputs(5937));
    layer2_outputs(4228) <= not(layer1_outputs(4073));
    layer2_outputs(4229) <= layer1_outputs(6817);
    layer2_outputs(4230) <= not(layer1_outputs(2709)) or (layer1_outputs(7662));
    layer2_outputs(4231) <= not((layer1_outputs(2631)) or (layer1_outputs(9166)));
    layer2_outputs(4232) <= layer1_outputs(3851);
    layer2_outputs(4233) <= layer1_outputs(2599);
    layer2_outputs(4234) <= not((layer1_outputs(312)) or (layer1_outputs(3630)));
    layer2_outputs(4235) <= layer1_outputs(7054);
    layer2_outputs(4236) <= (layer1_outputs(2035)) and (layer1_outputs(6278));
    layer2_outputs(4237) <= not(layer1_outputs(2941));
    layer2_outputs(4238) <= not((layer1_outputs(3300)) and (layer1_outputs(6161)));
    layer2_outputs(4239) <= (layer1_outputs(8825)) xor (layer1_outputs(6892));
    layer2_outputs(4240) <= not(layer1_outputs(7212)) or (layer1_outputs(7672));
    layer2_outputs(4241) <= (layer1_outputs(7324)) and not (layer1_outputs(9520));
    layer2_outputs(4242) <= layer1_outputs(3841);
    layer2_outputs(4243) <= (layer1_outputs(1075)) and (layer1_outputs(2175));
    layer2_outputs(4244) <= (layer1_outputs(7967)) and not (layer1_outputs(2621));
    layer2_outputs(4245) <= (layer1_outputs(1315)) xor (layer1_outputs(8398));
    layer2_outputs(4246) <= not((layer1_outputs(6319)) xor (layer1_outputs(3890)));
    layer2_outputs(4247) <= (layer1_outputs(1479)) and (layer1_outputs(4411));
    layer2_outputs(4248) <= '1';
    layer2_outputs(4249) <= not((layer1_outputs(956)) xor (layer1_outputs(6080)));
    layer2_outputs(4250) <= not(layer1_outputs(3462));
    layer2_outputs(4251) <= not(layer1_outputs(2369));
    layer2_outputs(4252) <= (layer1_outputs(1798)) and (layer1_outputs(6833));
    layer2_outputs(4253) <= layer1_outputs(1200);
    layer2_outputs(4254) <= (layer1_outputs(5897)) xor (layer1_outputs(1017));
    layer2_outputs(4255) <= (layer1_outputs(2420)) xor (layer1_outputs(6577));
    layer2_outputs(4256) <= (layer1_outputs(2881)) xor (layer1_outputs(8281));
    layer2_outputs(4257) <= (layer1_outputs(6974)) and not (layer1_outputs(4116));
    layer2_outputs(4258) <= layer1_outputs(2590);
    layer2_outputs(4259) <= (layer1_outputs(2710)) or (layer1_outputs(9454));
    layer2_outputs(4260) <= layer1_outputs(7646);
    layer2_outputs(4261) <= not(layer1_outputs(4711));
    layer2_outputs(4262) <= (layer1_outputs(7097)) xor (layer1_outputs(2937));
    layer2_outputs(4263) <= not(layer1_outputs(7980));
    layer2_outputs(4264) <= layer1_outputs(3154);
    layer2_outputs(4265) <= layer1_outputs(4180);
    layer2_outputs(4266) <= (layer1_outputs(4202)) or (layer1_outputs(3163));
    layer2_outputs(4267) <= not(layer1_outputs(10137));
    layer2_outputs(4268) <= not(layer1_outputs(7728));
    layer2_outputs(4269) <= not(layer1_outputs(5529));
    layer2_outputs(4270) <= (layer1_outputs(6019)) or (layer1_outputs(6571));
    layer2_outputs(4271) <= not(layer1_outputs(6788));
    layer2_outputs(4272) <= layer1_outputs(2466);
    layer2_outputs(4273) <= not(layer1_outputs(3852));
    layer2_outputs(4274) <= (layer1_outputs(6014)) and not (layer1_outputs(1120));
    layer2_outputs(4275) <= not(layer1_outputs(3722));
    layer2_outputs(4276) <= layer1_outputs(5305);
    layer2_outputs(4277) <= (layer1_outputs(430)) xor (layer1_outputs(4803));
    layer2_outputs(4278) <= layer1_outputs(6421);
    layer2_outputs(4279) <= not(layer1_outputs(5436));
    layer2_outputs(4280) <= layer1_outputs(1596);
    layer2_outputs(4281) <= layer1_outputs(6312);
    layer2_outputs(4282) <= not((layer1_outputs(5973)) and (layer1_outputs(7724)));
    layer2_outputs(4283) <= not(layer1_outputs(4172));
    layer2_outputs(4284) <= not(layer1_outputs(9050));
    layer2_outputs(4285) <= (layer1_outputs(1801)) and (layer1_outputs(3671));
    layer2_outputs(4286) <= not(layer1_outputs(2966));
    layer2_outputs(4287) <= not((layer1_outputs(3046)) or (layer1_outputs(9958)));
    layer2_outputs(4288) <= layer1_outputs(10059);
    layer2_outputs(4289) <= not((layer1_outputs(7805)) or (layer1_outputs(4241)));
    layer2_outputs(4290) <= (layer1_outputs(9007)) or (layer1_outputs(726));
    layer2_outputs(4291) <= layer1_outputs(6434);
    layer2_outputs(4292) <= (layer1_outputs(3092)) xor (layer1_outputs(3556));
    layer2_outputs(4293) <= layer1_outputs(2450);
    layer2_outputs(4294) <= (layer1_outputs(811)) or (layer1_outputs(4405));
    layer2_outputs(4295) <= layer1_outputs(2585);
    layer2_outputs(4296) <= not((layer1_outputs(7491)) and (layer1_outputs(4313)));
    layer2_outputs(4297) <= not(layer1_outputs(9416));
    layer2_outputs(4298) <= (layer1_outputs(2209)) xor (layer1_outputs(5200));
    layer2_outputs(4299) <= (layer1_outputs(4426)) xor (layer1_outputs(548));
    layer2_outputs(4300) <= not(layer1_outputs(2417));
    layer2_outputs(4301) <= not(layer1_outputs(1172));
    layer2_outputs(4302) <= layer1_outputs(542);
    layer2_outputs(4303) <= (layer1_outputs(9435)) and (layer1_outputs(2422));
    layer2_outputs(4304) <= (layer1_outputs(5840)) or (layer1_outputs(9527));
    layer2_outputs(4305) <= (layer1_outputs(5001)) xor (layer1_outputs(7517));
    layer2_outputs(4306) <= layer1_outputs(2697);
    layer2_outputs(4307) <= not((layer1_outputs(4585)) and (layer1_outputs(3017)));
    layer2_outputs(4308) <= not(layer1_outputs(6449));
    layer2_outputs(4309) <= layer1_outputs(6895);
    layer2_outputs(4310) <= (layer1_outputs(5221)) xor (layer1_outputs(2640));
    layer2_outputs(4311) <= not((layer1_outputs(8462)) xor (layer1_outputs(9982)));
    layer2_outputs(4312) <= not(layer1_outputs(1202));
    layer2_outputs(4313) <= layer1_outputs(3783);
    layer2_outputs(4314) <= (layer1_outputs(8871)) and (layer1_outputs(3954));
    layer2_outputs(4315) <= not(layer1_outputs(4265)) or (layer1_outputs(5271));
    layer2_outputs(4316) <= (layer1_outputs(10039)) and not (layer1_outputs(267));
    layer2_outputs(4317) <= (layer1_outputs(1592)) xor (layer1_outputs(902));
    layer2_outputs(4318) <= not(layer1_outputs(4106));
    layer2_outputs(4319) <= not((layer1_outputs(9042)) xor (layer1_outputs(1700)));
    layer2_outputs(4320) <= not(layer1_outputs(5403));
    layer2_outputs(4321) <= layer1_outputs(1164);
    layer2_outputs(4322) <= layer1_outputs(6891);
    layer2_outputs(4323) <= (layer1_outputs(1847)) and not (layer1_outputs(4496));
    layer2_outputs(4324) <= layer1_outputs(768);
    layer2_outputs(4325) <= (layer1_outputs(1322)) and not (layer1_outputs(4666));
    layer2_outputs(4326) <= not(layer1_outputs(4757));
    layer2_outputs(4327) <= not(layer1_outputs(6742)) or (layer1_outputs(7330));
    layer2_outputs(4328) <= (layer1_outputs(2656)) or (layer1_outputs(8437));
    layer2_outputs(4329) <= not(layer1_outputs(8432));
    layer2_outputs(4330) <= not(layer1_outputs(4957));
    layer2_outputs(4331) <= not(layer1_outputs(233));
    layer2_outputs(4332) <= layer1_outputs(5572);
    layer2_outputs(4333) <= not(layer1_outputs(1889));
    layer2_outputs(4334) <= not((layer1_outputs(4292)) or (layer1_outputs(3883)));
    layer2_outputs(4335) <= (layer1_outputs(4966)) or (layer1_outputs(9106));
    layer2_outputs(4336) <= not(layer1_outputs(7427));
    layer2_outputs(4337) <= not(layer1_outputs(2521));
    layer2_outputs(4338) <= not(layer1_outputs(169));
    layer2_outputs(4339) <= layer1_outputs(655);
    layer2_outputs(4340) <= not(layer1_outputs(8650));
    layer2_outputs(4341) <= (layer1_outputs(6)) and (layer1_outputs(7559));
    layer2_outputs(4342) <= layer1_outputs(14);
    layer2_outputs(4343) <= not((layer1_outputs(6408)) or (layer1_outputs(2574)));
    layer2_outputs(4344) <= (layer1_outputs(5808)) or (layer1_outputs(9880));
    layer2_outputs(4345) <= layer1_outputs(7744);
    layer2_outputs(4346) <= (layer1_outputs(5926)) and not (layer1_outputs(1655));
    layer2_outputs(4347) <= not(layer1_outputs(7289));
    layer2_outputs(4348) <= (layer1_outputs(2117)) and not (layer1_outputs(3214));
    layer2_outputs(4349) <= (layer1_outputs(7484)) and (layer1_outputs(4952));
    layer2_outputs(4350) <= not(layer1_outputs(7689));
    layer2_outputs(4351) <= (layer1_outputs(1240)) and not (layer1_outputs(5561));
    layer2_outputs(4352) <= layer1_outputs(3403);
    layer2_outputs(4353) <= not(layer1_outputs(3741));
    layer2_outputs(4354) <= layer1_outputs(4014);
    layer2_outputs(4355) <= not((layer1_outputs(8920)) xor (layer1_outputs(2099)));
    layer2_outputs(4356) <= layer1_outputs(9043);
    layer2_outputs(4357) <= (layer1_outputs(6424)) xor (layer1_outputs(6431));
    layer2_outputs(4358) <= not(layer1_outputs(7955)) or (layer1_outputs(8020));
    layer2_outputs(4359) <= not(layer1_outputs(3751));
    layer2_outputs(4360) <= (layer1_outputs(6244)) xor (layer1_outputs(4212));
    layer2_outputs(4361) <= (layer1_outputs(2965)) and not (layer1_outputs(3450));
    layer2_outputs(4362) <= not(layer1_outputs(419));
    layer2_outputs(4363) <= not((layer1_outputs(5578)) xor (layer1_outputs(1966)));
    layer2_outputs(4364) <= layer1_outputs(1854);
    layer2_outputs(4365) <= (layer1_outputs(6478)) or (layer1_outputs(5956));
    layer2_outputs(4366) <= not(layer1_outputs(4584));
    layer2_outputs(4367) <= layer1_outputs(4060);
    layer2_outputs(4368) <= not((layer1_outputs(780)) xor (layer1_outputs(4099)));
    layer2_outputs(4369) <= not(layer1_outputs(3126)) or (layer1_outputs(6484));
    layer2_outputs(4370) <= (layer1_outputs(8104)) and not (layer1_outputs(9945));
    layer2_outputs(4371) <= not(layer1_outputs(6945));
    layer2_outputs(4372) <= not((layer1_outputs(3692)) or (layer1_outputs(5298)));
    layer2_outputs(4373) <= (layer1_outputs(2026)) or (layer1_outputs(753));
    layer2_outputs(4374) <= (layer1_outputs(5094)) xor (layer1_outputs(7218));
    layer2_outputs(4375) <= not((layer1_outputs(6035)) xor (layer1_outputs(1373)));
    layer2_outputs(4376) <= not(layer1_outputs(1444));
    layer2_outputs(4377) <= not(layer1_outputs(6445));
    layer2_outputs(4378) <= layer1_outputs(4418);
    layer2_outputs(4379) <= layer1_outputs(6293);
    layer2_outputs(4380) <= not((layer1_outputs(1313)) xor (layer1_outputs(7928)));
    layer2_outputs(4381) <= layer1_outputs(1362);
    layer2_outputs(4382) <= layer1_outputs(10178);
    layer2_outputs(4383) <= layer1_outputs(8030);
    layer2_outputs(4384) <= not(layer1_outputs(10102));
    layer2_outputs(4385) <= layer1_outputs(2293);
    layer2_outputs(4386) <= (layer1_outputs(492)) or (layer1_outputs(9271));
    layer2_outputs(4387) <= not((layer1_outputs(9247)) or (layer1_outputs(3039)));
    layer2_outputs(4388) <= not(layer1_outputs(124));
    layer2_outputs(4389) <= layer1_outputs(9231);
    layer2_outputs(4390) <= (layer1_outputs(9898)) xor (layer1_outputs(5211));
    layer2_outputs(4391) <= (layer1_outputs(7600)) and not (layer1_outputs(9871));
    layer2_outputs(4392) <= (layer1_outputs(885)) xor (layer1_outputs(4634));
    layer2_outputs(4393) <= (layer1_outputs(8285)) and not (layer1_outputs(1196));
    layer2_outputs(4394) <= layer1_outputs(4900);
    layer2_outputs(4395) <= not(layer1_outputs(7082));
    layer2_outputs(4396) <= layer1_outputs(9285);
    layer2_outputs(4397) <= layer1_outputs(9559);
    layer2_outputs(4398) <= (layer1_outputs(2643)) or (layer1_outputs(10012));
    layer2_outputs(4399) <= (layer1_outputs(2336)) and not (layer1_outputs(6582));
    layer2_outputs(4400) <= not(layer1_outputs(1)) or (layer1_outputs(3143));
    layer2_outputs(4401) <= layer1_outputs(5812);
    layer2_outputs(4402) <= not(layer1_outputs(8913));
    layer2_outputs(4403) <= not(layer1_outputs(7135));
    layer2_outputs(4404) <= not(layer1_outputs(1261));
    layer2_outputs(4405) <= layer1_outputs(9008);
    layer2_outputs(4406) <= layer1_outputs(6674);
    layer2_outputs(4407) <= not(layer1_outputs(7911)) or (layer1_outputs(3345));
    layer2_outputs(4408) <= not(layer1_outputs(6119));
    layer2_outputs(4409) <= not(layer1_outputs(6410));
    layer2_outputs(4410) <= layer1_outputs(2075);
    layer2_outputs(4411) <= (layer1_outputs(2448)) xor (layer1_outputs(3663));
    layer2_outputs(4412) <= not(layer1_outputs(5851));
    layer2_outputs(4413) <= not(layer1_outputs(1549));
    layer2_outputs(4414) <= layer1_outputs(9738);
    layer2_outputs(4415) <= '0';
    layer2_outputs(4416) <= not(layer1_outputs(1526));
    layer2_outputs(4417) <= layer1_outputs(8958);
    layer2_outputs(4418) <= not((layer1_outputs(6555)) and (layer1_outputs(1064)));
    layer2_outputs(4419) <= layer1_outputs(8137);
    layer2_outputs(4420) <= not(layer1_outputs(9733)) or (layer1_outputs(7074));
    layer2_outputs(4421) <= layer1_outputs(6512);
    layer2_outputs(4422) <= layer1_outputs(6756);
    layer2_outputs(4423) <= layer1_outputs(5307);
    layer2_outputs(4424) <= layer1_outputs(6571);
    layer2_outputs(4425) <= not(layer1_outputs(10107)) or (layer1_outputs(8012));
    layer2_outputs(4426) <= not(layer1_outputs(9159));
    layer2_outputs(4427) <= layer1_outputs(9804);
    layer2_outputs(4428) <= not((layer1_outputs(9860)) or (layer1_outputs(3286)));
    layer2_outputs(4429) <= not(layer1_outputs(10103)) or (layer1_outputs(4507));
    layer2_outputs(4430) <= not((layer1_outputs(2177)) or (layer1_outputs(8942)));
    layer2_outputs(4431) <= not(layer1_outputs(2549));
    layer2_outputs(4432) <= not(layer1_outputs(7345));
    layer2_outputs(4433) <= layer1_outputs(5900);
    layer2_outputs(4434) <= not(layer1_outputs(4371));
    layer2_outputs(4435) <= (layer1_outputs(6163)) and not (layer1_outputs(140));
    layer2_outputs(4436) <= '0';
    layer2_outputs(4437) <= layer1_outputs(2455);
    layer2_outputs(4438) <= '0';
    layer2_outputs(4439) <= not((layer1_outputs(4617)) xor (layer1_outputs(45)));
    layer2_outputs(4440) <= not((layer1_outputs(5759)) and (layer1_outputs(5434)));
    layer2_outputs(4441) <= not((layer1_outputs(5046)) xor (layer1_outputs(3637)));
    layer2_outputs(4442) <= not((layer1_outputs(9824)) xor (layer1_outputs(1642)));
    layer2_outputs(4443) <= not((layer1_outputs(237)) xor (layer1_outputs(8013)));
    layer2_outputs(4444) <= not(layer1_outputs(7854));
    layer2_outputs(4445) <= layer1_outputs(9375);
    layer2_outputs(4446) <= not((layer1_outputs(1608)) xor (layer1_outputs(95)));
    layer2_outputs(4447) <= layer1_outputs(689);
    layer2_outputs(4448) <= not(layer1_outputs(875));
    layer2_outputs(4449) <= not(layer1_outputs(7456)) or (layer1_outputs(9433));
    layer2_outputs(4450) <= not(layer1_outputs(7936));
    layer2_outputs(4451) <= not((layer1_outputs(9954)) and (layer1_outputs(9930)));
    layer2_outputs(4452) <= not(layer1_outputs(9218));
    layer2_outputs(4453) <= layer1_outputs(233);
    layer2_outputs(4454) <= not(layer1_outputs(290));
    layer2_outputs(4455) <= not((layer1_outputs(4671)) or (layer1_outputs(10134)));
    layer2_outputs(4456) <= not(layer1_outputs(3035));
    layer2_outputs(4457) <= (layer1_outputs(8179)) and (layer1_outputs(9661));
    layer2_outputs(4458) <= not(layer1_outputs(2677));
    layer2_outputs(4459) <= layer1_outputs(3471);
    layer2_outputs(4460) <= (layer1_outputs(1968)) or (layer1_outputs(7048));
    layer2_outputs(4461) <= (layer1_outputs(5082)) xor (layer1_outputs(354));
    layer2_outputs(4462) <= layer1_outputs(6879);
    layer2_outputs(4463) <= not(layer1_outputs(8639));
    layer2_outputs(4464) <= layer1_outputs(10196);
    layer2_outputs(4465) <= (layer1_outputs(1956)) and (layer1_outputs(3513));
    layer2_outputs(4466) <= layer1_outputs(7930);
    layer2_outputs(4467) <= layer1_outputs(8453);
    layer2_outputs(4468) <= not((layer1_outputs(3659)) and (layer1_outputs(4797)));
    layer2_outputs(4469) <= (layer1_outputs(6931)) and not (layer1_outputs(7196));
    layer2_outputs(4470) <= layer1_outputs(2591);
    layer2_outputs(4471) <= layer1_outputs(6082);
    layer2_outputs(4472) <= not(layer1_outputs(1575)) or (layer1_outputs(8100));
    layer2_outputs(4473) <= not(layer1_outputs(3656));
    layer2_outputs(4474) <= (layer1_outputs(3555)) xor (layer1_outputs(4565));
    layer2_outputs(4475) <= not(layer1_outputs(448));
    layer2_outputs(4476) <= (layer1_outputs(7749)) and (layer1_outputs(301));
    layer2_outputs(4477) <= layer1_outputs(5285);
    layer2_outputs(4478) <= layer1_outputs(8342);
    layer2_outputs(4479) <= '0';
    layer2_outputs(4480) <= (layer1_outputs(3342)) and (layer1_outputs(9575));
    layer2_outputs(4481) <= (layer1_outputs(559)) xor (layer1_outputs(8322));
    layer2_outputs(4482) <= not((layer1_outputs(607)) or (layer1_outputs(107)));
    layer2_outputs(4483) <= not(layer1_outputs(2254));
    layer2_outputs(4484) <= not(layer1_outputs(1600));
    layer2_outputs(4485) <= not(layer1_outputs(4895)) or (layer1_outputs(1243));
    layer2_outputs(4486) <= not(layer1_outputs(2468));
    layer2_outputs(4487) <= not(layer1_outputs(2193));
    layer2_outputs(4488) <= layer1_outputs(9333);
    layer2_outputs(4489) <= (layer1_outputs(1614)) and not (layer1_outputs(651));
    layer2_outputs(4490) <= not((layer1_outputs(3472)) and (layer1_outputs(6977)));
    layer2_outputs(4491) <= layer1_outputs(8458);
    layer2_outputs(4492) <= layer1_outputs(7763);
    layer2_outputs(4493) <= not(layer1_outputs(6996));
    layer2_outputs(4494) <= not(layer1_outputs(1885)) or (layer1_outputs(8576));
    layer2_outputs(4495) <= not((layer1_outputs(509)) and (layer1_outputs(615)));
    layer2_outputs(4496) <= not((layer1_outputs(7671)) or (layer1_outputs(7447)));
    layer2_outputs(4497) <= (layer1_outputs(8151)) and not (layer1_outputs(7394));
    layer2_outputs(4498) <= not((layer1_outputs(8121)) and (layer1_outputs(2457)));
    layer2_outputs(4499) <= not(layer1_outputs(8344)) or (layer1_outputs(697));
    layer2_outputs(4500) <= not(layer1_outputs(1433));
    layer2_outputs(4501) <= not(layer1_outputs(1784));
    layer2_outputs(4502) <= layer1_outputs(6319);
    layer2_outputs(4503) <= layer1_outputs(6635);
    layer2_outputs(4504) <= not(layer1_outputs(7855));
    layer2_outputs(4505) <= (layer1_outputs(1463)) and (layer1_outputs(6152));
    layer2_outputs(4506) <= (layer1_outputs(6083)) xor (layer1_outputs(9260));
    layer2_outputs(4507) <= not(layer1_outputs(8575));
    layer2_outputs(4508) <= not((layer1_outputs(9193)) and (layer1_outputs(5617)));
    layer2_outputs(4509) <= not(layer1_outputs(5976));
    layer2_outputs(4510) <= (layer1_outputs(2059)) and not (layer1_outputs(7090));
    layer2_outputs(4511) <= not(layer1_outputs(1266));
    layer2_outputs(4512) <= layer1_outputs(2294);
    layer2_outputs(4513) <= layer1_outputs(726);
    layer2_outputs(4514) <= not(layer1_outputs(3364));
    layer2_outputs(4515) <= layer1_outputs(4973);
    layer2_outputs(4516) <= (layer1_outputs(4587)) and (layer1_outputs(8923));
    layer2_outputs(4517) <= not((layer1_outputs(7929)) xor (layer1_outputs(3147)));
    layer2_outputs(4518) <= not(layer1_outputs(5006));
    layer2_outputs(4519) <= not(layer1_outputs(4360));
    layer2_outputs(4520) <= not(layer1_outputs(8177));
    layer2_outputs(4521) <= layer1_outputs(4862);
    layer2_outputs(4522) <= not(layer1_outputs(8782));
    layer2_outputs(4523) <= layer1_outputs(4588);
    layer2_outputs(4524) <= not(layer1_outputs(365)) or (layer1_outputs(3266));
    layer2_outputs(4525) <= (layer1_outputs(3447)) and (layer1_outputs(3911));
    layer2_outputs(4526) <= layer1_outputs(8757);
    layer2_outputs(4527) <= (layer1_outputs(6897)) and not (layer1_outputs(6176));
    layer2_outputs(4528) <= not(layer1_outputs(5328)) or (layer1_outputs(9894));
    layer2_outputs(4529) <= layer1_outputs(4556);
    layer2_outputs(4530) <= not(layer1_outputs(4363));
    layer2_outputs(4531) <= (layer1_outputs(10223)) or (layer1_outputs(1893));
    layer2_outputs(4532) <= not((layer1_outputs(3350)) xor (layer1_outputs(4451)));
    layer2_outputs(4533) <= (layer1_outputs(850)) and not (layer1_outputs(5863));
    layer2_outputs(4534) <= not(layer1_outputs(3799));
    layer2_outputs(4535) <= not(layer1_outputs(4683)) or (layer1_outputs(6619));
    layer2_outputs(4536) <= not(layer1_outputs(3583));
    layer2_outputs(4537) <= (layer1_outputs(6575)) xor (layer1_outputs(5994));
    layer2_outputs(4538) <= not(layer1_outputs(2022));
    layer2_outputs(4539) <= not(layer1_outputs(2296));
    layer2_outputs(4540) <= not(layer1_outputs(1696));
    layer2_outputs(4541) <= layer1_outputs(10144);
    layer2_outputs(4542) <= not(layer1_outputs(3431));
    layer2_outputs(4543) <= not(layer1_outputs(9650));
    layer2_outputs(4544) <= layer1_outputs(2714);
    layer2_outputs(4545) <= (layer1_outputs(6989)) and not (layer1_outputs(5724));
    layer2_outputs(4546) <= not(layer1_outputs(7298));
    layer2_outputs(4547) <= (layer1_outputs(6467)) xor (layer1_outputs(1002));
    layer2_outputs(4548) <= not((layer1_outputs(309)) xor (layer1_outputs(1566)));
    layer2_outputs(4549) <= layer1_outputs(7199);
    layer2_outputs(4550) <= not(layer1_outputs(669));
    layer2_outputs(4551) <= not((layer1_outputs(7867)) or (layer1_outputs(537)));
    layer2_outputs(4552) <= not((layer1_outputs(9409)) and (layer1_outputs(3669)));
    layer2_outputs(4553) <= layer1_outputs(3030);
    layer2_outputs(4554) <= layer1_outputs(5932);
    layer2_outputs(4555) <= layer1_outputs(1546);
    layer2_outputs(4556) <= layer1_outputs(6610);
    layer2_outputs(4557) <= not(layer1_outputs(4461));
    layer2_outputs(4558) <= not(layer1_outputs(516));
    layer2_outputs(4559) <= (layer1_outputs(7615)) xor (layer1_outputs(7917));
    layer2_outputs(4560) <= (layer1_outputs(3829)) xor (layer1_outputs(5092));
    layer2_outputs(4561) <= not(layer1_outputs(5083));
    layer2_outputs(4562) <= (layer1_outputs(3071)) or (layer1_outputs(8065));
    layer2_outputs(4563) <= layer1_outputs(3706);
    layer2_outputs(4564) <= not(layer1_outputs(10237));
    layer2_outputs(4565) <= (layer1_outputs(8618)) and not (layer1_outputs(10070));
    layer2_outputs(4566) <= layer1_outputs(6991);
    layer2_outputs(4567) <= not(layer1_outputs(4879));
    layer2_outputs(4568) <= (layer1_outputs(3170)) xor (layer1_outputs(5072));
    layer2_outputs(4569) <= layer1_outputs(2771);
    layer2_outputs(4570) <= (layer1_outputs(8822)) xor (layer1_outputs(7112));
    layer2_outputs(4571) <= layer1_outputs(8081);
    layer2_outputs(4572) <= not(layer1_outputs(2333)) or (layer1_outputs(2138));
    layer2_outputs(4573) <= not(layer1_outputs(1689)) or (layer1_outputs(3643));
    layer2_outputs(4574) <= not(layer1_outputs(2196));
    layer2_outputs(4575) <= not(layer1_outputs(245));
    layer2_outputs(4576) <= layer1_outputs(6867);
    layer2_outputs(4577) <= layer1_outputs(6900);
    layer2_outputs(4578) <= layer1_outputs(243);
    layer2_outputs(4579) <= not((layer1_outputs(195)) xor (layer1_outputs(3143)));
    layer2_outputs(4580) <= (layer1_outputs(9082)) xor (layer1_outputs(177));
    layer2_outputs(4581) <= not(layer1_outputs(6375)) or (layer1_outputs(3862));
    layer2_outputs(4582) <= layer1_outputs(9588);
    layer2_outputs(4583) <= (layer1_outputs(6500)) or (layer1_outputs(5330));
    layer2_outputs(4584) <= not(layer1_outputs(5320));
    layer2_outputs(4585) <= (layer1_outputs(4322)) and not (layer1_outputs(4469));
    layer2_outputs(4586) <= layer1_outputs(6445);
    layer2_outputs(4587) <= not(layer1_outputs(4633));
    layer2_outputs(4588) <= (layer1_outputs(8595)) and not (layer1_outputs(6182));
    layer2_outputs(4589) <= not((layer1_outputs(3470)) or (layer1_outputs(10145)));
    layer2_outputs(4590) <= not(layer1_outputs(5035));
    layer2_outputs(4591) <= not(layer1_outputs(3095));
    layer2_outputs(4592) <= not((layer1_outputs(7354)) and (layer1_outputs(3114)));
    layer2_outputs(4593) <= (layer1_outputs(352)) or (layer1_outputs(9583));
    layer2_outputs(4594) <= layer1_outputs(7879);
    layer2_outputs(4595) <= (layer1_outputs(6249)) and not (layer1_outputs(5633));
    layer2_outputs(4596) <= not(layer1_outputs(3407)) or (layer1_outputs(1994));
    layer2_outputs(4597) <= (layer1_outputs(3508)) xor (layer1_outputs(1595));
    layer2_outputs(4598) <= not(layer1_outputs(8438));
    layer2_outputs(4599) <= (layer1_outputs(9439)) and not (layer1_outputs(1365));
    layer2_outputs(4600) <= not((layer1_outputs(4065)) and (layer1_outputs(2134)));
    layer2_outputs(4601) <= (layer1_outputs(678)) and not (layer1_outputs(2086));
    layer2_outputs(4602) <= (layer1_outputs(1933)) or (layer1_outputs(3263));
    layer2_outputs(4603) <= not(layer1_outputs(7210));
    layer2_outputs(4604) <= layer1_outputs(8134);
    layer2_outputs(4605) <= (layer1_outputs(5788)) or (layer1_outputs(4564));
    layer2_outputs(4606) <= not(layer1_outputs(3107));
    layer2_outputs(4607) <= (layer1_outputs(4934)) or (layer1_outputs(423));
    layer2_outputs(4608) <= not((layer1_outputs(3704)) xor (layer1_outputs(7413)));
    layer2_outputs(4609) <= layer1_outputs(1160);
    layer2_outputs(4610) <= not(layer1_outputs(5613)) or (layer1_outputs(3008));
    layer2_outputs(4611) <= (layer1_outputs(4302)) or (layer1_outputs(7374));
    layer2_outputs(4612) <= not(layer1_outputs(5673));
    layer2_outputs(4613) <= not(layer1_outputs(8591));
    layer2_outputs(4614) <= (layer1_outputs(5943)) xor (layer1_outputs(8768));
    layer2_outputs(4615) <= not(layer1_outputs(6259));
    layer2_outputs(4616) <= (layer1_outputs(5079)) and not (layer1_outputs(3856));
    layer2_outputs(4617) <= not((layer1_outputs(1305)) and (layer1_outputs(10184)));
    layer2_outputs(4618) <= not(layer1_outputs(4332));
    layer2_outputs(4619) <= not((layer1_outputs(7940)) xor (layer1_outputs(10027)));
    layer2_outputs(4620) <= not((layer1_outputs(158)) xor (layer1_outputs(4719)));
    layer2_outputs(4621) <= '0';
    layer2_outputs(4622) <= not((layer1_outputs(2720)) and (layer1_outputs(9049)));
    layer2_outputs(4623) <= (layer1_outputs(3357)) xor (layer1_outputs(9237));
    layer2_outputs(4624) <= not(layer1_outputs(6700));
    layer2_outputs(4625) <= layer1_outputs(2583);
    layer2_outputs(4626) <= layer1_outputs(1999);
    layer2_outputs(4627) <= not(layer1_outputs(5008)) or (layer1_outputs(8582));
    layer2_outputs(4628) <= not(layer1_outputs(4894));
    layer2_outputs(4629) <= not(layer1_outputs(6282)) or (layer1_outputs(8949));
    layer2_outputs(4630) <= (layer1_outputs(6968)) or (layer1_outputs(7961));
    layer2_outputs(4631) <= (layer1_outputs(5629)) or (layer1_outputs(5711));
    layer2_outputs(4632) <= not(layer1_outputs(410));
    layer2_outputs(4633) <= not(layer1_outputs(6504));
    layer2_outputs(4634) <= not(layer1_outputs(10206)) or (layer1_outputs(9613));
    layer2_outputs(4635) <= layer1_outputs(5289);
    layer2_outputs(4636) <= not(layer1_outputs(6621)) or (layer1_outputs(5345));
    layer2_outputs(4637) <= '1';
    layer2_outputs(4638) <= not(layer1_outputs(2119)) or (layer1_outputs(2435));
    layer2_outputs(4639) <= (layer1_outputs(6760)) xor (layer1_outputs(8279));
    layer2_outputs(4640) <= (layer1_outputs(7964)) and not (layer1_outputs(771));
    layer2_outputs(4641) <= not(layer1_outputs(5896)) or (layer1_outputs(6079));
    layer2_outputs(4642) <= not(layer1_outputs(3615));
    layer2_outputs(4643) <= not(layer1_outputs(9268));
    layer2_outputs(4644) <= not((layer1_outputs(2900)) and (layer1_outputs(4694)));
    layer2_outputs(4645) <= not((layer1_outputs(8410)) and (layer1_outputs(1953)));
    layer2_outputs(4646) <= not(layer1_outputs(1661));
    layer2_outputs(4647) <= not(layer1_outputs(4717));
    layer2_outputs(4648) <= layer1_outputs(592);
    layer2_outputs(4649) <= not((layer1_outputs(3376)) and (layer1_outputs(6417)));
    layer2_outputs(4650) <= (layer1_outputs(5777)) xor (layer1_outputs(2195));
    layer2_outputs(4651) <= (layer1_outputs(4285)) and (layer1_outputs(8828));
    layer2_outputs(4652) <= layer1_outputs(10202);
    layer2_outputs(4653) <= not((layer1_outputs(2405)) and (layer1_outputs(2162)));
    layer2_outputs(4654) <= layer1_outputs(10221);
    layer2_outputs(4655) <= not(layer1_outputs(5587));
    layer2_outputs(4656) <= layer1_outputs(5020);
    layer2_outputs(4657) <= not(layer1_outputs(2698));
    layer2_outputs(4658) <= not(layer1_outputs(6769)) or (layer1_outputs(6232));
    layer2_outputs(4659) <= layer1_outputs(4802);
    layer2_outputs(4660) <= (layer1_outputs(10094)) and not (layer1_outputs(838));
    layer2_outputs(4661) <= not(layer1_outputs(7757));
    layer2_outputs(4662) <= (layer1_outputs(8875)) xor (layer1_outputs(6116));
    layer2_outputs(4663) <= not(layer1_outputs(1014)) or (layer1_outputs(8413));
    layer2_outputs(4664) <= not(layer1_outputs(5301)) or (layer1_outputs(8066));
    layer2_outputs(4665) <= not((layer1_outputs(7141)) xor (layer1_outputs(2981)));
    layer2_outputs(4666) <= not(layer1_outputs(1591));
    layer2_outputs(4667) <= not(layer1_outputs(5807));
    layer2_outputs(4668) <= not(layer1_outputs(845));
    layer2_outputs(4669) <= not(layer1_outputs(4017)) or (layer1_outputs(3026));
    layer2_outputs(4670) <= layer1_outputs(2452);
    layer2_outputs(4671) <= not(layer1_outputs(9461));
    layer2_outputs(4672) <= not(layer1_outputs(1811)) or (layer1_outputs(2797));
    layer2_outputs(4673) <= not(layer1_outputs(4845));
    layer2_outputs(4674) <= not(layer1_outputs(663)) or (layer1_outputs(9116));
    layer2_outputs(4675) <= not((layer1_outputs(7651)) xor (layer1_outputs(79)));
    layer2_outputs(4676) <= not((layer1_outputs(4345)) xor (layer1_outputs(7875)));
    layer2_outputs(4677) <= not((layer1_outputs(8490)) or (layer1_outputs(7098)));
    layer2_outputs(4678) <= not(layer1_outputs(2118));
    layer2_outputs(4679) <= layer1_outputs(254);
    layer2_outputs(4680) <= not(layer1_outputs(10051));
    layer2_outputs(4681) <= (layer1_outputs(6207)) xor (layer1_outputs(8110));
    layer2_outputs(4682) <= (layer1_outputs(9619)) xor (layer1_outputs(3528));
    layer2_outputs(4683) <= '1';
    layer2_outputs(4684) <= layer1_outputs(5381);
    layer2_outputs(4685) <= not(layer1_outputs(2347));
    layer2_outputs(4686) <= not(layer1_outputs(10223));
    layer2_outputs(4687) <= not(layer1_outputs(8566));
    layer2_outputs(4688) <= (layer1_outputs(1823)) or (layer1_outputs(2091));
    layer2_outputs(4689) <= layer1_outputs(4955);
    layer2_outputs(4690) <= not(layer1_outputs(7348)) or (layer1_outputs(2672));
    layer2_outputs(4691) <= not(layer1_outputs(6224));
    layer2_outputs(4692) <= not((layer1_outputs(2267)) xor (layer1_outputs(3875)));
    layer2_outputs(4693) <= not(layer1_outputs(2536));
    layer2_outputs(4694) <= layer1_outputs(9313);
    layer2_outputs(4695) <= not(layer1_outputs(2618)) or (layer1_outputs(948));
    layer2_outputs(4696) <= not((layer1_outputs(1496)) and (layer1_outputs(8356)));
    layer2_outputs(4697) <= layer1_outputs(4110);
    layer2_outputs(4698) <= layer1_outputs(6011);
    layer2_outputs(4699) <= layer1_outputs(351);
    layer2_outputs(4700) <= (layer1_outputs(3652)) xor (layer1_outputs(4553));
    layer2_outputs(4701) <= not((layer1_outputs(1141)) and (layer1_outputs(4669)));
    layer2_outputs(4702) <= (layer1_outputs(1043)) and not (layer1_outputs(372));
    layer2_outputs(4703) <= not(layer1_outputs(5122));
    layer2_outputs(4704) <= not(layer1_outputs(8147));
    layer2_outputs(4705) <= not(layer1_outputs(3752));
    layer2_outputs(4706) <= '1';
    layer2_outputs(4707) <= not((layer1_outputs(10061)) xor (layer1_outputs(2483)));
    layer2_outputs(4708) <= (layer1_outputs(8995)) and not (layer1_outputs(7912));
    layer2_outputs(4709) <= not(layer1_outputs(5209));
    layer2_outputs(4710) <= (layer1_outputs(668)) or (layer1_outputs(10238));
    layer2_outputs(4711) <= not(layer1_outputs(9324));
    layer2_outputs(4712) <= not(layer1_outputs(2085));
    layer2_outputs(4713) <= layer1_outputs(9606);
    layer2_outputs(4714) <= not(layer1_outputs(9864));
    layer2_outputs(4715) <= not(layer1_outputs(9119));
    layer2_outputs(4716) <= (layer1_outputs(8980)) and (layer1_outputs(4189));
    layer2_outputs(4717) <= not((layer1_outputs(2895)) or (layer1_outputs(7166)));
    layer2_outputs(4718) <= layer1_outputs(662);
    layer2_outputs(4719) <= not(layer1_outputs(9766));
    layer2_outputs(4720) <= (layer1_outputs(2244)) xor (layer1_outputs(6597));
    layer2_outputs(4721) <= not((layer1_outputs(4262)) xor (layer1_outputs(1008)));
    layer2_outputs(4722) <= (layer1_outputs(882)) xor (layer1_outputs(2961));
    layer2_outputs(4723) <= layer1_outputs(6924);
    layer2_outputs(4724) <= (layer1_outputs(4858)) xor (layer1_outputs(8015));
    layer2_outputs(4725) <= layer1_outputs(918);
    layer2_outputs(4726) <= (layer1_outputs(8303)) and not (layer1_outputs(4638));
    layer2_outputs(4727) <= not(layer1_outputs(1534));
    layer2_outputs(4728) <= layer1_outputs(7442);
    layer2_outputs(4729) <= layer1_outputs(5101);
    layer2_outputs(4730) <= not(layer1_outputs(5334));
    layer2_outputs(4731) <= not(layer1_outputs(9193));
    layer2_outputs(4732) <= layer1_outputs(7459);
    layer2_outputs(4733) <= not(layer1_outputs(6987));
    layer2_outputs(4734) <= not(layer1_outputs(4386));
    layer2_outputs(4735) <= not(layer1_outputs(6548));
    layer2_outputs(4736) <= not(layer1_outputs(8325)) or (layer1_outputs(3291));
    layer2_outputs(4737) <= not(layer1_outputs(7755));
    layer2_outputs(4738) <= not(layer1_outputs(6664));
    layer2_outputs(4739) <= not(layer1_outputs(2567));
    layer2_outputs(4740) <= layer1_outputs(736);
    layer2_outputs(4741) <= layer1_outputs(1432);
    layer2_outputs(4742) <= (layer1_outputs(933)) xor (layer1_outputs(8529));
    layer2_outputs(4743) <= not((layer1_outputs(3893)) and (layer1_outputs(650)));
    layer2_outputs(4744) <= not((layer1_outputs(4786)) xor (layer1_outputs(1095)));
    layer2_outputs(4745) <= layer1_outputs(4092);
    layer2_outputs(4746) <= layer1_outputs(375);
    layer2_outputs(4747) <= (layer1_outputs(4833)) and not (layer1_outputs(1161));
    layer2_outputs(4748) <= not(layer1_outputs(4965)) or (layer1_outputs(8784));
    layer2_outputs(4749) <= layer1_outputs(7281);
    layer2_outputs(4750) <= not((layer1_outputs(8244)) and (layer1_outputs(4532)));
    layer2_outputs(4751) <= (layer1_outputs(9280)) and (layer1_outputs(6673));
    layer2_outputs(4752) <= not(layer1_outputs(10135)) or (layer1_outputs(4004));
    layer2_outputs(4753) <= layer1_outputs(1936);
    layer2_outputs(4754) <= not((layer1_outputs(3712)) xor (layer1_outputs(4748)));
    layer2_outputs(4755) <= not(layer1_outputs(7862));
    layer2_outputs(4756) <= not(layer1_outputs(4019)) or (layer1_outputs(470));
    layer2_outputs(4757) <= not(layer1_outputs(7268));
    layer2_outputs(4758) <= (layer1_outputs(7423)) xor (layer1_outputs(5978));
    layer2_outputs(4759) <= layer1_outputs(6480);
    layer2_outputs(4760) <= not(layer1_outputs(381));
    layer2_outputs(4761) <= not(layer1_outputs(5448)) or (layer1_outputs(6743));
    layer2_outputs(4762) <= not((layer1_outputs(3125)) xor (layer1_outputs(1111)));
    layer2_outputs(4763) <= not((layer1_outputs(5220)) xor (layer1_outputs(3076)));
    layer2_outputs(4764) <= layer1_outputs(7706);
    layer2_outputs(4765) <= not(layer1_outputs(1176)) or (layer1_outputs(5491));
    layer2_outputs(4766) <= layer1_outputs(8035);
    layer2_outputs(4767) <= (layer1_outputs(2736)) or (layer1_outputs(6713));
    layer2_outputs(4768) <= not((layer1_outputs(5552)) or (layer1_outputs(9335)));
    layer2_outputs(4769) <= not(layer1_outputs(8168)) or (layer1_outputs(8761));
    layer2_outputs(4770) <= layer1_outputs(6360);
    layer2_outputs(4771) <= (layer1_outputs(5898)) and (layer1_outputs(4916));
    layer2_outputs(4772) <= not((layer1_outputs(8167)) or (layer1_outputs(8747)));
    layer2_outputs(4773) <= not(layer1_outputs(3647));
    layer2_outputs(4774) <= layer1_outputs(5590);
    layer2_outputs(4775) <= (layer1_outputs(5458)) and not (layer1_outputs(1012));
    layer2_outputs(4776) <= layer1_outputs(9853);
    layer2_outputs(4777) <= layer1_outputs(5044);
    layer2_outputs(4778) <= layer1_outputs(6302);
    layer2_outputs(4779) <= layer1_outputs(9528);
    layer2_outputs(4780) <= layer1_outputs(6711);
    layer2_outputs(4781) <= not(layer1_outputs(2056)) or (layer1_outputs(9703));
    layer2_outputs(4782) <= (layer1_outputs(9597)) xor (layer1_outputs(2011));
    layer2_outputs(4783) <= not((layer1_outputs(3237)) xor (layer1_outputs(4897)));
    layer2_outputs(4784) <= not(layer1_outputs(9672));
    layer2_outputs(4785) <= not(layer1_outputs(3857));
    layer2_outputs(4786) <= layer1_outputs(7005);
    layer2_outputs(4787) <= '0';
    layer2_outputs(4788) <= not(layer1_outputs(139));
    layer2_outputs(4789) <= layer1_outputs(1700);
    layer2_outputs(4790) <= layer1_outputs(9035);
    layer2_outputs(4791) <= not(layer1_outputs(5997));
    layer2_outputs(4792) <= not(layer1_outputs(7706));
    layer2_outputs(4793) <= layer1_outputs(136);
    layer2_outputs(4794) <= layer1_outputs(8390);
    layer2_outputs(4795) <= not(layer1_outputs(7223)) or (layer1_outputs(4100));
    layer2_outputs(4796) <= (layer1_outputs(1108)) or (layer1_outputs(7050));
    layer2_outputs(4797) <= not(layer1_outputs(7877));
    layer2_outputs(4798) <= not((layer1_outputs(9272)) or (layer1_outputs(2202)));
    layer2_outputs(4799) <= (layer1_outputs(7472)) and not (layer1_outputs(5650));
    layer2_outputs(4800) <= layer1_outputs(9454);
    layer2_outputs(4801) <= layer1_outputs(3548);
    layer2_outputs(4802) <= layer1_outputs(6775);
    layer2_outputs(4803) <= not(layer1_outputs(9498)) or (layer1_outputs(3898));
    layer2_outputs(4804) <= not(layer1_outputs(246));
    layer2_outputs(4805) <= not(layer1_outputs(5489));
    layer2_outputs(4806) <= layer1_outputs(2615);
    layer2_outputs(4807) <= layer1_outputs(8252);
    layer2_outputs(4808) <= (layer1_outputs(3929)) xor (layer1_outputs(8877));
    layer2_outputs(4809) <= (layer1_outputs(8851)) and not (layer1_outputs(6587));
    layer2_outputs(4810) <= not(layer1_outputs(7384)) or (layer1_outputs(1748));
    layer2_outputs(4811) <= not(layer1_outputs(6709));
    layer2_outputs(4812) <= not((layer1_outputs(3137)) and (layer1_outputs(9339)));
    layer2_outputs(4813) <= not(layer1_outputs(9375)) or (layer1_outputs(6953));
    layer2_outputs(4814) <= layer1_outputs(8960);
    layer2_outputs(4815) <= layer1_outputs(3391);
    layer2_outputs(4816) <= not(layer1_outputs(5540)) or (layer1_outputs(1348));
    layer2_outputs(4817) <= layer1_outputs(4649);
    layer2_outputs(4818) <= not(layer1_outputs(8941)) or (layer1_outputs(9291));
    layer2_outputs(4819) <= '1';
    layer2_outputs(4820) <= not(layer1_outputs(4376));
    layer2_outputs(4821) <= not(layer1_outputs(8624));
    layer2_outputs(4822) <= layer1_outputs(8750);
    layer2_outputs(4823) <= not((layer1_outputs(10229)) xor (layer1_outputs(3719)));
    layer2_outputs(4824) <= not((layer1_outputs(6403)) or (layer1_outputs(882)));
    layer2_outputs(4825) <= not(layer1_outputs(8843));
    layer2_outputs(4826) <= not(layer1_outputs(3792));
    layer2_outputs(4827) <= layer1_outputs(2801);
    layer2_outputs(4828) <= (layer1_outputs(9298)) xor (layer1_outputs(6018));
    layer2_outputs(4829) <= (layer1_outputs(36)) xor (layer1_outputs(9871));
    layer2_outputs(4830) <= layer1_outputs(9091);
    layer2_outputs(4831) <= not((layer1_outputs(6758)) and (layer1_outputs(6640)));
    layer2_outputs(4832) <= (layer1_outputs(6123)) and not (layer1_outputs(566));
    layer2_outputs(4833) <= layer1_outputs(2541);
    layer2_outputs(4834) <= not(layer1_outputs(5532));
    layer2_outputs(4835) <= layer1_outputs(104);
    layer2_outputs(4836) <= not(layer1_outputs(3526));
    layer2_outputs(4837) <= not(layer1_outputs(1779));
    layer2_outputs(4838) <= layer1_outputs(9360);
    layer2_outputs(4839) <= layer1_outputs(6285);
    layer2_outputs(4840) <= layer1_outputs(6361);
    layer2_outputs(4841) <= not(layer1_outputs(5618));
    layer2_outputs(4842) <= not(layer1_outputs(2462)) or (layer1_outputs(5781));
    layer2_outputs(4843) <= layer1_outputs(5273);
    layer2_outputs(4844) <= not(layer1_outputs(4071)) or (layer1_outputs(4972));
    layer2_outputs(4845) <= layer1_outputs(6028);
    layer2_outputs(4846) <= layer1_outputs(264);
    layer2_outputs(4847) <= layer1_outputs(3144);
    layer2_outputs(4848) <= '0';
    layer2_outputs(4849) <= not(layer1_outputs(8245));
    layer2_outputs(4850) <= layer1_outputs(8710);
    layer2_outputs(4851) <= not(layer1_outputs(1308)) or (layer1_outputs(8196));
    layer2_outputs(4852) <= (layer1_outputs(2723)) xor (layer1_outputs(5948));
    layer2_outputs(4853) <= not((layer1_outputs(3658)) or (layer1_outputs(3358)));
    layer2_outputs(4854) <= layer1_outputs(9129);
    layer2_outputs(4855) <= layer1_outputs(5007);
    layer2_outputs(4856) <= layer1_outputs(1107);
    layer2_outputs(4857) <= layer1_outputs(8132);
    layer2_outputs(4858) <= not(layer1_outputs(1182));
    layer2_outputs(4859) <= layer1_outputs(3891);
    layer2_outputs(4860) <= not(layer1_outputs(6965));
    layer2_outputs(4861) <= (layer1_outputs(488)) and not (layer1_outputs(9726));
    layer2_outputs(4862) <= not(layer1_outputs(9393));
    layer2_outputs(4863) <= not((layer1_outputs(5531)) xor (layer1_outputs(5891)));
    layer2_outputs(4864) <= not((layer1_outputs(6852)) xor (layer1_outputs(6181)));
    layer2_outputs(4865) <= not(layer1_outputs(87));
    layer2_outputs(4866) <= layer1_outputs(464);
    layer2_outputs(4867) <= (layer1_outputs(7334)) xor (layer1_outputs(7162));
    layer2_outputs(4868) <= not(layer1_outputs(10073));
    layer2_outputs(4869) <= not(layer1_outputs(4760));
    layer2_outputs(4870) <= not(layer1_outputs(3398));
    layer2_outputs(4871) <= not(layer1_outputs(7643)) or (layer1_outputs(2986));
    layer2_outputs(4872) <= not(layer1_outputs(10232));
    layer2_outputs(4873) <= not(layer1_outputs(3502));
    layer2_outputs(4874) <= '1';
    layer2_outputs(4875) <= layer1_outputs(7981);
    layer2_outputs(4876) <= not(layer1_outputs(9808));
    layer2_outputs(4877) <= layer1_outputs(5250);
    layer2_outputs(4878) <= (layer1_outputs(4186)) or (layer1_outputs(1066));
    layer2_outputs(4879) <= (layer1_outputs(3146)) and not (layer1_outputs(3249));
    layer2_outputs(4880) <= '0';
    layer2_outputs(4881) <= not(layer1_outputs(3087));
    layer2_outputs(4882) <= layer1_outputs(9434);
    layer2_outputs(4883) <= not(layer1_outputs(6398));
    layer2_outputs(4884) <= (layer1_outputs(7434)) or (layer1_outputs(938));
    layer2_outputs(4885) <= not(layer1_outputs(9793));
    layer2_outputs(4886) <= not(layer1_outputs(4501));
    layer2_outputs(4887) <= not(layer1_outputs(6087));
    layer2_outputs(4888) <= not(layer1_outputs(38));
    layer2_outputs(4889) <= layer1_outputs(2916);
    layer2_outputs(4890) <= not(layer1_outputs(4771));
    layer2_outputs(4891) <= not(layer1_outputs(5326));
    layer2_outputs(4892) <= not(layer1_outputs(5622));
    layer2_outputs(4893) <= layer1_outputs(5915);
    layer2_outputs(4894) <= layer1_outputs(868);
    layer2_outputs(4895) <= not(layer1_outputs(2346));
    layer2_outputs(4896) <= (layer1_outputs(5063)) and not (layer1_outputs(8137));
    layer2_outputs(4897) <= (layer1_outputs(2857)) xor (layer1_outputs(4361));
    layer2_outputs(4898) <= (layer1_outputs(4234)) or (layer1_outputs(7235));
    layer2_outputs(4899) <= not(layer1_outputs(9236));
    layer2_outputs(4900) <= layer1_outputs(9379);
    layer2_outputs(4901) <= not(layer1_outputs(9752));
    layer2_outputs(4902) <= not((layer1_outputs(2283)) or (layer1_outputs(2403)));
    layer2_outputs(4903) <= layer1_outputs(4704);
    layer2_outputs(4904) <= layer1_outputs(4972);
    layer2_outputs(4905) <= not(layer1_outputs(1156));
    layer2_outputs(4906) <= (layer1_outputs(309)) and not (layer1_outputs(8778));
    layer2_outputs(4907) <= not((layer1_outputs(4851)) and (layer1_outputs(3673)));
    layer2_outputs(4908) <= not((layer1_outputs(8007)) xor (layer1_outputs(9433)));
    layer2_outputs(4909) <= layer1_outputs(9866);
    layer2_outputs(4910) <= layer1_outputs(4517);
    layer2_outputs(4911) <= not(layer1_outputs(291)) or (layer1_outputs(9496));
    layer2_outputs(4912) <= not(layer1_outputs(70));
    layer2_outputs(4913) <= layer1_outputs(10218);
    layer2_outputs(4914) <= not(layer1_outputs(6907));
    layer2_outputs(4915) <= not(layer1_outputs(144));
    layer2_outputs(4916) <= layer1_outputs(8220);
    layer2_outputs(4917) <= not(layer1_outputs(9857));
    layer2_outputs(4918) <= not(layer1_outputs(6347));
    layer2_outputs(4919) <= not(layer1_outputs(5663));
    layer2_outputs(4920) <= (layer1_outputs(5283)) and not (layer1_outputs(7094));
    layer2_outputs(4921) <= not((layer1_outputs(4000)) and (layer1_outputs(1040)));
    layer2_outputs(4922) <= (layer1_outputs(4410)) and not (layer1_outputs(9591));
    layer2_outputs(4923) <= (layer1_outputs(2881)) and not (layer1_outputs(3753));
    layer2_outputs(4924) <= (layer1_outputs(6799)) and not (layer1_outputs(950));
    layer2_outputs(4925) <= (layer1_outputs(9975)) and not (layer1_outputs(8159));
    layer2_outputs(4926) <= layer1_outputs(6160);
    layer2_outputs(4927) <= not(layer1_outputs(9419));
    layer2_outputs(4928) <= not(layer1_outputs(9283));
    layer2_outputs(4929) <= (layer1_outputs(8703)) or (layer1_outputs(5163));
    layer2_outputs(4930) <= not((layer1_outputs(3210)) and (layer1_outputs(2538)));
    layer2_outputs(4931) <= not(layer1_outputs(6971)) or (layer1_outputs(7906));
    layer2_outputs(4932) <= not(layer1_outputs(3136));
    layer2_outputs(4933) <= not(layer1_outputs(8126)) or (layer1_outputs(132));
    layer2_outputs(4934) <= layer1_outputs(9640);
    layer2_outputs(4935) <= not(layer1_outputs(59)) or (layer1_outputs(1752));
    layer2_outputs(4936) <= not(layer1_outputs(6114)) or (layer1_outputs(4715));
    layer2_outputs(4937) <= not(layer1_outputs(1744));
    layer2_outputs(4938) <= (layer1_outputs(2848)) xor (layer1_outputs(9033));
    layer2_outputs(4939) <= not(layer1_outputs(1806));
    layer2_outputs(4940) <= (layer1_outputs(1648)) or (layer1_outputs(6562));
    layer2_outputs(4941) <= (layer1_outputs(4978)) xor (layer1_outputs(8481));
    layer2_outputs(4942) <= layer1_outputs(6383);
    layer2_outputs(4943) <= layer1_outputs(547);
    layer2_outputs(4944) <= layer1_outputs(7691);
    layer2_outputs(4945) <= not((layer1_outputs(987)) xor (layer1_outputs(8706)));
    layer2_outputs(4946) <= (layer1_outputs(6518)) or (layer1_outputs(2674));
    layer2_outputs(4947) <= not(layer1_outputs(7525));
    layer2_outputs(4948) <= layer1_outputs(5031);
    layer2_outputs(4949) <= not(layer1_outputs(5867)) or (layer1_outputs(762));
    layer2_outputs(4950) <= '0';
    layer2_outputs(4951) <= not(layer1_outputs(6547));
    layer2_outputs(4952) <= (layer1_outputs(9457)) and (layer1_outputs(8393));
    layer2_outputs(4953) <= '1';
    layer2_outputs(4954) <= layer1_outputs(6094);
    layer2_outputs(4955) <= (layer1_outputs(7277)) and not (layer1_outputs(3175));
    layer2_outputs(4956) <= not(layer1_outputs(421));
    layer2_outputs(4957) <= (layer1_outputs(90)) and not (layer1_outputs(2500));
    layer2_outputs(4958) <= (layer1_outputs(235)) and not (layer1_outputs(509));
    layer2_outputs(4959) <= not(layer1_outputs(8431)) or (layer1_outputs(5798));
    layer2_outputs(4960) <= not(layer1_outputs(1380)) or (layer1_outputs(1564));
    layer2_outputs(4961) <= (layer1_outputs(458)) and not (layer1_outputs(1740));
    layer2_outputs(4962) <= (layer1_outputs(6043)) and (layer1_outputs(8970));
    layer2_outputs(4963) <= not(layer1_outputs(1345)) or (layer1_outputs(4615));
    layer2_outputs(4964) <= not(layer1_outputs(6747));
    layer2_outputs(4965) <= not(layer1_outputs(586));
    layer2_outputs(4966) <= (layer1_outputs(8631)) and not (layer1_outputs(2825));
    layer2_outputs(4967) <= not(layer1_outputs(6961));
    layer2_outputs(4968) <= (layer1_outputs(9304)) and not (layer1_outputs(4872));
    layer2_outputs(4969) <= not(layer1_outputs(8418)) or (layer1_outputs(58));
    layer2_outputs(4970) <= layer1_outputs(4348);
    layer2_outputs(4971) <= not(layer1_outputs(6332));
    layer2_outputs(4972) <= layer1_outputs(8855);
    layer2_outputs(4973) <= layer1_outputs(6944);
    layer2_outputs(4974) <= layer1_outputs(4278);
    layer2_outputs(4975) <= layer1_outputs(5343);
    layer2_outputs(4976) <= layer1_outputs(6487);
    layer2_outputs(4977) <= not(layer1_outputs(1585));
    layer2_outputs(4978) <= not(layer1_outputs(915)) or (layer1_outputs(6105));
    layer2_outputs(4979) <= layer1_outputs(7575);
    layer2_outputs(4980) <= not(layer1_outputs(7422));
    layer2_outputs(4981) <= not((layer1_outputs(1714)) xor (layer1_outputs(1697)));
    layer2_outputs(4982) <= layer1_outputs(1764);
    layer2_outputs(4983) <= not(layer1_outputs(5822)) or (layer1_outputs(8180));
    layer2_outputs(4984) <= layer1_outputs(10225);
    layer2_outputs(4985) <= (layer1_outputs(4406)) xor (layer1_outputs(439));
    layer2_outputs(4986) <= (layer1_outputs(9722)) and not (layer1_outputs(1708));
    layer2_outputs(4987) <= not(layer1_outputs(7901));
    layer2_outputs(4988) <= layer1_outputs(8479);
    layer2_outputs(4989) <= not((layer1_outputs(6250)) xor (layer1_outputs(6443)));
    layer2_outputs(4990) <= not(layer1_outputs(1220));
    layer2_outputs(4991) <= not((layer1_outputs(4921)) or (layer1_outputs(9381)));
    layer2_outputs(4992) <= (layer1_outputs(7840)) or (layer1_outputs(1613));
    layer2_outputs(4993) <= layer1_outputs(3316);
    layer2_outputs(4994) <= not(layer1_outputs(5212)) or (layer1_outputs(10046));
    layer2_outputs(4995) <= not((layer1_outputs(9639)) xor (layer1_outputs(6152)));
    layer2_outputs(4996) <= (layer1_outputs(6699)) xor (layer1_outputs(1360));
    layer2_outputs(4997) <= (layer1_outputs(1609)) or (layer1_outputs(1028));
    layer2_outputs(4998) <= layer1_outputs(7222);
    layer2_outputs(4999) <= (layer1_outputs(10060)) and (layer1_outputs(9021));
    layer2_outputs(5000) <= layer1_outputs(1975);
    layer2_outputs(5001) <= not(layer1_outputs(4433));
    layer2_outputs(5002) <= not(layer1_outputs(824));
    layer2_outputs(5003) <= not((layer1_outputs(4506)) or (layer1_outputs(3971)));
    layer2_outputs(5004) <= (layer1_outputs(7463)) and not (layer1_outputs(9140));
    layer2_outputs(5005) <= (layer1_outputs(5624)) xor (layer1_outputs(2628));
    layer2_outputs(5006) <= not(layer1_outputs(5157));
    layer2_outputs(5007) <= not(layer1_outputs(1388));
    layer2_outputs(5008) <= not((layer1_outputs(6915)) or (layer1_outputs(104)));
    layer2_outputs(5009) <= not((layer1_outputs(6887)) and (layer1_outputs(1298)));
    layer2_outputs(5010) <= not(layer1_outputs(3250));
    layer2_outputs(5011) <= layer1_outputs(8741);
    layer2_outputs(5012) <= not(layer1_outputs(9312));
    layer2_outputs(5013) <= (layer1_outputs(1896)) and not (layer1_outputs(3892));
    layer2_outputs(5014) <= (layer1_outputs(6815)) xor (layer1_outputs(4894));
    layer2_outputs(5015) <= layer1_outputs(7779);
    layer2_outputs(5016) <= not(layer1_outputs(6179));
    layer2_outputs(5017) <= not(layer1_outputs(9317));
    layer2_outputs(5018) <= not(layer1_outputs(9567)) or (layer1_outputs(5739));
    layer2_outputs(5019) <= not(layer1_outputs(4084));
    layer2_outputs(5020) <= not(layer1_outputs(9780));
    layer2_outputs(5021) <= (layer1_outputs(6710)) and (layer1_outputs(1932));
    layer2_outputs(5022) <= layer1_outputs(11);
    layer2_outputs(5023) <= layer1_outputs(7509);
    layer2_outputs(5024) <= (layer1_outputs(1182)) and not (layer1_outputs(9579));
    layer2_outputs(5025) <= layer1_outputs(7325);
    layer2_outputs(5026) <= layer1_outputs(6765);
    layer2_outputs(5027) <= layer1_outputs(3675);
    layer2_outputs(5028) <= (layer1_outputs(858)) or (layer1_outputs(9564));
    layer2_outputs(5029) <= layer1_outputs(5193);
    layer2_outputs(5030) <= not((layer1_outputs(204)) and (layer1_outputs(682)));
    layer2_outputs(5031) <= not(layer1_outputs(9094));
    layer2_outputs(5032) <= layer1_outputs(3298);
    layer2_outputs(5033) <= not(layer1_outputs(6888)) or (layer1_outputs(9231));
    layer2_outputs(5034) <= (layer1_outputs(7574)) and not (layer1_outputs(1545));
    layer2_outputs(5035) <= not(layer1_outputs(7252));
    layer2_outputs(5036) <= not((layer1_outputs(5240)) or (layer1_outputs(10057)));
    layer2_outputs(5037) <= (layer1_outputs(6947)) xor (layer1_outputs(334));
    layer2_outputs(5038) <= (layer1_outputs(5813)) and not (layer1_outputs(5521));
    layer2_outputs(5039) <= not(layer1_outputs(10092));
    layer2_outputs(5040) <= not(layer1_outputs(1343));
    layer2_outputs(5041) <= (layer1_outputs(2407)) and not (layer1_outputs(3262));
    layer2_outputs(5042) <= not(layer1_outputs(4829));
    layer2_outputs(5043) <= not(layer1_outputs(7913)) or (layer1_outputs(5224));
    layer2_outputs(5044) <= not(layer1_outputs(8705));
    layer2_outputs(5045) <= not(layer1_outputs(4257)) or (layer1_outputs(6196));
    layer2_outputs(5046) <= layer1_outputs(8937);
    layer2_outputs(5047) <= layer1_outputs(9628);
    layer2_outputs(5048) <= layer1_outputs(6463);
    layer2_outputs(5049) <= layer1_outputs(2591);
    layer2_outputs(5050) <= (layer1_outputs(9212)) xor (layer1_outputs(4581));
    layer2_outputs(5051) <= layer1_outputs(5742);
    layer2_outputs(5052) <= (layer1_outputs(7646)) and not (layer1_outputs(4475));
    layer2_outputs(5053) <= not(layer1_outputs(10105));
    layer2_outputs(5054) <= layer1_outputs(8284);
    layer2_outputs(5055) <= (layer1_outputs(2554)) and (layer1_outputs(7953));
    layer2_outputs(5056) <= layer1_outputs(2063);
    layer2_outputs(5057) <= layer1_outputs(3692);
    layer2_outputs(5058) <= layer1_outputs(8399);
    layer2_outputs(5059) <= (layer1_outputs(4927)) and not (layer1_outputs(8628));
    layer2_outputs(5060) <= not((layer1_outputs(2799)) and (layer1_outputs(3058)));
    layer2_outputs(5061) <= not((layer1_outputs(2344)) or (layer1_outputs(5866)));
    layer2_outputs(5062) <= not((layer1_outputs(3212)) or (layer1_outputs(1364)));
    layer2_outputs(5063) <= (layer1_outputs(10028)) xor (layer1_outputs(1154));
    layer2_outputs(5064) <= layer1_outputs(5182);
    layer2_outputs(5065) <= not((layer1_outputs(522)) and (layer1_outputs(2669)));
    layer2_outputs(5066) <= layer1_outputs(5768);
    layer2_outputs(5067) <= not((layer1_outputs(3633)) or (layer1_outputs(4913)));
    layer2_outputs(5068) <= not(layer1_outputs(191));
    layer2_outputs(5069) <= layer1_outputs(231);
    layer2_outputs(5070) <= layer1_outputs(7010);
    layer2_outputs(5071) <= (layer1_outputs(1133)) or (layer1_outputs(910));
    layer2_outputs(5072) <= not((layer1_outputs(7903)) xor (layer1_outputs(4238)));
    layer2_outputs(5073) <= not(layer1_outputs(4225));
    layer2_outputs(5074) <= layer1_outputs(2331);
    layer2_outputs(5075) <= layer1_outputs(6822);
    layer2_outputs(5076) <= not((layer1_outputs(676)) or (layer1_outputs(4820)));
    layer2_outputs(5077) <= not(layer1_outputs(3954));
    layer2_outputs(5078) <= layer1_outputs(9207);
    layer2_outputs(5079) <= not((layer1_outputs(5581)) xor (layer1_outputs(6629)));
    layer2_outputs(5080) <= not(layer1_outputs(4381)) or (layer1_outputs(7243));
    layer2_outputs(5081) <= not(layer1_outputs(3737));
    layer2_outputs(5082) <= layer1_outputs(1953);
    layer2_outputs(5083) <= not(layer1_outputs(4941));
    layer2_outputs(5084) <= layer1_outputs(1719);
    layer2_outputs(5085) <= not((layer1_outputs(9307)) or (layer1_outputs(2522)));
    layer2_outputs(5086) <= not((layer1_outputs(10092)) or (layer1_outputs(3259)));
    layer2_outputs(5087) <= layer1_outputs(1128);
    layer2_outputs(5088) <= (layer1_outputs(1076)) and not (layer1_outputs(4213));
    layer2_outputs(5089) <= layer1_outputs(453);
    layer2_outputs(5090) <= not(layer1_outputs(7437)) or (layer1_outputs(8390));
    layer2_outputs(5091) <= (layer1_outputs(2921)) xor (layer1_outputs(4018));
    layer2_outputs(5092) <= (layer1_outputs(908)) and not (layer1_outputs(1023));
    layer2_outputs(5093) <= not(layer1_outputs(7945));
    layer2_outputs(5094) <= not(layer1_outputs(4621));
    layer2_outputs(5095) <= not(layer1_outputs(3460)) or (layer1_outputs(3212));
    layer2_outputs(5096) <= layer1_outputs(501);
    layer2_outputs(5097) <= not((layer1_outputs(7086)) and (layer1_outputs(9617)));
    layer2_outputs(5098) <= layer1_outputs(6054);
    layer2_outputs(5099) <= not((layer1_outputs(9718)) xor (layer1_outputs(1328)));
    layer2_outputs(5100) <= layer1_outputs(9403);
    layer2_outputs(5101) <= not(layer1_outputs(5021));
    layer2_outputs(5102) <= not(layer1_outputs(9891));
    layer2_outputs(5103) <= (layer1_outputs(4984)) and not (layer1_outputs(8434));
    layer2_outputs(5104) <= (layer1_outputs(4896)) and not (layer1_outputs(2392));
    layer2_outputs(5105) <= not(layer1_outputs(2690));
    layer2_outputs(5106) <= (layer1_outputs(6383)) or (layer1_outputs(5952));
    layer2_outputs(5107) <= layer1_outputs(6502);
    layer2_outputs(5108) <= (layer1_outputs(6591)) and not (layer1_outputs(7675));
    layer2_outputs(5109) <= not((layer1_outputs(778)) xor (layer1_outputs(967)));
    layer2_outputs(5110) <= layer1_outputs(9234);
    layer2_outputs(5111) <= (layer1_outputs(4502)) or (layer1_outputs(1629));
    layer2_outputs(5112) <= (layer1_outputs(5676)) xor (layer1_outputs(632));
    layer2_outputs(5113) <= not(layer1_outputs(2187)) or (layer1_outputs(564));
    layer2_outputs(5114) <= not(layer1_outputs(6602)) or (layer1_outputs(37));
    layer2_outputs(5115) <= not((layer1_outputs(5265)) xor (layer1_outputs(9734)));
    layer2_outputs(5116) <= not(layer1_outputs(3253));
    layer2_outputs(5117) <= not(layer1_outputs(8303));
    layer2_outputs(5118) <= not((layer1_outputs(2760)) or (layer1_outputs(3741)));
    layer2_outputs(5119) <= layer1_outputs(2192);
    layer2_outputs(5120) <= not(layer1_outputs(10013));
    layer2_outputs(5121) <= not(layer1_outputs(9539)) or (layer1_outputs(6934));
    layer2_outputs(5122) <= layer1_outputs(4409);
    layer2_outputs(5123) <= not((layer1_outputs(716)) and (layer1_outputs(3812)));
    layer2_outputs(5124) <= (layer1_outputs(10226)) or (layer1_outputs(864));
    layer2_outputs(5125) <= layer1_outputs(5548);
    layer2_outputs(5126) <= (layer1_outputs(577)) xor (layer1_outputs(8292));
    layer2_outputs(5127) <= not((layer1_outputs(8513)) and (layer1_outputs(3517)));
    layer2_outputs(5128) <= not((layer1_outputs(4756)) or (layer1_outputs(3248)));
    layer2_outputs(5129) <= (layer1_outputs(4510)) xor (layer1_outputs(2605));
    layer2_outputs(5130) <= layer1_outputs(358);
    layer2_outputs(5131) <= (layer1_outputs(6090)) and not (layer1_outputs(9700));
    layer2_outputs(5132) <= (layer1_outputs(5302)) or (layer1_outputs(2211));
    layer2_outputs(5133) <= layer1_outputs(4967);
    layer2_outputs(5134) <= not((layer1_outputs(6889)) xor (layer1_outputs(1481)));
    layer2_outputs(5135) <= layer1_outputs(9957);
    layer2_outputs(5136) <= not(layer1_outputs(3348));
    layer2_outputs(5137) <= not(layer1_outputs(10029));
    layer2_outputs(5138) <= layer1_outputs(6180);
    layer2_outputs(5139) <= not(layer1_outputs(6261));
    layer2_outputs(5140) <= not(layer1_outputs(2464));
    layer2_outputs(5141) <= layer1_outputs(4885);
    layer2_outputs(5142) <= layer1_outputs(5529);
    layer2_outputs(5143) <= not(layer1_outputs(5866));
    layer2_outputs(5144) <= (layer1_outputs(320)) and not (layer1_outputs(1248));
    layer2_outputs(5145) <= not(layer1_outputs(9981));
    layer2_outputs(5146) <= not((layer1_outputs(2230)) and (layer1_outputs(428)));
    layer2_outputs(5147) <= not(layer1_outputs(31)) or (layer1_outputs(6619));
    layer2_outputs(5148) <= not(layer1_outputs(6223));
    layer2_outputs(5149) <= layer1_outputs(5368);
    layer2_outputs(5150) <= layer1_outputs(3986);
    layer2_outputs(5151) <= layer1_outputs(2031);
    layer2_outputs(5152) <= layer1_outputs(3938);
    layer2_outputs(5153) <= not((layer1_outputs(445)) or (layer1_outputs(8739)));
    layer2_outputs(5154) <= layer1_outputs(5633);
    layer2_outputs(5155) <= (layer1_outputs(8808)) and not (layer1_outputs(6541));
    layer2_outputs(5156) <= layer1_outputs(9179);
    layer2_outputs(5157) <= not(layer1_outputs(7124)) or (layer1_outputs(1848));
    layer2_outputs(5158) <= not(layer1_outputs(1906));
    layer2_outputs(5159) <= layer1_outputs(6649);
    layer2_outputs(5160) <= layer1_outputs(9792);
    layer2_outputs(5161) <= (layer1_outputs(10137)) xor (layer1_outputs(6554));
    layer2_outputs(5162) <= not(layer1_outputs(5191));
    layer2_outputs(5163) <= layer1_outputs(9971);
    layer2_outputs(5164) <= not(layer1_outputs(4511));
    layer2_outputs(5165) <= (layer1_outputs(8005)) xor (layer1_outputs(2044));
    layer2_outputs(5166) <= not(layer1_outputs(4405));
    layer2_outputs(5167) <= not(layer1_outputs(8649));
    layer2_outputs(5168) <= (layer1_outputs(10233)) xor (layer1_outputs(3426));
    layer2_outputs(5169) <= layer1_outputs(1197);
    layer2_outputs(5170) <= (layer1_outputs(9589)) and not (layer1_outputs(1196));
    layer2_outputs(5171) <= (layer1_outputs(3710)) or (layer1_outputs(1604));
    layer2_outputs(5172) <= '1';
    layer2_outputs(5173) <= not(layer1_outputs(3652)) or (layer1_outputs(7351));
    layer2_outputs(5174) <= (layer1_outputs(4352)) or (layer1_outputs(1136));
    layer2_outputs(5175) <= not(layer1_outputs(8550)) or (layer1_outputs(10212));
    layer2_outputs(5176) <= not((layer1_outputs(8052)) and (layer1_outputs(7835)));
    layer2_outputs(5177) <= not(layer1_outputs(7976));
    layer2_outputs(5178) <= '0';
    layer2_outputs(5179) <= not((layer1_outputs(4624)) xor (layer1_outputs(4754)));
    layer2_outputs(5180) <= layer1_outputs(8122);
    layer2_outputs(5181) <= layer1_outputs(1921);
    layer2_outputs(5182) <= not(layer1_outputs(9383));
    layer2_outputs(5183) <= not((layer1_outputs(2528)) or (layer1_outputs(7555)));
    layer2_outputs(5184) <= (layer1_outputs(9406)) and (layer1_outputs(391));
    layer2_outputs(5185) <= not(layer1_outputs(3545));
    layer2_outputs(5186) <= not(layer1_outputs(5612));
    layer2_outputs(5187) <= not(layer1_outputs(829));
    layer2_outputs(5188) <= (layer1_outputs(4572)) and not (layer1_outputs(7147));
    layer2_outputs(5189) <= layer1_outputs(2686);
    layer2_outputs(5190) <= not(layer1_outputs(2700));
    layer2_outputs(5191) <= layer1_outputs(7937);
    layer2_outputs(5192) <= not(layer1_outputs(3062));
    layer2_outputs(5193) <= '1';
    layer2_outputs(5194) <= not(layer1_outputs(9453)) or (layer1_outputs(9146));
    layer2_outputs(5195) <= not((layer1_outputs(7178)) or (layer1_outputs(6362)));
    layer2_outputs(5196) <= layer1_outputs(351);
    layer2_outputs(5197) <= not(layer1_outputs(476)) or (layer1_outputs(9584));
    layer2_outputs(5198) <= (layer1_outputs(1)) or (layer1_outputs(5623));
    layer2_outputs(5199) <= (layer1_outputs(398)) and not (layer1_outputs(2200));
    layer2_outputs(5200) <= not(layer1_outputs(9762));
    layer2_outputs(5201) <= not((layer1_outputs(5813)) and (layer1_outputs(6050)));
    layer2_outputs(5202) <= layer1_outputs(4348);
    layer2_outputs(5203) <= not(layer1_outputs(8974)) or (layer1_outputs(5748));
    layer2_outputs(5204) <= (layer1_outputs(3596)) xor (layer1_outputs(8016));
    layer2_outputs(5205) <= layer1_outputs(2647);
    layer2_outputs(5206) <= (layer1_outputs(8496)) xor (layer1_outputs(5970));
    layer2_outputs(5207) <= layer1_outputs(7497);
    layer2_outputs(5208) <= not(layer1_outputs(9134)) or (layer1_outputs(4906));
    layer2_outputs(5209) <= layer1_outputs(5076);
    layer2_outputs(5210) <= not(layer1_outputs(1985));
    layer2_outputs(5211) <= not(layer1_outputs(1004));
    layer2_outputs(5212) <= layer1_outputs(6729);
    layer2_outputs(5213) <= layer1_outputs(440);
    layer2_outputs(5214) <= '1';
    layer2_outputs(5215) <= not(layer1_outputs(5446));
    layer2_outputs(5216) <= not(layer1_outputs(6685));
    layer2_outputs(5217) <= not(layer1_outputs(9654)) or (layer1_outputs(6509));
    layer2_outputs(5218) <= layer1_outputs(5753);
    layer2_outputs(5219) <= not(layer1_outputs(4455)) or (layer1_outputs(2800));
    layer2_outputs(5220) <= not(layer1_outputs(6647));
    layer2_outputs(5221) <= (layer1_outputs(8732)) or (layer1_outputs(1944));
    layer2_outputs(5222) <= (layer1_outputs(8593)) and (layer1_outputs(5154));
    layer2_outputs(5223) <= layer1_outputs(4114);
    layer2_outputs(5224) <= (layer1_outputs(4631)) and (layer1_outputs(9494));
    layer2_outputs(5225) <= (layer1_outputs(2305)) and (layer1_outputs(2758));
    layer2_outputs(5226) <= not((layer1_outputs(9595)) and (layer1_outputs(9142)));
    layer2_outputs(5227) <= (layer1_outputs(3477)) xor (layer1_outputs(4192));
    layer2_outputs(5228) <= not((layer1_outputs(6831)) and (layer1_outputs(4724)));
    layer2_outputs(5229) <= (layer1_outputs(2772)) xor (layer1_outputs(5709));
    layer2_outputs(5230) <= (layer1_outputs(8049)) or (layer1_outputs(4864));
    layer2_outputs(5231) <= layer1_outputs(7511);
    layer2_outputs(5232) <= not(layer1_outputs(982));
    layer2_outputs(5233) <= not((layer1_outputs(6782)) or (layer1_outputs(6107)));
    layer2_outputs(5234) <= (layer1_outputs(8535)) and not (layer1_outputs(1138));
    layer2_outputs(5235) <= not(layer1_outputs(2916));
    layer2_outputs(5236) <= (layer1_outputs(6637)) and (layer1_outputs(3990));
    layer2_outputs(5237) <= layer1_outputs(9952);
    layer2_outputs(5238) <= layer1_outputs(5927);
    layer2_outputs(5239) <= layer1_outputs(2524);
    layer2_outputs(5240) <= not(layer1_outputs(7044));
    layer2_outputs(5241) <= layer1_outputs(3100);
    layer2_outputs(5242) <= '0';
    layer2_outputs(5243) <= (layer1_outputs(2859)) and not (layer1_outputs(6644));
    layer2_outputs(5244) <= (layer1_outputs(5085)) xor (layer1_outputs(9830));
    layer2_outputs(5245) <= layer1_outputs(5176);
    layer2_outputs(5246) <= layer1_outputs(6055);
    layer2_outputs(5247) <= not(layer1_outputs(2869));
    layer2_outputs(5248) <= (layer1_outputs(8831)) and not (layer1_outputs(9786));
    layer2_outputs(5249) <= (layer1_outputs(8415)) and not (layer1_outputs(1916));
    layer2_outputs(5250) <= not(layer1_outputs(10033));
    layer2_outputs(5251) <= not(layer1_outputs(1794));
    layer2_outputs(5252) <= (layer1_outputs(3903)) and not (layer1_outputs(9999));
    layer2_outputs(5253) <= not((layer1_outputs(4834)) or (layer1_outputs(3433)));
    layer2_outputs(5254) <= layer1_outputs(3367);
    layer2_outputs(5255) <= not(layer1_outputs(9437)) or (layer1_outputs(4788));
    layer2_outputs(5256) <= (layer1_outputs(7297)) and (layer1_outputs(8067));
    layer2_outputs(5257) <= (layer1_outputs(4161)) and not (layer1_outputs(5022));
    layer2_outputs(5258) <= layer1_outputs(9233);
    layer2_outputs(5259) <= not(layer1_outputs(1231));
    layer2_outputs(5260) <= (layer1_outputs(1341)) or (layer1_outputs(8525));
    layer2_outputs(5261) <= not((layer1_outputs(7262)) xor (layer1_outputs(8066)));
    layer2_outputs(5262) <= (layer1_outputs(7667)) or (layer1_outputs(8554));
    layer2_outputs(5263) <= layer1_outputs(4112);
    layer2_outputs(5264) <= (layer1_outputs(1325)) xor (layer1_outputs(6656));
    layer2_outputs(5265) <= layer1_outputs(7175);
    layer2_outputs(5266) <= layer1_outputs(6452);
    layer2_outputs(5267) <= (layer1_outputs(4580)) and not (layer1_outputs(8697));
    layer2_outputs(5268) <= not(layer1_outputs(7670)) or (layer1_outputs(5953));
    layer2_outputs(5269) <= not(layer1_outputs(4359));
    layer2_outputs(5270) <= not(layer1_outputs(9280)) or (layer1_outputs(8503));
    layer2_outputs(5271) <= not((layer1_outputs(1630)) xor (layer1_outputs(6415)));
    layer2_outputs(5272) <= not(layer1_outputs(6020)) or (layer1_outputs(6964));
    layer2_outputs(5273) <= layer1_outputs(5592);
    layer2_outputs(5274) <= layer1_outputs(7608);
    layer2_outputs(5275) <= layer1_outputs(8534);
    layer2_outputs(5276) <= layer1_outputs(2499);
    layer2_outputs(5277) <= '1';
    layer2_outputs(5278) <= layer1_outputs(298);
    layer2_outputs(5279) <= (layer1_outputs(5535)) xor (layer1_outputs(1812));
    layer2_outputs(5280) <= not(layer1_outputs(3773));
    layer2_outputs(5281) <= not(layer1_outputs(9184)) or (layer1_outputs(4645));
    layer2_outputs(5282) <= not(layer1_outputs(8543));
    layer2_outputs(5283) <= not((layer1_outputs(6211)) or (layer1_outputs(8315)));
    layer2_outputs(5284) <= not((layer1_outputs(5292)) and (layer1_outputs(3427)));
    layer2_outputs(5285) <= (layer1_outputs(3517)) and not (layer1_outputs(6214));
    layer2_outputs(5286) <= not((layer1_outputs(432)) and (layer1_outputs(703)));
    layer2_outputs(5287) <= not(layer1_outputs(7787));
    layer2_outputs(5288) <= (layer1_outputs(836)) and not (layer1_outputs(6504));
    layer2_outputs(5289) <= not(layer1_outputs(8202));
    layer2_outputs(5290) <= layer1_outputs(6341);
    layer2_outputs(5291) <= layer1_outputs(4646);
    layer2_outputs(5292) <= (layer1_outputs(3731)) xor (layer1_outputs(719));
    layer2_outputs(5293) <= not((layer1_outputs(6954)) xor (layer1_outputs(997)));
    layer2_outputs(5294) <= not(layer1_outputs(9266));
    layer2_outputs(5295) <= layer1_outputs(8707);
    layer2_outputs(5296) <= not(layer1_outputs(2887));
    layer2_outputs(5297) <= layer1_outputs(1251);
    layer2_outputs(5298) <= layer1_outputs(4940);
    layer2_outputs(5299) <= (layer1_outputs(8593)) xor (layer1_outputs(5421));
    layer2_outputs(5300) <= not(layer1_outputs(8182));
    layer2_outputs(5301) <= not(layer1_outputs(4618)) or (layer1_outputs(5635));
    layer2_outputs(5302) <= layer1_outputs(9117);
    layer2_outputs(5303) <= layer1_outputs(2884);
    layer2_outputs(5304) <= (layer1_outputs(9082)) or (layer1_outputs(7985));
    layer2_outputs(5305) <= (layer1_outputs(5877)) xor (layer1_outputs(9519));
    layer2_outputs(5306) <= not((layer1_outputs(6790)) and (layer1_outputs(8466)));
    layer2_outputs(5307) <= (layer1_outputs(5473)) xor (layer1_outputs(1844));
    layer2_outputs(5308) <= not(layer1_outputs(1835));
    layer2_outputs(5309) <= not(layer1_outputs(6306));
    layer2_outputs(5310) <= layer1_outputs(6797);
    layer2_outputs(5311) <= not(layer1_outputs(6201));
    layer2_outputs(5312) <= not(layer1_outputs(1211));
    layer2_outputs(5313) <= layer1_outputs(2420);
    layer2_outputs(5314) <= not(layer1_outputs(2613));
    layer2_outputs(5315) <= not((layer1_outputs(5865)) or (layer1_outputs(6340)));
    layer2_outputs(5316) <= not((layer1_outputs(6003)) xor (layer1_outputs(3474)));
    layer2_outputs(5317) <= not(layer1_outputs(9684));
    layer2_outputs(5318) <= not((layer1_outputs(9868)) xor (layer1_outputs(7069)));
    layer2_outputs(5319) <= (layer1_outputs(592)) xor (layer1_outputs(1272));
    layer2_outputs(5320) <= layer1_outputs(8731);
    layer2_outputs(5321) <= (layer1_outputs(2749)) and not (layer1_outputs(4674));
    layer2_outputs(5322) <= layer1_outputs(9424);
    layer2_outputs(5323) <= layer1_outputs(397);
    layer2_outputs(5324) <= layer1_outputs(5510);
    layer2_outputs(5325) <= not((layer1_outputs(3028)) xor (layer1_outputs(5070)));
    layer2_outputs(5326) <= not(layer1_outputs(2681));
    layer2_outputs(5327) <= not(layer1_outputs(5363));
    layer2_outputs(5328) <= layer1_outputs(9088);
    layer2_outputs(5329) <= not((layer1_outputs(621)) and (layer1_outputs(9835)));
    layer2_outputs(5330) <= not(layer1_outputs(7451));
    layer2_outputs(5331) <= layer1_outputs(6826);
    layer2_outputs(5332) <= not(layer1_outputs(10191)) or (layer1_outputs(10136));
    layer2_outputs(5333) <= layer1_outputs(1676);
    layer2_outputs(5334) <= layer1_outputs(7711);
    layer2_outputs(5335) <= layer1_outputs(4942);
    layer2_outputs(5336) <= not((layer1_outputs(9594)) or (layer1_outputs(9458)));
    layer2_outputs(5337) <= not(layer1_outputs(3999));
    layer2_outputs(5338) <= not(layer1_outputs(517)) or (layer1_outputs(9605));
    layer2_outputs(5339) <= not(layer1_outputs(7022)) or (layer1_outputs(4295));
    layer2_outputs(5340) <= not(layer1_outputs(6843));
    layer2_outputs(5341) <= not(layer1_outputs(7089)) or (layer1_outputs(5195));
    layer2_outputs(5342) <= not(layer1_outputs(2190));
    layer2_outputs(5343) <= not(layer1_outputs(7982)) or (layer1_outputs(5505));
    layer2_outputs(5344) <= not((layer1_outputs(10171)) xor (layer1_outputs(9799)));
    layer2_outputs(5345) <= not(layer1_outputs(1822)) or (layer1_outputs(3780));
    layer2_outputs(5346) <= layer1_outputs(6251);
    layer2_outputs(5347) <= not(layer1_outputs(4890));
    layer2_outputs(5348) <= not(layer1_outputs(5275));
    layer2_outputs(5349) <= not((layer1_outputs(9460)) or (layer1_outputs(5923)));
    layer2_outputs(5350) <= layer1_outputs(5193);
    layer2_outputs(5351) <= layer1_outputs(6884);
    layer2_outputs(5352) <= not(layer1_outputs(6568));
    layer2_outputs(5353) <= not((layer1_outputs(3330)) and (layer1_outputs(5570)));
    layer2_outputs(5354) <= '0';
    layer2_outputs(5355) <= layer1_outputs(3190);
    layer2_outputs(5356) <= not(layer1_outputs(3290));
    layer2_outputs(5357) <= layer1_outputs(8655);
    layer2_outputs(5358) <= not(layer1_outputs(8086));
    layer2_outputs(5359) <= not(layer1_outputs(5189));
    layer2_outputs(5360) <= '0';
    layer2_outputs(5361) <= not(layer1_outputs(1110));
    layer2_outputs(5362) <= not(layer1_outputs(3515));
    layer2_outputs(5363) <= not(layer1_outputs(912));
    layer2_outputs(5364) <= layer1_outputs(9540);
    layer2_outputs(5365) <= layer1_outputs(923);
    layer2_outputs(5366) <= not(layer1_outputs(6444)) or (layer1_outputs(8687));
    layer2_outputs(5367) <= (layer1_outputs(2880)) and (layer1_outputs(8596));
    layer2_outputs(5368) <= not((layer1_outputs(9523)) or (layer1_outputs(8553)));
    layer2_outputs(5369) <= layer1_outputs(9863);
    layer2_outputs(5370) <= layer1_outputs(2416);
    layer2_outputs(5371) <= not(layer1_outputs(2904)) or (layer1_outputs(4066));
    layer2_outputs(5372) <= not(layer1_outputs(587));
    layer2_outputs(5373) <= not((layer1_outputs(267)) and (layer1_outputs(1691)));
    layer2_outputs(5374) <= (layer1_outputs(2734)) xor (layer1_outputs(10201));
    layer2_outputs(5375) <= not(layer1_outputs(6988));
    layer2_outputs(5376) <= not(layer1_outputs(6253));
    layer2_outputs(5377) <= not(layer1_outputs(8456)) or (layer1_outputs(10211));
    layer2_outputs(5378) <= not((layer1_outputs(9016)) xor (layer1_outputs(8632)));
    layer2_outputs(5379) <= layer1_outputs(408);
    layer2_outputs(5380) <= layer1_outputs(8560);
    layer2_outputs(5381) <= not(layer1_outputs(2564));
    layer2_outputs(5382) <= layer1_outputs(1437);
    layer2_outputs(5383) <= not(layer1_outputs(1448));
    layer2_outputs(5384) <= '0';
    layer2_outputs(5385) <= layer1_outputs(343);
    layer2_outputs(5386) <= layer1_outputs(6237);
    layer2_outputs(5387) <= not(layer1_outputs(2934));
    layer2_outputs(5388) <= not((layer1_outputs(2135)) and (layer1_outputs(8710)));
    layer2_outputs(5389) <= (layer1_outputs(1244)) or (layer1_outputs(6496));
    layer2_outputs(5390) <= (layer1_outputs(7140)) xor (layer1_outputs(5128));
    layer2_outputs(5391) <= '1';
    layer2_outputs(5392) <= layer1_outputs(4067);
    layer2_outputs(5393) <= (layer1_outputs(9894)) and (layer1_outputs(9067));
    layer2_outputs(5394) <= not(layer1_outputs(1198));
    layer2_outputs(5395) <= not(layer1_outputs(9112));
    layer2_outputs(5396) <= not(layer1_outputs(5108)) or (layer1_outputs(3068));
    layer2_outputs(5397) <= not(layer1_outputs(7775));
    layer2_outputs(5398) <= not((layer1_outputs(1080)) or (layer1_outputs(7746)));
    layer2_outputs(5399) <= layer1_outputs(7385);
    layer2_outputs(5400) <= not((layer1_outputs(4567)) xor (layer1_outputs(1000)));
    layer2_outputs(5401) <= not(layer1_outputs(6550));
    layer2_outputs(5402) <= not((layer1_outputs(9968)) xor (layer1_outputs(6251)));
    layer2_outputs(5403) <= not(layer1_outputs(9632)) or (layer1_outputs(114));
    layer2_outputs(5404) <= (layer1_outputs(2756)) and not (layer1_outputs(553));
    layer2_outputs(5405) <= not((layer1_outputs(8204)) and (layer1_outputs(9890)));
    layer2_outputs(5406) <= (layer1_outputs(7980)) xor (layer1_outputs(4220));
    layer2_outputs(5407) <= (layer1_outputs(6831)) and not (layer1_outputs(6629));
    layer2_outputs(5408) <= layer1_outputs(3817);
    layer2_outputs(5409) <= not((layer1_outputs(4971)) xor (layer1_outputs(9322)));
    layer2_outputs(5410) <= '0';
    layer2_outputs(5411) <= not(layer1_outputs(3577));
    layer2_outputs(5412) <= (layer1_outputs(8454)) and not (layer1_outputs(8097));
    layer2_outputs(5413) <= not(layer1_outputs(2886));
    layer2_outputs(5414) <= not(layer1_outputs(6701));
    layer2_outputs(5415) <= not(layer1_outputs(1544)) or (layer1_outputs(8070));
    layer2_outputs(5416) <= (layer1_outputs(3820)) and not (layer1_outputs(2815));
    layer2_outputs(5417) <= not(layer1_outputs(9573));
    layer2_outputs(5418) <= not(layer1_outputs(1377));
    layer2_outputs(5419) <= layer1_outputs(1847);
    layer2_outputs(5420) <= '0';
    layer2_outputs(5421) <= layer1_outputs(6256);
    layer2_outputs(5422) <= not(layer1_outputs(987));
    layer2_outputs(5423) <= not(layer1_outputs(6595)) or (layer1_outputs(4070));
    layer2_outputs(5424) <= layer1_outputs(8664);
    layer2_outputs(5425) <= not((layer1_outputs(8366)) or (layer1_outputs(4850)));
    layer2_outputs(5426) <= not(layer1_outputs(9926));
    layer2_outputs(5427) <= layer1_outputs(5153);
    layer2_outputs(5428) <= not((layer1_outputs(8620)) or (layer1_outputs(1760)));
    layer2_outputs(5429) <= (layer1_outputs(5634)) and (layer1_outputs(6072));
    layer2_outputs(5430) <= layer1_outputs(8143);
    layer2_outputs(5431) <= (layer1_outputs(8469)) and not (layer1_outputs(7056));
    layer2_outputs(5432) <= layer1_outputs(3202);
    layer2_outputs(5433) <= not(layer1_outputs(5993));
    layer2_outputs(5434) <= layer1_outputs(3769);
    layer2_outputs(5435) <= not(layer1_outputs(5148));
    layer2_outputs(5436) <= not(layer1_outputs(9029));
    layer2_outputs(5437) <= (layer1_outputs(8318)) xor (layer1_outputs(1757));
    layer2_outputs(5438) <= layer1_outputs(10005);
    layer2_outputs(5439) <= not(layer1_outputs(4602));
    layer2_outputs(5440) <= (layer1_outputs(1565)) and not (layer1_outputs(5046));
    layer2_outputs(5441) <= layer1_outputs(758);
    layer2_outputs(5442) <= (layer1_outputs(8655)) and (layer1_outputs(122));
    layer2_outputs(5443) <= not(layer1_outputs(1744));
    layer2_outputs(5444) <= not(layer1_outputs(4288));
    layer2_outputs(5445) <= layer1_outputs(3727);
    layer2_outputs(5446) <= layer1_outputs(6746);
    layer2_outputs(5447) <= layer1_outputs(2223);
    layer2_outputs(5448) <= not(layer1_outputs(9273)) or (layer1_outputs(1249));
    layer2_outputs(5449) <= (layer1_outputs(9305)) xor (layer1_outputs(5261));
    layer2_outputs(5450) <= not(layer1_outputs(8586));
    layer2_outputs(5451) <= layer1_outputs(4364);
    layer2_outputs(5452) <= layer1_outputs(5849);
    layer2_outputs(5453) <= layer1_outputs(7611);
    layer2_outputs(5454) <= layer1_outputs(734);
    layer2_outputs(5455) <= (layer1_outputs(4061)) and (layer1_outputs(8218));
    layer2_outputs(5456) <= not((layer1_outputs(9581)) xor (layer1_outputs(178)));
    layer2_outputs(5457) <= layer1_outputs(6132);
    layer2_outputs(5458) <= not((layer1_outputs(415)) xor (layer1_outputs(6970)));
    layer2_outputs(5459) <= (layer1_outputs(876)) and (layer1_outputs(7996));
    layer2_outputs(5460) <= not((layer1_outputs(7317)) xor (layer1_outputs(1618)));
    layer2_outputs(5461) <= layer1_outputs(3808);
    layer2_outputs(5462) <= layer1_outputs(6551);
    layer2_outputs(5463) <= layer1_outputs(7185);
    layer2_outputs(5464) <= layer1_outputs(8984);
    layer2_outputs(5465) <= layer1_outputs(7224);
    layer2_outputs(5466) <= not((layer1_outputs(6242)) or (layer1_outputs(3734)));
    layer2_outputs(5467) <= (layer1_outputs(331)) and not (layer1_outputs(7892));
    layer2_outputs(5468) <= (layer1_outputs(5170)) xor (layer1_outputs(765));
    layer2_outputs(5469) <= layer1_outputs(10163);
    layer2_outputs(5470) <= not(layer1_outputs(1872)) or (layer1_outputs(5998));
    layer2_outputs(5471) <= not(layer1_outputs(7549));
    layer2_outputs(5472) <= (layer1_outputs(8361)) xor (layer1_outputs(6920));
    layer2_outputs(5473) <= (layer1_outputs(5779)) and not (layer1_outputs(8769));
    layer2_outputs(5474) <= layer1_outputs(2344);
    layer2_outputs(5475) <= layer1_outputs(5641);
    layer2_outputs(5476) <= (layer1_outputs(6292)) or (layer1_outputs(9995));
    layer2_outputs(5477) <= not((layer1_outputs(9472)) xor (layer1_outputs(8582)));
    layer2_outputs(5478) <= (layer1_outputs(4542)) or (layer1_outputs(2278));
    layer2_outputs(5479) <= layer1_outputs(1278);
    layer2_outputs(5480) <= '0';
    layer2_outputs(5481) <= layer1_outputs(5043);
    layer2_outputs(5482) <= layer1_outputs(6508);
    layer2_outputs(5483) <= not(layer1_outputs(7287)) or (layer1_outputs(1194));
    layer2_outputs(5484) <= (layer1_outputs(6650)) and not (layer1_outputs(5950));
    layer2_outputs(5485) <= not(layer1_outputs(2979)) or (layer1_outputs(6201));
    layer2_outputs(5486) <= (layer1_outputs(3871)) or (layer1_outputs(9283));
    layer2_outputs(5487) <= not((layer1_outputs(1418)) or (layer1_outputs(2065)));
    layer2_outputs(5488) <= not((layer1_outputs(7590)) and (layer1_outputs(5404)));
    layer2_outputs(5489) <= layer1_outputs(6092);
    layer2_outputs(5490) <= not(layer1_outputs(4849));
    layer2_outputs(5491) <= not(layer1_outputs(8154)) or (layer1_outputs(5903));
    layer2_outputs(5492) <= (layer1_outputs(2521)) or (layer1_outputs(995));
    layer2_outputs(5493) <= not(layer1_outputs(1713)) or (layer1_outputs(3331));
    layer2_outputs(5494) <= layer1_outputs(4080);
    layer2_outputs(5495) <= layer1_outputs(4882);
    layer2_outputs(5496) <= layer1_outputs(9387);
    layer2_outputs(5497) <= layer1_outputs(7144);
    layer2_outputs(5498) <= not(layer1_outputs(1777));
    layer2_outputs(5499) <= (layer1_outputs(6737)) and not (layer1_outputs(8672));
    layer2_outputs(5500) <= layer1_outputs(3262);
    layer2_outputs(5501) <= not(layer1_outputs(243));
    layer2_outputs(5502) <= layer1_outputs(578);
    layer2_outputs(5503) <= not(layer1_outputs(2726));
    layer2_outputs(5504) <= (layer1_outputs(5636)) xor (layer1_outputs(5565));
    layer2_outputs(5505) <= layer1_outputs(9672);
    layer2_outputs(5506) <= not(layer1_outputs(9128));
    layer2_outputs(5507) <= layer1_outputs(8995);
    layer2_outputs(5508) <= not(layer1_outputs(505)) or (layer1_outputs(4013));
    layer2_outputs(5509) <= not(layer1_outputs(1343));
    layer2_outputs(5510) <= layer1_outputs(5026);
    layer2_outputs(5511) <= not(layer1_outputs(5389)) or (layer1_outputs(9501));
    layer2_outputs(5512) <= not(layer1_outputs(7797));
    layer2_outputs(5513) <= layer1_outputs(2153);
    layer2_outputs(5514) <= not(layer1_outputs(646));
    layer2_outputs(5515) <= not((layer1_outputs(9179)) or (layer1_outputs(729)));
    layer2_outputs(5516) <= not(layer1_outputs(2830));
    layer2_outputs(5517) <= not((layer1_outputs(1269)) and (layer1_outputs(4390)));
    layer2_outputs(5518) <= not(layer1_outputs(3436));
    layer2_outputs(5519) <= not(layer1_outputs(219));
    layer2_outputs(5520) <= layer1_outputs(3373);
    layer2_outputs(5521) <= not((layer1_outputs(3180)) or (layer1_outputs(2477)));
    layer2_outputs(5522) <= layer1_outputs(1416);
    layer2_outputs(5523) <= not(layer1_outputs(7275));
    layer2_outputs(5524) <= not(layer1_outputs(3551));
    layer2_outputs(5525) <= layer1_outputs(1065);
    layer2_outputs(5526) <= layer1_outputs(7234);
    layer2_outputs(5527) <= layer1_outputs(4859);
    layer2_outputs(5528) <= not(layer1_outputs(7461));
    layer2_outputs(5529) <= not(layer1_outputs(4494));
    layer2_outputs(5530) <= not(layer1_outputs(5585));
    layer2_outputs(5531) <= layer1_outputs(5116);
    layer2_outputs(5532) <= (layer1_outputs(2241)) and not (layer1_outputs(1055));
    layer2_outputs(5533) <= layer1_outputs(1950);
    layer2_outputs(5534) <= not(layer1_outputs(1046));
    layer2_outputs(5535) <= not(layer1_outputs(2838));
    layer2_outputs(5536) <= (layer1_outputs(2176)) xor (layer1_outputs(4745));
    layer2_outputs(5537) <= layer1_outputs(6353);
    layer2_outputs(5538) <= not(layer1_outputs(5795));
    layer2_outputs(5539) <= (layer1_outputs(53)) or (layer1_outputs(6275));
    layer2_outputs(5540) <= (layer1_outputs(336)) xor (layer1_outputs(7720));
    layer2_outputs(5541) <= not(layer1_outputs(6177)) or (layer1_outputs(7504));
    layer2_outputs(5542) <= layer1_outputs(5329);
    layer2_outputs(5543) <= not(layer1_outputs(4550));
    layer2_outputs(5544) <= not(layer1_outputs(4091));
    layer2_outputs(5545) <= (layer1_outputs(9238)) xor (layer1_outputs(4351));
    layer2_outputs(5546) <= not(layer1_outputs(10108));
    layer2_outputs(5547) <= layer1_outputs(9048);
    layer2_outputs(5548) <= (layer1_outputs(8651)) or (layer1_outputs(8945));
    layer2_outputs(5549) <= not((layer1_outputs(2826)) and (layer1_outputs(4881)));
    layer2_outputs(5550) <= (layer1_outputs(3318)) or (layer1_outputs(3752));
    layer2_outputs(5551) <= layer1_outputs(9759);
    layer2_outputs(5552) <= '1';
    layer2_outputs(5553) <= layer1_outputs(9462);
    layer2_outputs(5554) <= layer1_outputs(7775);
    layer2_outputs(5555) <= (layer1_outputs(4684)) and (layer1_outputs(5388));
    layer2_outputs(5556) <= layer1_outputs(2493);
    layer2_outputs(5557) <= layer1_outputs(226);
    layer2_outputs(5558) <= layer1_outputs(8504);
    layer2_outputs(5559) <= not((layer1_outputs(3444)) or (layer1_outputs(5832)));
    layer2_outputs(5560) <= not(layer1_outputs(3895));
    layer2_outputs(5561) <= layer1_outputs(5188);
    layer2_outputs(5562) <= (layer1_outputs(8536)) xor (layer1_outputs(7117));
    layer2_outputs(5563) <= not(layer1_outputs(5335));
    layer2_outputs(5564) <= layer1_outputs(9831);
    layer2_outputs(5565) <= layer1_outputs(5030);
    layer2_outputs(5566) <= not(layer1_outputs(1270)) or (layer1_outputs(9078));
    layer2_outputs(5567) <= '0';
    layer2_outputs(5568) <= not(layer1_outputs(1546));
    layer2_outputs(5569) <= not(layer1_outputs(8115));
    layer2_outputs(5570) <= layer1_outputs(8607);
    layer2_outputs(5571) <= not(layer1_outputs(7440));
    layer2_outputs(5572) <= not((layer1_outputs(7060)) xor (layer1_outputs(3685)));
    layer2_outputs(5573) <= not((layer1_outputs(10209)) xor (layer1_outputs(9240)));
    layer2_outputs(5574) <= layer1_outputs(4957);
    layer2_outputs(5575) <= not(layer1_outputs(8656)) or (layer1_outputs(1030));
    layer2_outputs(5576) <= not(layer1_outputs(2088));
    layer2_outputs(5577) <= (layer1_outputs(2633)) and not (layer1_outputs(7734));
    layer2_outputs(5578) <= not((layer1_outputs(8370)) or (layer1_outputs(511)));
    layer2_outputs(5579) <= layer1_outputs(2418);
    layer2_outputs(5580) <= not((layer1_outputs(5205)) and (layer1_outputs(7368)));
    layer2_outputs(5581) <= not((layer1_outputs(8743)) xor (layer1_outputs(1073)));
    layer2_outputs(5582) <= not(layer1_outputs(9990));
    layer2_outputs(5583) <= not(layer1_outputs(4420)) or (layer1_outputs(8292));
    layer2_outputs(5584) <= not(layer1_outputs(7211)) or (layer1_outputs(5670));
    layer2_outputs(5585) <= not(layer1_outputs(1674));
    layer2_outputs(5586) <= not(layer1_outputs(4661));
    layer2_outputs(5587) <= not(layer1_outputs(5421));
    layer2_outputs(5588) <= (layer1_outputs(3539)) and not (layer1_outputs(10095));
    layer2_outputs(5589) <= not((layer1_outputs(7412)) xor (layer1_outputs(3021)));
    layer2_outputs(5590) <= (layer1_outputs(7922)) and (layer1_outputs(2266));
    layer2_outputs(5591) <= not(layer1_outputs(3709));
    layer2_outputs(5592) <= not(layer1_outputs(3198));
    layer2_outputs(5593) <= not(layer1_outputs(6210));
    layer2_outputs(5594) <= layer1_outputs(9594);
    layer2_outputs(5595) <= (layer1_outputs(10014)) and (layer1_outputs(3244));
    layer2_outputs(5596) <= layer1_outputs(7584);
    layer2_outputs(5597) <= (layer1_outputs(8110)) and not (layer1_outputs(1562));
    layer2_outputs(5598) <= layer1_outputs(1129);
    layer2_outputs(5599) <= layer1_outputs(188);
    layer2_outputs(5600) <= layer1_outputs(195);
    layer2_outputs(5601) <= (layer1_outputs(308)) and (layer1_outputs(8933));
    layer2_outputs(5602) <= not(layer1_outputs(7267));
    layer2_outputs(5603) <= layer1_outputs(9829);
    layer2_outputs(5604) <= (layer1_outputs(1342)) and not (layer1_outputs(818));
    layer2_outputs(5605) <= (layer1_outputs(1992)) xor (layer1_outputs(6435));
    layer2_outputs(5606) <= layer1_outputs(4034);
    layer2_outputs(5607) <= layer1_outputs(3527);
    layer2_outputs(5608) <= not(layer1_outputs(9079));
    layer2_outputs(5609) <= not(layer1_outputs(7498));
    layer2_outputs(5610) <= layer1_outputs(2971);
    layer2_outputs(5611) <= not(layer1_outputs(8053));
    layer2_outputs(5612) <= not(layer1_outputs(827));
    layer2_outputs(5613) <= not(layer1_outputs(867));
    layer2_outputs(5614) <= layer1_outputs(8326);
    layer2_outputs(5615) <= layer1_outputs(9848);
    layer2_outputs(5616) <= not(layer1_outputs(4121));
    layer2_outputs(5617) <= not(layer1_outputs(8394));
    layer2_outputs(5618) <= (layer1_outputs(1344)) or (layer1_outputs(4049));
    layer2_outputs(5619) <= layer1_outputs(640);
    layer2_outputs(5620) <= not(layer1_outputs(6053));
    layer2_outputs(5621) <= layer1_outputs(2680);
    layer2_outputs(5622) <= not(layer1_outputs(9976));
    layer2_outputs(5623) <= not(layer1_outputs(746));
    layer2_outputs(5624) <= (layer1_outputs(4249)) xor (layer1_outputs(8926));
    layer2_outputs(5625) <= not(layer1_outputs(569));
    layer2_outputs(5626) <= layer1_outputs(3977);
    layer2_outputs(5627) <= not(layer1_outputs(6169)) or (layer1_outputs(5571));
    layer2_outputs(5628) <= not(layer1_outputs(7400));
    layer2_outputs(5629) <= not((layer1_outputs(3011)) xor (layer1_outputs(2729)));
    layer2_outputs(5630) <= not((layer1_outputs(2757)) xor (layer1_outputs(3393)));
    layer2_outputs(5631) <= layer1_outputs(1337);
    layer2_outputs(5632) <= layer1_outputs(6365);
    layer2_outputs(5633) <= not(layer1_outputs(10205));
    layer2_outputs(5634) <= not((layer1_outputs(3830)) or (layer1_outputs(7640)));
    layer2_outputs(5635) <= not(layer1_outputs(6669));
    layer2_outputs(5636) <= not(layer1_outputs(420));
    layer2_outputs(5637) <= not(layer1_outputs(5040));
    layer2_outputs(5638) <= layer1_outputs(7848);
    layer2_outputs(5639) <= not(layer1_outputs(6204));
    layer2_outputs(5640) <= not((layer1_outputs(356)) or (layer1_outputs(5296)));
    layer2_outputs(5641) <= not(layer1_outputs(2784)) or (layer1_outputs(9148));
    layer2_outputs(5642) <= layer1_outputs(7689);
    layer2_outputs(5643) <= layer1_outputs(6721);
    layer2_outputs(5644) <= layer1_outputs(4283);
    layer2_outputs(5645) <= layer1_outputs(402);
    layer2_outputs(5646) <= not(layer1_outputs(8539));
    layer2_outputs(5647) <= layer1_outputs(6708);
    layer2_outputs(5648) <= not(layer1_outputs(332));
    layer2_outputs(5649) <= not(layer1_outputs(9788));
    layer2_outputs(5650) <= not(layer1_outputs(8853));
    layer2_outputs(5651) <= not((layer1_outputs(4210)) xor (layer1_outputs(6664)));
    layer2_outputs(5652) <= layer1_outputs(4708);
    layer2_outputs(5653) <= not(layer1_outputs(8211));
    layer2_outputs(5654) <= layer1_outputs(2958);
    layer2_outputs(5655) <= not(layer1_outputs(9000));
    layer2_outputs(5656) <= layer1_outputs(6796);
    layer2_outputs(5657) <= layer1_outputs(820);
    layer2_outputs(5658) <= not((layer1_outputs(9422)) or (layer1_outputs(8093)));
    layer2_outputs(5659) <= layer1_outputs(2168);
    layer2_outputs(5660) <= layer1_outputs(6497);
    layer2_outputs(5661) <= layer1_outputs(3976);
    layer2_outputs(5662) <= not(layer1_outputs(2303));
    layer2_outputs(5663) <= not(layer1_outputs(2587));
    layer2_outputs(5664) <= layer1_outputs(3228);
    layer2_outputs(5665) <= not((layer1_outputs(1715)) or (layer1_outputs(5737)));
    layer2_outputs(5666) <= (layer1_outputs(6617)) and (layer1_outputs(5481));
    layer2_outputs(5667) <= (layer1_outputs(2329)) and (layer1_outputs(1622));
    layer2_outputs(5668) <= not(layer1_outputs(6455));
    layer2_outputs(5669) <= (layer1_outputs(7051)) xor (layer1_outputs(5041));
    layer2_outputs(5670) <= (layer1_outputs(8082)) and not (layer1_outputs(5909));
    layer2_outputs(5671) <= layer1_outputs(7582);
    layer2_outputs(5672) <= not(layer1_outputs(1324));
    layer2_outputs(5673) <= not(layer1_outputs(8778)) or (layer1_outputs(685));
    layer2_outputs(5674) <= (layer1_outputs(4081)) or (layer1_outputs(3757));
    layer2_outputs(5675) <= not((layer1_outputs(9370)) or (layer1_outputs(9937)));
    layer2_outputs(5676) <= (layer1_outputs(1027)) and not (layer1_outputs(3273));
    layer2_outputs(5677) <= not((layer1_outputs(6438)) xor (layer1_outputs(9530)));
    layer2_outputs(5678) <= not(layer1_outputs(5111));
    layer2_outputs(5679) <= (layer1_outputs(6115)) and (layer1_outputs(1467));
    layer2_outputs(5680) <= not(layer1_outputs(9360));
    layer2_outputs(5681) <= not(layer1_outputs(2991));
    layer2_outputs(5682) <= not(layer1_outputs(484));
    layer2_outputs(5683) <= (layer1_outputs(2492)) and not (layer1_outputs(2363));
    layer2_outputs(5684) <= not(layer1_outputs(4330));
    layer2_outputs(5685) <= not(layer1_outputs(5413));
    layer2_outputs(5686) <= not(layer1_outputs(253));
    layer2_outputs(5687) <= not((layer1_outputs(8259)) and (layer1_outputs(2706)));
    layer2_outputs(5688) <= (layer1_outputs(1146)) and not (layer1_outputs(6643));
    layer2_outputs(5689) <= layer1_outputs(2402);
    layer2_outputs(5690) <= not(layer1_outputs(9290));
    layer2_outputs(5691) <= layer1_outputs(9557);
    layer2_outputs(5692) <= (layer1_outputs(7499)) and (layer1_outputs(1752));
    layer2_outputs(5693) <= (layer1_outputs(9511)) and not (layer1_outputs(4332));
    layer2_outputs(5694) <= not(layer1_outputs(2543));
    layer2_outputs(5695) <= layer1_outputs(1100);
    layer2_outputs(5696) <= layer1_outputs(2268);
    layer2_outputs(5697) <= layer1_outputs(4337);
    layer2_outputs(5698) <= (layer1_outputs(6574)) xor (layer1_outputs(3273));
    layer2_outputs(5699) <= not(layer1_outputs(1403));
    layer2_outputs(5700) <= not(layer1_outputs(2661));
    layer2_outputs(5701) <= layer1_outputs(1287);
    layer2_outputs(5702) <= not(layer1_outputs(7739));
    layer2_outputs(5703) <= layer1_outputs(6811);
    layer2_outputs(5704) <= not(layer1_outputs(27));
    layer2_outputs(5705) <= not(layer1_outputs(3645));
    layer2_outputs(5706) <= (layer1_outputs(1501)) and not (layer1_outputs(8298));
    layer2_outputs(5707) <= not(layer1_outputs(9713));
    layer2_outputs(5708) <= layer1_outputs(1014);
    layer2_outputs(5709) <= not(layer1_outputs(561)) or (layer1_outputs(9019));
    layer2_outputs(5710) <= layer1_outputs(8171);
    layer2_outputs(5711) <= not(layer1_outputs(2083));
    layer2_outputs(5712) <= (layer1_outputs(2)) xor (layer1_outputs(6103));
    layer2_outputs(5713) <= not(layer1_outputs(3278));
    layer2_outputs(5714) <= layer1_outputs(10129);
    layer2_outputs(5715) <= layer1_outputs(9957);
    layer2_outputs(5716) <= layer1_outputs(8152);
    layer2_outputs(5717) <= layer1_outputs(1086);
    layer2_outputs(5718) <= (layer1_outputs(5673)) xor (layer1_outputs(7902));
    layer2_outputs(5719) <= not(layer1_outputs(3617));
    layer2_outputs(5720) <= (layer1_outputs(3748)) and not (layer1_outputs(3315));
    layer2_outputs(5721) <= (layer1_outputs(1785)) or (layer1_outputs(4716));
    layer2_outputs(5722) <= layer1_outputs(6703);
    layer2_outputs(5723) <= not(layer1_outputs(9935));
    layer2_outputs(5724) <= not((layer1_outputs(3934)) or (layer1_outputs(1383)));
    layer2_outputs(5725) <= layer1_outputs(928);
    layer2_outputs(5726) <= (layer1_outputs(6121)) xor (layer1_outputs(8844));
    layer2_outputs(5727) <= not(layer1_outputs(9423));
    layer2_outputs(5728) <= '1';
    layer2_outputs(5729) <= not(layer1_outputs(2192));
    layer2_outputs(5730) <= (layer1_outputs(8402)) or (layer1_outputs(452));
    layer2_outputs(5731) <= not(layer1_outputs(8772)) or (layer1_outputs(3705));
    layer2_outputs(5732) <= not(layer1_outputs(4176));
    layer2_outputs(5733) <= layer1_outputs(3600);
    layer2_outputs(5734) <= not((layer1_outputs(482)) xor (layer1_outputs(8884)));
    layer2_outputs(5735) <= not(layer1_outputs(8813));
    layer2_outputs(5736) <= not((layer1_outputs(5360)) or (layer1_outputs(10153)));
    layer2_outputs(5737) <= not(layer1_outputs(2762));
    layer2_outputs(5738) <= not(layer1_outputs(9316));
    layer2_outputs(5739) <= not((layer1_outputs(1242)) xor (layer1_outputs(9876)));
    layer2_outputs(5740) <= layer1_outputs(414);
    layer2_outputs(5741) <= not(layer1_outputs(9481)) or (layer1_outputs(7284));
    layer2_outputs(5742) <= layer1_outputs(9746);
    layer2_outputs(5743) <= (layer1_outputs(9195)) and not (layer1_outputs(3987));
    layer2_outputs(5744) <= (layer1_outputs(5077)) and (layer1_outputs(9751));
    layer2_outputs(5745) <= layer1_outputs(8339);
    layer2_outputs(5746) <= not(layer1_outputs(3308));
    layer2_outputs(5747) <= not(layer1_outputs(713));
    layer2_outputs(5748) <= not((layer1_outputs(8808)) xor (layer1_outputs(1123)));
    layer2_outputs(5749) <= not(layer1_outputs(10077));
    layer2_outputs(5750) <= not(layer1_outputs(5350));
    layer2_outputs(5751) <= not(layer1_outputs(2621));
    layer2_outputs(5752) <= layer1_outputs(198);
    layer2_outputs(5753) <= not((layer1_outputs(1009)) or (layer1_outputs(9724)));
    layer2_outputs(5754) <= (layer1_outputs(7749)) and (layer1_outputs(794));
    layer2_outputs(5755) <= (layer1_outputs(29)) and (layer1_outputs(4479));
    layer2_outputs(5756) <= not(layer1_outputs(4237));
    layer2_outputs(5757) <= not(layer1_outputs(900));
    layer2_outputs(5758) <= not(layer1_outputs(904));
    layer2_outputs(5759) <= layer1_outputs(10224);
    layer2_outputs(5760) <= (layer1_outputs(6606)) or (layer1_outputs(3688));
    layer2_outputs(5761) <= not(layer1_outputs(174));
    layer2_outputs(5762) <= layer1_outputs(1833);
    layer2_outputs(5763) <= not(layer1_outputs(1149)) or (layer1_outputs(5019));
    layer2_outputs(5764) <= layer1_outputs(5620);
    layer2_outputs(5765) <= layer1_outputs(1939);
    layer2_outputs(5766) <= (layer1_outputs(4875)) and not (layer1_outputs(1510));
    layer2_outputs(5767) <= not((layer1_outputs(2241)) xor (layer1_outputs(8925)));
    layer2_outputs(5768) <= not(layer1_outputs(8233));
    layer2_outputs(5769) <= not(layer1_outputs(10011));
    layer2_outputs(5770) <= layer1_outputs(7988);
    layer2_outputs(5771) <= '1';
    layer2_outputs(5772) <= not(layer1_outputs(8764));
    layer2_outputs(5773) <= not(layer1_outputs(2998));
    layer2_outputs(5774) <= (layer1_outputs(2984)) and not (layer1_outputs(4699));
    layer2_outputs(5775) <= (layer1_outputs(7618)) or (layer1_outputs(2888));
    layer2_outputs(5776) <= (layer1_outputs(5972)) and not (layer1_outputs(8931));
    layer2_outputs(5777) <= layer1_outputs(3213);
    layer2_outputs(5778) <= layer1_outputs(9692);
    layer2_outputs(5779) <= not((layer1_outputs(6701)) or (layer1_outputs(5281)));
    layer2_outputs(5780) <= layer1_outputs(4249);
    layer2_outputs(5781) <= not(layer1_outputs(8284)) or (layer1_outputs(8883));
    layer2_outputs(5782) <= (layer1_outputs(4605)) and not (layer1_outputs(8146));
    layer2_outputs(5783) <= layer1_outputs(4074);
    layer2_outputs(5784) <= not(layer1_outputs(4174)) or (layer1_outputs(8054));
    layer2_outputs(5785) <= not(layer1_outputs(7165));
    layer2_outputs(5786) <= (layer1_outputs(4043)) and (layer1_outputs(3010));
    layer2_outputs(5787) <= layer1_outputs(166);
    layer2_outputs(5788) <= not(layer1_outputs(4785));
    layer2_outputs(5789) <= layer1_outputs(2458);
    layer2_outputs(5790) <= not((layer1_outputs(8612)) or (layer1_outputs(234)));
    layer2_outputs(5791) <= (layer1_outputs(820)) and not (layer1_outputs(8460));
    layer2_outputs(5792) <= not(layer1_outputs(5534));
    layer2_outputs(5793) <= not(layer1_outputs(1087));
    layer2_outputs(5794) <= not(layer1_outputs(9487)) or (layer1_outputs(1236));
    layer2_outputs(5795) <= layer1_outputs(168);
    layer2_outputs(5796) <= not(layer1_outputs(7493));
    layer2_outputs(5797) <= not(layer1_outputs(568));
    layer2_outputs(5798) <= (layer1_outputs(2386)) and not (layer1_outputs(8634));
    layer2_outputs(5799) <= not(layer1_outputs(6490)) or (layer1_outputs(752));
    layer2_outputs(5800) <= not((layer1_outputs(8337)) and (layer1_outputs(2429)));
    layer2_outputs(5801) <= not(layer1_outputs(2612));
    layer2_outputs(5802) <= layer1_outputs(2334);
    layer2_outputs(5803) <= not(layer1_outputs(2183));
    layer2_outputs(5804) <= not(layer1_outputs(7839));
    layer2_outputs(5805) <= (layer1_outputs(6306)) and not (layer1_outputs(567));
    layer2_outputs(5806) <= not((layer1_outputs(3739)) and (layer1_outputs(9441)));
    layer2_outputs(5807) <= layer1_outputs(2993);
    layer2_outputs(5808) <= not(layer1_outputs(2410)) or (layer1_outputs(8026));
    layer2_outputs(5809) <= not((layer1_outputs(3000)) xor (layer1_outputs(8162)));
    layer2_outputs(5810) <= not(layer1_outputs(3549));
    layer2_outputs(5811) <= not(layer1_outputs(2473));
    layer2_outputs(5812) <= not(layer1_outputs(436)) or (layer1_outputs(8610));
    layer2_outputs(5813) <= not(layer1_outputs(899));
    layer2_outputs(5814) <= layer1_outputs(7323);
    layer2_outputs(5815) <= '1';
    layer2_outputs(5816) <= (layer1_outputs(3803)) xor (layer1_outputs(9418));
    layer2_outputs(5817) <= layer1_outputs(9993);
    layer2_outputs(5818) <= layer1_outputs(198);
    layer2_outputs(5819) <= not(layer1_outputs(6038));
    layer2_outputs(5820) <= (layer1_outputs(10022)) and not (layer1_outputs(7667));
    layer2_outputs(5821) <= not(layer1_outputs(5591)) or (layer1_outputs(3102));
    layer2_outputs(5822) <= not(layer1_outputs(3295)) or (layer1_outputs(5317));
    layer2_outputs(5823) <= (layer1_outputs(4597)) and (layer1_outputs(4857));
    layer2_outputs(5824) <= layer1_outputs(327);
    layer2_outputs(5825) <= not((layer1_outputs(4624)) xor (layer1_outputs(5061)));
    layer2_outputs(5826) <= not(layer1_outputs(2087));
    layer2_outputs(5827) <= layer1_outputs(7718);
    layer2_outputs(5828) <= (layer1_outputs(3056)) and (layer1_outputs(6593));
    layer2_outputs(5829) <= layer1_outputs(8159);
    layer2_outputs(5830) <= layer1_outputs(899);
    layer2_outputs(5831) <= layer1_outputs(8188);
    layer2_outputs(5832) <= not(layer1_outputs(3372)) or (layer1_outputs(6044));
    layer2_outputs(5833) <= not(layer1_outputs(7375)) or (layer1_outputs(5141));
    layer2_outputs(5834) <= (layer1_outputs(746)) or (layer1_outputs(9281));
    layer2_outputs(5835) <= not(layer1_outputs(4735));
    layer2_outputs(5836) <= not(layer1_outputs(9880));
    layer2_outputs(5837) <= not(layer1_outputs(1171));
    layer2_outputs(5838) <= (layer1_outputs(5666)) or (layer1_outputs(3172));
    layer2_outputs(5839) <= not(layer1_outputs(3490));
    layer2_outputs(5840) <= layer1_outputs(3599);
    layer2_outputs(5841) <= (layer1_outputs(2503)) and not (layer1_outputs(9456));
    layer2_outputs(5842) <= not(layer1_outputs(8438));
    layer2_outputs(5843) <= not(layer1_outputs(8136));
    layer2_outputs(5844) <= not(layer1_outputs(97));
    layer2_outputs(5845) <= layer1_outputs(8099);
    layer2_outputs(5846) <= not(layer1_outputs(6820)) or (layer1_outputs(1772));
    layer2_outputs(5847) <= not(layer1_outputs(947));
    layer2_outputs(5848) <= layer1_outputs(9765);
    layer2_outputs(5849) <= not((layer1_outputs(2456)) xor (layer1_outputs(1792)));
    layer2_outputs(5850) <= not(layer1_outputs(8464));
    layer2_outputs(5851) <= (layer1_outputs(78)) and (layer1_outputs(5990));
    layer2_outputs(5852) <= '1';
    layer2_outputs(5853) <= not((layer1_outputs(8440)) xor (layer1_outputs(3192)));
    layer2_outputs(5854) <= not(layer1_outputs(9984));
    layer2_outputs(5855) <= layer1_outputs(4344);
    layer2_outputs(5856) <= (layer1_outputs(2596)) and not (layer1_outputs(5272));
    layer2_outputs(5857) <= not(layer1_outputs(10005));
    layer2_outputs(5858) <= not(layer1_outputs(4401)) or (layer1_outputs(3336));
    layer2_outputs(5859) <= not((layer1_outputs(107)) or (layer1_outputs(6303)));
    layer2_outputs(5860) <= not((layer1_outputs(6715)) xor (layer1_outputs(722)));
    layer2_outputs(5861) <= (layer1_outputs(2025)) and not (layer1_outputs(5797));
    layer2_outputs(5862) <= not(layer1_outputs(7181));
    layer2_outputs(5863) <= not((layer1_outputs(4200)) xor (layer1_outputs(6019)));
    layer2_outputs(5864) <= layer1_outputs(3173);
    layer2_outputs(5865) <= not(layer1_outputs(3155));
    layer2_outputs(5866) <= not(layer1_outputs(1834));
    layer2_outputs(5867) <= not(layer1_outputs(8785));
    layer2_outputs(5868) <= not((layer1_outputs(6304)) and (layer1_outputs(3264)));
    layer2_outputs(5869) <= layer1_outputs(8313);
    layer2_outputs(5870) <= not((layer1_outputs(1385)) and (layer1_outputs(2019)));
    layer2_outputs(5871) <= (layer1_outputs(8025)) and (layer1_outputs(2684));
    layer2_outputs(5872) <= not(layer1_outputs(9690));
    layer2_outputs(5873) <= not(layer1_outputs(2424));
    layer2_outputs(5874) <= not(layer1_outputs(300));
    layer2_outputs(5875) <= not(layer1_outputs(5803)) or (layer1_outputs(7721));
    layer2_outputs(5876) <= layer1_outputs(4430);
    layer2_outputs(5877) <= not(layer1_outputs(9707));
    layer2_outputs(5878) <= not(layer1_outputs(765)) or (layer1_outputs(3522));
    layer2_outputs(5879) <= (layer1_outputs(1513)) xor (layer1_outputs(2404));
    layer2_outputs(5880) <= not(layer1_outputs(6457));
    layer2_outputs(5881) <= (layer1_outputs(8227)) and not (layer1_outputs(555));
    layer2_outputs(5882) <= layer1_outputs(1165);
    layer2_outputs(5883) <= not(layer1_outputs(3225));
    layer2_outputs(5884) <= (layer1_outputs(1384)) and not (layer1_outputs(8008));
    layer2_outputs(5885) <= not(layer1_outputs(8269)) or (layer1_outputs(1863));
    layer2_outputs(5886) <= not((layer1_outputs(9875)) xor (layer1_outputs(5089)));
    layer2_outputs(5887) <= not(layer1_outputs(2744)) or (layer1_outputs(255));
    layer2_outputs(5888) <= layer1_outputs(3446);
    layer2_outputs(5889) <= (layer1_outputs(7115)) or (layer1_outputs(8865));
    layer2_outputs(5890) <= (layer1_outputs(6018)) or (layer1_outputs(4558));
    layer2_outputs(5891) <= layer1_outputs(9518);
    layer2_outputs(5892) <= not((layer1_outputs(958)) xor (layer1_outputs(348)));
    layer2_outputs(5893) <= not((layer1_outputs(1000)) or (layer1_outputs(3933)));
    layer2_outputs(5894) <= not(layer1_outputs(8106));
    layer2_outputs(5895) <= not(layer1_outputs(4520));
    layer2_outputs(5896) <= not(layer1_outputs(7598));
    layer2_outputs(5897) <= not((layer1_outputs(1894)) or (layer1_outputs(1022)));
    layer2_outputs(5898) <= layer1_outputs(8935);
    layer2_outputs(5899) <= layer1_outputs(4020);
    layer2_outputs(5900) <= layer1_outputs(595);
    layer2_outputs(5901) <= layer1_outputs(6933);
    layer2_outputs(5902) <= layer1_outputs(4039);
    layer2_outputs(5903) <= not(layer1_outputs(5783));
    layer2_outputs(5904) <= not((layer1_outputs(9689)) xor (layer1_outputs(916)));
    layer2_outputs(5905) <= not(layer1_outputs(8469));
    layer2_outputs(5906) <= (layer1_outputs(1165)) or (layer1_outputs(7311));
    layer2_outputs(5907) <= '1';
    layer2_outputs(5908) <= not((layer1_outputs(3180)) or (layer1_outputs(9492)));
    layer2_outputs(5909) <= layer1_outputs(3693);
    layer2_outputs(5910) <= (layer1_outputs(3808)) or (layer1_outputs(7827));
    layer2_outputs(5911) <= layer1_outputs(1928);
    layer2_outputs(5912) <= layer1_outputs(9359);
    layer2_outputs(5913) <= not(layer1_outputs(3555));
    layer2_outputs(5914) <= layer1_outputs(7543);
    layer2_outputs(5915) <= (layer1_outputs(6422)) and not (layer1_outputs(1299));
    layer2_outputs(5916) <= not(layer1_outputs(9442)) or (layer1_outputs(9909));
    layer2_outputs(5917) <= layer1_outputs(4960);
    layer2_outputs(5918) <= (layer1_outputs(7247)) xor (layer1_outputs(5785));
    layer2_outputs(5919) <= not(layer1_outputs(4726));
    layer2_outputs(5920) <= layer1_outputs(6611);
    layer2_outputs(5921) <= layer1_outputs(9261);
    layer2_outputs(5922) <= not((layer1_outputs(3795)) xor (layer1_outputs(1270)));
    layer2_outputs(5923) <= not(layer1_outputs(1389));
    layer2_outputs(5924) <= (layer1_outputs(3467)) xor (layer1_outputs(7381));
    layer2_outputs(5925) <= not(layer1_outputs(5337)) or (layer1_outputs(3794));
    layer2_outputs(5926) <= layer1_outputs(2261);
    layer2_outputs(5927) <= layer1_outputs(9578);
    layer2_outputs(5928) <= not(layer1_outputs(8689)) or (layer1_outputs(4289));
    layer2_outputs(5929) <= (layer1_outputs(4493)) and not (layer1_outputs(1453));
    layer2_outputs(5930) <= layer1_outputs(3021);
    layer2_outputs(5931) <= not(layer1_outputs(5226));
    layer2_outputs(5932) <= '1';
    layer2_outputs(5933) <= not((layer1_outputs(5594)) or (layer1_outputs(8713)));
    layer2_outputs(5934) <= layer1_outputs(1707);
    layer2_outputs(5935) <= not(layer1_outputs(6197));
    layer2_outputs(5936) <= (layer1_outputs(3595)) and not (layer1_outputs(273));
    layer2_outputs(5937) <= (layer1_outputs(6475)) and (layer1_outputs(1507));
    layer2_outputs(5938) <= not((layer1_outputs(4768)) xor (layer1_outputs(4218)));
    layer2_outputs(5939) <= layer1_outputs(8051);
    layer2_outputs(5940) <= not(layer1_outputs(4610));
    layer2_outputs(5941) <= layer1_outputs(2583);
    layer2_outputs(5942) <= layer1_outputs(6599);
    layer2_outputs(5943) <= layer1_outputs(2517);
    layer2_outputs(5944) <= (layer1_outputs(3493)) or (layer1_outputs(2225));
    layer2_outputs(5945) <= not((layer1_outputs(5056)) and (layer1_outputs(1670)));
    layer2_outputs(5946) <= (layer1_outputs(3847)) and not (layer1_outputs(106));
    layer2_outputs(5947) <= '1';
    layer2_outputs(5948) <= (layer1_outputs(1793)) and not (layer1_outputs(4115));
    layer2_outputs(5949) <= not((layer1_outputs(2243)) or (layer1_outputs(9605)));
    layer2_outputs(5950) <= not(layer1_outputs(9874));
    layer2_outputs(5951) <= layer1_outputs(4850);
    layer2_outputs(5952) <= layer1_outputs(4082);
    layer2_outputs(5953) <= (layer1_outputs(77)) and not (layer1_outputs(3375));
    layer2_outputs(5954) <= layer1_outputs(5357);
    layer2_outputs(5955) <= not(layer1_outputs(1273));
    layer2_outputs(5956) <= layer1_outputs(7663);
    layer2_outputs(5957) <= (layer1_outputs(5389)) and not (layer1_outputs(9941));
    layer2_outputs(5958) <= layer1_outputs(3379);
    layer2_outputs(5959) <= layer1_outputs(2533);
    layer2_outputs(5960) <= (layer1_outputs(7779)) and (layer1_outputs(3070));
    layer2_outputs(5961) <= layer1_outputs(1787);
    layer2_outputs(5962) <= not(layer1_outputs(2777));
    layer2_outputs(5963) <= not(layer1_outputs(766));
    layer2_outputs(5964) <= not(layer1_outputs(9651)) or (layer1_outputs(3620));
    layer2_outputs(5965) <= not(layer1_outputs(7065));
    layer2_outputs(5966) <= not(layer1_outputs(4184));
    layer2_outputs(5967) <= (layer1_outputs(1878)) and (layer1_outputs(5815));
    layer2_outputs(5968) <= not((layer1_outputs(6718)) and (layer1_outputs(3309)));
    layer2_outputs(5969) <= not(layer1_outputs(5150));
    layer2_outputs(5970) <= layer1_outputs(4084);
    layer2_outputs(5971) <= not(layer1_outputs(8654));
    layer2_outputs(5972) <= not(layer1_outputs(2232)) or (layer1_outputs(7927));
    layer2_outputs(5973) <= not(layer1_outputs(5683)) or (layer1_outputs(150));
    layer2_outputs(5974) <= not(layer1_outputs(25));
    layer2_outputs(5975) <= not(layer1_outputs(9833)) or (layer1_outputs(9138));
    layer2_outputs(5976) <= layer1_outputs(1374);
    layer2_outputs(5977) <= (layer1_outputs(109)) and (layer1_outputs(2753));
    layer2_outputs(5978) <= not(layer1_outputs(2838));
    layer2_outputs(5979) <= (layer1_outputs(5881)) and (layer1_outputs(9822));
    layer2_outputs(5980) <= layer1_outputs(5438);
    layer2_outputs(5981) <= not(layer1_outputs(5433));
    layer2_outputs(5982) <= layer1_outputs(7814);
    layer2_outputs(5983) <= layer1_outputs(5819);
    layer2_outputs(5984) <= (layer1_outputs(1722)) and not (layer1_outputs(9845));
    layer2_outputs(5985) <= not(layer1_outputs(8881)) or (layer1_outputs(4836));
    layer2_outputs(5986) <= not((layer1_outputs(2567)) or (layer1_outputs(6205)));
    layer2_outputs(5987) <= layer1_outputs(1885);
    layer2_outputs(5988) <= (layer1_outputs(2049)) and (layer1_outputs(4371));
    layer2_outputs(5989) <= (layer1_outputs(8482)) and (layer1_outputs(3898));
    layer2_outputs(5990) <= not((layer1_outputs(8666)) and (layer1_outputs(6635)));
    layer2_outputs(5991) <= not(layer1_outputs(2755));
    layer2_outputs(5992) <= (layer1_outputs(8530)) and not (layer1_outputs(8503));
    layer2_outputs(5993) <= not((layer1_outputs(1652)) xor (layer1_outputs(2072)));
    layer2_outputs(5994) <= (layer1_outputs(7772)) and not (layer1_outputs(732));
    layer2_outputs(5995) <= not(layer1_outputs(1283));
    layer2_outputs(5996) <= layer1_outputs(2895);
    layer2_outputs(5997) <= '1';
    layer2_outputs(5998) <= layer1_outputs(8032);
    layer2_outputs(5999) <= not(layer1_outputs(7531));
    layer2_outputs(6000) <= (layer1_outputs(9735)) and not (layer1_outputs(10203));
    layer2_outputs(6001) <= layer1_outputs(9213);
    layer2_outputs(6002) <= not(layer1_outputs(4198));
    layer2_outputs(6003) <= layer1_outputs(932);
    layer2_outputs(6004) <= not(layer1_outputs(7367));
    layer2_outputs(6005) <= (layer1_outputs(7451)) and (layer1_outputs(9160));
    layer2_outputs(6006) <= not(layer1_outputs(9794));
    layer2_outputs(6007) <= layer1_outputs(7951);
    layer2_outputs(6008) <= (layer1_outputs(8888)) and not (layer1_outputs(468));
    layer2_outputs(6009) <= not(layer1_outputs(2641));
    layer2_outputs(6010) <= not(layer1_outputs(636)) or (layer1_outputs(8382));
    layer2_outputs(6011) <= not(layer1_outputs(3451));
    layer2_outputs(6012) <= not(layer1_outputs(9064));
    layer2_outputs(6013) <= (layer1_outputs(7576)) or (layer1_outputs(4055));
    layer2_outputs(6014) <= layer1_outputs(5410);
    layer2_outputs(6015) <= layer1_outputs(5782);
    layer2_outputs(6016) <= layer1_outputs(4353);
    layer2_outputs(6017) <= (layer1_outputs(9187)) and not (layer1_outputs(7548));
    layer2_outputs(6018) <= layer1_outputs(2253);
    layer2_outputs(6019) <= layer1_outputs(3823);
    layer2_outputs(6020) <= not(layer1_outputs(2979));
    layer2_outputs(6021) <= not(layer1_outputs(9582));
    layer2_outputs(6022) <= not(layer1_outputs(6012));
    layer2_outputs(6023) <= (layer1_outputs(4114)) and (layer1_outputs(6297));
    layer2_outputs(6024) <= not((layer1_outputs(4219)) xor (layer1_outputs(2980)));
    layer2_outputs(6025) <= not((layer1_outputs(9190)) xor (layer1_outputs(8804)));
    layer2_outputs(6026) <= not(layer1_outputs(6036));
    layer2_outputs(6027) <= not(layer1_outputs(8961));
    layer2_outputs(6028) <= not((layer1_outputs(2294)) xor (layer1_outputs(7680)));
    layer2_outputs(6029) <= layer1_outputs(3791);
    layer2_outputs(6030) <= not(layer1_outputs(7152));
    layer2_outputs(6031) <= (layer1_outputs(1130)) and (layer1_outputs(3320));
    layer2_outputs(6032) <= '1';
    layer2_outputs(6033) <= not(layer1_outputs(4735)) or (layer1_outputs(8158));
    layer2_outputs(6034) <= layer1_outputs(5939);
    layer2_outputs(6035) <= not(layer1_outputs(626));
    layer2_outputs(6036) <= layer1_outputs(6189);
    layer2_outputs(6037) <= layer1_outputs(8360);
    layer2_outputs(6038) <= layer1_outputs(9569);
    layer2_outputs(6039) <= layer1_outputs(5016);
    layer2_outputs(6040) <= layer1_outputs(9669);
    layer2_outputs(6041) <= layer1_outputs(9609);
    layer2_outputs(6042) <= not(layer1_outputs(9990));
    layer2_outputs(6043) <= layer1_outputs(3529);
    layer2_outputs(6044) <= not((layer1_outputs(4221)) xor (layer1_outputs(7136)));
    layer2_outputs(6045) <= not(layer1_outputs(402));
    layer2_outputs(6046) <= layer1_outputs(2540);
    layer2_outputs(6047) <= not(layer1_outputs(9876));
    layer2_outputs(6048) <= not(layer1_outputs(565)) or (layer1_outputs(9349));
    layer2_outputs(6049) <= not(layer1_outputs(7342));
    layer2_outputs(6050) <= (layer1_outputs(7597)) xor (layer1_outputs(9347));
    layer2_outputs(6051) <= layer1_outputs(8989);
    layer2_outputs(6052) <= (layer1_outputs(6525)) and not (layer1_outputs(3857));
    layer2_outputs(6053) <= layer1_outputs(6133);
    layer2_outputs(6054) <= layer1_outputs(9914);
    layer2_outputs(6055) <= layer1_outputs(2132);
    layer2_outputs(6056) <= not((layer1_outputs(9615)) and (layer1_outputs(9757)));
    layer2_outputs(6057) <= not((layer1_outputs(3726)) or (layer1_outputs(5497)));
    layer2_outputs(6058) <= not(layer1_outputs(10194));
    layer2_outputs(6059) <= layer1_outputs(4177);
    layer2_outputs(6060) <= (layer1_outputs(4458)) xor (layer1_outputs(1430));
    layer2_outputs(6061) <= layer1_outputs(444);
    layer2_outputs(6062) <= layer1_outputs(845);
    layer2_outputs(6063) <= layer1_outputs(2047);
    layer2_outputs(6064) <= (layer1_outputs(3160)) and (layer1_outputs(5455));
    layer2_outputs(6065) <= layer1_outputs(409);
    layer2_outputs(6066) <= (layer1_outputs(3105)) and not (layer1_outputs(9777));
    layer2_outputs(6067) <= layer1_outputs(9438);
    layer2_outputs(6068) <= not(layer1_outputs(4557));
    layer2_outputs(6069) <= not(layer1_outputs(7018)) or (layer1_outputs(7270));
    layer2_outputs(6070) <= not(layer1_outputs(6900)) or (layer1_outputs(4546));
    layer2_outputs(6071) <= (layer1_outputs(8958)) and (layer1_outputs(7990));
    layer2_outputs(6072) <= layer1_outputs(9538);
    layer2_outputs(6073) <= not(layer1_outputs(8877)) or (layer1_outputs(2849));
    layer2_outputs(6074) <= not((layer1_outputs(5359)) and (layer1_outputs(8420)));
    layer2_outputs(6075) <= not(layer1_outputs(1007));
    layer2_outputs(6076) <= (layer1_outputs(1511)) and (layer1_outputs(7239));
    layer2_outputs(6077) <= (layer1_outputs(4882)) xor (layer1_outputs(9468));
    layer2_outputs(6078) <= layer1_outputs(2017);
    layer2_outputs(6079) <= not(layer1_outputs(2094));
    layer2_outputs(6080) <= not(layer1_outputs(5558)) or (layer1_outputs(6059));
    layer2_outputs(6081) <= not((layer1_outputs(5705)) or (layer1_outputs(4492)));
    layer2_outputs(6082) <= layer1_outputs(5028);
    layer2_outputs(6083) <= (layer1_outputs(3307)) and (layer1_outputs(8868));
    layer2_outputs(6084) <= layer1_outputs(29);
    layer2_outputs(6085) <= not((layer1_outputs(5966)) xor (layer1_outputs(3360)));
    layer2_outputs(6086) <= not((layer1_outputs(9463)) xor (layer1_outputs(5419)));
    layer2_outputs(6087) <= not(layer1_outputs(3939));
    layer2_outputs(6088) <= (layer1_outputs(1722)) and not (layer1_outputs(4022));
    layer2_outputs(6089) <= (layer1_outputs(8921)) or (layer1_outputs(6593));
    layer2_outputs(6090) <= (layer1_outputs(1181)) and not (layer1_outputs(4937));
    layer2_outputs(6091) <= not(layer1_outputs(3147)) or (layer1_outputs(4797));
    layer2_outputs(6092) <= (layer1_outputs(2903)) and not (layer1_outputs(2513));
    layer2_outputs(6093) <= not(layer1_outputs(3497));
    layer2_outputs(6094) <= not(layer1_outputs(4775));
    layer2_outputs(6095) <= not(layer1_outputs(4328));
    layer2_outputs(6096) <= (layer1_outputs(4682)) and (layer1_outputs(3217));
    layer2_outputs(6097) <= not((layer1_outputs(5675)) or (layer1_outputs(200)));
    layer2_outputs(6098) <= not(layer1_outputs(6088));
    layer2_outputs(6099) <= layer1_outputs(8552);
    layer2_outputs(6100) <= not((layer1_outputs(1898)) and (layer1_outputs(4453)));
    layer2_outputs(6101) <= not(layer1_outputs(2966));
    layer2_outputs(6102) <= layer1_outputs(3457);
    layer2_outputs(6103) <= (layer1_outputs(4752)) and not (layer1_outputs(3113));
    layer2_outputs(6104) <= layer1_outputs(5371);
    layer2_outputs(6105) <= not(layer1_outputs(4635));
    layer2_outputs(6106) <= (layer1_outputs(9951)) or (layer1_outputs(8409));
    layer2_outputs(6107) <= not(layer1_outputs(1408));
    layer2_outputs(6108) <= not(layer1_outputs(861));
    layer2_outputs(6109) <= not((layer1_outputs(7244)) and (layer1_outputs(5458)));
    layer2_outputs(6110) <= layer1_outputs(5175);
    layer2_outputs(6111) <= not(layer1_outputs(4338));
    layer2_outputs(6112) <= (layer1_outputs(4567)) or (layer1_outputs(1031));
    layer2_outputs(6113) <= layer1_outputs(6001);
    layer2_outputs(6114) <= (layer1_outputs(7710)) and (layer1_outputs(877));
    layer2_outputs(6115) <= layer1_outputs(5135);
    layer2_outputs(6116) <= layer1_outputs(5724);
    layer2_outputs(6117) <= not((layer1_outputs(1439)) or (layer1_outputs(3397)));
    layer2_outputs(6118) <= not(layer1_outputs(2038));
    layer2_outputs(6119) <= not(layer1_outputs(6056)) or (layer1_outputs(6612));
    layer2_outputs(6120) <= not((layer1_outputs(7255)) or (layer1_outputs(3751)));
    layer2_outputs(6121) <= (layer1_outputs(389)) and (layer1_outputs(5035));
    layer2_outputs(6122) <= not((layer1_outputs(5766)) and (layer1_outputs(1986)));
    layer2_outputs(6123) <= not(layer1_outputs(8319));
    layer2_outputs(6124) <= not(layer1_outputs(2143));
    layer2_outputs(6125) <= not(layer1_outputs(713));
    layer2_outputs(6126) <= layer1_outputs(2390);
    layer2_outputs(6127) <= not(layer1_outputs(435));
    layer2_outputs(6128) <= not(layer1_outputs(2573));
    layer2_outputs(6129) <= layer1_outputs(9338);
    layer2_outputs(6130) <= not((layer1_outputs(7318)) and (layer1_outputs(1384)));
    layer2_outputs(6131) <= (layer1_outputs(7356)) and not (layer1_outputs(3992));
    layer2_outputs(6132) <= not(layer1_outputs(3760));
    layer2_outputs(6133) <= layer1_outputs(5000);
    layer2_outputs(6134) <= not(layer1_outputs(853)) or (layer1_outputs(8413));
    layer2_outputs(6135) <= layer1_outputs(1024);
    layer2_outputs(6136) <= not(layer1_outputs(6976));
    layer2_outputs(6137) <= not(layer1_outputs(494));
    layer2_outputs(6138) <= not((layer1_outputs(985)) xor (layer1_outputs(1466)));
    layer2_outputs(6139) <= layer1_outputs(261);
    layer2_outputs(6140) <= not(layer1_outputs(3573));
    layer2_outputs(6141) <= (layer1_outputs(8282)) and not (layer1_outputs(3186));
    layer2_outputs(6142) <= layer1_outputs(7743);
    layer2_outputs(6143) <= not(layer1_outputs(7656));
    layer2_outputs(6144) <= layer1_outputs(5984);
    layer2_outputs(6145) <= not(layer1_outputs(805));
    layer2_outputs(6146) <= layer1_outputs(9796);
    layer2_outputs(6147) <= layer1_outputs(6534);
    layer2_outputs(6148) <= (layer1_outputs(4166)) and not (layer1_outputs(42));
    layer2_outputs(6149) <= not(layer1_outputs(2115));
    layer2_outputs(6150) <= not(layer1_outputs(3199));
    layer2_outputs(6151) <= layer1_outputs(8375);
    layer2_outputs(6152) <= not(layer1_outputs(7456));
    layer2_outputs(6153) <= layer1_outputs(7890);
    layer2_outputs(6154) <= not(layer1_outputs(7444));
    layer2_outputs(6155) <= '1';
    layer2_outputs(6156) <= not(layer1_outputs(2035));
    layer2_outputs(6157) <= not(layer1_outputs(4932)) or (layer1_outputs(2892));
    layer2_outputs(6158) <= (layer1_outputs(10150)) and not (layer1_outputs(4293));
    layer2_outputs(6159) <= not(layer1_outputs(1078));
    layer2_outputs(6160) <= not((layer1_outputs(8938)) xor (layer1_outputs(1142)));
    layer2_outputs(6161) <= layer1_outputs(9122);
    layer2_outputs(6162) <= layer1_outputs(6582);
    layer2_outputs(6163) <= layer1_outputs(4989);
    layer2_outputs(6164) <= (layer1_outputs(7904)) xor (layer1_outputs(1019));
    layer2_outputs(6165) <= (layer1_outputs(9452)) or (layer1_outputs(8476));
    layer2_outputs(6166) <= not(layer1_outputs(3351)) or (layer1_outputs(8371));
    layer2_outputs(6167) <= (layer1_outputs(1849)) and (layer1_outputs(5387));
    layer2_outputs(6168) <= layer1_outputs(7066);
    layer2_outputs(6169) <= layer1_outputs(238);
    layer2_outputs(6170) <= not(layer1_outputs(2088)) or (layer1_outputs(4036));
    layer2_outputs(6171) <= not((layer1_outputs(2974)) or (layer1_outputs(5039)));
    layer2_outputs(6172) <= layer1_outputs(6523);
    layer2_outputs(6173) <= not(layer1_outputs(5467));
    layer2_outputs(6174) <= '0';
    layer2_outputs(6175) <= (layer1_outputs(4500)) or (layer1_outputs(1523));
    layer2_outputs(6176) <= layer1_outputs(7822);
    layer2_outputs(6177) <= layer1_outputs(6931);
    layer2_outputs(6178) <= (layer1_outputs(7471)) or (layer1_outputs(3022));
    layer2_outputs(6179) <= not((layer1_outputs(6763)) xor (layer1_outputs(2475)));
    layer2_outputs(6180) <= (layer1_outputs(9831)) and not (layer1_outputs(8991));
    layer2_outputs(6181) <= not((layer1_outputs(1284)) and (layer1_outputs(1581)));
    layer2_outputs(6182) <= not(layer1_outputs(7477));
    layer2_outputs(6183) <= not((layer1_outputs(6119)) or (layer1_outputs(5963)));
    layer2_outputs(6184) <= not(layer1_outputs(4397));
    layer2_outputs(6185) <= not(layer1_outputs(5878));
    layer2_outputs(6186) <= layer1_outputs(5514);
    layer2_outputs(6187) <= not(layer1_outputs(1643));
    layer2_outputs(6188) <= layer1_outputs(3503);
    layer2_outputs(6189) <= not(layer1_outputs(6318));
    layer2_outputs(6190) <= (layer1_outputs(8694)) and not (layer1_outputs(4556));
    layer2_outputs(6191) <= not((layer1_outputs(7118)) or (layer1_outputs(6054)));
    layer2_outputs(6192) <= layer1_outputs(8779);
    layer2_outputs(6193) <= not(layer1_outputs(4264));
    layer2_outputs(6194) <= not(layer1_outputs(5825));
    layer2_outputs(6195) <= (layer1_outputs(2097)) xor (layer1_outputs(5488));
    layer2_outputs(6196) <= not((layer1_outputs(6786)) and (layer1_outputs(407)));
    layer2_outputs(6197) <= not((layer1_outputs(2748)) xor (layer1_outputs(3448)));
    layer2_outputs(6198) <= not(layer1_outputs(7125));
    layer2_outputs(6199) <= layer1_outputs(7756);
    layer2_outputs(6200) <= (layer1_outputs(1818)) and not (layer1_outputs(8133));
    layer2_outputs(6201) <= (layer1_outputs(6543)) xor (layer1_outputs(1364));
    layer2_outputs(6202) <= not((layer1_outputs(1499)) or (layer1_outputs(1025)));
    layer2_outputs(6203) <= not(layer1_outputs(1376));
    layer2_outputs(6204) <= (layer1_outputs(5220)) and not (layer1_outputs(9030));
    layer2_outputs(6205) <= not(layer1_outputs(183));
    layer2_outputs(6206) <= not(layer1_outputs(6535));
    layer2_outputs(6207) <= not(layer1_outputs(5282));
    layer2_outputs(6208) <= not(layer1_outputs(9277)) or (layer1_outputs(8923));
    layer2_outputs(6209) <= layer1_outputs(328);
    layer2_outputs(6210) <= layer1_outputs(6088);
    layer2_outputs(6211) <= not((layer1_outputs(9575)) and (layer1_outputs(4743)));
    layer2_outputs(6212) <= layer1_outputs(2405);
    layer2_outputs(6213) <= layer1_outputs(115);
    layer2_outputs(6214) <= not((layer1_outputs(4878)) xor (layer1_outputs(8164)));
    layer2_outputs(6215) <= (layer1_outputs(9593)) or (layer1_outputs(10115));
    layer2_outputs(6216) <= not((layer1_outputs(400)) xor (layer1_outputs(4739)));
    layer2_outputs(6217) <= layer1_outputs(3737);
    layer2_outputs(6218) <= layer1_outputs(1400);
    layer2_outputs(6219) <= not(layer1_outputs(333));
    layer2_outputs(6220) <= layer1_outputs(1715);
    layer2_outputs(6221) <= (layer1_outputs(4090)) xor (layer1_outputs(9514));
    layer2_outputs(6222) <= not(layer1_outputs(663));
    layer2_outputs(6223) <= (layer1_outputs(6469)) xor (layer1_outputs(1740));
    layer2_outputs(6224) <= layer1_outputs(8776);
    layer2_outputs(6225) <= not(layer1_outputs(2484));
    layer2_outputs(6226) <= layer1_outputs(6717);
    layer2_outputs(6227) <= not(layer1_outputs(5187));
    layer2_outputs(6228) <= layer1_outputs(3033);
    layer2_outputs(6229) <= layer1_outputs(2899);
    layer2_outputs(6230) <= not((layer1_outputs(5761)) xor (layer1_outputs(7516)));
    layer2_outputs(6231) <= not((layer1_outputs(8730)) and (layer1_outputs(1123)));
    layer2_outputs(6232) <= layer1_outputs(5464);
    layer2_outputs(6233) <= not((layer1_outputs(6076)) and (layer1_outputs(6973)));
    layer2_outputs(6234) <= layer1_outputs(1521);
    layer2_outputs(6235) <= not(layer1_outputs(8111)) or (layer1_outputs(10068));
    layer2_outputs(6236) <= not(layer1_outputs(798));
    layer2_outputs(6237) <= not(layer1_outputs(2391)) or (layer1_outputs(8547));
    layer2_outputs(6238) <= layer1_outputs(8166);
    layer2_outputs(6239) <= (layer1_outputs(4232)) and not (layer1_outputs(386));
    layer2_outputs(6240) <= layer1_outputs(4192);
    layer2_outputs(6241) <= layer1_outputs(5760);
    layer2_outputs(6242) <= not(layer1_outputs(7438));
    layer2_outputs(6243) <= not((layer1_outputs(4146)) and (layer1_outputs(273)));
    layer2_outputs(6244) <= not(layer1_outputs(4214));
    layer2_outputs(6245) <= (layer1_outputs(8062)) and (layer1_outputs(7654));
    layer2_outputs(6246) <= layer1_outputs(6193);
    layer2_outputs(6247) <= not((layer1_outputs(9966)) xor (layer1_outputs(5649)));
    layer2_outputs(6248) <= '1';
    layer2_outputs(6249) <= (layer1_outputs(5869)) and not (layer1_outputs(8436));
    layer2_outputs(6250) <= not(layer1_outputs(3667)) or (layer1_outputs(2415));
    layer2_outputs(6251) <= (layer1_outputs(1219)) xor (layer1_outputs(10056));
    layer2_outputs(6252) <= not(layer1_outputs(8119));
    layer2_outputs(6253) <= not(layer1_outputs(8275)) or (layer1_outputs(7481));
    layer2_outputs(6254) <= not(layer1_outputs(590));
    layer2_outputs(6255) <= not(layer1_outputs(9805));
    layer2_outputs(6256) <= layer1_outputs(2067);
    layer2_outputs(6257) <= (layer1_outputs(7725)) or (layer1_outputs(4717));
    layer2_outputs(6258) <= layer1_outputs(758);
    layer2_outputs(6259) <= (layer1_outputs(8074)) and not (layer1_outputs(6356));
    layer2_outputs(6260) <= (layer1_outputs(8215)) and (layer1_outputs(1332));
    layer2_outputs(6261) <= not(layer1_outputs(8251));
    layer2_outputs(6262) <= not(layer1_outputs(2376));
    layer2_outputs(6263) <= layer1_outputs(2337);
    layer2_outputs(6264) <= layer1_outputs(7190);
    layer2_outputs(6265) <= layer1_outputs(7924);
    layer2_outputs(6266) <= (layer1_outputs(1516)) xor (layer1_outputs(2926));
    layer2_outputs(6267) <= (layer1_outputs(4820)) xor (layer1_outputs(2114));
    layer2_outputs(6268) <= (layer1_outputs(5400)) and (layer1_outputs(8581));
    layer2_outputs(6269) <= not(layer1_outputs(3463));
    layer2_outputs(6270) <= not(layer1_outputs(3806));
    layer2_outputs(6271) <= (layer1_outputs(8352)) and not (layer1_outputs(4235));
    layer2_outputs(6272) <= (layer1_outputs(127)) xor (layer1_outputs(8816));
    layer2_outputs(6273) <= (layer1_outputs(5310)) xor (layer1_outputs(2996));
    layer2_outputs(6274) <= layer1_outputs(3828);
    layer2_outputs(6275) <= not((layer1_outputs(1753)) and (layer1_outputs(216)));
    layer2_outputs(6276) <= layer1_outputs(1757);
    layer2_outputs(6277) <= not(layer1_outputs(5948));
    layer2_outputs(6278) <= layer1_outputs(879);
    layer2_outputs(6279) <= not(layer1_outputs(5313));
    layer2_outputs(6280) <= not((layer1_outputs(1525)) and (layer1_outputs(8427)));
    layer2_outputs(6281) <= layer1_outputs(9552);
    layer2_outputs(6282) <= layer1_outputs(2438);
    layer2_outputs(6283) <= not(layer1_outputs(5660));
    layer2_outputs(6284) <= layer1_outputs(4734);
    layer2_outputs(6285) <= not(layer1_outputs(878));
    layer2_outputs(6286) <= (layer1_outputs(3853)) xor (layer1_outputs(8201));
    layer2_outputs(6287) <= not(layer1_outputs(6273));
    layer2_outputs(6288) <= (layer1_outputs(2551)) and not (layer1_outputs(3597));
    layer2_outputs(6289) <= (layer1_outputs(7614)) and not (layer1_outputs(8677));
    layer2_outputs(6290) <= layer1_outputs(812);
    layer2_outputs(6291) <= layer1_outputs(9493);
    layer2_outputs(6292) <= not((layer1_outputs(8332)) xor (layer1_outputs(2759)));
    layer2_outputs(6293) <= not(layer1_outputs(1038)) or (layer1_outputs(6207));
    layer2_outputs(6294) <= layer1_outputs(933);
    layer2_outputs(6295) <= not(layer1_outputs(3097));
    layer2_outputs(6296) <= not(layer1_outputs(2615));
    layer2_outputs(6297) <= (layer1_outputs(8374)) xor (layer1_outputs(6323));
    layer2_outputs(6298) <= not(layer1_outputs(6146));
    layer2_outputs(6299) <= not(layer1_outputs(9552));
    layer2_outputs(6300) <= not(layer1_outputs(4359));
    layer2_outputs(6301) <= (layer1_outputs(1906)) or (layer1_outputs(1635));
    layer2_outputs(6302) <= '1';
    layer2_outputs(6303) <= layer1_outputs(3011);
    layer2_outputs(6304) <= layer1_outputs(8484);
    layer2_outputs(6305) <= layer1_outputs(9163);
    layer2_outputs(6306) <= not(layer1_outputs(4970));
    layer2_outputs(6307) <= not(layer1_outputs(137));
    layer2_outputs(6308) <= (layer1_outputs(7252)) and not (layer1_outputs(9198));
    layer2_outputs(6309) <= layer1_outputs(10096);
    layer2_outputs(6310) <= (layer1_outputs(3971)) and (layer1_outputs(9323));
    layer2_outputs(6311) <= not(layer1_outputs(2604)) or (layer1_outputs(2637));
    layer2_outputs(6312) <= not(layer1_outputs(4392)) or (layer1_outputs(2280));
    layer2_outputs(6313) <= not(layer1_outputs(8446));
    layer2_outputs(6314) <= not(layer1_outputs(8636));
    layer2_outputs(6315) <= (layer1_outputs(2210)) and not (layer1_outputs(8364));
    layer2_outputs(6316) <= layer1_outputs(7309);
    layer2_outputs(6317) <= (layer1_outputs(3165)) or (layer1_outputs(5121));
    layer2_outputs(6318) <= layer1_outputs(2974);
    layer2_outputs(6319) <= layer1_outputs(2310);
    layer2_outputs(6320) <= layer1_outputs(7158);
    layer2_outputs(6321) <= (layer1_outputs(5413)) and (layer1_outputs(7872));
    layer2_outputs(6322) <= not(layer1_outputs(6156));
    layer2_outputs(6323) <= not(layer1_outputs(1506));
    layer2_outputs(6324) <= not(layer1_outputs(3715));
    layer2_outputs(6325) <= layer1_outputs(1518);
    layer2_outputs(6326) <= (layer1_outputs(9274)) and not (layer1_outputs(4161));
    layer2_outputs(6327) <= not((layer1_outputs(1307)) xor (layer1_outputs(3005)));
    layer2_outputs(6328) <= not(layer1_outputs(4659));
    layer2_outputs(6329) <= (layer1_outputs(1828)) and not (layer1_outputs(204));
    layer2_outputs(6330) <= not((layer1_outputs(7394)) or (layer1_outputs(6163)));
    layer2_outputs(6331) <= (layer1_outputs(743)) xor (layer1_outputs(4880));
    layer2_outputs(6332) <= (layer1_outputs(9910)) or (layer1_outputs(9100));
    layer2_outputs(6333) <= not(layer1_outputs(9307)) or (layer1_outputs(4832));
    layer2_outputs(6334) <= (layer1_outputs(7112)) or (layer1_outputs(1282));
    layer2_outputs(6335) <= (layer1_outputs(253)) xor (layer1_outputs(7789));
    layer2_outputs(6336) <= not((layer1_outputs(8206)) xor (layer1_outputs(9743)));
    layer2_outputs(6337) <= not(layer1_outputs(3761));
    layer2_outputs(6338) <= (layer1_outputs(7293)) and not (layer1_outputs(4662));
    layer2_outputs(6339) <= layer1_outputs(4123);
    layer2_outputs(6340) <= layer1_outputs(7353);
    layer2_outputs(6341) <= not((layer1_outputs(232)) xor (layer1_outputs(8709)));
    layer2_outputs(6342) <= layer1_outputs(489);
    layer2_outputs(6343) <= layer1_outputs(6987);
    layer2_outputs(6344) <= layer1_outputs(5671);
    layer2_outputs(6345) <= not(layer1_outputs(4487));
    layer2_outputs(6346) <= (layer1_outputs(9411)) and (layer1_outputs(2077));
    layer2_outputs(6347) <= not(layer1_outputs(381));
    layer2_outputs(6348) <= not(layer1_outputs(5783));
    layer2_outputs(6349) <= layer1_outputs(4846);
    layer2_outputs(6350) <= layer1_outputs(830);
    layer2_outputs(6351) <= not(layer1_outputs(3666)) or (layer1_outputs(7959));
    layer2_outputs(6352) <= not(layer1_outputs(5088));
    layer2_outputs(6353) <= not((layer1_outputs(5388)) or (layer1_outputs(2783)));
    layer2_outputs(6354) <= not(layer1_outputs(6608)) or (layer1_outputs(5164));
    layer2_outputs(6355) <= not(layer1_outputs(230));
    layer2_outputs(6356) <= not(layer1_outputs(9823)) or (layer1_outputs(7040));
    layer2_outputs(6357) <= '0';
    layer2_outputs(6358) <= not(layer1_outputs(1967));
    layer2_outputs(6359) <= not(layer1_outputs(128));
    layer2_outputs(6360) <= (layer1_outputs(2801)) and not (layer1_outputs(4570));
    layer2_outputs(6361) <= not((layer1_outputs(8271)) or (layer1_outputs(6882)));
    layer2_outputs(6362) <= (layer1_outputs(8326)) or (layer1_outputs(4657));
    layer2_outputs(6363) <= not(layer1_outputs(4002));
    layer2_outputs(6364) <= (layer1_outputs(9489)) and not (layer1_outputs(1851));
    layer2_outputs(6365) <= not(layer1_outputs(110));
    layer2_outputs(6366) <= layer1_outputs(9257);
    layer2_outputs(6367) <= not((layer1_outputs(8627)) or (layer1_outputs(7356)));
    layer2_outputs(6368) <= (layer1_outputs(10062)) and not (layer1_outputs(5237));
    layer2_outputs(6369) <= not(layer1_outputs(6394));
    layer2_outputs(6370) <= layer1_outputs(8090);
    layer2_outputs(6371) <= layer1_outputs(4935);
    layer2_outputs(6372) <= '1';
    layer2_outputs(6373) <= not(layer1_outputs(1267)) or (layer1_outputs(4277));
    layer2_outputs(6374) <= not(layer1_outputs(8505)) or (layer1_outputs(3588));
    layer2_outputs(6375) <= layer1_outputs(4435);
    layer2_outputs(6376) <= layer1_outputs(5762);
    layer2_outputs(6377) <= not(layer1_outputs(6368));
    layer2_outputs(6378) <= not(layer1_outputs(8831));
    layer2_outputs(6379) <= layer1_outputs(7022);
    layer2_outputs(6380) <= (layer1_outputs(2523)) and not (layer1_outputs(8804));
    layer2_outputs(6381) <= not(layer1_outputs(9156));
    layer2_outputs(6382) <= not(layer1_outputs(1539));
    layer2_outputs(6383) <= layer1_outputs(277);
    layer2_outputs(6384) <= layer1_outputs(5067);
    layer2_outputs(6385) <= not(layer1_outputs(9003));
    layer2_outputs(6386) <= layer1_outputs(3464);
    layer2_outputs(6387) <= layer1_outputs(2722);
    layer2_outputs(6388) <= (layer1_outputs(4219)) and not (layer1_outputs(9652));
    layer2_outputs(6389) <= not(layer1_outputs(7773)) or (layer1_outputs(8213));
    layer2_outputs(6390) <= layer1_outputs(85);
    layer2_outputs(6391) <= not(layer1_outputs(9377));
    layer2_outputs(6392) <= not(layer1_outputs(6485)) or (layer1_outputs(6847));
    layer2_outputs(6393) <= (layer1_outputs(7071)) xor (layer1_outputs(8522));
    layer2_outputs(6394) <= not(layer1_outputs(9986)) or (layer1_outputs(3188));
    layer2_outputs(6395) <= not(layer1_outputs(2925));
    layer2_outputs(6396) <= not((layer1_outputs(7373)) or (layer1_outputs(3868)));
    layer2_outputs(6397) <= (layer1_outputs(7280)) and not (layer1_outputs(2796));
    layer2_outputs(6398) <= layer1_outputs(6184);
    layer2_outputs(6399) <= layer1_outputs(8570);
    layer2_outputs(6400) <= (layer1_outputs(7978)) and not (layer1_outputs(5438));
    layer2_outputs(6401) <= not((layer1_outputs(2803)) or (layer1_outputs(1109)));
    layer2_outputs(6402) <= (layer1_outputs(2889)) or (layer1_outputs(244));
    layer2_outputs(6403) <= layer1_outputs(2149);
    layer2_outputs(6404) <= not(layer1_outputs(7024));
    layer2_outputs(6405) <= (layer1_outputs(8147)) and not (layer1_outputs(4115));
    layer2_outputs(6406) <= layer1_outputs(2139);
    layer2_outputs(6407) <= (layer1_outputs(8922)) and (layer1_outputs(3197));
    layer2_outputs(6408) <= not(layer1_outputs(3860)) or (layer1_outputs(8508));
    layer2_outputs(6409) <= not(layer1_outputs(5349));
    layer2_outputs(6410) <= layer1_outputs(5081);
    layer2_outputs(6411) <= not(layer1_outputs(9698));
    layer2_outputs(6412) <= not((layer1_outputs(9558)) xor (layer1_outputs(8672)));
    layer2_outputs(6413) <= not(layer1_outputs(2218));
    layer2_outputs(6414) <= not(layer1_outputs(3628));
    layer2_outputs(6415) <= layer1_outputs(146);
    layer2_outputs(6416) <= not(layer1_outputs(9937)) or (layer1_outputs(9872));
    layer2_outputs(6417) <= (layer1_outputs(9197)) xor (layer1_outputs(3302));
    layer2_outputs(6418) <= not(layer1_outputs(4518));
    layer2_outputs(6419) <= layer1_outputs(6811);
    layer2_outputs(6420) <= layer1_outputs(9303);
    layer2_outputs(6421) <= layer1_outputs(4186);
    layer2_outputs(6422) <= not((layer1_outputs(6195)) and (layer1_outputs(5546)));
    layer2_outputs(6423) <= (layer1_outputs(8268)) and (layer1_outputs(2005));
    layer2_outputs(6424) <= layer1_outputs(9123);
    layer2_outputs(6425) <= layer1_outputs(612);
    layer2_outputs(6426) <= not(layer1_outputs(4156)) or (layer1_outputs(5258));
    layer2_outputs(6427) <= not(layer1_outputs(9720)) or (layer1_outputs(7932));
    layer2_outputs(6428) <= not(layer1_outputs(7934)) or (layer1_outputs(5427));
    layer2_outputs(6429) <= layer1_outputs(9115);
    layer2_outputs(6430) <= layer1_outputs(3370);
    layer2_outputs(6431) <= not(layer1_outputs(4001));
    layer2_outputs(6432) <= not((layer1_outputs(10186)) xor (layer1_outputs(3475)));
    layer2_outputs(6433) <= not((layer1_outputs(5888)) and (layer1_outputs(7791)));
    layer2_outputs(6434) <= not(layer1_outputs(2696));
    layer2_outputs(6435) <= '1';
    layer2_outputs(6436) <= (layer1_outputs(8378)) or (layer1_outputs(9991));
    layer2_outputs(6437) <= (layer1_outputs(1509)) and not (layer1_outputs(4267));
    layer2_outputs(6438) <= layer1_outputs(7482);
    layer2_outputs(6439) <= not(layer1_outputs(2325));
    layer2_outputs(6440) <= (layer1_outputs(9425)) or (layer1_outputs(6055));
    layer2_outputs(6441) <= layer1_outputs(4044);
    layer2_outputs(6442) <= not(layer1_outputs(1320));
    layer2_outputs(6443) <= layer1_outputs(3124);
    layer2_outputs(6444) <= not((layer1_outputs(1393)) xor (layer1_outputs(3289)));
    layer2_outputs(6445) <= layer1_outputs(5541);
    layer2_outputs(6446) <= (layer1_outputs(8060)) or (layer1_outputs(4907));
    layer2_outputs(6447) <= (layer1_outputs(3243)) xor (layer1_outputs(6874));
    layer2_outputs(6448) <= layer1_outputs(9555);
    layer2_outputs(6449) <= (layer1_outputs(9535)) and not (layer1_outputs(7679));
    layer2_outputs(6450) <= not(layer1_outputs(5449));
    layer2_outputs(6451) <= (layer1_outputs(8787)) xor (layer1_outputs(3363));
    layer2_outputs(6452) <= not((layer1_outputs(8187)) and (layer1_outputs(3548)));
    layer2_outputs(6453) <= (layer1_outputs(1298)) or (layer1_outputs(6974));
    layer2_outputs(6454) <= not(layer1_outputs(5045));
    layer2_outputs(6455) <= layer1_outputs(1584);
    layer2_outputs(6456) <= not((layer1_outputs(8898)) and (layer1_outputs(7904)));
    layer2_outputs(6457) <= layer1_outputs(1361);
    layer2_outputs(6458) <= (layer1_outputs(34)) and (layer1_outputs(7322));
    layer2_outputs(6459) <= not(layer1_outputs(7878)) or (layer1_outputs(4920));
    layer2_outputs(6460) <= (layer1_outputs(3569)) or (layer1_outputs(2184));
    layer2_outputs(6461) <= not(layer1_outputs(9269));
    layer2_outputs(6462) <= not((layer1_outputs(7839)) xor (layer1_outputs(2779)));
    layer2_outputs(6463) <= not((layer1_outputs(10128)) or (layer1_outputs(6042)));
    layer2_outputs(6464) <= not(layer1_outputs(7100));
    layer2_outputs(6465) <= not(layer1_outputs(7752));
    layer2_outputs(6466) <= not(layer1_outputs(5379));
    layer2_outputs(6467) <= layer1_outputs(547);
    layer2_outputs(6468) <= (layer1_outputs(2099)) xor (layer1_outputs(5791));
    layer2_outputs(6469) <= layer1_outputs(6353);
    layer2_outputs(6470) <= not(layer1_outputs(3816));
    layer2_outputs(6471) <= layer1_outputs(696);
    layer2_outputs(6472) <= (layer1_outputs(9714)) and not (layer1_outputs(4103));
    layer2_outputs(6473) <= (layer1_outputs(9495)) and not (layer1_outputs(6499));
    layer2_outputs(6474) <= layer1_outputs(4297);
    layer2_outputs(6475) <= (layer1_outputs(9946)) and not (layer1_outputs(2496));
    layer2_outputs(6476) <= (layer1_outputs(3962)) or (layer1_outputs(5791));
    layer2_outputs(6477) <= not(layer1_outputs(9145));
    layer2_outputs(6478) <= layer1_outputs(9257);
    layer2_outputs(6479) <= '1';
    layer2_outputs(6480) <= (layer1_outputs(5909)) and not (layer1_outputs(9149));
    layer2_outputs(6481) <= layer1_outputs(8684);
    layer2_outputs(6482) <= not((layer1_outputs(4648)) xor (layer1_outputs(4101)));
    layer2_outputs(6483) <= not(layer1_outputs(7470));
    layer2_outputs(6484) <= (layer1_outputs(8318)) and (layer1_outputs(2870));
    layer2_outputs(6485) <= layer1_outputs(2081);
    layer2_outputs(6486) <= layer1_outputs(4578);
    layer2_outputs(6487) <= not(layer1_outputs(5367));
    layer2_outputs(6488) <= not(layer1_outputs(4));
    layer2_outputs(6489) <= (layer1_outputs(7239)) xor (layer1_outputs(9993));
    layer2_outputs(6490) <= (layer1_outputs(8019)) and not (layer1_outputs(3112));
    layer2_outputs(6491) <= not((layer1_outputs(7459)) or (layer1_outputs(2406)));
    layer2_outputs(6492) <= (layer1_outputs(73)) or (layer1_outputs(7262));
    layer2_outputs(6493) <= layer1_outputs(6740);
    layer2_outputs(6494) <= not(layer1_outputs(724));
    layer2_outputs(6495) <= not(layer1_outputs(2003));
    layer2_outputs(6496) <= not((layer1_outputs(9579)) xor (layer1_outputs(675)));
    layer2_outputs(6497) <= not(layer1_outputs(9444));
    layer2_outputs(6498) <= layer1_outputs(2688);
    layer2_outputs(6499) <= not(layer1_outputs(382));
    layer2_outputs(6500) <= (layer1_outputs(1800)) and not (layer1_outputs(2098));
    layer2_outputs(6501) <= '1';
    layer2_outputs(6502) <= (layer1_outputs(767)) or (layer1_outputs(24));
    layer2_outputs(6503) <= not(layer1_outputs(2744)) or (layer1_outputs(4533));
    layer2_outputs(6504) <= not(layer1_outputs(781));
    layer2_outputs(6505) <= (layer1_outputs(8231)) and (layer1_outputs(6953));
    layer2_outputs(6506) <= (layer1_outputs(8380)) and (layer1_outputs(2687));
    layer2_outputs(6507) <= layer1_outputs(56);
    layer2_outputs(6508) <= layer1_outputs(751);
    layer2_outputs(6509) <= not(layer1_outputs(744));
    layer2_outputs(6510) <= not(layer1_outputs(3730));
    layer2_outputs(6511) <= layer1_outputs(7116);
    layer2_outputs(6512) <= (layer1_outputs(1493)) xor (layer1_outputs(1904));
    layer2_outputs(6513) <= not(layer1_outputs(10149));
    layer2_outputs(6514) <= '1';
    layer2_outputs(6515) <= layer1_outputs(7357);
    layer2_outputs(6516) <= layer1_outputs(9066);
    layer2_outputs(6517) <= (layer1_outputs(3387)) or (layer1_outputs(7246));
    layer2_outputs(6518) <= not(layer1_outputs(5225));
    layer2_outputs(6519) <= not((layer1_outputs(1678)) xor (layer1_outputs(3421)));
    layer2_outputs(6520) <= not(layer1_outputs(22));
    layer2_outputs(6521) <= (layer1_outputs(3099)) and (layer1_outputs(9165));
    layer2_outputs(6522) <= not(layer1_outputs(8017)) or (layer1_outputs(4677));
    layer2_outputs(6523) <= not((layer1_outputs(2708)) or (layer1_outputs(9479)));
    layer2_outputs(6524) <= not((layer1_outputs(5594)) and (layer1_outputs(2778)));
    layer2_outputs(6525) <= (layer1_outputs(7630)) or (layer1_outputs(2014));
    layer2_outputs(6526) <= layer1_outputs(3264);
    layer2_outputs(6527) <= not(layer1_outputs(4011));
    layer2_outputs(6528) <= layer1_outputs(9377);
    layer2_outputs(6529) <= (layer1_outputs(5689)) or (layer1_outputs(6343));
    layer2_outputs(6530) <= not((layer1_outputs(2877)) or (layer1_outputs(1605)));
    layer2_outputs(6531) <= not(layer1_outputs(2702));
    layer2_outputs(6532) <= (layer1_outputs(2864)) and (layer1_outputs(9612));
    layer2_outputs(6533) <= layer1_outputs(7344);
    layer2_outputs(6534) <= layer1_outputs(518);
    layer2_outputs(6535) <= not(layer1_outputs(9005)) or (layer1_outputs(10183));
    layer2_outputs(6536) <= layer1_outputs(638);
    layer2_outputs(6537) <= not(layer1_outputs(3994));
    layer2_outputs(6538) <= (layer1_outputs(3714)) and not (layer1_outputs(6688));
    layer2_outputs(6539) <= not((layer1_outputs(7442)) or (layer1_outputs(7898)));
    layer2_outputs(6540) <= layer1_outputs(10040);
    layer2_outputs(6541) <= not(layer1_outputs(9985)) or (layer1_outputs(8644));
    layer2_outputs(6542) <= layer1_outputs(8907);
    layer2_outputs(6543) <= layer1_outputs(5145);
    layer2_outputs(6544) <= layer1_outputs(7046);
    layer2_outputs(6545) <= not((layer1_outputs(2892)) or (layer1_outputs(3597)));
    layer2_outputs(6546) <= layer1_outputs(5957);
    layer2_outputs(6547) <= not(layer1_outputs(4819));
    layer2_outputs(6548) <= layer1_outputs(3101);
    layer2_outputs(6549) <= not(layer1_outputs(395));
    layer2_outputs(6550) <= (layer1_outputs(9928)) and not (layer1_outputs(2824));
    layer2_outputs(6551) <= not(layer1_outputs(7907));
    layer2_outputs(6552) <= not(layer1_outputs(6680));
    layer2_outputs(6553) <= layer1_outputs(8499);
    layer2_outputs(6554) <= layer1_outputs(608);
    layer2_outputs(6555) <= layer1_outputs(7626);
    layer2_outputs(6556) <= not(layer1_outputs(9234));
    layer2_outputs(6557) <= not(layer1_outputs(5931));
    layer2_outputs(6558) <= (layer1_outputs(2383)) xor (layer1_outputs(6142));
    layer2_outputs(6559) <= layer1_outputs(2728);
    layer2_outputs(6560) <= (layer1_outputs(5925)) and (layer1_outputs(4663));
    layer2_outputs(6561) <= '1';
    layer2_outputs(6562) <= not(layer1_outputs(251));
    layer2_outputs(6563) <= not((layer1_outputs(3575)) and (layer1_outputs(2359)));
    layer2_outputs(6564) <= not(layer1_outputs(1881));
    layer2_outputs(6565) <= not(layer1_outputs(6387)) or (layer1_outputs(7737));
    layer2_outputs(6566) <= layer1_outputs(4950);
    layer2_outputs(6567) <= '1';
    layer2_outputs(6568) <= not((layer1_outputs(5669)) or (layer1_outputs(9450)));
    layer2_outputs(6569) <= (layer1_outputs(2588)) and not (layer1_outputs(9642));
    layer2_outputs(6570) <= (layer1_outputs(5205)) or (layer1_outputs(3016));
    layer2_outputs(6571) <= (layer1_outputs(7050)) and (layer1_outputs(9866));
    layer2_outputs(6572) <= layer1_outputs(6499);
    layer2_outputs(6573) <= not((layer1_outputs(8669)) and (layer1_outputs(6469)));
    layer2_outputs(6574) <= not(layer1_outputs(7443));
    layer2_outputs(6575) <= not((layer1_outputs(1553)) or (layer1_outputs(2430)));
    layer2_outputs(6576) <= layer1_outputs(8840);
    layer2_outputs(6577) <= layer1_outputs(153);
    layer2_outputs(6578) <= layer1_outputs(8634);
    layer2_outputs(6579) <= not(layer1_outputs(87));
    layer2_outputs(6580) <= '0';
    layer2_outputs(6581) <= layer1_outputs(3070);
    layer2_outputs(6582) <= not(layer1_outputs(6371));
    layer2_outputs(6583) <= not((layer1_outputs(7036)) and (layer1_outputs(3179)));
    layer2_outputs(6584) <= (layer1_outputs(1729)) or (layer1_outputs(9677));
    layer2_outputs(6585) <= layer1_outputs(1960);
    layer2_outputs(6586) <= (layer1_outputs(5551)) xor (layer1_outputs(4275));
    layer2_outputs(6587) <= not((layer1_outputs(7089)) and (layer1_outputs(8401)));
    layer2_outputs(6588) <= not(layer1_outputs(2870)) or (layer1_outputs(4826));
    layer2_outputs(6589) <= not((layer1_outputs(7121)) and (layer1_outputs(7961)));
    layer2_outputs(6590) <= not(layer1_outputs(3054));
    layer2_outputs(6591) <= not(layer1_outputs(4125));
    layer2_outputs(6592) <= (layer1_outputs(2040)) or (layer1_outputs(5873));
    layer2_outputs(6593) <= not(layer1_outputs(9756));
    layer2_outputs(6594) <= not(layer1_outputs(4943)) or (layer1_outputs(3201));
    layer2_outputs(6595) <= not(layer1_outputs(2045));
    layer2_outputs(6596) <= not((layer1_outputs(1308)) and (layer1_outputs(5525)));
    layer2_outputs(6597) <= not((layer1_outputs(2967)) and (layer1_outputs(3088)));
    layer2_outputs(6598) <= not(layer1_outputs(2918));
    layer2_outputs(6599) <= not(layer1_outputs(8172));
    layer2_outputs(6600) <= (layer1_outputs(5291)) and not (layer1_outputs(5));
    layer2_outputs(6601) <= not((layer1_outputs(3488)) and (layer1_outputs(6876)));
    layer2_outputs(6602) <= layer1_outputs(1926);
    layer2_outputs(6603) <= (layer1_outputs(9742)) and not (layer1_outputs(2854));
    layer2_outputs(6604) <= not((layer1_outputs(2531)) or (layer1_outputs(8142)));
    layer2_outputs(6605) <= (layer1_outputs(5776)) or (layer1_outputs(8098));
    layer2_outputs(6606) <= not((layer1_outputs(4358)) and (layer1_outputs(8290)));
    layer2_outputs(6607) <= not(layer1_outputs(3579));
    layer2_outputs(6608) <= not((layer1_outputs(2182)) and (layer1_outputs(8506)));
    layer2_outputs(6609) <= not(layer1_outputs(1370));
    layer2_outputs(6610) <= not(layer1_outputs(1467));
    layer2_outputs(6611) <= not((layer1_outputs(633)) xor (layer1_outputs(7029)));
    layer2_outputs(6612) <= not(layer1_outputs(7369));
    layer2_outputs(6613) <= (layer1_outputs(6374)) and (layer1_outputs(5538));
    layer2_outputs(6614) <= layer1_outputs(1875);
    layer2_outputs(6615) <= not(layer1_outputs(4973)) or (layer1_outputs(4708));
    layer2_outputs(6616) <= layer1_outputs(1892);
    layer2_outputs(6617) <= not((layer1_outputs(2144)) or (layer1_outputs(6327)));
    layer2_outputs(6618) <= (layer1_outputs(10071)) and not (layer1_outputs(5460));
    layer2_outputs(6619) <= not(layer1_outputs(7785)) or (layer1_outputs(1081));
    layer2_outputs(6620) <= not(layer1_outputs(3945));
    layer2_outputs(6621) <= not(layer1_outputs(8331));
    layer2_outputs(6622) <= layer1_outputs(613);
    layer2_outputs(6623) <= (layer1_outputs(6648)) and (layer1_outputs(6600));
    layer2_outputs(6624) <= not((layer1_outputs(8910)) xor (layer1_outputs(1144)));
    layer2_outputs(6625) <= layer1_outputs(2537);
    layer2_outputs(6626) <= not(layer1_outputs(487));
    layer2_outputs(6627) <= not(layer1_outputs(3016));
    layer2_outputs(6628) <= layer1_outputs(2231);
    layer2_outputs(6629) <= not((layer1_outputs(767)) or (layer1_outputs(9886)));
    layer2_outputs(6630) <= layer1_outputs(2623);
    layer2_outputs(6631) <= not(layer1_outputs(995));
    layer2_outputs(6632) <= (layer1_outputs(297)) xor (layer1_outputs(9536));
    layer2_outputs(6633) <= not(layer1_outputs(4279)) or (layer1_outputs(9361));
    layer2_outputs(6634) <= layer1_outputs(936);
    layer2_outputs(6635) <= not(layer1_outputs(700));
    layer2_outputs(6636) <= layer1_outputs(4128);
    layer2_outputs(6637) <= (layer1_outputs(6143)) and not (layer1_outputs(2482));
    layer2_outputs(6638) <= not(layer1_outputs(10215));
    layer2_outputs(6639) <= not(layer1_outputs(7703));
    layer2_outputs(6640) <= layer1_outputs(976);
    layer2_outputs(6641) <= not(layer1_outputs(4809));
    layer2_outputs(6642) <= (layer1_outputs(2267)) and not (layer1_outputs(7746));
    layer2_outputs(6643) <= not(layer1_outputs(1404));
    layer2_outputs(6644) <= not((layer1_outputs(254)) and (layer1_outputs(45)));
    layer2_outputs(6645) <= layer1_outputs(601);
    layer2_outputs(6646) <= (layer1_outputs(72)) or (layer1_outputs(9859));
    layer2_outputs(6647) <= (layer1_outputs(7401)) and not (layer1_outputs(8746));
    layer2_outputs(6648) <= not(layer1_outputs(7743));
    layer2_outputs(6649) <= not(layer1_outputs(6566));
    layer2_outputs(6650) <= not(layer1_outputs(4445));
    layer2_outputs(6651) <= not(layer1_outputs(4063));
    layer2_outputs(6652) <= not(layer1_outputs(2781)) or (layer1_outputs(4065));
    layer2_outputs(6653) <= not(layer1_outputs(2326));
    layer2_outputs(6654) <= (layer1_outputs(535)) or (layer1_outputs(4688));
    layer2_outputs(6655) <= layer1_outputs(4031);
    layer2_outputs(6656) <= not(layer1_outputs(9916)) or (layer1_outputs(3403));
    layer2_outputs(6657) <= layer1_outputs(527);
    layer2_outputs(6658) <= layer1_outputs(405);
    layer2_outputs(6659) <= (layer1_outputs(6601)) and (layer1_outputs(8879));
    layer2_outputs(6660) <= (layer1_outputs(117)) and (layer1_outputs(6122));
    layer2_outputs(6661) <= not((layer1_outputs(5072)) and (layer1_outputs(8182)));
    layer2_outputs(6662) <= not((layer1_outputs(722)) xor (layer1_outputs(8854)));
    layer2_outputs(6663) <= layer1_outputs(8510);
    layer2_outputs(6664) <= layer1_outputs(8417);
    layer2_outputs(6665) <= not((layer1_outputs(5735)) and (layer1_outputs(3319)));
    layer2_outputs(6666) <= not(layer1_outputs(1896));
    layer2_outputs(6667) <= layer1_outputs(1679);
    layer2_outputs(6668) <= (layer1_outputs(8597)) and (layer1_outputs(5394));
    layer2_outputs(6669) <= layer1_outputs(5565);
    layer2_outputs(6670) <= layer1_outputs(937);
    layer2_outputs(6671) <= not(layer1_outputs(9342));
    layer2_outputs(6672) <= not((layer1_outputs(4203)) and (layer1_outputs(862)));
    layer2_outputs(6673) <= not(layer1_outputs(8908)) or (layer1_outputs(1940));
    layer2_outputs(6674) <= not(layer1_outputs(4267));
    layer2_outputs(6675) <= layer1_outputs(7314);
    layer2_outputs(6676) <= layer1_outputs(4067);
    layer2_outputs(6677) <= not(layer1_outputs(8053));
    layer2_outputs(6678) <= (layer1_outputs(7450)) and not (layer1_outputs(5372));
    layer2_outputs(6679) <= layer1_outputs(1810);
    layer2_outputs(6680) <= layer1_outputs(4180);
    layer2_outputs(6681) <= (layer1_outputs(2902)) and not (layer1_outputs(7377));
    layer2_outputs(6682) <= (layer1_outputs(5158)) and not (layer1_outputs(3442));
    layer2_outputs(6683) <= not(layer1_outputs(9394));
    layer2_outputs(6684) <= not(layer1_outputs(1051)) or (layer1_outputs(4269));
    layer2_outputs(6685) <= layer1_outputs(6455);
    layer2_outputs(6686) <= (layer1_outputs(2234)) xor (layer1_outputs(2759));
    layer2_outputs(6687) <= not((layer1_outputs(8763)) xor (layer1_outputs(6750)));
    layer2_outputs(6688) <= not(layer1_outputs(7899));
    layer2_outputs(6689) <= not(layer1_outputs(1939)) or (layer1_outputs(4033));
    layer2_outputs(6690) <= (layer1_outputs(6230)) and (layer1_outputs(4586));
    layer2_outputs(6691) <= not((layer1_outputs(279)) or (layer1_outputs(3323)));
    layer2_outputs(6692) <= layer1_outputs(5068);
    layer2_outputs(6693) <= '1';
    layer2_outputs(6694) <= not(layer1_outputs(6546));
    layer2_outputs(6695) <= layer1_outputs(2082);
    layer2_outputs(6696) <= (layer1_outputs(5168)) or (layer1_outputs(2617));
    layer2_outputs(6697) <= (layer1_outputs(1157)) and (layer1_outputs(377));
    layer2_outputs(6698) <= (layer1_outputs(5287)) xor (layer1_outputs(800));
    layer2_outputs(6699) <= not(layer1_outputs(4580));
    layer2_outputs(6700) <= not(layer1_outputs(8727));
    layer2_outputs(6701) <= layer1_outputs(4423);
    layer2_outputs(6702) <= layer1_outputs(896);
    layer2_outputs(6703) <= layer1_outputs(3405);
    layer2_outputs(6704) <= layer1_outputs(2494);
    layer2_outputs(6705) <= layer1_outputs(8827);
    layer2_outputs(6706) <= (layer1_outputs(5012)) and not (layer1_outputs(1062));
    layer2_outputs(6707) <= not(layer1_outputs(8524));
    layer2_outputs(6708) <= (layer1_outputs(782)) xor (layer1_outputs(7919));
    layer2_outputs(6709) <= (layer1_outputs(8950)) and not (layer1_outputs(7119));
    layer2_outputs(6710) <= not(layer1_outputs(5986));
    layer2_outputs(6711) <= not(layer1_outputs(182));
    layer2_outputs(6712) <= (layer1_outputs(8657)) xor (layer1_outputs(2284));
    layer2_outputs(6713) <= not(layer1_outputs(2969));
    layer2_outputs(6714) <= not(layer1_outputs(185)) or (layer1_outputs(9014));
    layer2_outputs(6715) <= not((layer1_outputs(1692)) or (layer1_outputs(6452)));
    layer2_outputs(6716) <= layer1_outputs(814);
    layer2_outputs(6717) <= layer1_outputs(8660);
    layer2_outputs(6718) <= not((layer1_outputs(2319)) and (layer1_outputs(9508)));
    layer2_outputs(6719) <= (layer1_outputs(964)) and not (layer1_outputs(7338));
    layer2_outputs(6720) <= not((layer1_outputs(727)) or (layer1_outputs(7764)));
    layer2_outputs(6721) <= (layer1_outputs(8906)) xor (layer1_outputs(2072));
    layer2_outputs(6722) <= layer1_outputs(7241);
    layer2_outputs(6723) <= not((layer1_outputs(382)) and (layer1_outputs(8752)));
    layer2_outputs(6724) <= (layer1_outputs(6372)) xor (layer1_outputs(10103));
    layer2_outputs(6725) <= (layer1_outputs(9901)) and (layer1_outputs(2273));
    layer2_outputs(6726) <= not(layer1_outputs(426));
    layer2_outputs(6727) <= (layer1_outputs(278)) and not (layer1_outputs(3429));
    layer2_outputs(6728) <= not(layer1_outputs(258));
    layer2_outputs(6729) <= (layer1_outputs(5267)) and (layer1_outputs(2195));
    layer2_outputs(6730) <= layer1_outputs(5804);
    layer2_outputs(6731) <= (layer1_outputs(9525)) or (layer1_outputs(903));
    layer2_outputs(6732) <= layer1_outputs(7149);
    layer2_outputs(6733) <= layer1_outputs(3435);
    layer2_outputs(6734) <= not(layer1_outputs(2364));
    layer2_outputs(6735) <= not(layer1_outputs(4958)) or (layer1_outputs(9286));
    layer2_outputs(6736) <= not(layer1_outputs(2886));
    layer2_outputs(6737) <= layer1_outputs(2994);
    layer2_outputs(6738) <= not(layer1_outputs(8961));
    layer2_outputs(6739) <= not(layer1_outputs(9145));
    layer2_outputs(6740) <= not(layer1_outputs(1446)) or (layer1_outputs(4525));
    layer2_outputs(6741) <= layer1_outputs(8271);
    layer2_outputs(6742) <= (layer1_outputs(2467)) and (layer1_outputs(3055));
    layer2_outputs(6743) <= layer1_outputs(7288);
    layer2_outputs(6744) <= layer1_outputs(6118);
    layer2_outputs(6745) <= layer1_outputs(711);
    layer2_outputs(6746) <= layer1_outputs(7074);
    layer2_outputs(6747) <= layer1_outputs(8293);
    layer2_outputs(6748) <= layer1_outputs(10130);
    layer2_outputs(6749) <= not(layer1_outputs(1624));
    layer2_outputs(6750) <= not(layer1_outputs(1519)) or (layer1_outputs(9982));
    layer2_outputs(6751) <= (layer1_outputs(3586)) and (layer1_outputs(7047));
    layer2_outputs(6752) <= not((layer1_outputs(5123)) and (layer1_outputs(1128)));
    layer2_outputs(6753) <= (layer1_outputs(5825)) xor (layer1_outputs(628));
    layer2_outputs(6754) <= layer1_outputs(3983);
    layer2_outputs(6755) <= layer1_outputs(8037);
    layer2_outputs(6756) <= layer1_outputs(1245);
    layer2_outputs(6757) <= not((layer1_outputs(6530)) xor (layer1_outputs(4414)));
    layer2_outputs(6758) <= not(layer1_outputs(3141));
    layer2_outputs(6759) <= not(layer1_outputs(699));
    layer2_outputs(6760) <= layer1_outputs(5449);
    layer2_outputs(6761) <= layer1_outputs(7454);
    layer2_outputs(6762) <= not(layer1_outputs(5930));
    layer2_outputs(6763) <= not(layer1_outputs(438));
    layer2_outputs(6764) <= not((layer1_outputs(3024)) or (layer1_outputs(9315)));
    layer2_outputs(6765) <= not(layer1_outputs(8868));
    layer2_outputs(6766) <= not((layer1_outputs(1977)) or (layer1_outputs(6907)));
    layer2_outputs(6767) <= layer1_outputs(4712);
    layer2_outputs(6768) <= layer1_outputs(1371);
    layer2_outputs(6769) <= (layer1_outputs(5921)) xor (layer1_outputs(4796));
    layer2_outputs(6770) <= (layer1_outputs(9186)) xor (layer1_outputs(9941));
    layer2_outputs(6771) <= not(layer1_outputs(4934)) or (layer1_outputs(5215));
    layer2_outputs(6772) <= not(layer1_outputs(10114));
    layer2_outputs(6773) <= not((layer1_outputs(2674)) xor (layer1_outputs(10139)));
    layer2_outputs(6774) <= (layer1_outputs(1710)) xor (layer1_outputs(4976));
    layer2_outputs(6775) <= (layer1_outputs(7697)) and not (layer1_outputs(8565));
    layer2_outputs(6776) <= not(layer1_outputs(4225));
    layer2_outputs(6777) <= not(layer1_outputs(4759));
    layer2_outputs(6778) <= layer1_outputs(8718);
    layer2_outputs(6779) <= not((layer1_outputs(2341)) or (layer1_outputs(7925)));
    layer2_outputs(6780) <= not(layer1_outputs(5416));
    layer2_outputs(6781) <= layer1_outputs(5918);
    layer2_outputs(6782) <= layer1_outputs(6563);
    layer2_outputs(6783) <= layer1_outputs(3472);
    layer2_outputs(6784) <= layer1_outputs(444);
    layer2_outputs(6785) <= not((layer1_outputs(5047)) xor (layer1_outputs(6814)));
    layer2_outputs(6786) <= (layer1_outputs(5525)) or (layer1_outputs(9339));
    layer2_outputs(6787) <= (layer1_outputs(523)) and not (layer1_outputs(742));
    layer2_outputs(6788) <= layer1_outputs(6087);
    layer2_outputs(6789) <= not(layer1_outputs(1662));
    layer2_outputs(6790) <= not(layer1_outputs(6655)) or (layer1_outputs(8447));
    layer2_outputs(6791) <= (layer1_outputs(4426)) and not (layer1_outputs(9015));
    layer2_outputs(6792) <= not((layer1_outputs(8685)) and (layer1_outputs(8861)));
    layer2_outputs(6793) <= not(layer1_outputs(8699));
    layer2_outputs(6794) <= not(layer1_outputs(7662));
    layer2_outputs(6795) <= not((layer1_outputs(3533)) and (layer1_outputs(8599)));
    layer2_outputs(6796) <= not((layer1_outputs(7469)) xor (layer1_outputs(316)));
    layer2_outputs(6797) <= not((layer1_outputs(6601)) xor (layer1_outputs(9453)));
    layer2_outputs(6798) <= not(layer1_outputs(5465));
    layer2_outputs(6799) <= not((layer1_outputs(8696)) xor (layer1_outputs(5138)));
    layer2_outputs(6800) <= not((layer1_outputs(5002)) or (layer1_outputs(9203)));
    layer2_outputs(6801) <= not(layer1_outputs(1590)) or (layer1_outputs(4777));
    layer2_outputs(6802) <= not(layer1_outputs(8845));
    layer2_outputs(6803) <= layer1_outputs(2579);
    layer2_outputs(6804) <= not((layer1_outputs(4227)) and (layer1_outputs(5850)));
    layer2_outputs(6805) <= (layer1_outputs(4002)) or (layer1_outputs(7801));
    layer2_outputs(6806) <= not(layer1_outputs(1129));
    layer2_outputs(6807) <= layer1_outputs(2542);
    layer2_outputs(6808) <= '1';
    layer2_outputs(6809) <= (layer1_outputs(9630)) and not (layer1_outputs(6725));
    layer2_outputs(6810) <= not(layer1_outputs(481));
    layer2_outputs(6811) <= (layer1_outputs(46)) xor (layer1_outputs(581));
    layer2_outputs(6812) <= layer1_outputs(6872);
    layer2_outputs(6813) <= layer1_outputs(658);
    layer2_outputs(6814) <= '1';
    layer2_outputs(6815) <= not(layer1_outputs(8886));
    layer2_outputs(6816) <= (layer1_outputs(7505)) xor (layer1_outputs(460));
    layer2_outputs(6817) <= not((layer1_outputs(8228)) xor (layer1_outputs(9020)));
    layer2_outputs(6818) <= layer1_outputs(3464);
    layer2_outputs(6819) <= not(layer1_outputs(9712)) or (layer1_outputs(3665));
    layer2_outputs(6820) <= not(layer1_outputs(2331));
    layer2_outputs(6821) <= not(layer1_outputs(4953));
    layer2_outputs(6822) <= layer1_outputs(1233);
    layer2_outputs(6823) <= not(layer1_outputs(7204));
    layer2_outputs(6824) <= (layer1_outputs(98)) or (layer1_outputs(8421));
    layer2_outputs(6825) <= not(layer1_outputs(3879));
    layer2_outputs(6826) <= (layer1_outputs(6456)) and not (layer1_outputs(5742));
    layer2_outputs(6827) <= not((layer1_outputs(6967)) and (layer1_outputs(9484)));
    layer2_outputs(6828) <= not(layer1_outputs(6114));
    layer2_outputs(6829) <= not((layer1_outputs(7392)) and (layer1_outputs(6730)));
    layer2_outputs(6830) <= layer1_outputs(4480);
    layer2_outputs(6831) <= layer1_outputs(4566);
    layer2_outputs(6832) <= not(layer1_outputs(1654));
    layer2_outputs(6833) <= (layer1_outputs(8842)) or (layer1_outputs(9192));
    layer2_outputs(6834) <= (layer1_outputs(4402)) or (layer1_outputs(8262));
    layer2_outputs(6835) <= not(layer1_outputs(9270));
    layer2_outputs(6836) <= layer1_outputs(1074);
    layer2_outputs(6837) <= not(layer1_outputs(10083));
    layer2_outputs(6838) <= not(layer1_outputs(9852));
    layer2_outputs(6839) <= not(layer1_outputs(9911)) or (layer1_outputs(9356));
    layer2_outputs(6840) <= layer1_outputs(9635);
    layer2_outputs(6841) <= not(layer1_outputs(2995));
    layer2_outputs(6842) <= not((layer1_outputs(5387)) xor (layer1_outputs(3824)));
    layer2_outputs(6843) <= not(layer1_outputs(3353));
    layer2_outputs(6844) <= not(layer1_outputs(1659));
    layer2_outputs(6845) <= not(layer1_outputs(1617));
    layer2_outputs(6846) <= layer1_outputs(6871);
    layer2_outputs(6847) <= not(layer1_outputs(8895));
    layer2_outputs(6848) <= not(layer1_outputs(10239));
    layer2_outputs(6849) <= not(layer1_outputs(8034)) or (layer1_outputs(5677));
    layer2_outputs(6850) <= not((layer1_outputs(2126)) or (layer1_outputs(837)));
    layer2_outputs(6851) <= not(layer1_outputs(9545));
    layer2_outputs(6852) <= layer1_outputs(5196);
    layer2_outputs(6853) <= layer1_outputs(7383);
    layer2_outputs(6854) <= not(layer1_outputs(6460)) or (layer1_outputs(4214));
    layer2_outputs(6855) <= layer1_outputs(9788);
    layer2_outputs(6856) <= not(layer1_outputs(5606));
    layer2_outputs(6857) <= layer1_outputs(3351);
    layer2_outputs(6858) <= not(layer1_outputs(129));
    layer2_outputs(6859) <= (layer1_outputs(9547)) and not (layer1_outputs(7147));
    layer2_outputs(6860) <= (layer1_outputs(3304)) xor (layer1_outputs(10067));
    layer2_outputs(6861) <= layer1_outputs(4966);
    layer2_outputs(6862) <= layer1_outputs(9053);
    layer2_outputs(6863) <= layer1_outputs(5153);
    layer2_outputs(6864) <= (layer1_outputs(10000)) and not (layer1_outputs(4059));
    layer2_outputs(6865) <= not((layer1_outputs(3623)) xor (layer1_outputs(1469)));
    layer2_outputs(6866) <= not(layer1_outputs(1218)) or (layer1_outputs(4854));
    layer2_outputs(6867) <= layer1_outputs(8673);
    layer2_outputs(6868) <= layer1_outputs(1781);
    layer2_outputs(6869) <= layer1_outputs(7952);
    layer2_outputs(6870) <= (layer1_outputs(8356)) xor (layer1_outputs(4709));
    layer2_outputs(6871) <= layer1_outputs(3359);
    layer2_outputs(6872) <= (layer1_outputs(8404)) and not (layer1_outputs(5896));
    layer2_outputs(6873) <= (layer1_outputs(8203)) and not (layer1_outputs(9000));
    layer2_outputs(6874) <= (layer1_outputs(6603)) and not (layer1_outputs(1960));
    layer2_outputs(6875) <= layer1_outputs(5043);
    layer2_outputs(6876) <= layer1_outputs(6741);
    layer2_outputs(6877) <= '0';
    layer2_outputs(6878) <= not(layer1_outputs(5773));
    layer2_outputs(6879) <= layer1_outputs(4977);
    layer2_outputs(6880) <= not((layer1_outputs(6795)) and (layer1_outputs(6489)));
    layer2_outputs(6881) <= not(layer1_outputs(6495));
    layer2_outputs(6882) <= layer1_outputs(1232);
    layer2_outputs(6883) <= layer1_outputs(6024);
    layer2_outputs(6884) <= layer1_outputs(3749);
    layer2_outputs(6885) <= not((layer1_outputs(4303)) xor (layer1_outputs(9404)));
    layer2_outputs(6886) <= layer1_outputs(6103);
    layer2_outputs(6887) <= not((layer1_outputs(8680)) and (layer1_outputs(568)));
    layer2_outputs(6888) <= layer1_outputs(6397);
    layer2_outputs(6889) <= not(layer1_outputs(6691)) or (layer1_outputs(6509));
    layer2_outputs(6890) <= (layer1_outputs(5917)) and not (layer1_outputs(1178));
    layer2_outputs(6891) <= layer1_outputs(3782);
    layer2_outputs(6892) <= (layer1_outputs(1502)) and not (layer1_outputs(2173));
    layer2_outputs(6893) <= not(layer1_outputs(9293)) or (layer1_outputs(557));
    layer2_outputs(6894) <= not(layer1_outputs(1365)) or (layer1_outputs(5029));
    layer2_outputs(6895) <= not(layer1_outputs(945)) or (layer1_outputs(4449));
    layer2_outputs(6896) <= not(layer1_outputs(5021));
    layer2_outputs(6897) <= (layer1_outputs(2821)) and not (layer1_outputs(6653));
    layer2_outputs(6898) <= (layer1_outputs(6982)) and (layer1_outputs(6966));
    layer2_outputs(6899) <= (layer1_outputs(7647)) and not (layer1_outputs(9752));
    layer2_outputs(6900) <= (layer1_outputs(5664)) and not (layer1_outputs(4910));
    layer2_outputs(6901) <= not(layer1_outputs(7788));
    layer2_outputs(6902) <= not(layer1_outputs(6523)) or (layer1_outputs(1607));
    layer2_outputs(6903) <= not(layer1_outputs(2127));
    layer2_outputs(6904) <= (layer1_outputs(126)) xor (layer1_outputs(3415));
    layer2_outputs(6905) <= layer1_outputs(3773);
    layer2_outputs(6906) <= not(layer1_outputs(3599)) or (layer1_outputs(578));
    layer2_outputs(6907) <= (layer1_outputs(10120)) or (layer1_outputs(7302));
    layer2_outputs(6908) <= not(layer1_outputs(9562));
    layer2_outputs(6909) <= (layer1_outputs(9417)) and not (layer1_outputs(9837));
    layer2_outputs(6910) <= not(layer1_outputs(2459));
    layer2_outputs(6911) <= layer1_outputs(3509);
    layer2_outputs(6912) <= not((layer1_outputs(7851)) xor (layer1_outputs(4747)));
    layer2_outputs(6913) <= not(layer1_outputs(5333));
    layer2_outputs(6914) <= not((layer1_outputs(10066)) and (layer1_outputs(8818)));
    layer2_outputs(6915) <= (layer1_outputs(227)) and not (layer1_outputs(1414));
    layer2_outputs(6916) <= not((layer1_outputs(8583)) xor (layer1_outputs(3775)));
    layer2_outputs(6917) <= layer1_outputs(652);
    layer2_outputs(6918) <= (layer1_outputs(2155)) and not (layer1_outputs(1266));
    layer2_outputs(6919) <= not(layer1_outputs(8834));
    layer2_outputs(6920) <= layer1_outputs(8787);
    layer2_outputs(6921) <= not(layer1_outputs(4276));
    layer2_outputs(6922) <= not(layer1_outputs(1079));
    layer2_outputs(6923) <= layer1_outputs(8569);
    layer2_outputs(6924) <= not((layer1_outputs(5891)) xor (layer1_outputs(6946)));
    layer2_outputs(6925) <= not(layer1_outputs(652)) or (layer1_outputs(8533));
    layer2_outputs(6926) <= layer1_outputs(983);
    layer2_outputs(6927) <= not((layer1_outputs(8722)) or (layer1_outputs(9748)));
    layer2_outputs(6928) <= (layer1_outputs(4697)) xor (layer1_outputs(6990));
    layer2_outputs(6929) <= '0';
    layer2_outputs(6930) <= not((layer1_outputs(749)) or (layer1_outputs(4732)));
    layer2_outputs(6931) <= not((layer1_outputs(2137)) xor (layer1_outputs(10126)));
    layer2_outputs(6932) <= not(layer1_outputs(3835));
    layer2_outputs(6933) <= not(layer1_outputs(4463));
    layer2_outputs(6934) <= not(layer1_outputs(1815));
    layer2_outputs(6935) <= not(layer1_outputs(6516));
    layer2_outputs(6936) <= layer1_outputs(5763);
    layer2_outputs(6937) <= not(layer1_outputs(3995));
    layer2_outputs(6938) <= layer1_outputs(5826);
    layer2_outputs(6939) <= layer1_outputs(3510);
    layer2_outputs(6940) <= not(layer1_outputs(7360)) or (layer1_outputs(7475));
    layer2_outputs(6941) <= not(layer1_outputs(6647));
    layer2_outputs(6942) <= (layer1_outputs(631)) xor (layer1_outputs(5494));
    layer2_outputs(6943) <= not(layer1_outputs(3609));
    layer2_outputs(6944) <= not(layer1_outputs(668));
    layer2_outputs(6945) <= not(layer1_outputs(531));
    layer2_outputs(6946) <= not(layer1_outputs(9027));
    layer2_outputs(6947) <= not(layer1_outputs(6772));
    layer2_outputs(6948) <= layer1_outputs(8755);
    layer2_outputs(6949) <= (layer1_outputs(7480)) or (layer1_outputs(7362));
    layer2_outputs(6950) <= (layer1_outputs(9438)) and (layer1_outputs(10043));
    layer2_outputs(6951) <= layer1_outputs(4229);
    layer2_outputs(6952) <= not(layer1_outputs(3915));
    layer2_outputs(6953) <= not((layer1_outputs(5218)) xor (layer1_outputs(44)));
    layer2_outputs(6954) <= not(layer1_outputs(3875));
    layer2_outputs(6955) <= layer1_outputs(1005);
    layer2_outputs(6956) <= not(layer1_outputs(7207)) or (layer1_outputs(539));
    layer2_outputs(6957) <= (layer1_outputs(2248)) and not (layer1_outputs(9584));
    layer2_outputs(6958) <= not(layer1_outputs(4384));
    layer2_outputs(6959) <= layer1_outputs(3648);
    layer2_outputs(6960) <= not((layer1_outputs(2861)) xor (layer1_outputs(707)));
    layer2_outputs(6961) <= (layer1_outputs(9795)) xor (layer1_outputs(4012));
    layer2_outputs(6962) <= layer1_outputs(7255);
    layer2_outputs(6963) <= layer1_outputs(4910);
    layer2_outputs(6964) <= not(layer1_outputs(7254));
    layer2_outputs(6965) <= (layer1_outputs(8226)) or (layer1_outputs(9604));
    layer2_outputs(6966) <= (layer1_outputs(3365)) xor (layer1_outputs(6410));
    layer2_outputs(6967) <= (layer1_outputs(9813)) xor (layer1_outputs(3484));
    layer2_outputs(6968) <= '1';
    layer2_outputs(6969) <= not(layer1_outputs(7753)) or (layer1_outputs(3883));
    layer2_outputs(6970) <= (layer1_outputs(3633)) and (layer1_outputs(8407));
    layer2_outputs(6971) <= not(layer1_outputs(3152));
    layer2_outputs(6972) <= not(layer1_outputs(1356));
    layer2_outputs(6973) <= layer1_outputs(4428);
    layer2_outputs(6974) <= (layer1_outputs(393)) and not (layer1_outputs(9664));
    layer2_outputs(6975) <= not(layer1_outputs(5796));
    layer2_outputs(6976) <= not(layer1_outputs(540));
    layer2_outputs(6977) <= layer1_outputs(4536);
    layer2_outputs(6978) <= layer1_outputs(2489);
    layer2_outputs(6979) <= not((layer1_outputs(7122)) or (layer1_outputs(5892)));
    layer2_outputs(6980) <= (layer1_outputs(7635)) and not (layer1_outputs(3718));
    layer2_outputs(6981) <= not(layer1_outputs(9701));
    layer2_outputs(6982) <= not(layer1_outputs(7754));
    layer2_outputs(6983) <= (layer1_outputs(1761)) and not (layer1_outputs(4678));
    layer2_outputs(6984) <= layer1_outputs(8948);
    layer2_outputs(6985) <= not((layer1_outputs(3738)) xor (layer1_outputs(3988)));
    layer2_outputs(6986) <= not(layer1_outputs(2320));
    layer2_outputs(6987) <= layer1_outputs(5889);
    layer2_outputs(6988) <= layer1_outputs(4588);
    layer2_outputs(6989) <= layer1_outputs(4014);
    layer2_outputs(6990) <= not(layer1_outputs(8693)) or (layer1_outputs(8547));
    layer2_outputs(6991) <= not(layer1_outputs(6845));
    layer2_outputs(6992) <= (layer1_outputs(732)) or (layer1_outputs(5236));
    layer2_outputs(6993) <= not((layer1_outputs(4450)) and (layer1_outputs(3701)));
    layer2_outputs(6994) <= not(layer1_outputs(6401)) or (layer1_outputs(2941));
    layer2_outputs(6995) <= not(layer1_outputs(8765));
    layer2_outputs(6996) <= layer1_outputs(2480);
    layer2_outputs(6997) <= layer1_outputs(4626);
    layer2_outputs(6998) <= layer1_outputs(1770);
    layer2_outputs(6999) <= not((layer1_outputs(2832)) xor (layer1_outputs(4998)));
    layer2_outputs(7000) <= (layer1_outputs(6787)) and not (layer1_outputs(9940));
    layer2_outputs(7001) <= layer1_outputs(895);
    layer2_outputs(7002) <= not(layer1_outputs(5606));
    layer2_outputs(7003) <= not(layer1_outputs(3434));
    layer2_outputs(7004) <= not(layer1_outputs(5066));
    layer2_outputs(7005) <= layer1_outputs(6572);
    layer2_outputs(7006) <= layer1_outputs(1331);
    layer2_outputs(7007) <= (layer1_outputs(4554)) and not (layer1_outputs(2076));
    layer2_outputs(7008) <= layer1_outputs(2573);
    layer2_outputs(7009) <= layer1_outputs(857);
    layer2_outputs(7010) <= not(layer1_outputs(8930));
    layer2_outputs(7011) <= not((layer1_outputs(5392)) xor (layer1_outputs(9924)));
    layer2_outputs(7012) <= not((layer1_outputs(2508)) xor (layer1_outputs(7925)));
    layer2_outputs(7013) <= not(layer1_outputs(3501)) or (layer1_outputs(2302));
    layer2_outputs(7014) <= not(layer1_outputs(7227));
    layer2_outputs(7015) <= not(layer1_outputs(8421)) or (layer1_outputs(9140));
    layer2_outputs(7016) <= not(layer1_outputs(9617)) or (layer1_outputs(1162));
    layer2_outputs(7017) <= layer1_outputs(4645);
    layer2_outputs(7018) <= not(layer1_outputs(4309));
    layer2_outputs(7019) <= not(layer1_outputs(2169)) or (layer1_outputs(4856));
    layer2_outputs(7020) <= not(layer1_outputs(9535));
    layer2_outputs(7021) <= not(layer1_outputs(8441)) or (layer1_outputs(2655));
    layer2_outputs(7022) <= not(layer1_outputs(4253));
    layer2_outputs(7023) <= not(layer1_outputs(3534));
    layer2_outputs(7024) <= (layer1_outputs(7758)) and not (layer1_outputs(3705));
    layer2_outputs(7025) <= layer1_outputs(1466);
    layer2_outputs(7026) <= (layer1_outputs(7570)) or (layer1_outputs(7738));
    layer2_outputs(7027) <= not(layer1_outputs(257));
    layer2_outputs(7028) <= not(layer1_outputs(9821));
    layer2_outputs(7029) <= (layer1_outputs(8376)) and (layer1_outputs(923));
    layer2_outputs(7030) <= '0';
    layer2_outputs(7031) <= not(layer1_outputs(6053));
    layer2_outputs(7032) <= (layer1_outputs(4933)) and not (layer1_outputs(7842));
    layer2_outputs(7033) <= layer1_outputs(9964);
    layer2_outputs(7034) <= layer1_outputs(5390);
    layer2_outputs(7035) <= not((layer1_outputs(6668)) and (layer1_outputs(5334)));
    layer2_outputs(7036) <= not(layer1_outputs(2301)) or (layer1_outputs(1269));
    layer2_outputs(7037) <= layer1_outputs(8946);
    layer2_outputs(7038) <= not(layer1_outputs(9403));
    layer2_outputs(7039) <= not(layer1_outputs(9017));
    layer2_outputs(7040) <= not(layer1_outputs(3749));
    layer2_outputs(7041) <= layer1_outputs(6442);
    layer2_outputs(7042) <= not(layer1_outputs(8621));
    layer2_outputs(7043) <= not(layer1_outputs(4370)) or (layer1_outputs(2669));
    layer2_outputs(7044) <= not(layer1_outputs(2574));
    layer2_outputs(7045) <= not((layer1_outputs(9900)) xor (layer1_outputs(8757)));
    layer2_outputs(7046) <= not(layer1_outputs(6340));
    layer2_outputs(7047) <= layer1_outputs(789);
    layer2_outputs(7048) <= layer1_outputs(6226);
    layer2_outputs(7049) <= (layer1_outputs(4539)) xor (layer1_outputs(7759));
    layer2_outputs(7050) <= not(layer1_outputs(6878));
    layer2_outputs(7051) <= not(layer1_outputs(3781));
    layer2_outputs(7052) <= layer1_outputs(6236);
    layer2_outputs(7053) <= not((layer1_outputs(1443)) xor (layer1_outputs(9567)));
    layer2_outputs(7054) <= layer1_outputs(2541);
    layer2_outputs(7055) <= (layer1_outputs(5280)) or (layer1_outputs(1119));
    layer2_outputs(7056) <= (layer1_outputs(4478)) and not (layer1_outputs(7799));
    layer2_outputs(7057) <= not(layer1_outputs(4054));
    layer2_outputs(7058) <= (layer1_outputs(5504)) and (layer1_outputs(8102));
    layer2_outputs(7059) <= not(layer1_outputs(515));
    layer2_outputs(7060) <= not(layer1_outputs(4644)) or (layer1_outputs(459));
    layer2_outputs(7061) <= layer1_outputs(30);
    layer2_outputs(7062) <= not((layer1_outputs(3538)) xor (layer1_outputs(897)));
    layer2_outputs(7063) <= not(layer1_outputs(2576));
    layer2_outputs(7064) <= layer1_outputs(294);
    layer2_outputs(7065) <= not((layer1_outputs(9999)) or (layer1_outputs(7258)));
    layer2_outputs(7066) <= not(layer1_outputs(7986));
    layer2_outputs(7067) <= layer1_outputs(10214);
    layer2_outputs(7068) <= not(layer1_outputs(6506));
    layer2_outputs(7069) <= (layer1_outputs(7079)) and (layer1_outputs(8452));
    layer2_outputs(7070) <= not((layer1_outputs(4220)) and (layer1_outputs(5441)));
    layer2_outputs(7071) <= (layer1_outputs(8893)) xor (layer1_outputs(5340));
    layer2_outputs(7072) <= (layer1_outputs(3045)) and not (layer1_outputs(2780));
    layer2_outputs(7073) <= not(layer1_outputs(3721));
    layer2_outputs(7074) <= not(layer1_outputs(6046));
    layer2_outputs(7075) <= not(layer1_outputs(9580));
    layer2_outputs(7076) <= not((layer1_outputs(6035)) xor (layer1_outputs(4514)));
    layer2_outputs(7077) <= not(layer1_outputs(2379));
    layer2_outputs(7078) <= not(layer1_outputs(6144));
    layer2_outputs(7079) <= layer1_outputs(1383);
    layer2_outputs(7080) <= not((layer1_outputs(4112)) or (layer1_outputs(3067)));
    layer2_outputs(7081) <= not(layer1_outputs(1216));
    layer2_outputs(7082) <= not((layer1_outputs(6963)) or (layer1_outputs(9664)));
    layer2_outputs(7083) <= layer1_outputs(5014);
    layer2_outputs(7084) <= not((layer1_outputs(7998)) and (layer1_outputs(7562)));
    layer2_outputs(7085) <= (layer1_outputs(4062)) xor (layer1_outputs(9484));
    layer2_outputs(7086) <= not((layer1_outputs(3632)) and (layer1_outputs(632)));
    layer2_outputs(7087) <= (layer1_outputs(8795)) and not (layer1_outputs(9557));
    layer2_outputs(7088) <= not(layer1_outputs(6367));
    layer2_outputs(7089) <= not(layer1_outputs(2715));
    layer2_outputs(7090) <= (layer1_outputs(3287)) and not (layer1_outputs(2321));
    layer2_outputs(7091) <= (layer1_outputs(3725)) xor (layer1_outputs(3753));
    layer2_outputs(7092) <= not(layer1_outputs(9266));
    layer2_outputs(7093) <= not(layer1_outputs(396));
    layer2_outputs(7094) <= layer1_outputs(3845);
    layer2_outputs(7095) <= (layer1_outputs(5640)) and (layer1_outputs(6240));
    layer2_outputs(7096) <= layer1_outputs(2775);
    layer2_outputs(7097) <= layer1_outputs(6255);
    layer2_outputs(7098) <= layer1_outputs(939);
    layer2_outputs(7099) <= not(layer1_outputs(1094));
    layer2_outputs(7100) <= (layer1_outputs(4557)) xor (layer1_outputs(8181));
    layer2_outputs(7101) <= not(layer1_outputs(6755));
    layer2_outputs(7102) <= not(layer1_outputs(3846)) or (layer1_outputs(2602));
    layer2_outputs(7103) <= not(layer1_outputs(3758));
    layer2_outputs(7104) <= (layer1_outputs(3077)) xor (layer1_outputs(4571));
    layer2_outputs(7105) <= (layer1_outputs(1177)) and (layer1_outputs(1221));
    layer2_outputs(7106) <= not(layer1_outputs(7028));
    layer2_outputs(7107) <= (layer1_outputs(5258)) and not (layer1_outputs(3374));
    layer2_outputs(7108) <= not((layer1_outputs(1289)) or (layer1_outputs(372)));
    layer2_outputs(7109) <= not((layer1_outputs(1783)) and (layer1_outputs(4481)));
    layer2_outputs(7110) <= (layer1_outputs(1230)) xor (layer1_outputs(8103));
    layer2_outputs(7111) <= not(layer1_outputs(1168));
    layer2_outputs(7112) <= layer1_outputs(2570);
    layer2_outputs(7113) <= (layer1_outputs(9912)) and not (layer1_outputs(5860));
    layer2_outputs(7114) <= not((layer1_outputs(9921)) and (layer1_outputs(2545)));
    layer2_outputs(7115) <= (layer1_outputs(1281)) xor (layer1_outputs(6925));
    layer2_outputs(7116) <= (layer1_outputs(7339)) and not (layer1_outputs(2280));
    layer2_outputs(7117) <= not(layer1_outputs(6813));
    layer2_outputs(7118) <= layer1_outputs(552);
    layer2_outputs(7119) <= layer1_outputs(2156);
    layer2_outputs(7120) <= layer1_outputs(2205);
    layer2_outputs(7121) <= not(layer1_outputs(5036));
    layer2_outputs(7122) <= not(layer1_outputs(7142));
    layer2_outputs(7123) <= (layer1_outputs(259)) and (layer1_outputs(3058));
    layer2_outputs(7124) <= not(layer1_outputs(3776));
    layer2_outputs(7125) <= not(layer1_outputs(4736));
    layer2_outputs(7126) <= (layer1_outputs(7606)) or (layer1_outputs(4335));
    layer2_outputs(7127) <= (layer1_outputs(4308)) or (layer1_outputs(6109));
    layer2_outputs(7128) <= (layer1_outputs(2328)) xor (layer1_outputs(8896));
    layer2_outputs(7129) <= '0';
    layer2_outputs(7130) <= layer1_outputs(2764);
    layer2_outputs(7131) <= not(layer1_outputs(1671)) or (layer1_outputs(3657));
    layer2_outputs(7132) <= (layer1_outputs(9662)) and not (layer1_outputs(5897));
    layer2_outputs(7133) <= not((layer1_outputs(5920)) xor (layer1_outputs(1322)));
    layer2_outputs(7134) <= not(layer1_outputs(3311));
    layer2_outputs(7135) <= (layer1_outputs(4570)) and not (layer1_outputs(2283));
    layer2_outputs(7136) <= not(layer1_outputs(7233));
    layer2_outputs(7137) <= layer1_outputs(5076);
    layer2_outputs(7138) <= not(layer1_outputs(3800));
    layer2_outputs(7139) <= (layer1_outputs(4006)) and not (layer1_outputs(620));
    layer2_outputs(7140) <= (layer1_outputs(6867)) and not (layer1_outputs(4140));
    layer2_outputs(7141) <= layer1_outputs(5323);
    layer2_outputs(7142) <= not((layer1_outputs(2603)) or (layer1_outputs(2233)));
    layer2_outputs(7143) <= not(layer1_outputs(7637)) or (layer1_outputs(770));
    layer2_outputs(7144) <= layer1_outputs(1458);
    layer2_outputs(7145) <= not(layer1_outputs(3493)) or (layer1_outputs(7323));
    layer2_outputs(7146) <= not((layer1_outputs(3491)) or (layer1_outputs(5296)));
    layer2_outputs(7147) <= not((layer1_outputs(5463)) xor (layer1_outputs(9774)));
    layer2_outputs(7148) <= not(layer1_outputs(8183));
    layer2_outputs(7149) <= not(layer1_outputs(329));
    layer2_outputs(7150) <= '0';
    layer2_outputs(7151) <= layer1_outputs(9186);
    layer2_outputs(7152) <= not((layer1_outputs(9572)) xor (layer1_outputs(8058)));
    layer2_outputs(7153) <= not(layer1_outputs(6435));
    layer2_outputs(7154) <= layer1_outputs(1774);
    layer2_outputs(7155) <= layer1_outputs(8223);
    layer2_outputs(7156) <= layer1_outputs(8338);
    layer2_outputs(7157) <= layer1_outputs(4127);
    layer2_outputs(7158) <= not((layer1_outputs(2891)) and (layer1_outputs(3247)));
    layer2_outputs(7159) <= (layer1_outputs(6262)) and (layer1_outputs(3596));
    layer2_outputs(7160) <= (layer1_outputs(991)) and not (layer1_outputs(483));
    layer2_outputs(7161) <= not(layer1_outputs(5317));
    layer2_outputs(7162) <= '0';
    layer2_outputs(7163) <= not(layer1_outputs(2045));
    layer2_outputs(7164) <= not(layer1_outputs(5835));
    layer2_outputs(7165) <= (layer1_outputs(2580)) and not (layer1_outputs(1058));
    layer2_outputs(7166) <= (layer1_outputs(5988)) and (layer1_outputs(1102));
    layer2_outputs(7167) <= not(layer1_outputs(6981)) or (layer1_outputs(8957));
    layer2_outputs(7168) <= not(layer1_outputs(4604));
    layer2_outputs(7169) <= not(layer1_outputs(4781));
    layer2_outputs(7170) <= (layer1_outputs(3463)) and not (layer1_outputs(5923));
    layer2_outputs(7171) <= not(layer1_outputs(3787));
    layer2_outputs(7172) <= not(layer1_outputs(4905));
    layer2_outputs(7173) <= layer1_outputs(6600);
    layer2_outputs(7174) <= not(layer1_outputs(6267));
    layer2_outputs(7175) <= not(layer1_outputs(4283));
    layer2_outputs(7176) <= (layer1_outputs(4610)) and (layer1_outputs(2107));
    layer2_outputs(7177) <= not(layer1_outputs(8708));
    layer2_outputs(7178) <= not(layer1_outputs(5206));
    layer2_outputs(7179) <= layer1_outputs(6982);
    layer2_outputs(7180) <= (layer1_outputs(8953)) and not (layer1_outputs(5650));
    layer2_outputs(7181) <= not(layer1_outputs(9144));
    layer2_outputs(7182) <= layer1_outputs(4689);
    layer2_outputs(7183) <= not(layer1_outputs(9376));
    layer2_outputs(7184) <= layer1_outputs(10064);
    layer2_outputs(7185) <= not(layer1_outputs(8613));
    layer2_outputs(7186) <= (layer1_outputs(855)) xor (layer1_outputs(9362));
    layer2_outputs(7187) <= not((layer1_outputs(6178)) xor (layer1_outputs(3052)));
    layer2_outputs(7188) <= not((layer1_outputs(10034)) and (layer1_outputs(348)));
    layer2_outputs(7189) <= layer1_outputs(4763);
    layer2_outputs(7190) <= not(layer1_outputs(5691));
    layer2_outputs(7191) <= layer1_outputs(170);
    layer2_outputs(7192) <= (layer1_outputs(3629)) and (layer1_outputs(9637));
    layer2_outputs(7193) <= (layer1_outputs(8157)) xor (layer1_outputs(7490));
    layer2_outputs(7194) <= not(layer1_outputs(9745)) or (layer1_outputs(7581));
    layer2_outputs(7195) <= not((layer1_outputs(8031)) xor (layer1_outputs(2481)));
    layer2_outputs(7196) <= not(layer1_outputs(9189));
    layer2_outputs(7197) <= not(layer1_outputs(4992));
    layer2_outputs(7198) <= layer1_outputs(9412);
    layer2_outputs(7199) <= (layer1_outputs(8257)) and not (layer1_outputs(7268));
    layer2_outputs(7200) <= layer1_outputs(1375);
    layer2_outputs(7201) <= layer1_outputs(3442);
    layer2_outputs(7202) <= not(layer1_outputs(2268));
    layer2_outputs(7203) <= layer1_outputs(2277);
    layer2_outputs(7204) <= (layer1_outputs(10189)) or (layer1_outputs(7791));
    layer2_outputs(7205) <= not(layer1_outputs(162));
    layer2_outputs(7206) <= (layer1_outputs(3868)) xor (layer1_outputs(3900));
    layer2_outputs(7207) <= (layer1_outputs(9043)) or (layer1_outputs(4620));
    layer2_outputs(7208) <= not(layer1_outputs(5688));
    layer2_outputs(7209) <= '1';
    layer2_outputs(7210) <= (layer1_outputs(1092)) or (layer1_outputs(6836));
    layer2_outputs(7211) <= not(layer1_outputs(9276));
    layer2_outputs(7212) <= (layer1_outputs(7049)) and not (layer1_outputs(9944));
    layer2_outputs(7213) <= layer1_outputs(8063);
    layer2_outputs(7214) <= not((layer1_outputs(6097)) and (layer1_outputs(5034)));
    layer2_outputs(7215) <= not(layer1_outputs(4812)) or (layer1_outputs(9437));
    layer2_outputs(7216) <= not(layer1_outputs(9455));
    layer2_outputs(7217) <= (layer1_outputs(4722)) xor (layer1_outputs(702));
    layer2_outputs(7218) <= layer1_outputs(5555);
    layer2_outputs(7219) <= not((layer1_outputs(5603)) and (layer1_outputs(155)));
    layer2_outputs(7220) <= (layer1_outputs(2154)) and (layer1_outputs(2610));
    layer2_outputs(7221) <= (layer1_outputs(8334)) xor (layer1_outputs(3049));
    layer2_outputs(7222) <= not(layer1_outputs(810));
    layer2_outputs(7223) <= not(layer1_outputs(7858));
    layer2_outputs(7224) <= '1';
    layer2_outputs(7225) <= not(layer1_outputs(1156));
    layer2_outputs(7226) <= not(layer1_outputs(8810));
    layer2_outputs(7227) <= (layer1_outputs(5032)) and (layer1_outputs(9985));
    layer2_outputs(7228) <= not(layer1_outputs(4320));
    layer2_outputs(7229) <= (layer1_outputs(4808)) xor (layer1_outputs(6073));
    layer2_outputs(7230) <= not(layer1_outputs(9069));
    layer2_outputs(7231) <= not(layer1_outputs(6590)) or (layer1_outputs(4188));
    layer2_outputs(7232) <= not(layer1_outputs(9022));
    layer2_outputs(7233) <= layer1_outputs(6805);
    layer2_outputs(7234) <= not(layer1_outputs(5352));
    layer2_outputs(7235) <= layer1_outputs(4277);
    layer2_outputs(7236) <= layer1_outputs(3591);
    layer2_outputs(7237) <= (layer1_outputs(7313)) and (layer1_outputs(5983));
    layer2_outputs(7238) <= not(layer1_outputs(2644));
    layer2_outputs(7239) <= not(layer1_outputs(4054));
    layer2_outputs(7240) <= not((layer1_outputs(2747)) or (layer1_outputs(5075)));
    layer2_outputs(7241) <= not((layer1_outputs(1637)) or (layer1_outputs(5837)));
    layer2_outputs(7242) <= (layer1_outputs(8508)) and not (layer1_outputs(3256));
    layer2_outputs(7243) <= not(layer1_outputs(646));
    layer2_outputs(7244) <= layer1_outputs(2556);
    layer2_outputs(7245) <= (layer1_outputs(2909)) xor (layer1_outputs(1907));
    layer2_outputs(7246) <= not((layer1_outputs(3952)) or (layer1_outputs(5024)));
    layer2_outputs(7247) <= layer1_outputs(9656);
    layer2_outputs(7248) <= (layer1_outputs(4982)) or (layer1_outputs(4176));
    layer2_outputs(7249) <= not(layer1_outputs(2316));
    layer2_outputs(7250) <= '0';
    layer2_outputs(7251) <= not(layer1_outputs(834));
    layer2_outputs(7252) <= not(layer1_outputs(2291));
    layer2_outputs(7253) <= not(layer1_outputs(891));
    layer2_outputs(7254) <= not(layer1_outputs(10191));
    layer2_outputs(7255) <= not(layer1_outputs(8243));
    layer2_outputs(7256) <= layer1_outputs(5409);
    layer2_outputs(7257) <= (layer1_outputs(3695)) and (layer1_outputs(9885));
    layer2_outputs(7258) <= not(layer1_outputs(1260));
    layer2_outputs(7259) <= layer1_outputs(9350);
    layer2_outputs(7260) <= not(layer1_outputs(4895));
    layer2_outputs(7261) <= not(layer1_outputs(2823)) or (layer1_outputs(2737));
    layer2_outputs(7262) <= not(layer1_outputs(4123));
    layer2_outputs(7263) <= layer1_outputs(5500);
    layer2_outputs(7264) <= layer1_outputs(3573);
    layer2_outputs(7265) <= not(layer1_outputs(1582)) or (layer1_outputs(3996));
    layer2_outputs(7266) <= (layer1_outputs(5544)) and not (layer1_outputs(7276));
    layer2_outputs(7267) <= not(layer1_outputs(6876)) or (layer1_outputs(3382));
    layer2_outputs(7268) <= (layer1_outputs(238)) and not (layer1_outputs(3584));
    layer2_outputs(7269) <= (layer1_outputs(1964)) and not (layer1_outputs(3834));
    layer2_outputs(7270) <= (layer1_outputs(4347)) xor (layer1_outputs(1506));
    layer2_outputs(7271) <= not(layer1_outputs(1612));
    layer2_outputs(7272) <= (layer1_outputs(5243)) and not (layer1_outputs(9080));
    layer2_outputs(7273) <= layer1_outputs(8960);
    layer2_outputs(7274) <= not(layer1_outputs(20));
    layer2_outputs(7275) <= not(layer1_outputs(5218));
    layer2_outputs(7276) <= layer1_outputs(3450);
    layer2_outputs(7277) <= (layer1_outputs(2129)) and not (layer1_outputs(9724));
    layer2_outputs(7278) <= not(layer1_outputs(7823));
    layer2_outputs(7279) <= not(layer1_outputs(6810)) or (layer1_outputs(7228));
    layer2_outputs(7280) <= not(layer1_outputs(5593));
    layer2_outputs(7281) <= (layer1_outputs(2683)) xor (layer1_outputs(7733));
    layer2_outputs(7282) <= not(layer1_outputs(6967));
    layer2_outputs(7283) <= layer1_outputs(8716);
    layer2_outputs(7284) <= (layer1_outputs(9749)) or (layer1_outputs(270));
    layer2_outputs(7285) <= not(layer1_outputs(4787));
    layer2_outputs(7286) <= (layer1_outputs(228)) xor (layer1_outputs(4375));
    layer2_outputs(7287) <= (layer1_outputs(3506)) and not (layer1_outputs(9485));
    layer2_outputs(7288) <= (layer1_outputs(8675)) and not (layer1_outputs(2358));
    layer2_outputs(7289) <= not(layer1_outputs(4918)) or (layer1_outputs(3476));
    layer2_outputs(7290) <= not(layer1_outputs(5364)) or (layer1_outputs(5346));
    layer2_outputs(7291) <= not(layer1_outputs(755));
    layer2_outputs(7292) <= layer1_outputs(2894);
    layer2_outputs(7293) <= (layer1_outputs(2925)) xor (layer1_outputs(4745));
    layer2_outputs(7294) <= layer1_outputs(6498);
    layer2_outputs(7295) <= layer1_outputs(8696);
    layer2_outputs(7296) <= layer1_outputs(6768);
    layer2_outputs(7297) <= (layer1_outputs(6625)) and not (layer1_outputs(2377));
    layer2_outputs(7298) <= layer1_outputs(3639);
    layer2_outputs(7299) <= not(layer1_outputs(9608));
    layer2_outputs(7300) <= not((layer1_outputs(5509)) xor (layer1_outputs(1085)));
    layer2_outputs(7301) <= layer1_outputs(8093);
    layer2_outputs(7302) <= not(layer1_outputs(6794));
    layer2_outputs(7303) <= not(layer1_outputs(773));
    layer2_outputs(7304) <= not(layer1_outputs(4750));
    layer2_outputs(7305) <= not(layer1_outputs(6308));
    layer2_outputs(7306) <= (layer1_outputs(4453)) xor (layer1_outputs(5729));
    layer2_outputs(7307) <= layer1_outputs(1411);
    layer2_outputs(7308) <= (layer1_outputs(8688)) and not (layer1_outputs(4981));
    layer2_outputs(7309) <= layer1_outputs(1429);
    layer2_outputs(7310) <= not((layer1_outputs(3193)) and (layer1_outputs(1390)));
    layer2_outputs(7311) <= not(layer1_outputs(7448));
    layer2_outputs(7312) <= layer1_outputs(3476);
    layer2_outputs(7313) <= not(layer1_outputs(8882));
    layer2_outputs(7314) <= not(layer1_outputs(7744));
    layer2_outputs(7315) <= not(layer1_outputs(10020));
    layer2_outputs(7316) <= not((layer1_outputs(5790)) or (layer1_outputs(5652)));
    layer2_outputs(7317) <= layer1_outputs(6534);
    layer2_outputs(7318) <= not(layer1_outputs(125));
    layer2_outputs(7319) <= not(layer1_outputs(3195));
    layer2_outputs(7320) <= not(layer1_outputs(1965));
    layer2_outputs(7321) <= (layer1_outputs(9634)) and (layer1_outputs(6442));
    layer2_outputs(7322) <= layer1_outputs(5116);
    layer2_outputs(7323) <= not(layer1_outputs(3191));
    layer2_outputs(7324) <= layer1_outputs(9268);
    layer2_outputs(7325) <= (layer1_outputs(9320)) xor (layer1_outputs(9297));
    layer2_outputs(7326) <= not(layer1_outputs(8334)) or (layer1_outputs(3008));
    layer2_outputs(7327) <= not(layer1_outputs(1613));
    layer2_outputs(7328) <= (layer1_outputs(1726)) and not (layer1_outputs(9218));
    layer2_outputs(7329) <= not(layer1_outputs(6586)) or (layer1_outputs(8601));
    layer2_outputs(7330) <= not(layer1_outputs(4572)) or (layer1_outputs(3071));
    layer2_outputs(7331) <= (layer1_outputs(5027)) xor (layer1_outputs(7577));
    layer2_outputs(7332) <= layer1_outputs(212);
    layer2_outputs(7333) <= (layer1_outputs(6159)) and not (layer1_outputs(1018));
    layer2_outputs(7334) <= not((layer1_outputs(2123)) or (layer1_outputs(1158)));
    layer2_outputs(7335) <= layer1_outputs(7642);
    layer2_outputs(7336) <= not(layer1_outputs(8504)) or (layer1_outputs(7718));
    layer2_outputs(7337) <= layer1_outputs(5029);
    layer2_outputs(7338) <= not((layer1_outputs(2948)) and (layer1_outputs(1478)));
    layer2_outputs(7339) <= (layer1_outputs(161)) and (layer1_outputs(8448));
    layer2_outputs(7340) <= (layer1_outputs(1693)) and (layer1_outputs(4243));
    layer2_outputs(7341) <= (layer1_outputs(7140)) and not (layer1_outputs(7427));
    layer2_outputs(7342) <= layer1_outputs(5336);
    layer2_outputs(7343) <= (layer1_outputs(9714)) xor (layer1_outputs(6510));
    layer2_outputs(7344) <= not(layer1_outputs(4988)) or (layer1_outputs(3936));
    layer2_outputs(7345) <= not(layer1_outputs(4113));
    layer2_outputs(7346) <= not(layer1_outputs(9202));
    layer2_outputs(7347) <= layer1_outputs(1684);
    layer2_outputs(7348) <= layer1_outputs(2257);
    layer2_outputs(7349) <= not(layer1_outputs(9713));
    layer2_outputs(7350) <= not(layer1_outputs(8247)) or (layer1_outputs(2549));
    layer2_outputs(7351) <= (layer1_outputs(2620)) or (layer1_outputs(9706));
    layer2_outputs(7352) <= not(layer1_outputs(1070));
    layer2_outputs(7353) <= (layer1_outputs(3511)) xor (layer1_outputs(7141));
    layer2_outputs(7354) <= (layer1_outputs(5519)) xor (layer1_outputs(3818));
    layer2_outputs(7355) <= not((layer1_outputs(8024)) xor (layer1_outputs(7033)));
    layer2_outputs(7356) <= not(layer1_outputs(8700));
    layer2_outputs(7357) <= (layer1_outputs(3094)) and (layer1_outputs(4893));
    layer2_outputs(7358) <= (layer1_outputs(1619)) and not (layer1_outputs(3409));
    layer2_outputs(7359) <= not(layer1_outputs(3307));
    layer2_outputs(7360) <= not((layer1_outputs(687)) xor (layer1_outputs(4499)));
    layer2_outputs(7361) <= layer1_outputs(2193);
    layer2_outputs(7362) <= not(layer1_outputs(9319));
    layer2_outputs(7363) <= not(layer1_outputs(2812));
    layer2_outputs(7364) <= not(layer1_outputs(6634));
    layer2_outputs(7365) <= (layer1_outputs(5545)) or (layer1_outputs(3214));
    layer2_outputs(7366) <= layer1_outputs(9554);
    layer2_outputs(7367) <= not((layer1_outputs(4945)) xor (layer1_outputs(365)));
    layer2_outputs(7368) <= not(layer1_outputs(10138));
    layer2_outputs(7369) <= layer1_outputs(4424);
    layer2_outputs(7370) <= (layer1_outputs(1682)) xor (layer1_outputs(6428));
    layer2_outputs(7371) <= not(layer1_outputs(1026));
    layer2_outputs(7372) <= not(layer1_outputs(255));
    layer2_outputs(7373) <= not(layer1_outputs(4603));
    layer2_outputs(7374) <= (layer1_outputs(5061)) and not (layer1_outputs(8979));
    layer2_outputs(7375) <= not((layer1_outputs(8994)) xor (layer1_outputs(10122)));
    layer2_outputs(7376) <= not(layer1_outputs(5087)) or (layer1_outputs(7171));
    layer2_outputs(7377) <= layer1_outputs(7389);
    layer2_outputs(7378) <= not((layer1_outputs(2029)) xor (layer1_outputs(8343)));
    layer2_outputs(7379) <= not((layer1_outputs(8109)) or (layer1_outputs(1277)));
    layer2_outputs(7380) <= layer1_outputs(8306);
    layer2_outputs(7381) <= layer1_outputs(1579);
    layer2_outputs(7382) <= layer1_outputs(8780);
    layer2_outputs(7383) <= layer1_outputs(5731);
    layer2_outputs(7384) <= layer1_outputs(807);
    layer2_outputs(7385) <= not((layer1_outputs(9213)) xor (layer1_outputs(8937)));
    layer2_outputs(7386) <= not(layer1_outputs(941));
    layer2_outputs(7387) <= not(layer1_outputs(137));
    layer2_outputs(7388) <= not((layer1_outputs(7361)) or (layer1_outputs(5102)));
    layer2_outputs(7389) <= not(layer1_outputs(627));
    layer2_outputs(7390) <= layer1_outputs(4698);
    layer2_outputs(7391) <= not(layer1_outputs(3210)) or (layer1_outputs(6239));
    layer2_outputs(7392) <= (layer1_outputs(5841)) and not (layer1_outputs(2950));
    layer2_outputs(7393) <= not(layer1_outputs(9041));
    layer2_outputs(7394) <= layer1_outputs(2715);
    layer2_outputs(7395) <= not(layer1_outputs(7174));
    layer2_outputs(7396) <= not(layer1_outputs(8355));
    layer2_outputs(7397) <= (layer1_outputs(7767)) xor (layer1_outputs(5924));
    layer2_outputs(7398) <= layer1_outputs(1982);
    layer2_outputs(7399) <= not((layer1_outputs(462)) xor (layer1_outputs(1187)));
    layer2_outputs(7400) <= not((layer1_outputs(7577)) or (layer1_outputs(3774)));
    layer2_outputs(7401) <= not(layer1_outputs(10199));
    layer2_outputs(7402) <= not(layer1_outputs(9118)) or (layer1_outputs(4442));
    layer2_outputs(7403) <= layer1_outputs(1830);
    layer2_outputs(7404) <= layer1_outputs(4037);
    layer2_outputs(7405) <= (layer1_outputs(4963)) and not (layer1_outputs(7173));
    layer2_outputs(7406) <= not((layer1_outputs(2629)) or (layer1_outputs(5494)));
    layer2_outputs(7407) <= layer1_outputs(1797);
    layer2_outputs(7408) <= layer1_outputs(9025);
    layer2_outputs(7409) <= not(layer1_outputs(8880));
    layer2_outputs(7410) <= not((layer1_outputs(3930)) and (layer1_outputs(1698)));
    layer2_outputs(7411) <= not((layer1_outputs(6642)) xor (layer1_outputs(424)));
    layer2_outputs(7412) <= (layer1_outputs(454)) and (layer1_outputs(5126));
    layer2_outputs(7413) <= not(layer1_outputs(5241)) or (layer1_outputs(4055));
    layer2_outputs(7414) <= layer1_outputs(4406);
    layer2_outputs(7415) <= (layer1_outputs(1845)) xor (layer1_outputs(541));
    layer2_outputs(7416) <= layer1_outputs(2794);
    layer2_outputs(7417) <= not(layer1_outputs(5101));
    layer2_outputs(7418) <= not(layer1_outputs(139));
    layer2_outputs(7419) <= (layer1_outputs(8178)) xor (layer1_outputs(3109));
    layer2_outputs(7420) <= not(layer1_outputs(4162)) or (layer1_outputs(4149));
    layer2_outputs(7421) <= not((layer1_outputs(8562)) xor (layer1_outputs(3735)));
    layer2_outputs(7422) <= not(layer1_outputs(7766));
    layer2_outputs(7423) <= layer1_outputs(2636);
    layer2_outputs(7424) <= (layer1_outputs(4027)) and not (layer1_outputs(7528));
    layer2_outputs(7425) <= not(layer1_outputs(1214)) or (layer1_outputs(2004));
    layer2_outputs(7426) <= layer1_outputs(6908);
    layer2_outputs(7427) <= (layer1_outputs(3918)) xor (layer1_outputs(3014));
    layer2_outputs(7428) <= not((layer1_outputs(326)) and (layer1_outputs(325)));
    layer2_outputs(7429) <= (layer1_outputs(4380)) and not (layer1_outputs(1224));
    layer2_outputs(7430) <= (layer1_outputs(1931)) and not (layer1_outputs(5910));
    layer2_outputs(7431) <= not(layer1_outputs(2520)) or (layer1_outputs(9352));
    layer2_outputs(7432) <= (layer1_outputs(5134)) and (layer1_outputs(6762));
    layer2_outputs(7433) <= (layer1_outputs(4195)) and not (layer1_outputs(527));
    layer2_outputs(7434) <= not(layer1_outputs(3399)) or (layer1_outputs(6245));
    layer2_outputs(7435) <= not((layer1_outputs(8802)) and (layer1_outputs(434)));
    layer2_outputs(7436) <= (layer1_outputs(6855)) or (layer1_outputs(3591));
    layer2_outputs(7437) <= (layer1_outputs(7500)) xor (layer1_outputs(9793));
    layer2_outputs(7438) <= not(layer1_outputs(3465));
    layer2_outputs(7439) <= (layer1_outputs(5362)) and not (layer1_outputs(2912));
    layer2_outputs(7440) <= not(layer1_outputs(7633));
    layer2_outputs(7441) <= layer1_outputs(3779);
    layer2_outputs(7442) <= layer1_outputs(5033);
    layer2_outputs(7443) <= layer1_outputs(7821);
    layer2_outputs(7444) <= not(layer1_outputs(66)) or (layer1_outputs(6308));
    layer2_outputs(7445) <= not(layer1_outputs(2032));
    layer2_outputs(7446) <= not(layer1_outputs(9903));
    layer2_outputs(7447) <= not((layer1_outputs(8885)) and (layer1_outputs(7327)));
    layer2_outputs(7448) <= layer1_outputs(3585);
    layer2_outputs(7449) <= not(layer1_outputs(4964)) or (layer1_outputs(4083));
    layer2_outputs(7450) <= layer1_outputs(8656);
    layer2_outputs(7451) <= layer1_outputs(9784);
    layer2_outputs(7452) <= not((layer1_outputs(455)) and (layer1_outputs(5372)));
    layer2_outputs(7453) <= layer1_outputs(259);
    layer2_outputs(7454) <= not((layer1_outputs(7314)) xor (layer1_outputs(7282)));
    layer2_outputs(7455) <= not(layer1_outputs(27));
    layer2_outputs(7456) <= not(layer1_outputs(4924)) or (layer1_outputs(3816));
    layer2_outputs(7457) <= (layer1_outputs(3665)) and not (layer1_outputs(10231));
    layer2_outputs(7458) <= layer1_outputs(9807);
    layer2_outputs(7459) <= layer1_outputs(8139);
    layer2_outputs(7460) <= not(layer1_outputs(3459));
    layer2_outputs(7461) <= (layer1_outputs(6607)) and (layer1_outputs(10033));
    layer2_outputs(7462) <= not(layer1_outputs(1453)) or (layer1_outputs(8348));
    layer2_outputs(7463) <= (layer1_outputs(6960)) and (layer1_outputs(8285));
    layer2_outputs(7464) <= not(layer1_outputs(7101));
    layer2_outputs(7465) <= layer1_outputs(8528);
    layer2_outputs(7466) <= (layer1_outputs(5765)) and not (layer1_outputs(7015));
    layer2_outputs(7467) <= not(layer1_outputs(5336));
    layer2_outputs(7468) <= (layer1_outputs(9271)) xor (layer1_outputs(7039));
    layer2_outputs(7469) <= (layer1_outputs(573)) and not (layer1_outputs(3208));
    layer2_outputs(7470) <= not(layer1_outputs(2809));
    layer2_outputs(7471) <= not(layer1_outputs(2536));
    layer2_outputs(7472) <= not((layer1_outputs(6233)) and (layer1_outputs(7844)));
    layer2_outputs(7473) <= layer1_outputs(4632);
    layer2_outputs(7474) <= layer1_outputs(78);
    layer2_outputs(7475) <= not(layer1_outputs(2249));
    layer2_outputs(7476) <= layer1_outputs(10208);
    layer2_outputs(7477) <= (layer1_outputs(4350)) or (layer1_outputs(1927));
    layer2_outputs(7478) <= not((layer1_outputs(9928)) and (layer1_outputs(8109)));
    layer2_outputs(7479) <= not(layer1_outputs(1134)) or (layer1_outputs(10131));
    layer2_outputs(7480) <= (layer1_outputs(436)) xor (layer1_outputs(9658));
    layer2_outputs(7481) <= layer1_outputs(7483);
    layer2_outputs(7482) <= layer1_outputs(5922);
    layer2_outputs(7483) <= not(layer1_outputs(772));
    layer2_outputs(7484) <= not(layer1_outputs(5437));
    layer2_outputs(7485) <= layer1_outputs(9429);
    layer2_outputs(7486) <= layer1_outputs(4985);
    layer2_outputs(7487) <= layer1_outputs(3976);
    layer2_outputs(7488) <= not(layer1_outputs(388));
    layer2_outputs(7489) <= (layer1_outputs(5182)) and not (layer1_outputs(2041));
    layer2_outputs(7490) <= not(layer1_outputs(2642));
    layer2_outputs(7491) <= layer1_outputs(7215);
    layer2_outputs(7492) <= not(layer1_outputs(3956));
    layer2_outputs(7493) <= not(layer1_outputs(6986)) or (layer1_outputs(7548));
    layer2_outputs(7494) <= layer1_outputs(6229);
    layer2_outputs(7495) <= not((layer1_outputs(2825)) or (layer1_outputs(5332)));
    layer2_outputs(7496) <= not(layer1_outputs(815));
    layer2_outputs(7497) <= not((layer1_outputs(2701)) or (layer1_outputs(5995)));
    layer2_outputs(7498) <= layer1_outputs(4024);
    layer2_outputs(7499) <= not(layer1_outputs(838));
    layer2_outputs(7500) <= not(layer1_outputs(6717));
    layer2_outputs(7501) <= not(layer1_outputs(1987));
    layer2_outputs(7502) <= not(layer1_outputs(602));
    layer2_outputs(7503) <= (layer1_outputs(8423)) and (layer1_outputs(6284));
    layer2_outputs(7504) <= layer1_outputs(8546);
    layer2_outputs(7505) <= (layer1_outputs(10050)) and (layer1_outputs(1408));
    layer2_outputs(7506) <= (layer1_outputs(3324)) and (layer1_outputs(4491));
    layer2_outputs(7507) <= layer1_outputs(1071);
    layer2_outputs(7508) <= not(layer1_outputs(3344));
    layer2_outputs(7509) <= layer1_outputs(6542);
    layer2_outputs(7510) <= '1';
    layer2_outputs(7511) <= not((layer1_outputs(6812)) or (layer1_outputs(1187)));
    layer2_outputs(7512) <= (layer1_outputs(6470)) and not (layer1_outputs(3969));
    layer2_outputs(7513) <= not(layer1_outputs(4535));
    layer2_outputs(7514) <= layer1_outputs(1837);
    layer2_outputs(7515) <= layer1_outputs(7013);
    layer2_outputs(7516) <= not((layer1_outputs(6015)) or (layer1_outputs(965)));
    layer2_outputs(7517) <= not(layer1_outputs(8011));
    layer2_outputs(7518) <= layer1_outputs(10118);
    layer2_outputs(7519) <= layer1_outputs(614);
    layer2_outputs(7520) <= layer1_outputs(3458);
    layer2_outputs(7521) <= not(layer1_outputs(4531)) or (layer1_outputs(7009));
    layer2_outputs(7522) <= layer1_outputs(5432);
    layer2_outputs(7523) <= layer1_outputs(583);
    layer2_outputs(7524) <= (layer1_outputs(7521)) and not (layer1_outputs(3794));
    layer2_outputs(7525) <= not((layer1_outputs(7970)) xor (layer1_outputs(6074)));
    layer2_outputs(7526) <= not((layer1_outputs(5705)) xor (layer1_outputs(3280)));
    layer2_outputs(7527) <= layer1_outputs(2121);
    layer2_outputs(7528) <= (layer1_outputs(5848)) and (layer1_outputs(1494));
    layer2_outputs(7529) <= (layer1_outputs(61)) and not (layer1_outputs(3156));
    layer2_outputs(7530) <= layer1_outputs(9102);
    layer2_outputs(7531) <= (layer1_outputs(7482)) and (layer1_outputs(1603));
    layer2_outputs(7532) <= layer1_outputs(471);
    layer2_outputs(7533) <= layer1_outputs(1601);
    layer2_outputs(7534) <= layer1_outputs(4155);
    layer2_outputs(7535) <= layer1_outputs(5119);
    layer2_outputs(7536) <= not(layer1_outputs(5148));
    layer2_outputs(7537) <= layer1_outputs(8982);
    layer2_outputs(7538) <= layer1_outputs(9430);
    layer2_outputs(7539) <= layer1_outputs(9973);
    layer2_outputs(7540) <= (layer1_outputs(4785)) or (layer1_outputs(5974));
    layer2_outputs(7541) <= not((layer1_outputs(3418)) xor (layer1_outputs(2926)));
    layer2_outputs(7542) <= not((layer1_outputs(7417)) xor (layer1_outputs(5685)));
    layer2_outputs(7543) <= not(layer1_outputs(5194)) or (layer1_outputs(3347));
    layer2_outputs(7544) <= layer1_outputs(8406);
    layer2_outputs(7545) <= not((layer1_outputs(777)) and (layer1_outputs(9834)));
    layer2_outputs(7546) <= not(layer1_outputs(2555)) or (layer1_outputs(8209));
    layer2_outputs(7547) <= not(layer1_outputs(6234));
    layer2_outputs(7548) <= layer1_outputs(10030);
    layer2_outputs(7549) <= layer1_outputs(4823);
    layer2_outputs(7550) <= (layer1_outputs(413)) or (layer1_outputs(4228));
    layer2_outputs(7551) <= not((layer1_outputs(6206)) or (layer1_outputs(5254)));
    layer2_outputs(7552) <= layer1_outputs(41);
    layer2_outputs(7553) <= not((layer1_outputs(4087)) xor (layer1_outputs(3681)));
    layer2_outputs(7554) <= not(layer1_outputs(5601));
    layer2_outputs(7555) <= layer1_outputs(7569);
    layer2_outputs(7556) <= (layer1_outputs(8638)) xor (layer1_outputs(1065));
    layer2_outputs(7557) <= not(layer1_outputs(7277));
    layer2_outputs(7558) <= not(layer1_outputs(5495));
    layer2_outputs(7559) <= (layer1_outputs(2760)) or (layer1_outputs(8249));
    layer2_outputs(7560) <= not(layer1_outputs(5930));
    layer2_outputs(7561) <= layer1_outputs(2648);
    layer2_outputs(7562) <= not(layer1_outputs(1430));
    layer2_outputs(7563) <= not(layer1_outputs(4510));
    layer2_outputs(7564) <= not(layer1_outputs(7331)) or (layer1_outputs(7994));
    layer2_outputs(7565) <= not((layer1_outputs(3769)) xor (layer1_outputs(8389)));
    layer2_outputs(7566) <= (layer1_outputs(8819)) or (layer1_outputs(1237));
    layer2_outputs(7567) <= layer1_outputs(1366);
    layer2_outputs(7568) <= not(layer1_outputs(10157));
    layer2_outputs(7569) <= layer1_outputs(8856);
    layer2_outputs(7570) <= not((layer1_outputs(5445)) xor (layer1_outputs(4154)));
    layer2_outputs(7571) <= layer1_outputs(10123);
    layer2_outputs(7572) <= (layer1_outputs(7166)) or (layer1_outputs(2898));
    layer2_outputs(7573) <= (layer1_outputs(4047)) xor (layer1_outputs(8726));
    layer2_outputs(7574) <= not(layer1_outputs(10050)) or (layer1_outputs(4209));
    layer2_outputs(7575) <= '0';
    layer2_outputs(7576) <= not(layer1_outputs(666));
    layer2_outputs(7577) <= not(layer1_outputs(9147));
    layer2_outputs(7578) <= layer1_outputs(8439);
    layer2_outputs(7579) <= not(layer1_outputs(427));
    layer2_outputs(7580) <= layer1_outputs(969);
    layer2_outputs(7581) <= not((layer1_outputs(5526)) xor (layer1_outputs(1633)));
    layer2_outputs(7582) <= layer1_outputs(5370);
    layer2_outputs(7583) <= (layer1_outputs(1675)) and not (layer1_outputs(3696));
    layer2_outputs(7584) <= layer1_outputs(40);
    layer2_outputs(7585) <= not(layer1_outputs(2470));
    layer2_outputs(7586) <= layer1_outputs(6579);
    layer2_outputs(7587) <= layer1_outputs(4460);
    layer2_outputs(7588) <= not(layer1_outputs(10032));
    layer2_outputs(7589) <= layer1_outputs(6078);
    layer2_outputs(7590) <= layer1_outputs(4559);
    layer2_outputs(7591) <= not(layer1_outputs(4634));
    layer2_outputs(7592) <= layer1_outputs(3145);
    layer2_outputs(7593) <= layer1_outputs(3216);
    layer2_outputs(7594) <= not(layer1_outputs(3437));
    layer2_outputs(7595) <= not(layer1_outputs(9154));
    layer2_outputs(7596) <= not(layer1_outputs(262));
    layer2_outputs(7597) <= layer1_outputs(6277);
    layer2_outputs(7598) <= (layer1_outputs(2570)) xor (layer1_outputs(10070));
    layer2_outputs(7599) <= not(layer1_outputs(5326)) or (layer1_outputs(2575));
    layer2_outputs(7600) <= not(layer1_outputs(8520)) or (layer1_outputs(8337));
    layer2_outputs(7601) <= layer1_outputs(981);
    layer2_outputs(7602) <= not(layer1_outputs(7368));
    layer2_outputs(7603) <= (layer1_outputs(8427)) and not (layer1_outputs(4356));
    layer2_outputs(7604) <= layer1_outputs(7864);
    layer2_outputs(7605) <= (layer1_outputs(1931)) xor (layer1_outputs(1755));
    layer2_outputs(7606) <= not(layer1_outputs(7257));
    layer2_outputs(7607) <= not(layer1_outputs(617)) or (layer1_outputs(6845));
    layer2_outputs(7608) <= not((layer1_outputs(7983)) or (layer1_outputs(4662)));
    layer2_outputs(7609) <= not((layer1_outputs(7092)) and (layer1_outputs(4534)));
    layer2_outputs(7610) <= layer1_outputs(3656);
    layer2_outputs(7611) <= layer1_outputs(10006);
    layer2_outputs(7612) <= not((layer1_outputs(2381)) xor (layer1_outputs(1275)));
    layer2_outputs(7613) <= (layer1_outputs(5697)) and not (layer1_outputs(8153));
    layer2_outputs(7614) <= not(layer1_outputs(2893));
    layer2_outputs(7615) <= not((layer1_outputs(1596)) xor (layer1_outputs(455)));
    layer2_outputs(7616) <= not(layer1_outputs(7222));
    layer2_outputs(7617) <= not(layer1_outputs(10148));
    layer2_outputs(7618) <= not(layer1_outputs(2058));
    layer2_outputs(7619) <= not((layer1_outputs(3641)) xor (layer1_outputs(6833)));
    layer2_outputs(7620) <= (layer1_outputs(91)) or (layer1_outputs(1235));
    layer2_outputs(7621) <= not((layer1_outputs(6590)) xor (layer1_outputs(5289)));
    layer2_outputs(7622) <= layer1_outputs(8999);
    layer2_outputs(7623) <= (layer1_outputs(8384)) and not (layer1_outputs(2020));
    layer2_outputs(7624) <= '0';
    layer2_outputs(7625) <= not(layer1_outputs(9136)) or (layer1_outputs(6498));
    layer2_outputs(7626) <= layer1_outputs(6637);
    layer2_outputs(7627) <= not(layer1_outputs(909));
    layer2_outputs(7628) <= not(layer1_outputs(2113));
    layer2_outputs(7629) <= (layer1_outputs(10099)) and not (layer1_outputs(3861));
    layer2_outputs(7630) <= layer1_outputs(8512);
    layer2_outputs(7631) <= not((layer1_outputs(8262)) or (layer1_outputs(2499)));
    layer2_outputs(7632) <= (layer1_outputs(1047)) and not (layer1_outputs(6844));
    layer2_outputs(7633) <= layer1_outputs(5799);
    layer2_outputs(7634) <= layer1_outputs(5078);
    layer2_outputs(7635) <= not(layer1_outputs(6860));
    layer2_outputs(7636) <= (layer1_outputs(3516)) and (layer1_outputs(7093));
    layer2_outputs(7637) <= (layer1_outputs(8215)) xor (layer1_outputs(4026));
    layer2_outputs(7638) <= (layer1_outputs(4578)) and not (layer1_outputs(4761));
    layer2_outputs(7639) <= not((layer1_outputs(7006)) or (layer1_outputs(8912)));
    layer2_outputs(7640) <= layer1_outputs(5130);
    layer2_outputs(7641) <= not(layer1_outputs(8050));
    layer2_outputs(7642) <= not(layer1_outputs(7306));
    layer2_outputs(7643) <= not((layer1_outputs(3161)) xor (layer1_outputs(7198)));
    layer2_outputs(7644) <= layer1_outputs(9545);
    layer2_outputs(7645) <= layer1_outputs(9697);
    layer2_outputs(7646) <= not(layer1_outputs(9199)) or (layer1_outputs(2685));
    layer2_outputs(7647) <= not(layer1_outputs(7958)) or (layer1_outputs(7920));
    layer2_outputs(7648) <= layer1_outputs(8847);
    layer2_outputs(7649) <= layer1_outputs(7230);
    layer2_outputs(7650) <= not(layer1_outputs(4995)) or (layer1_outputs(6263));
    layer2_outputs(7651) <= not(layer1_outputs(4987));
    layer2_outputs(7652) <= not(layer1_outputs(1413)) or (layer1_outputs(2234));
    layer2_outputs(7653) <= not(layer1_outputs(2396)) or (layer1_outputs(4814));
    layer2_outputs(7654) <= layer1_outputs(2407);
    layer2_outputs(7655) <= layer1_outputs(6086);
    layer2_outputs(7656) <= (layer1_outputs(6427)) xor (layer1_outputs(2887));
    layer2_outputs(7657) <= layer1_outputs(6545);
    layer2_outputs(7658) <= layer1_outputs(8425);
    layer2_outputs(7659) <= layer1_outputs(182);
    layer2_outputs(7660) <= layer1_outputs(1945);
    layer2_outputs(7661) <= layer1_outputs(6765);
    layer2_outputs(7662) <= (layer1_outputs(2964)) and not (layer1_outputs(3138));
    layer2_outputs(7663) <= layer1_outputs(1228);
    layer2_outputs(7664) <= layer1_outputs(7139);
    layer2_outputs(7665) <= not(layer1_outputs(6626));
    layer2_outputs(7666) <= layer1_outputs(8988);
    layer2_outputs(7667) <= not((layer1_outputs(10159)) and (layer1_outputs(3823)));
    layer2_outputs(7668) <= layer1_outputs(5162);
    layer2_outputs(7669) <= not(layer1_outputs(2685)) or (layer1_outputs(5864));
    layer2_outputs(7670) <= (layer1_outputs(5711)) and not (layer1_outputs(8729));
    layer2_outputs(7671) <= not(layer1_outputs(7630)) or (layer1_outputs(1254));
    layer2_outputs(7672) <= (layer1_outputs(5304)) xor (layer1_outputs(4792));
    layer2_outputs(7673) <= layer1_outputs(5319);
    layer2_outputs(7674) <= not(layer1_outputs(1832));
    layer2_outputs(7675) <= not(layer1_outputs(565)) or (layer1_outputs(3099));
    layer2_outputs(7676) <= not((layer1_outputs(1415)) and (layer1_outputs(3313)));
    layer2_outputs(7677) <= not(layer1_outputs(1389));
    layer2_outputs(7678) <= not(layer1_outputs(8523));
    layer2_outputs(7679) <= not((layer1_outputs(4197)) or (layer1_outputs(4774)));
    layer2_outputs(7680) <= (layer1_outputs(5201)) or (layer1_outputs(6894));
    layer2_outputs(7681) <= (layer1_outputs(3505)) and (layer1_outputs(5559));
    layer2_outputs(7682) <= layer1_outputs(135);
    layer2_outputs(7683) <= layer1_outputs(10181);
    layer2_outputs(7684) <= not((layer1_outputs(3889)) or (layer1_outputs(7755)));
    layer2_outputs(7685) <= not(layer1_outputs(3660)) or (layer1_outputs(9686));
    layer2_outputs(7686) <= not(layer1_outputs(484));
    layer2_outputs(7687) <= not(layer1_outputs(10111)) or (layer1_outputs(2328));
    layer2_outputs(7688) <= layer1_outputs(2706);
    layer2_outputs(7689) <= (layer1_outputs(889)) xor (layer1_outputs(6909));
    layer2_outputs(7690) <= not(layer1_outputs(448));
    layer2_outputs(7691) <= not(layer1_outputs(6998)) or (layer1_outputs(4680));
    layer2_outputs(7692) <= not(layer1_outputs(9955));
    layer2_outputs(7693) <= not(layer1_outputs(700)) or (layer1_outputs(4124));
    layer2_outputs(7694) <= not(layer1_outputs(2831));
    layer2_outputs(7695) <= not(layer1_outputs(4539)) or (layer1_outputs(9089));
    layer2_outputs(7696) <= not(layer1_outputs(9821)) or (layer1_outputs(1112));
    layer2_outputs(7697) <= not(layer1_outputs(3296));
    layer2_outputs(7698) <= not((layer1_outputs(1693)) or (layer1_outputs(7243)));
    layer2_outputs(7699) <= not((layer1_outputs(2137)) xor (layer1_outputs(7969)));
    layer2_outputs(7700) <= not((layer1_outputs(9101)) xor (layer1_outputs(2395)));
    layer2_outputs(7701) <= not(layer1_outputs(10174));
    layer2_outputs(7702) <= not(layer1_outputs(1616));
    layer2_outputs(7703) <= not(layer1_outputs(8899));
    layer2_outputs(7704) <= (layer1_outputs(2781)) and (layer1_outputs(5344));
    layer2_outputs(7705) <= (layer1_outputs(2563)) and (layer1_outputs(1247));
    layer2_outputs(7706) <= layer1_outputs(8498);
    layer2_outputs(7707) <= (layer1_outputs(7216)) or (layer1_outputs(6733));
    layer2_outputs(7708) <= not(layer1_outputs(9987));
    layer2_outputs(7709) <= not(layer1_outputs(2819));
    layer2_outputs(7710) <= (layer1_outputs(3602)) and (layer1_outputs(4472));
    layer2_outputs(7711) <= '0';
    layer2_outputs(7712) <= (layer1_outputs(9926)) and (layer1_outputs(1701));
    layer2_outputs(7713) <= not((layer1_outputs(725)) xor (layer1_outputs(3086)));
    layer2_outputs(7714) <= (layer1_outputs(7431)) xor (layer1_outputs(7187));
    layer2_outputs(7715) <= not(layer1_outputs(3319));
    layer2_outputs(7716) <= layer1_outputs(575);
    layer2_outputs(7717) <= not(layer1_outputs(7760));
    layer2_outputs(7718) <= not((layer1_outputs(8310)) xor (layer1_outputs(6513)));
    layer2_outputs(7719) <= layer1_outputs(6196);
    layer2_outputs(7720) <= layer1_outputs(8826);
    layer2_outputs(7721) <= not(layer1_outputs(474));
    layer2_outputs(7722) <= not((layer1_outputs(5563)) or (layer1_outputs(7478)));
    layer2_outputs(7723) <= not((layer1_outputs(8386)) and (layer1_outputs(7676)));
    layer2_outputs(7724) <= not(layer1_outputs(166));
    layer2_outputs(7725) <= not(layer1_outputs(9908));
    layer2_outputs(7726) <= layer1_outputs(7281);
    layer2_outputs(7727) <= layer1_outputs(8760);
    layer2_outputs(7728) <= layer1_outputs(288);
    layer2_outputs(7729) <= layer1_outputs(5612);
    layer2_outputs(7730) <= (layer1_outputs(6260)) and (layer1_outputs(7374));
    layer2_outputs(7731) <= not(layer1_outputs(9172));
    layer2_outputs(7732) <= not(layer1_outputs(949)) or (layer1_outputs(4339));
    layer2_outputs(7733) <= not((layer1_outputs(1559)) or (layer1_outputs(9952)));
    layer2_outputs(7734) <= not(layer1_outputs(6995));
    layer2_outputs(7735) <= not((layer1_outputs(6771)) xor (layer1_outputs(8963)));
    layer2_outputs(7736) <= layer1_outputs(8760);
    layer2_outputs(7737) <= (layer1_outputs(8023)) xor (layer1_outputs(7861));
    layer2_outputs(7738) <= not(layer1_outputs(4233));
    layer2_outputs(7739) <= not((layer1_outputs(6935)) xor (layer1_outputs(8551)));
    layer2_outputs(7740) <= not(layer1_outputs(1950));
    layer2_outputs(7741) <= not(layer1_outputs(7317));
    layer2_outputs(7742) <= not((layer1_outputs(2339)) or (layer1_outputs(8747)));
    layer2_outputs(7743) <= layer1_outputs(5048);
    layer2_outputs(7744) <= not((layer1_outputs(3871)) and (layer1_outputs(8521)));
    layer2_outputs(7745) <= (layer1_outputs(9448)) and not (layer1_outputs(2670));
    layer2_outputs(7746) <= (layer1_outputs(9345)) xor (layer1_outputs(8096));
    layer2_outputs(7747) <= (layer1_outputs(6792)) and not (layer1_outputs(3703));
    layer2_outputs(7748) <= not((layer1_outputs(6652)) xor (layer1_outputs(5256)));
    layer2_outputs(7749) <= layer1_outputs(9204);
    layer2_outputs(7750) <= (layer1_outputs(1468)) and not (layer1_outputs(2714));
    layer2_outputs(7751) <= layer1_outputs(6810);
    layer2_outputs(7752) <= not(layer1_outputs(5456)) or (layer1_outputs(4185));
    layer2_outputs(7753) <= (layer1_outputs(5422)) and not (layer1_outputs(9335));
    layer2_outputs(7754) <= layer1_outputs(7901);
    layer2_outputs(7755) <= (layer1_outputs(1956)) and not (layer1_outputs(9731));
    layer2_outputs(7756) <= not(layer1_outputs(2920)) or (layer1_outputs(7541));
    layer2_outputs(7757) <= (layer1_outputs(7382)) and not (layer1_outputs(407));
    layer2_outputs(7758) <= (layer1_outputs(2816)) xor (layer1_outputs(7591));
    layer2_outputs(7759) <= (layer1_outputs(9500)) or (layer1_outputs(8798));
    layer2_outputs(7760) <= not(layer1_outputs(3218));
    layer2_outputs(7761) <= layer1_outputs(9897);
    layer2_outputs(7762) <= (layer1_outputs(3111)) or (layer1_outputs(2560));
    layer2_outputs(7763) <= not(layer1_outputs(2946)) or (layer1_outputs(5637));
    layer2_outputs(7764) <= (layer1_outputs(5425)) and not (layer1_outputs(9516));
    layer2_outputs(7765) <= not(layer1_outputs(5831));
    layer2_outputs(7766) <= layer1_outputs(5213);
    layer2_outputs(7767) <= not(layer1_outputs(4940));
    layer2_outputs(7768) <= layer1_outputs(7732);
    layer2_outputs(7769) <= (layer1_outputs(5818)) and not (layer1_outputs(3921));
    layer2_outputs(7770) <= not((layer1_outputs(4191)) xor (layer1_outputs(1031)));
    layer2_outputs(7771) <= not(layer1_outputs(4515));
    layer2_outputs(7772) <= not(layer1_outputs(9755)) or (layer1_outputs(1631));
    layer2_outputs(7773) <= (layer1_outputs(8124)) xor (layer1_outputs(7885));
    layer2_outputs(7774) <= (layer1_outputs(8892)) or (layer1_outputs(6131));
    layer2_outputs(7775) <= not(layer1_outputs(10026)) or (layer1_outputs(4280));
    layer2_outputs(7776) <= (layer1_outputs(9171)) xor (layer1_outputs(133));
    layer2_outputs(7777) <= not(layer1_outputs(6038));
    layer2_outputs(7778) <= not(layer1_outputs(1882));
    layer2_outputs(7779) <= not((layer1_outputs(1555)) and (layer1_outputs(981)));
    layer2_outputs(7780) <= not((layer1_outputs(8869)) and (layer1_outputs(7546)));
    layer2_outputs(7781) <= (layer1_outputs(4432)) and not (layer1_outputs(3293));
    layer2_outputs(7782) <= not((layer1_outputs(8819)) or (layer1_outputs(3654)));
    layer2_outputs(7783) <= not(layer1_outputs(941));
    layer2_outputs(7784) <= layer1_outputs(7011);
    layer2_outputs(7785) <= (layer1_outputs(8274)) and (layer1_outputs(2565));
    layer2_outputs(7786) <= not(layer1_outputs(3708));
    layer2_outputs(7787) <= not(layer1_outputs(956));
    layer2_outputs(7788) <= not(layer1_outputs(8827));
    layer2_outputs(7789) <= not((layer1_outputs(852)) xor (layer1_outputs(7611)));
    layer2_outputs(7790) <= not(layer1_outputs(9500));
    layer2_outputs(7791) <= (layer1_outputs(2279)) xor (layer1_outputs(4616));
    layer2_outputs(7792) <= (layer1_outputs(6187)) or (layer1_outputs(9427));
    layer2_outputs(7793) <= layer1_outputs(8541);
    layer2_outputs(7794) <= not(layer1_outputs(116));
    layer2_outputs(7795) <= (layer1_outputs(8501)) and not (layer1_outputs(7433));
    layer2_outputs(7796) <= (layer1_outputs(5823)) and not (layer1_outputs(6677));
    layer2_outputs(7797) <= (layer1_outputs(815)) xor (layer1_outputs(6451));
    layer2_outputs(7798) <= not(layer1_outputs(4075)) or (layer1_outputs(6851));
    layer2_outputs(7799) <= (layer1_outputs(4729)) xor (layer1_outputs(649));
    layer2_outputs(7800) <= not((layer1_outputs(8204)) and (layer1_outputs(5982)));
    layer2_outputs(7801) <= (layer1_outputs(988)) xor (layer1_outputs(4914));
    layer2_outputs(7802) <= (layer1_outputs(7383)) xor (layer1_outputs(2068));
    layer2_outputs(7803) <= (layer1_outputs(3719)) and (layer1_outputs(7950));
    layer2_outputs(7804) <= layer1_outputs(7894);
    layer2_outputs(7805) <= not(layer1_outputs(5272));
    layer2_outputs(7806) <= not((layer1_outputs(8517)) or (layer1_outputs(2360)));
    layer2_outputs(7807) <= (layer1_outputs(110)) xor (layer1_outputs(5009));
    layer2_outputs(7808) <= not(layer1_outputs(5315)) or (layer1_outputs(2027));
    layer2_outputs(7809) <= layer1_outputs(8761);
    layer2_outputs(7810) <= (layer1_outputs(6883)) and (layer1_outputs(6875));
    layer2_outputs(7811) <= (layer1_outputs(7054)) xor (layer1_outputs(6074));
    layer2_outputs(7812) <= not((layer1_outputs(3115)) or (layer1_outputs(9882)));
    layer2_outputs(7813) <= not(layer1_outputs(1578));
    layer2_outputs(7814) <= not((layer1_outputs(7312)) and (layer1_outputs(2873)));
    layer2_outputs(7815) <= (layer1_outputs(1309)) and not (layer1_outputs(1153));
    layer2_outputs(7816) <= not(layer1_outputs(136));
    layer2_outputs(7817) <= (layer1_outputs(5797)) or (layer1_outputs(8091));
    layer2_outputs(7818) <= (layer1_outputs(1541)) xor (layer1_outputs(2228));
    layer2_outputs(7819) <= not(layer1_outputs(6735));
    layer2_outputs(7820) <= not(layer1_outputs(8376));
    layer2_outputs(7821) <= layer1_outputs(2066);
    layer2_outputs(7822) <= (layer1_outputs(7614)) and not (layer1_outputs(4800));
    layer2_outputs(7823) <= layer1_outputs(5345);
    layer2_outputs(7824) <= (layer1_outputs(9900)) and (layer1_outputs(9045));
    layer2_outputs(7825) <= not(layer1_outputs(3853));
    layer2_outputs(7826) <= layer1_outputs(5743);
    layer2_outputs(7827) <= (layer1_outputs(543)) xor (layer1_outputs(8567));
    layer2_outputs(7828) <= not((layer1_outputs(6578)) and (layer1_outputs(2474)));
    layer2_outputs(7829) <= (layer1_outputs(7946)) and (layer1_outputs(935));
    layer2_outputs(7830) <= not((layer1_outputs(9602)) xor (layer1_outputs(9251)));
    layer2_outputs(7831) <= not(layer1_outputs(7201));
    layer2_outputs(7832) <= not(layer1_outputs(8296));
    layer2_outputs(7833) <= layer1_outputs(6505);
    layer2_outputs(7834) <= not(layer1_outputs(6744));
    layer2_outputs(7835) <= (layer1_outputs(10221)) and not (layer1_outputs(9621));
    layer2_outputs(7836) <= (layer1_outputs(10179)) xor (layer1_outputs(193));
    layer2_outputs(7837) <= not(layer1_outputs(7556));
    layer2_outputs(7838) <= (layer1_outputs(9530)) xor (layer1_outputs(8489));
    layer2_outputs(7839) <= (layer1_outputs(217)) and (layer1_outputs(3073));
    layer2_outputs(7840) <= layer1_outputs(1378);
    layer2_outputs(7841) <= not(layer1_outputs(9504)) or (layer1_outputs(2221));
    layer2_outputs(7842) <= not(layer1_outputs(3912));
    layer2_outputs(7843) <= (layer1_outputs(8155)) xor (layer1_outputs(7721));
    layer2_outputs(7844) <= not(layer1_outputs(5447));
    layer2_outputs(7845) <= layer1_outputs(6130);
    layer2_outputs(7846) <= not(layer1_outputs(3822)) or (layer1_outputs(3354));
    layer2_outputs(7847) <= not((layer1_outputs(2901)) xor (layer1_outputs(643)));
    layer2_outputs(7848) <= not((layer1_outputs(3576)) or (layer1_outputs(9625)));
    layer2_outputs(7849) <= layer1_outputs(4951);
    layer2_outputs(7850) <= layer1_outputs(1763);
    layer2_outputs(7851) <= not((layer1_outputs(6375)) xor (layer1_outputs(9746)));
    layer2_outputs(7852) <= not(layer1_outputs(7973)) or (layer1_outputs(870));
    layer2_outputs(7853) <= not(layer1_outputs(8678));
    layer2_outputs(7854) <= not(layer1_outputs(3379)) or (layer1_outputs(1013));
    layer2_outputs(7855) <= layer1_outputs(7361);
    layer2_outputs(7856) <= layer1_outputs(9210);
    layer2_outputs(7857) <= not(layer1_outputs(1235));
    layer2_outputs(7858) <= not((layer1_outputs(4671)) or (layer1_outputs(9587)));
    layer2_outputs(7859) <= (layer1_outputs(4136)) and not (layer1_outputs(4538));
    layer2_outputs(7860) <= not(layer1_outputs(5854));
    layer2_outputs(7861) <= not((layer1_outputs(2278)) or (layer1_outputs(5517)));
    layer2_outputs(7862) <= not(layer1_outputs(9645));
    layer2_outputs(7863) <= not(layer1_outputs(4755));
    layer2_outputs(7864) <= layer1_outputs(6008);
    layer2_outputs(7865) <= not((layer1_outputs(9169)) and (layer1_outputs(9945)));
    layer2_outputs(7866) <= (layer1_outputs(1533)) and (layer1_outputs(8148));
    layer2_outputs(7867) <= layer1_outputs(1431);
    layer2_outputs(7868) <= not(layer1_outputs(4853)) or (layer1_outputs(7070));
    layer2_outputs(7869) <= (layer1_outputs(5959)) xor (layer1_outputs(6447));
    layer2_outputs(7870) <= not((layer1_outputs(7299)) or (layer1_outputs(6190)));
    layer2_outputs(7871) <= layer1_outputs(666);
    layer2_outputs(7872) <= (layer1_outputs(966)) xor (layer1_outputs(1461));
    layer2_outputs(7873) <= layer1_outputs(3438);
    layer2_outputs(7874) <= not(layer1_outputs(7163));
    layer2_outputs(7875) <= not((layer1_outputs(6149)) and (layer1_outputs(1813)));
    layer2_outputs(7876) <= not(layer1_outputs(3335));
    layer2_outputs(7877) <= layer1_outputs(2627);
    layer2_outputs(7878) <= (layer1_outputs(2042)) xor (layer1_outputs(9221));
    layer2_outputs(7879) <= (layer1_outputs(7519)) and (layer1_outputs(8537));
    layer2_outputs(7880) <= not(layer1_outputs(408));
    layer2_outputs(7881) <= layer1_outputs(9529);
    layer2_outputs(7882) <= layer1_outputs(9060);
    layer2_outputs(7883) <= layer1_outputs(2879);
    layer2_outputs(7884) <= layer1_outputs(8987);
    layer2_outputs(7885) <= layer1_outputs(1511);
    layer2_outputs(7886) <= layer1_outputs(7638);
    layer2_outputs(7887) <= (layer1_outputs(7781)) and not (layer1_outputs(1561));
    layer2_outputs(7888) <= (layer1_outputs(4094)) and not (layer1_outputs(5771));
    layer2_outputs(7889) <= not((layer1_outputs(1103)) and (layer1_outputs(6745)));
    layer2_outputs(7890) <= layer1_outputs(1202);
    layer2_outputs(7891) <= layer1_outputs(2639);
    layer2_outputs(7892) <= not(layer1_outputs(4540));
    layer2_outputs(7893) <= not(layer1_outputs(3781));
    layer2_outputs(7894) <= not((layer1_outputs(2104)) or (layer1_outputs(7362)));
    layer2_outputs(7895) <= not(layer1_outputs(6441));
    layer2_outputs(7896) <= layer1_outputs(1522);
    layer2_outputs(7897) <= (layer1_outputs(5386)) and (layer1_outputs(65));
    layer2_outputs(7898) <= not(layer1_outputs(6359));
    layer2_outputs(7899) <= not(layer1_outputs(2940));
    layer2_outputs(7900) <= not(layer1_outputs(2054));
    layer2_outputs(7901) <= not((layer1_outputs(1025)) or (layer1_outputs(3921)));
    layer2_outputs(7902) <= not(layer1_outputs(4921));
    layer2_outputs(7903) <= not(layer1_outputs(296));
    layer2_outputs(7904) <= not(layer1_outputs(2737));
    layer2_outputs(7905) <= (layer1_outputs(951)) and (layer1_outputs(4329));
    layer2_outputs(7906) <= (layer1_outputs(6890)) xor (layer1_outputs(5285));
    layer2_outputs(7907) <= not(layer1_outputs(9163));
    layer2_outputs(7908) <= not(layer1_outputs(459));
    layer2_outputs(7909) <= (layer1_outputs(1858)) and not (layer1_outputs(9206));
    layer2_outputs(7910) <= layer1_outputs(6857);
    layer2_outputs(7911) <= not(layer1_outputs(5952));
    layer2_outputs(7912) <= (layer1_outputs(789)) xor (layer1_outputs(5099));
    layer2_outputs(7913) <= not(layer1_outputs(634));
    layer2_outputs(7914) <= layer1_outputs(1569);
    layer2_outputs(7915) <= not(layer1_outputs(3114));
    layer2_outputs(7916) <= not((layer1_outputs(106)) and (layer1_outputs(7823)));
    layer2_outputs(7917) <= layer1_outputs(2160);
    layer2_outputs(7918) <= not((layer1_outputs(7881)) and (layer1_outputs(9386)));
    layer2_outputs(7919) <= layer1_outputs(5436);
    layer2_outputs(7920) <= layer1_outputs(4171);
    layer2_outputs(7921) <= not((layer1_outputs(5709)) or (layer1_outputs(9086)));
    layer2_outputs(7922) <= not(layer1_outputs(6241));
    layer2_outputs(7923) <= layer1_outputs(2543);
    layer2_outputs(7924) <= layer1_outputs(9699);
    layer2_outputs(7925) <= not((layer1_outputs(3420)) and (layer1_outputs(3348)));
    layer2_outputs(7926) <= not(layer1_outputs(6310)) or (layer1_outputs(6409));
    layer2_outputs(7927) <= layer1_outputs(4440);
    layer2_outputs(7928) <= layer1_outputs(9819);
    layer2_outputs(7929) <= not(layer1_outputs(5537)) or (layer1_outputs(3161));
    layer2_outputs(7930) <= layer1_outputs(2712);
    layer2_outputs(7931) <= not(layer1_outputs(6583));
    layer2_outputs(7932) <= layer1_outputs(6186);
    layer2_outputs(7933) <= (layer1_outputs(5335)) xor (layer1_outputs(2753));
    layer2_outputs(7934) <= layer1_outputs(5186);
    layer2_outputs(7935) <= layer1_outputs(6031);
    layer2_outputs(7936) <= (layer1_outputs(6870)) and not (layer1_outputs(6641));
    layer2_outputs(7937) <= layer1_outputs(3906);
    layer2_outputs(7938) <= not((layer1_outputs(7137)) and (layer1_outputs(5822)));
    layer2_outputs(7939) <= layer1_outputs(3618);
    layer2_outputs(7940) <= layer1_outputs(8849);
    layer2_outputs(7941) <= not(layer1_outputs(9167));
    layer2_outputs(7942) <= (layer1_outputs(3447)) and not (layer1_outputs(5938));
    layer2_outputs(7943) <= not(layer1_outputs(67));
    layer2_outputs(7944) <= not((layer1_outputs(9012)) xor (layer1_outputs(133)));
    layer2_outputs(7945) <= layer1_outputs(7686);
    layer2_outputs(7946) <= (layer1_outputs(7979)) and (layer1_outputs(3923));
    layer2_outputs(7947) <= not((layer1_outputs(5053)) xor (layer1_outputs(7987)));
    layer2_outputs(7948) <= layer1_outputs(6901);
    layer2_outputs(7949) <= layer1_outputs(5601);
    layer2_outputs(7950) <= not(layer1_outputs(5207));
    layer2_outputs(7951) <= not(layer1_outputs(535));
    layer2_outputs(7952) <= layer1_outputs(2787);
    layer2_outputs(7953) <= not(layer1_outputs(2095));
    layer2_outputs(7954) <= layer1_outputs(4883);
    layer2_outputs(7955) <= not(layer1_outputs(3234)) or (layer1_outputs(7806));
    layer2_outputs(7956) <= layer1_outputs(2404);
    layer2_outputs(7957) <= not(layer1_outputs(9512));
    layer2_outputs(7958) <= (layer1_outputs(7410)) and not (layer1_outputs(5163));
    layer2_outputs(7959) <= not(layer1_outputs(6243)) or (layer1_outputs(4476));
    layer2_outputs(7960) <= layer1_outputs(5422);
    layer2_outputs(7961) <= (layer1_outputs(8847)) or (layer1_outputs(1902));
    layer2_outputs(7962) <= not(layer1_outputs(5119));
    layer2_outputs(7963) <= not(layer1_outputs(5859));
    layer2_outputs(7964) <= not(layer1_outputs(6436));
    layer2_outputs(7965) <= layer1_outputs(5066);
    layer2_outputs(7966) <= (layer1_outputs(373)) or (layer1_outputs(5085));
    layer2_outputs(7967) <= not(layer1_outputs(3744)) or (layer1_outputs(2949));
    layer2_outputs(7968) <= not(layer1_outputs(2550));
    layer2_outputs(7969) <= layer1_outputs(6194);
    layer2_outputs(7970) <= layer1_outputs(1810);
    layer2_outputs(7971) <= not((layer1_outputs(8879)) xor (layer1_outputs(2024)));
    layer2_outputs(7972) <= not((layer1_outputs(8266)) or (layer1_outputs(1673)));
    layer2_outputs(7973) <= (layer1_outputs(5543)) and not (layer1_outputs(1349));
    layer2_outputs(7974) <= not((layer1_outputs(7894)) and (layer1_outputs(6446)));
    layer2_outputs(7975) <= layer1_outputs(2077);
    layer2_outputs(7976) <= not((layer1_outputs(7072)) or (layer1_outputs(915)));
    layer2_outputs(7977) <= layer1_outputs(8872);
    layer2_outputs(7978) <= '0';
    layer2_outputs(7979) <= not(layer1_outputs(5311));
    layer2_outputs(7980) <= not(layer1_outputs(7145));
    layer2_outputs(7981) <= not((layer1_outputs(3784)) and (layer1_outputs(3684)));
    layer2_outputs(7982) <= (layer1_outputs(9615)) xor (layer1_outputs(7695));
    layer2_outputs(7983) <= not(layer1_outputs(6786));
    layer2_outputs(7984) <= layer1_outputs(3922);
    layer2_outputs(7985) <= not((layer1_outputs(1450)) xor (layer1_outputs(4230)));
    layer2_outputs(7986) <= not(layer1_outputs(4672));
    layer2_outputs(7987) <= not(layer1_outputs(9045));
    layer2_outputs(7988) <= (layer1_outputs(8704)) or (layer1_outputs(8240));
    layer2_outputs(7989) <= layer1_outputs(4404);
    layer2_outputs(7990) <= not(layer1_outputs(5720));
    layer2_outputs(7991) <= (layer1_outputs(2839)) xor (layer1_outputs(9673));
    layer2_outputs(7992) <= layer1_outputs(2216);
    layer2_outputs(7993) <= layer1_outputs(7066);
    layer2_outputs(7994) <= layer1_outputs(3284);
    layer2_outputs(7995) <= (layer1_outputs(10085)) xor (layer1_outputs(5661));
    layer2_outputs(7996) <= not(layer1_outputs(6712)) or (layer1_outputs(4837));
    layer2_outputs(7997) <= not(layer1_outputs(8637));
    layer2_outputs(7998) <= (layer1_outputs(2166)) xor (layer1_outputs(9591));
    layer2_outputs(7999) <= layer1_outputs(604);
    layer2_outputs(8000) <= not((layer1_outputs(7197)) or (layer1_outputs(8119)));
    layer2_outputs(8001) <= (layer1_outputs(5377)) xor (layer1_outputs(507));
    layer2_outputs(8002) <= layer1_outputs(5512);
    layer2_outputs(8003) <= not(layer1_outputs(3043)) or (layer1_outputs(7931));
    layer2_outputs(8004) <= layer1_outputs(8795);
    layer2_outputs(8005) <= not(layer1_outputs(9178));
    layer2_outputs(8006) <= layer1_outputs(8561);
    layer2_outputs(8007) <= (layer1_outputs(5470)) xor (layer1_outputs(4146));
    layer2_outputs(8008) <= not((layer1_outputs(3165)) xor (layer1_outputs(3678)));
    layer2_outputs(8009) <= (layer1_outputs(10222)) or (layer1_outputs(7928));
    layer2_outputs(8010) <= (layer1_outputs(8056)) and not (layer1_outputs(4347));
    layer2_outputs(8011) <= layer1_outputs(6636);
    layer2_outputs(8012) <= not(layer1_outputs(295));
    layer2_outputs(8013) <= layer1_outputs(2105);
    layer2_outputs(8014) <= not(layer1_outputs(9512));
    layer2_outputs(8015) <= not(layer1_outputs(7253)) or (layer1_outputs(3408));
    layer2_outputs(8016) <= (layer1_outputs(3232)) xor (layer1_outputs(6503));
    layer2_outputs(8017) <= not(layer1_outputs(6699));
    layer2_outputs(8018) <= not(layer1_outputs(3894)) or (layer1_outputs(7993));
    layer2_outputs(8019) <= '1';
    layer2_outputs(8020) <= layer1_outputs(6770);
    layer2_outputs(8021) <= (layer1_outputs(7130)) and (layer1_outputs(2446));
    layer2_outputs(8022) <= not(layer1_outputs(3562));
    layer2_outputs(8023) <= layer1_outputs(5507);
    layer2_outputs(8024) <= not(layer1_outputs(1145));
    layer2_outputs(8025) <= layer1_outputs(6465);
    layer2_outputs(8026) <= layer1_outputs(3734);
    layer2_outputs(8027) <= layer1_outputs(9542);
    layer2_outputs(8028) <= layer1_outputs(496);
    layer2_outputs(8029) <= layer1_outputs(3239);
    layer2_outputs(8030) <= layer1_outputs(3097);
    layer2_outputs(8031) <= layer1_outputs(7557);
    layer2_outputs(8032) <= not(layer1_outputs(9302));
    layer2_outputs(8033) <= '1';
    layer2_outputs(8034) <= layer1_outputs(3929);
    layer2_outputs(8035) <= (layer1_outputs(8190)) xor (layer1_outputs(4766));
    layer2_outputs(8036) <= layer1_outputs(2079);
    layer2_outputs(8037) <= not(layer1_outputs(879));
    layer2_outputs(8038) <= (layer1_outputs(2324)) and (layer1_outputs(531));
    layer2_outputs(8039) <= (layer1_outputs(7168)) and not (layer1_outputs(2697));
    layer2_outputs(8040) <= (layer1_outputs(3200)) and not (layer1_outputs(2924));
    layer2_outputs(8041) <= not(layer1_outputs(6979));
    layer2_outputs(8042) <= layer1_outputs(2236);
    layer2_outputs(8043) <= not(layer1_outputs(1113));
    layer2_outputs(8044) <= (layer1_outputs(3299)) and not (layer1_outputs(9685));
    layer2_outputs(8045) <= not(layer1_outputs(7185));
    layer2_outputs(8046) <= (layer1_outputs(4159)) and not (layer1_outputs(3677));
    layer2_outputs(8047) <= not((layer1_outputs(6161)) xor (layer1_outputs(4903)));
    layer2_outputs(8048) <= layer1_outputs(3145);
    layer2_outputs(8049) <= layer1_outputs(1884);
    layer2_outputs(8050) <= not((layer1_outputs(2505)) xor (layer1_outputs(3261)));
    layer2_outputs(8051) <= not(layer1_outputs(7203));
    layer2_outputs(8052) <= (layer1_outputs(316)) and not (layer1_outputs(5328));
    layer2_outputs(8053) <= layer1_outputs(4513);
    layer2_outputs(8054) <= (layer1_outputs(4840)) and (layer1_outputs(2313));
    layer2_outputs(8055) <= layer1_outputs(5255);
    layer2_outputs(8056) <= not(layer1_outputs(5146));
    layer2_outputs(8057) <= layer1_outputs(341);
    layer2_outputs(8058) <= (layer1_outputs(8947)) xor (layer1_outputs(3032));
    layer2_outputs(8059) <= not(layer1_outputs(1047));
    layer2_outputs(8060) <= not(layer1_outputs(2345));
    layer2_outputs(8061) <= not(layer1_outputs(8451));
    layer2_outputs(8062) <= not(layer1_outputs(3532));
    layer2_outputs(8063) <= (layer1_outputs(3318)) and not (layer1_outputs(2126));
    layer2_outputs(8064) <= not(layer1_outputs(6594));
    layer2_outputs(8065) <= not(layer1_outputs(5757));
    layer2_outputs(8066) <= not((layer1_outputs(1576)) xor (layer1_outputs(970)));
    layer2_outputs(8067) <= layer1_outputs(9126);
    layer2_outputs(8068) <= layer1_outputs(9585);
    layer2_outputs(8069) <= not(layer1_outputs(93));
    layer2_outputs(8070) <= not(layer1_outputs(5604)) or (layer1_outputs(6208));
    layer2_outputs(8071) <= not((layer1_outputs(292)) or (layer1_outputs(5197)));
    layer2_outputs(8072) <= (layer1_outputs(4627)) and not (layer1_outputs(8813));
    layer2_outputs(8073) <= not(layer1_outputs(1473));
    layer2_outputs(8074) <= (layer1_outputs(2785)) or (layer1_outputs(7396));
    layer2_outputs(8075) <= not(layer1_outputs(9003));
    layer2_outputs(8076) <= not((layer1_outputs(1545)) xor (layer1_outputs(2585)));
    layer2_outputs(8077) <= (layer1_outputs(2911)) and not (layer1_outputs(6248));
    layer2_outputs(8078) <= layer1_outputs(5060);
    layer2_outputs(8079) <= layer1_outputs(992);
    layer2_outputs(8080) <= layer1_outputs(2219);
    layer2_outputs(8081) <= (layer1_outputs(7240)) and (layer1_outputs(2840));
    layer2_outputs(8082) <= not(layer1_outputs(396));
    layer2_outputs(8083) <= not(layer1_outputs(8805));
    layer2_outputs(8084) <= (layer1_outputs(2030)) and not (layer1_outputs(3343));
    layer2_outputs(8085) <= not(layer1_outputs(6654));
    layer2_outputs(8086) <= not((layer1_outputs(285)) or (layer1_outputs(2496)));
    layer2_outputs(8087) <= layer1_outputs(10222);
    layer2_outputs(8088) <= (layer1_outputs(2389)) and (layer1_outputs(8557));
    layer2_outputs(8089) <= not(layer1_outputs(2377)) or (layer1_outputs(2902));
    layer2_outputs(8090) <= layer1_outputs(5768);
    layer2_outputs(8091) <= layer1_outputs(1550);
    layer2_outputs(8092) <= (layer1_outputs(5166)) and not (layer1_outputs(2176));
    layer2_outputs(8093) <= not((layer1_outputs(7234)) or (layer1_outputs(101)));
    layer2_outputs(8094) <= not((layer1_outputs(2671)) xor (layer1_outputs(3135)));
    layer2_outputs(8095) <= not((layer1_outputs(4848)) xor (layer1_outputs(3483)));
    layer2_outputs(8096) <= (layer1_outputs(529)) and (layer1_outputs(4873));
    layer2_outputs(8097) <= not(layer1_outputs(8212));
    layer2_outputs(8098) <= not(layer1_outputs(3955)) or (layer1_outputs(8812));
    layer2_outputs(8099) <= not((layer1_outputs(7861)) xor (layer1_outputs(3370)));
    layer2_outputs(8100) <= (layer1_outputs(8647)) and not (layer1_outputs(6565));
    layer2_outputs(8101) <= not(layer1_outputs(4587));
    layer2_outputs(8102) <= not(layer1_outputs(1397));
    layer2_outputs(8103) <= (layer1_outputs(7944)) and not (layer1_outputs(598));
    layer2_outputs(8104) <= not(layer1_outputs(3295)) or (layer1_outputs(6697));
    layer2_outputs(8105) <= not(layer1_outputs(8939)) or (layer1_outputs(7795));
    layer2_outputs(8106) <= not(layer1_outputs(307));
    layer2_outputs(8107) <= not((layer1_outputs(1329)) and (layer1_outputs(986)));
    layer2_outputs(8108) <= not(layer1_outputs(1588)) or (layer1_outputs(901));
    layer2_outputs(8109) <= (layer1_outputs(2307)) xor (layer1_outputs(7917));
    layer2_outputs(8110) <= not((layer1_outputs(6530)) and (layer1_outputs(4997)));
    layer2_outputs(8111) <= not(layer1_outputs(9395)) or (layer1_outputs(2809));
    layer2_outputs(8112) <= not(layer1_outputs(1769)) or (layer1_outputs(3048));
    layer2_outputs(8113) <= not((layer1_outputs(8777)) xor (layer1_outputs(4158)));
    layer2_outputs(8114) <= not(layer1_outputs(7536));
    layer2_outputs(8115) <= (layer1_outputs(8889)) and not (layer1_outputs(6423));
    layer2_outputs(8116) <= layer1_outputs(4676);
    layer2_outputs(8117) <= not(layer1_outputs(9001));
    layer2_outputs(8118) <= (layer1_outputs(3047)) and not (layer1_outputs(8242));
    layer2_outputs(8119) <= not(layer1_outputs(901));
    layer2_outputs(8120) <= (layer1_outputs(2919)) or (layer1_outputs(3521));
    layer2_outputs(8121) <= layer1_outputs(2975);
    layer2_outputs(8122) <= layer1_outputs(10101);
    layer2_outputs(8123) <= (layer1_outputs(7123)) xor (layer1_outputs(9026));
    layer2_outputs(8124) <= not(layer1_outputs(7834));
    layer2_outputs(8125) <= not((layer1_outputs(5461)) xor (layer1_outputs(4552)));
    layer2_outputs(8126) <= (layer1_outputs(5308)) and (layer1_outputs(3616));
    layer2_outputs(8127) <= not(layer1_outputs(7303)) or (layer1_outputs(4899));
    layer2_outputs(8128) <= layer1_outputs(7378);
    layer2_outputs(8129) <= not(layer1_outputs(8373));
    layer2_outputs(8130) <= not((layer1_outputs(7651)) xor (layer1_outputs(3716)));
    layer2_outputs(8131) <= not((layer1_outputs(2769)) and (layer1_outputs(8157)));
    layer2_outputs(8132) <= not(layer1_outputs(9318));
    layer2_outputs(8133) <= layer1_outputs(8406);
    layer2_outputs(8134) <= (layer1_outputs(8205)) and (layer1_outputs(2860));
    layer2_outputs(8135) <= not(layer1_outputs(1346)) or (layer1_outputs(7380));
    layer2_outputs(8136) <= layer1_outputs(1678);
    layer2_outputs(8137) <= not(layer1_outputs(8140)) or (layer1_outputs(4991));
    layer2_outputs(8138) <= not(layer1_outputs(5672)) or (layer1_outputs(473));
    layer2_outputs(8139) <= (layer1_outputs(8925)) and (layer1_outputs(5616));
    layer2_outputs(8140) <= (layer1_outputs(5662)) or (layer1_outputs(435));
    layer2_outputs(8141) <= layer1_outputs(9609);
    layer2_outputs(8142) <= not(layer1_outputs(7468));
    layer2_outputs(8143) <= layer1_outputs(5967);
    layer2_outputs(8144) <= not((layer1_outputs(6975)) xor (layer1_outputs(6772)));
    layer2_outputs(8145) <= layer1_outputs(6901);
    layer2_outputs(8146) <= not(layer1_outputs(9624));
    layer2_outputs(8147) <= layer1_outputs(656);
    layer2_outputs(8148) <= not(layer1_outputs(703));
    layer2_outputs(8149) <= (layer1_outputs(8189)) and not (layer1_outputs(2132));
    layer2_outputs(8150) <= not(layer1_outputs(5392));
    layer2_outputs(8151) <= not((layer1_outputs(5004)) and (layer1_outputs(1567)));
    layer2_outputs(8152) <= layer1_outputs(9647);
    layer2_outputs(8153) <= (layer1_outputs(6697)) and not (layer1_outputs(8594));
    layer2_outputs(8154) <= layer1_outputs(8207);
    layer2_outputs(8155) <= layer1_outputs(10224);
    layer2_outputs(8156) <= layer1_outputs(5515);
    layer2_outputs(8157) <= not(layer1_outputs(5553)) or (layer1_outputs(2668));
    layer2_outputs(8158) <= not(layer1_outputs(4484));
    layer2_outputs(8159) <= layer1_outputs(3359);
    layer2_outputs(8160) <= not(layer1_outputs(2721));
    layer2_outputs(8161) <= not(layer1_outputs(5706));
    layer2_outputs(8162) <= not(layer1_outputs(2031));
    layer2_outputs(8163) <= layer1_outputs(5103);
    layer2_outputs(8164) <= layer1_outputs(2776);
    layer2_outputs(8165) <= not(layer1_outputs(7643));
    layer2_outputs(8166) <= '0';
    layer2_outputs(8167) <= (layer1_outputs(4604)) and not (layer1_outputs(4636));
    layer2_outputs(8168) <= layer1_outputs(6350);
    layer2_outputs(8169) <= (layer1_outputs(7647)) or (layer1_outputs(3697));
    layer2_outputs(8170) <= '1';
    layer2_outputs(8171) <= not((layer1_outputs(8551)) or (layer1_outputs(5694)));
    layer2_outputs(8172) <= '1';
    layer2_outputs(8173) <= not(layer1_outputs(4945));
    layer2_outputs(8174) <= layer1_outputs(4047);
    layer2_outputs(8175) <= not(layer1_outputs(3595));
    layer2_outputs(8176) <= not(layer1_outputs(9372));
    layer2_outputs(8177) <= layer1_outputs(1619);
    layer2_outputs(8178) <= layer1_outputs(3914);
    layer2_outputs(8179) <= not((layer1_outputs(5944)) xor (layer1_outputs(2571)));
    layer2_outputs(8180) <= not((layer1_outputs(32)) and (layer1_outputs(9854)));
    layer2_outputs(8181) <= layer1_outputs(1432);
    layer2_outputs(8182) <= (layer1_outputs(1603)) and (layer1_outputs(3455));
    layer2_outputs(8183) <= (layer1_outputs(7939)) and not (layer1_outputs(6904));
    layer2_outputs(8184) <= layer1_outputs(2122);
    layer2_outputs(8185) <= layer1_outputs(2036);
    layer2_outputs(8186) <= not(layer1_outputs(2905)) or (layer1_outputs(3878));
    layer2_outputs(8187) <= layer1_outputs(7659);
    layer2_outputs(8188) <= '0';
    layer2_outputs(8189) <= not((layer1_outputs(6466)) xor (layer1_outputs(3036)));
    layer2_outputs(8190) <= layer1_outputs(2542);
    layer2_outputs(8191) <= layer1_outputs(10113);
    layer2_outputs(8192) <= not(layer1_outputs(9775));
    layer2_outputs(8193) <= not((layer1_outputs(3410)) and (layer1_outputs(9332)));
    layer2_outputs(8194) <= layer1_outputs(2243);
    layer2_outputs(8195) <= not(layer1_outputs(769));
    layer2_outputs(8196) <= '0';
    layer2_outputs(8197) <= not(layer1_outputs(2696));
    layer2_outputs(8198) <= layer1_outputs(9735);
    layer2_outputs(8199) <= not((layer1_outputs(754)) and (layer1_outputs(5968)));
    layer2_outputs(8200) <= not((layer1_outputs(260)) or (layer1_outputs(8194)));
    layer2_outputs(8201) <= not(layer1_outputs(1768));
    layer2_outputs(8202) <= '1';
    layer2_outputs(8203) <= not(layer1_outputs(1116));
    layer2_outputs(8204) <= not(layer1_outputs(2380));
    layer2_outputs(8205) <= (layer1_outputs(5203)) and not (layer1_outputs(9016));
    layer2_outputs(8206) <= not((layer1_outputs(3943)) xor (layer1_outputs(1694)));
    layer2_outputs(8207) <= not(layer1_outputs(8142));
    layer2_outputs(8208) <= (layer1_outputs(963)) or (layer1_outputs(1482));
    layer2_outputs(8209) <= not((layer1_outputs(8340)) and (layer1_outputs(187)));
    layer2_outputs(8210) <= not(layer1_outputs(1010));
    layer2_outputs(8211) <= layer1_outputs(4976);
    layer2_outputs(8212) <= layer1_outputs(1477);
    layer2_outputs(8213) <= not(layer1_outputs(2276));
    layer2_outputs(8214) <= layer1_outputs(5733);
    layer2_outputs(8215) <= not(layer1_outputs(2229)) or (layer1_outputs(9544));
    layer2_outputs(8216) <= not(layer1_outputs(118));
    layer2_outputs(8217) <= not((layer1_outputs(485)) xor (layer1_outputs(3152)));
    layer2_outputs(8218) <= layer1_outputs(7269);
    layer2_outputs(8219) <= layer1_outputs(1743);
    layer2_outputs(8220) <= not(layer1_outputs(2772));
    layer2_outputs(8221) <= (layer1_outputs(8631)) or (layer1_outputs(2990));
    layer2_outputs(8222) <= not(layer1_outputs(5621));
    layer2_outputs(8223) <= (layer1_outputs(9325)) and (layer1_outputs(5232));
    layer2_outputs(8224) <= layer1_outputs(5545);
    layer2_outputs(8225) <= not(layer1_outputs(9925));
    layer2_outputs(8226) <= layer1_outputs(4888);
    layer2_outputs(8227) <= not(layer1_outputs(5713));
    layer2_outputs(8228) <= (layer1_outputs(8857)) or (layer1_outputs(7579));
    layer2_outputs(8229) <= layer1_outputs(7445);
    layer2_outputs(8230) <= (layer1_outputs(7824)) and not (layer1_outputs(8811));
    layer2_outputs(8231) <= layer1_outputs(5655);
    layer2_outputs(8232) <= (layer1_outputs(2566)) or (layer1_outputs(566));
    layer2_outputs(8233) <= layer1_outputs(343);
    layer2_outputs(8234) <= layer1_outputs(10094);
    layer2_outputs(8235) <= not(layer1_outputs(1788));
    layer2_outputs(8236) <= not(layer1_outputs(881));
    layer2_outputs(8237) <= not(layer1_outputs(5341)) or (layer1_outputs(9065));
    layer2_outputs(8238) <= not(layer1_outputs(998));
    layer2_outputs(8239) <= layer1_outputs(6909);
    layer2_outputs(8240) <= layer1_outputs(9616);
    layer2_outputs(8241) <= (layer1_outputs(9738)) or (layer1_outputs(8073));
    layer2_outputs(8242) <= (layer1_outputs(9898)) xor (layer1_outputs(2108));
    layer2_outputs(8243) <= not((layer1_outputs(6458)) and (layer1_outputs(4870)));
    layer2_outputs(8244) <= not((layer1_outputs(4898)) xor (layer1_outputs(9463)));
    layer2_outputs(8245) <= not(layer1_outputs(10162));
    layer2_outputs(8246) <= not(layer1_outputs(1829)) or (layer1_outputs(6802));
    layer2_outputs(8247) <= layer1_outputs(5752);
    layer2_outputs(8248) <= not(layer1_outputs(7842));
    layer2_outputs(8249) <= not(layer1_outputs(9634));
    layer2_outputs(8250) <= layer1_outputs(2390);
    layer2_outputs(8251) <= not(layer1_outputs(7621));
    layer2_outputs(8252) <= not((layer1_outputs(9446)) xor (layer1_outputs(1908)));
    layer2_outputs(8253) <= layer1_outputs(6102);
    layer2_outputs(8254) <= (layer1_outputs(5356)) or (layer1_outputs(5206));
    layer2_outputs(8255) <= not(layer1_outputs(1472));
    layer2_outputs(8256) <= (layer1_outputs(3941)) or (layer1_outputs(4187));
    layer2_outputs(8257) <= not(layer1_outputs(8214));
    layer2_outputs(8258) <= not(layer1_outputs(4890));
    layer2_outputs(8259) <= not(layer1_outputs(6448)) or (layer1_outputs(5268));
    layer2_outputs(8260) <= not(layer1_outputs(5659));
    layer2_outputs(8261) <= (layer1_outputs(2471)) xor (layer1_outputs(1747));
    layer2_outputs(8262) <= not(layer1_outputs(9351));
    layer2_outputs(8263) <= not(layer1_outputs(2422)) or (layer1_outputs(3231));
    layer2_outputs(8264) <= (layer1_outputs(1255)) or (layer1_outputs(4755));
    layer2_outputs(8265) <= (layer1_outputs(3167)) and not (layer1_outputs(1094));
    layer2_outputs(8266) <= not(layer1_outputs(2734));
    layer2_outputs(8267) <= (layer1_outputs(772)) and (layer1_outputs(9191));
    layer2_outputs(8268) <= not((layer1_outputs(6186)) xor (layer1_outputs(8270)));
    layer2_outputs(8269) <= not(layer1_outputs(6936));
    layer2_outputs(8270) <= (layer1_outputs(9320)) or (layer1_outputs(4749));
    layer2_outputs(8271) <= layer1_outputs(2972);
    layer2_outputs(8272) <= not((layer1_outputs(5204)) or (layer1_outputs(4774)));
    layer2_outputs(8273) <= not(layer1_outputs(5740));
    layer2_outputs(8274) <= (layer1_outputs(8955)) xor (layer1_outputs(3108));
    layer2_outputs(8275) <= layer1_outputs(10184);
    layer2_outputs(8276) <= (layer1_outputs(7593)) and not (layer1_outputs(6562));
    layer2_outputs(8277) <= layer1_outputs(9013);
    layer2_outputs(8278) <= layer1_outputs(2938);
    layer2_outputs(8279) <= (layer1_outputs(5290)) and not (layer1_outputs(4658));
    layer2_outputs(8280) <= not(layer1_outputs(2189));
    layer2_outputs(8281) <= not(layer1_outputs(2701));
    layer2_outputs(8282) <= layer1_outputs(8564);
    layer2_outputs(8283) <= '0';
    layer2_outputs(8284) <= layer1_outputs(6936);
    layer2_outputs(8285) <= layer1_outputs(3268);
    layer2_outputs(8286) <= layer1_outputs(7400);
    layer2_outputs(8287) <= not(layer1_outputs(1423));
    layer2_outputs(8288) <= layer1_outputs(3546);
    layer2_outputs(8289) <= (layer1_outputs(9915)) xor (layer1_outputs(44));
    layer2_outputs(8290) <= layer1_outputs(9288);
    layer2_outputs(8291) <= layer1_outputs(1353);
    layer2_outputs(8292) <= not(layer1_outputs(4694));
    layer2_outputs(8293) <= layer1_outputs(576);
    layer2_outputs(8294) <= (layer1_outputs(5955)) xor (layer1_outputs(6627));
    layer2_outputs(8295) <= layer1_outputs(1988);
    layer2_outputs(8296) <= not(layer1_outputs(9805));
    layer2_outputs(8297) <= not(layer1_outputs(244));
    layer2_outputs(8298) <= (layer1_outputs(5836)) and (layer1_outputs(6459));
    layer2_outputs(8299) <= not((layer1_outputs(1772)) xor (layer1_outputs(1229)));
    layer2_outputs(8300) <= layer1_outputs(823);
    layer2_outputs(8301) <= (layer1_outputs(1016)) or (layer1_outputs(1388));
    layer2_outputs(8302) <= (layer1_outputs(3159)) and not (layer1_outputs(9716));
    layer2_outputs(8303) <= not(layer1_outputs(2364));
    layer2_outputs(8304) <= (layer1_outputs(7088)) xor (layer1_outputs(9244));
    layer2_outputs(8305) <= layer1_outputs(9687);
    layer2_outputs(8306) <= layer1_outputs(2047);
    layer2_outputs(8307) <= layer1_outputs(1627);
    layer2_outputs(8308) <= not(layer1_outputs(5994)) or (layer1_outputs(601));
    layer2_outputs(8309) <= layer1_outputs(9471);
    layer2_outputs(8310) <= layer1_outputs(3968);
    layer2_outputs(8311) <= layer1_outputs(6250);
    layer2_outputs(8312) <= not(layer1_outputs(208)) or (layer1_outputs(7369));
    layer2_outputs(8313) <= (layer1_outputs(5862)) and (layer1_outputs(1359));
    layer2_outputs(8314) <= not((layer1_outputs(7161)) and (layer1_outputs(4110)));
    layer2_outputs(8315) <= (layer1_outputs(7437)) or (layer1_outputs(4981));
    layer2_outputs(8316) <= not(layer1_outputs(7148));
    layer2_outputs(8317) <= not(layer1_outputs(9086));
    layer2_outputs(8318) <= layer1_outputs(7897);
    layer2_outputs(8319) <= not(layer1_outputs(8725)) or (layer1_outputs(7878));
    layer2_outputs(8320) <= not(layer1_outputs(1451));
    layer2_outputs(8321) <= layer1_outputs(1066);
    layer2_outputs(8322) <= layer1_outputs(1655);
    layer2_outputs(8323) <= not((layer1_outputs(4685)) or (layer1_outputs(2765)));
    layer2_outputs(8324) <= not(layer1_outputs(8519));
    layer2_outputs(8325) <= layer1_outputs(3827);
    layer2_outputs(8326) <= layer1_outputs(6657);
    layer2_outputs(8327) <= (layer1_outputs(7162)) and not (layer1_outputs(1830));
    layer2_outputs(8328) <= not(layer1_outputs(10174));
    layer2_outputs(8329) <= layer1_outputs(3996);
    layer2_outputs(8330) <= layer1_outputs(8578);
    layer2_outputs(8331) <= (layer1_outputs(9948)) and (layer1_outputs(9174));
    layer2_outputs(8332) <= layer1_outputs(5566);
    layer2_outputs(8333) <= not(layer1_outputs(9054));
    layer2_outputs(8334) <= not(layer1_outputs(5611));
    layer2_outputs(8335) <= not(layer1_outputs(755));
    layer2_outputs(8336) <= (layer1_outputs(9947)) or (layer1_outputs(4273));
    layer2_outputs(8337) <= layer1_outputs(1857);
    layer2_outputs(8338) <= '1';
    layer2_outputs(8339) <= not((layer1_outputs(3394)) or (layer1_outputs(4664)));
    layer2_outputs(8340) <= not(layer1_outputs(4105));
    layer2_outputs(8341) <= '1';
    layer2_outputs(8342) <= not(layer1_outputs(1347)) or (layer1_outputs(7));
    layer2_outputs(8343) <= (layer1_outputs(3707)) xor (layer1_outputs(3649));
    layer2_outputs(8344) <= not((layer1_outputs(2528)) xor (layer1_outputs(2882)));
    layer2_outputs(8345) <= (layer1_outputs(7916)) and (layer1_outputs(9099));
    layer2_outputs(8346) <= not((layer1_outputs(2639)) xor (layer1_outputs(8291)));
    layer2_outputs(8347) <= not(layer1_outputs(3015)) or (layer1_outputs(8766));
    layer2_outputs(8348) <= layer1_outputs(1854);
    layer2_outputs(8349) <= layer1_outputs(9614);
    layer2_outputs(8350) <= not(layer1_outputs(705));
    layer2_outputs(8351) <= layer1_outputs(2411);
    layer2_outputs(8352) <= (layer1_outputs(1492)) and not (layer1_outputs(1524));
    layer2_outputs(8353) <= not(layer1_outputs(5065)) or (layer1_outputs(7209));
    layer2_outputs(8354) <= not(layer1_outputs(8458));
    layer2_outputs(8355) <= (layer1_outputs(6908)) and not (layer1_outputs(8720));
    layer2_outputs(8356) <= not((layer1_outputs(9860)) or (layer1_outputs(4397)));
    layer2_outputs(8357) <= (layer1_outputs(8463)) and not (layer1_outputs(6800));
    layer2_outputs(8358) <= layer1_outputs(10117);
    layer2_outputs(8359) <= layer1_outputs(6215);
    layer2_outputs(8360) <= (layer1_outputs(9878)) xor (layer1_outputs(7632));
    layer2_outputs(8361) <= not(layer1_outputs(6280));
    layer2_outputs(8362) <= layer1_outputs(2629);
    layer2_outputs(8363) <= layer1_outputs(2174);
    layer2_outputs(8364) <= not((layer1_outputs(4100)) and (layer1_outputs(4594)));
    layer2_outputs(8365) <= not(layer1_outputs(8131));
    layer2_outputs(8366) <= (layer1_outputs(9196)) and (layer1_outputs(2876));
    layer2_outputs(8367) <= not(layer1_outputs(2376)) or (layer1_outputs(1484));
    layer2_outputs(8368) <= (layer1_outputs(3945)) and (layer1_outputs(6458));
    layer2_outputs(8369) <= (layer1_outputs(6578)) and (layer1_outputs(4460));
    layer2_outputs(8370) <= layer1_outputs(7558);
    layer2_outputs(8371) <= (layer1_outputs(7615)) and not (layer1_outputs(6684));
    layer2_outputs(8372) <= (layer1_outputs(7554)) or (layer1_outputs(7247));
    layer2_outputs(8373) <= layer1_outputs(10003);
    layer2_outputs(8374) <= layer1_outputs(2945);
    layer2_outputs(8375) <= (layer1_outputs(7710)) xor (layer1_outputs(174));
    layer2_outputs(8376) <= not(layer1_outputs(4315));
    layer2_outputs(8377) <= not(layer1_outputs(108));
    layer2_outputs(8378) <= layer1_outputs(8962);
    layer2_outputs(8379) <= not(layer1_outputs(2942));
    layer2_outputs(8380) <= '1';
    layer2_outputs(8381) <= (layer1_outputs(8821)) and (layer1_outputs(9337));
    layer2_outputs(8382) <= (layer1_outputs(5754)) and not (layer1_outputs(4571));
    layer2_outputs(8383) <= layer1_outputs(9912);
    layer2_outputs(8384) <= (layer1_outputs(8976)) and not (layer1_outputs(1248));
    layer2_outputs(8385) <= not(layer1_outputs(8515)) or (layer1_outputs(4685));
    layer2_outputs(8386) <= not(layer1_outputs(6688));
    layer2_outputs(8387) <= not(layer1_outputs(2023));
    layer2_outputs(8388) <= not(layer1_outputs(8973));
    layer2_outputs(8389) <= layer1_outputs(5528);
    layer2_outputs(8390) <= not(layer1_outputs(7745));
    layer2_outputs(8391) <= not(layer1_outputs(9370));
    layer2_outputs(8392) <= (layer1_outputs(2764)) and not (layer1_outputs(6273));
    layer2_outputs(8393) <= layer1_outputs(26);
    layer2_outputs(8394) <= not(layer1_outputs(4720)) or (layer1_outputs(906));
    layer2_outputs(8395) <= not((layer1_outputs(8691)) xor (layer1_outputs(756)));
    layer2_outputs(8396) <= (layer1_outputs(2423)) or (layer1_outputs(9338));
    layer2_outputs(8397) <= not(layer1_outputs(4142));
    layer2_outputs(8398) <= not(layer1_outputs(952)) or (layer1_outputs(5861));
    layer2_outputs(8399) <= layer1_outputs(1717);
    layer2_outputs(8400) <= not(layer1_outputs(6359));
    layer2_outputs(8401) <= layer1_outputs(6563);
    layer2_outputs(8402) <= not(layer1_outputs(4848));
    layer2_outputs(8403) <= not(layer1_outputs(7703));
    layer2_outputs(8404) <= not(layer1_outputs(6309));
    layer2_outputs(8405) <= '1';
    layer2_outputs(8406) <= not(layer1_outputs(1572)) or (layer1_outputs(5682));
    layer2_outputs(8407) <= not(layer1_outputs(3859));
    layer2_outputs(8408) <= not((layer1_outputs(6125)) xor (layer1_outputs(491)));
    layer2_outputs(8409) <= not(layer1_outputs(6466)) or (layer1_outputs(8919));
    layer2_outputs(8410) <= not(layer1_outputs(414));
    layer2_outputs(8411) <= not(layer1_outputs(8534));
    layer2_outputs(8412) <= layer1_outputs(8116);
    layer2_outputs(8413) <= layer1_outputs(9931);
    layer2_outputs(8414) <= not(layer1_outputs(5622));
    layer2_outputs(8415) <= not(layer1_outputs(1929));
    layer2_outputs(8416) <= not(layer1_outputs(3622)) or (layer1_outputs(10036));
    layer2_outputs(8417) <= (layer1_outputs(220)) or (layer1_outputs(8873));
    layer2_outputs(8418) <= layer1_outputs(3762);
    layer2_outputs(8419) <= not(layer1_outputs(7445));
    layer2_outputs(8420) <= layer1_outputs(8751);
    layer2_outputs(8421) <= not(layer1_outputs(3698)) or (layer1_outputs(5080));
    layer2_outputs(8422) <= not((layer1_outputs(618)) and (layer1_outputs(4746)));
    layer2_outputs(8423) <= not(layer1_outputs(10187));
    layer2_outputs(8424) <= not(layer1_outputs(9959));
    layer2_outputs(8425) <= (layer1_outputs(4058)) or (layer1_outputs(9023));
    layer2_outputs(8426) <= not(layer1_outputs(6325));
    layer2_outputs(8427) <= (layer1_outputs(1334)) or (layer1_outputs(3064));
    layer2_outputs(8428) <= layer1_outputs(4029);
    layer2_outputs(8429) <= layer1_outputs(113);
    layer2_outputs(8430) <= (layer1_outputs(1922)) and not (layer1_outputs(4767));
    layer2_outputs(8431) <= layer1_outputs(10199);
    layer2_outputs(8432) <= not(layer1_outputs(7060));
    layer2_outputs(8433) <= not((layer1_outputs(8322)) and (layer1_outputs(9717)));
    layer2_outputs(8434) <= (layer1_outputs(10075)) or (layer1_outputs(782));
    layer2_outputs(8435) <= not((layer1_outputs(1872)) and (layer1_outputs(10138)));
    layer2_outputs(8436) <= not(layer1_outputs(4505));
    layer2_outputs(8437) <= layer1_outputs(6404);
    layer2_outputs(8438) <= (layer1_outputs(5502)) and not (layer1_outputs(2822));
    layer2_outputs(8439) <= not(layer1_outputs(9175));
    layer2_outputs(8440) <= (layer1_outputs(2816)) xor (layer1_outputs(2845));
    layer2_outputs(8441) <= layer1_outputs(5987);
    layer2_outputs(8442) <= not(layer1_outputs(4692));
    layer2_outputs(8443) <= layer1_outputs(9199);
    layer2_outputs(8444) <= not(layer1_outputs(2434)) or (layer1_outputs(8071));
    layer2_outputs(8445) <= not(layer1_outputs(1515)) or (layer1_outputs(4839));
    layer2_outputs(8446) <= layer1_outputs(5560);
    layer2_outputs(8447) <= not((layer1_outputs(7457)) and (layer1_outputs(5354)));
    layer2_outputs(8448) <= layer1_outputs(8230);
    layer2_outputs(8449) <= not(layer1_outputs(4650));
    layer2_outputs(8450) <= layer1_outputs(6780);
    layer2_outputs(8451) <= (layer1_outputs(3519)) or (layer1_outputs(8179));
    layer2_outputs(8452) <= (layer1_outputs(9481)) and not (layer1_outputs(7962));
    layer2_outputs(8453) <= not((layer1_outputs(9547)) xor (layer1_outputs(7770)));
    layer2_outputs(8454) <= not((layer1_outputs(3411)) xor (layer1_outputs(8103)));
    layer2_outputs(8455) <= not(layer1_outputs(7580));
    layer2_outputs(8456) <= not((layer1_outputs(8018)) and (layer1_outputs(2425)));
    layer2_outputs(8457) <= (layer1_outputs(8351)) or (layer1_outputs(7579));
    layer2_outputs(8458) <= layer1_outputs(3535);
    layer2_outputs(8459) <= layer1_outputs(3888);
    layer2_outputs(8460) <= not(layer1_outputs(9205));
    layer2_outputs(8461) <= layer1_outputs(3653);
    layer2_outputs(8462) <= not(layer1_outputs(4273));
    layer2_outputs(8463) <= not(layer1_outputs(4696));
    layer2_outputs(8464) <= layer1_outputs(6529);
    layer2_outputs(8465) <= not(layer1_outputs(2042));
    layer2_outputs(8466) <= not(layer1_outputs(5856));
    layer2_outputs(8467) <= not(layer1_outputs(8849));
    layer2_outputs(8468) <= layer1_outputs(4652);
    layer2_outputs(8469) <= layer1_outputs(3727);
    layer2_outputs(8470) <= (layer1_outputs(3828)) and not (layer1_outputs(2732));
    layer2_outputs(8471) <= layer1_outputs(362);
    layer2_outputs(8472) <= not(layer1_outputs(6796)) or (layer1_outputs(9497));
    layer2_outputs(8473) <= layer1_outputs(715);
    layer2_outputs(8474) <= not(layer1_outputs(1191));
    layer2_outputs(8475) <= not(layer1_outputs(5014));
    layer2_outputs(8476) <= (layer1_outputs(6777)) and (layer1_outputs(2102));
    layer2_outputs(8477) <= not(layer1_outputs(6494));
    layer2_outputs(8478) <= not((layer1_outputs(1106)) and (layer1_outputs(3864)));
    layer2_outputs(8479) <= not(layer1_outputs(7453)) or (layer1_outputs(9868));
    layer2_outputs(8480) <= (layer1_outputs(1816)) and (layer1_outputs(1917));
    layer2_outputs(8481) <= not((layer1_outputs(7052)) and (layer1_outputs(7194)));
    layer2_outputs(8482) <= not(layer1_outputs(7938)) or (layer1_outputs(7083));
    layer2_outputs(8483) <= not((layer1_outputs(8248)) xor (layer1_outputs(7683)));
    layer2_outputs(8484) <= (layer1_outputs(1242)) and (layer1_outputs(1532));
    layer2_outputs(8485) <= layer1_outputs(3091);
    layer2_outputs(8486) <= (layer1_outputs(5801)) or (layer1_outputs(4794));
    layer2_outputs(8487) <= not(layer1_outputs(8740)) or (layer1_outputs(1019));
    layer2_outputs(8488) <= (layer1_outputs(600)) xor (layer1_outputs(3449));
    layer2_outputs(8489) <= layer1_outputs(2692);
    layer2_outputs(8490) <= layer1_outputs(5471);
    layer2_outputs(8491) <= not(layer1_outputs(7267));
    layer2_outputs(8492) <= layer1_outputs(5812);
    layer2_outputs(8493) <= (layer1_outputs(7335)) and (layer1_outputs(8021));
    layer2_outputs(8494) <= not(layer1_outputs(996));
    layer2_outputs(8495) <= not(layer1_outputs(4120));
    layer2_outputs(8496) <= layer1_outputs(1959);
    layer2_outputs(8497) <= not(layer1_outputs(4216));
    layer2_outputs(8498) <= (layer1_outputs(3231)) xor (layer1_outputs(8345));
    layer2_outputs(8499) <= not((layer1_outputs(3211)) or (layer1_outputs(10190)));
    layer2_outputs(8500) <= not(layer1_outputs(4630));
    layer2_outputs(8501) <= not((layer1_outputs(7831)) and (layer1_outputs(4750)));
    layer2_outputs(8502) <= (layer1_outputs(1523)) and not (layer1_outputs(427));
    layer2_outputs(8503) <= not((layer1_outputs(9534)) or (layer1_outputs(8688)));
    layer2_outputs(8504) <= not(layer1_outputs(1500)) or (layer1_outputs(3728));
    layer2_outputs(8505) <= not(layer1_outputs(8812)) or (layer1_outputs(3352));
    layer2_outputs(8506) <= not(layer1_outputs(4817));
    layer2_outputs(8507) <= (layer1_outputs(4825)) xor (layer1_outputs(3051));
    layer2_outputs(8508) <= layer1_outputs(826);
    layer2_outputs(8509) <= not(layer1_outputs(7042));
    layer2_outputs(8510) <= not((layer1_outputs(1731)) or (layer1_outputs(5582)));
    layer2_outputs(8511) <= not(layer1_outputs(2111));
    layer2_outputs(8512) <= layer1_outputs(8715);
    layer2_outputs(8513) <= layer1_outputs(6681);
    layer2_outputs(8514) <= (layer1_outputs(5325)) and not (layer1_outputs(6288));
    layer2_outputs(8515) <= (layer1_outputs(8811)) and not (layer1_outputs(1952));
    layer2_outputs(8516) <= (layer1_outputs(745)) and not (layer1_outputs(5837));
    layer2_outputs(8517) <= layer1_outputs(8207);
    layer2_outputs(8518) <= not(layer1_outputs(823));
    layer2_outputs(8519) <= not(layer1_outputs(9119));
    layer2_outputs(8520) <= not((layer1_outputs(7967)) and (layer1_outputs(1316)));
    layer2_outputs(8521) <= layer1_outputs(1219);
    layer2_outputs(8522) <= not((layer1_outputs(1336)) and (layer1_outputs(1183)));
    layer2_outputs(8523) <= not(layer1_outputs(5787));
    layer2_outputs(8524) <= (layer1_outputs(7759)) and not (layer1_outputs(9671));
    layer2_outputs(8525) <= (layer1_outputs(6072)) and not (layer1_outputs(1067));
    layer2_outputs(8526) <= not(layer1_outputs(534));
    layer2_outputs(8527) <= not((layer1_outputs(7026)) or (layer1_outputs(2428)));
    layer2_outputs(8528) <= not((layer1_outputs(8529)) or (layer1_outputs(1333)));
    layer2_outputs(8529) <= not(layer1_outputs(4861));
    layer2_outputs(8530) <= layer1_outputs(5497);
    layer2_outputs(8531) <= not(layer1_outputs(9412)) or (layer1_outputs(4317));
    layer2_outputs(8532) <= '0';
    layer2_outputs(8533) <= layer1_outputs(939);
    layer2_outputs(8534) <= (layer1_outputs(1736)) and (layer1_outputs(8123));
    layer2_outputs(8535) <= not(layer1_outputs(5230));
    layer2_outputs(8536) <= (layer1_outputs(9625)) or (layer1_outputs(896));
    layer2_outputs(8537) <= (layer1_outputs(7462)) and not (layer1_outputs(807));
    layer2_outputs(8538) <= (layer1_outputs(5905)) xor (layer1_outputs(1366));
    layer2_outputs(8539) <= not((layer1_outputs(7077)) or (layer1_outputs(5698)));
    layer2_outputs(8540) <= not((layer1_outputs(5173)) and (layer1_outputs(6517)));
    layer2_outputs(8541) <= not((layer1_outputs(4252)) xor (layer1_outputs(5252)));
    layer2_outputs(8542) <= (layer1_outputs(8219)) and not (layer1_outputs(6891));
    layer2_outputs(8543) <= layer1_outputs(371);
    layer2_outputs(8544) <= not((layer1_outputs(8401)) and (layer1_outputs(2214)));
    layer2_outputs(8545) <= not((layer1_outputs(1460)) or (layer1_outputs(5209)));
    layer2_outputs(8546) <= not(layer1_outputs(6784));
    layer2_outputs(8547) <= layer1_outputs(5899);
    layer2_outputs(8548) <= (layer1_outputs(3334)) or (layer1_outputs(7802));
    layer2_outputs(8549) <= not(layer1_outputs(8623)) or (layer1_outputs(3905));
    layer2_outputs(8550) <= not(layer1_outputs(4808));
    layer2_outputs(8551) <= not(layer1_outputs(3553)) or (layer1_outputs(4690));
    layer2_outputs(8552) <= not(layer1_outputs(10226));
    layer2_outputs(8553) <= not(layer1_outputs(4279)) or (layer1_outputs(4555));
    layer2_outputs(8554) <= (layer1_outputs(1231)) and (layer1_outputs(3064));
    layer2_outputs(8555) <= not(layer1_outputs(9332));
    layer2_outputs(8556) <= layer1_outputs(6331);
    layer2_outputs(8557) <= not(layer1_outputs(1565));
    layer2_outputs(8558) <= not(layer1_outputs(3306));
    layer2_outputs(8559) <= layer1_outputs(8117);
    layer2_outputs(8560) <= layer1_outputs(759);
    layer2_outputs(8561) <= layer1_outputs(6212);
    layer2_outputs(8562) <= not(layer1_outputs(8357));
    layer2_outputs(8563) <= layer1_outputs(1109);
    layer2_outputs(8564) <= not(layer1_outputs(7564));
    layer2_outputs(8565) <= layer1_outputs(370);
    layer2_outputs(8566) <= (layer1_outputs(8040)) and not (layer1_outputs(3916));
    layer2_outputs(8567) <= layer1_outputs(3269);
    layer2_outputs(8568) <= not((layer1_outputs(8111)) xor (layer1_outputs(6586)));
    layer2_outputs(8569) <= '0';
    layer2_outputs(8570) <= layer1_outputs(739);
    layer2_outputs(8571) <= not((layer1_outputs(3683)) or (layer1_outputs(5739)));
    layer2_outputs(8572) <= layer1_outputs(944);
    layer2_outputs(8573) <= not(layer1_outputs(2791)) or (layer1_outputs(3031));
    layer2_outputs(8574) <= layer1_outputs(5223);
    layer2_outputs(8575) <= not((layer1_outputs(1140)) xor (layer1_outputs(10098)));
    layer2_outputs(8576) <= layer1_outputs(7572);
    layer2_outputs(8577) <= not(layer1_outputs(4109)) or (layer1_outputs(33));
    layer2_outputs(8578) <= layer1_outputs(4201);
    layer2_outputs(8579) <= (layer1_outputs(2394)) or (layer1_outputs(7120));
    layer2_outputs(8580) <= not(layer1_outputs(3205));
    layer2_outputs(8581) <= not(layer1_outputs(7192));
    layer2_outputs(8582) <= not(layer1_outputs(5792));
    layer2_outputs(8583) <= layer1_outputs(4113);
    layer2_outputs(8584) <= layer1_outputs(8786);
    layer2_outputs(8585) <= layer1_outputs(5599);
    layer2_outputs(8586) <= (layer1_outputs(7068)) xor (layer1_outputs(4651));
    layer2_outputs(8587) <= layer1_outputs(3970);
    layer2_outputs(8588) <= not(layer1_outputs(8712));
    layer2_outputs(8589) <= (layer1_outputs(2712)) and (layer1_outputs(1284));
    layer2_outputs(8590) <= not(layer1_outputs(9725)) or (layer1_outputs(2787));
    layer2_outputs(8591) <= (layer1_outputs(10182)) and not (layer1_outputs(1209));
    layer2_outputs(8592) <= not((layer1_outputs(10037)) and (layer1_outputs(2579)));
    layer2_outputs(8593) <= (layer1_outputs(5967)) and (layer1_outputs(4722));
    layer2_outputs(8594) <= not(layer1_outputs(4037)) or (layer1_outputs(7550));
    layer2_outputs(8595) <= not(layer1_outputs(2512));
    layer2_outputs(8596) <= (layer1_outputs(418)) xor (layer1_outputs(4300));
    layer2_outputs(8597) <= not(layer1_outputs(1749));
    layer2_outputs(8598) <= not(layer1_outputs(2789));
    layer2_outputs(8599) <= layer1_outputs(2140);
    layer2_outputs(8600) <= (layer1_outputs(8475)) and not (layer1_outputs(769));
    layer2_outputs(8601) <= not(layer1_outputs(5985));
    layer2_outputs(8602) <= not(layer1_outputs(2834));
    layer2_outputs(8603) <= not(layer1_outputs(141)) or (layer1_outputs(8931));
    layer2_outputs(8604) <= not((layer1_outputs(5588)) or (layer1_outputs(4929)));
    layer2_outputs(8605) <= layer1_outputs(3206);
    layer2_outputs(8606) <= not((layer1_outputs(10161)) and (layer1_outputs(4918)));
    layer2_outputs(8607) <= not(layer1_outputs(6627));
    layer2_outputs(8608) <= (layer1_outputs(4543)) and not (layer1_outputs(10118));
    layer2_outputs(8609) <= not(layer1_outputs(3952)) or (layer1_outputs(1889));
    layer2_outputs(8610) <= layer1_outputs(7031);
    layer2_outputs(8611) <= not(layer1_outputs(1735));
    layer2_outputs(8612) <= (layer1_outputs(230)) xor (layer1_outputs(2296));
    layer2_outputs(8613) <= not((layer1_outputs(9216)) or (layer1_outputs(3331)));
    layer2_outputs(8614) <= (layer1_outputs(9408)) and (layer1_outputs(8869));
    layer2_outputs(8615) <= layer1_outputs(5651);
    layer2_outputs(8616) <= layer1_outputs(10195);
    layer2_outputs(8617) <= not(layer1_outputs(683)) or (layer1_outputs(2837));
    layer2_outputs(8618) <= layer1_outputs(6365);
    layer2_outputs(8619) <= layer1_outputs(1990);
    layer2_outputs(8620) <= layer1_outputs(1976);
    layer2_outputs(8621) <= layer1_outputs(9683);
    layer2_outputs(8622) <= layer1_outputs(2249);
    layer2_outputs(8623) <= layer1_outputs(8502);
    layer2_outputs(8624) <= (layer1_outputs(9400)) or (layer1_outputs(7254));
    layer2_outputs(8625) <= (layer1_outputs(704)) or (layer1_outputs(6399));
    layer2_outputs(8626) <= layer1_outputs(1179);
    layer2_outputs(8627) <= (layer1_outputs(4357)) and not (layer1_outputs(9118));
    layer2_outputs(8628) <= layer1_outputs(9259);
    layer2_outputs(8629) <= not((layer1_outputs(9171)) xor (layer1_outputs(5093)));
    layer2_outputs(8630) <= layer1_outputs(5904);
    layer2_outputs(8631) <= not(layer1_outputs(3174));
    layer2_outputs(8632) <= layer1_outputs(6267);
    layer2_outputs(8633) <= not(layer1_outputs(972));
    layer2_outputs(8634) <= layer1_outputs(8403);
    layer2_outputs(8635) <= layer1_outputs(2835);
    layer2_outputs(8636) <= (layer1_outputs(7424)) xor (layer1_outputs(8129));
    layer2_outputs(8637) <= not(layer1_outputs(4380));
    layer2_outputs(8638) <= not(layer1_outputs(7820));
    layer2_outputs(8639) <= not(layer1_outputs(5349));
    layer2_outputs(8640) <= layer1_outputs(6401);
    layer2_outputs(8641) <= not(layer1_outputs(8766)) or (layer1_outputs(7131));
    layer2_outputs(8642) <= (layer1_outputs(9264)) and not (layer1_outputs(7349));
    layer2_outputs(8643) <= not(layer1_outputs(1462));
    layer2_outputs(8644) <= not(layer1_outputs(7155));
    layer2_outputs(8645) <= not(layer1_outputs(1151)) or (layer1_outputs(6014));
    layer2_outputs(8646) <= not(layer1_outputs(9896));
    layer2_outputs(8647) <= (layer1_outputs(9538)) and not (layer1_outputs(1042));
    layer2_outputs(8648) <= layer1_outputs(5942);
    layer2_outputs(8649) <= not(layer1_outputs(491)) or (layer1_outputs(7603));
    layer2_outputs(8650) <= not(layer1_outputs(6165));
    layer2_outputs(8651) <= not(layer1_outputs(4697));
    layer2_outputs(8652) <= layer1_outputs(5917);
    layer2_outputs(8653) <= layer1_outputs(5811);
    layer2_outputs(8654) <= (layer1_outputs(7432)) xor (layer1_outputs(6269));
    layer2_outputs(8655) <= layer1_outputs(4149);
    layer2_outputs(8656) <= not(layer1_outputs(4838));
    layer2_outputs(8657) <= not(layer1_outputs(7236));
    layer2_outputs(8658) <= not(layer1_outputs(9492));
    layer2_outputs(8659) <= not((layer1_outputs(1401)) or (layer1_outputs(909)));
    layer2_outputs(8660) <= layer1_outputs(5251);
    layer2_outputs(8661) <= layer1_outputs(1627);
    layer2_outputs(8662) <= (layer1_outputs(8949)) or (layer1_outputs(8722));
    layer2_outputs(8663) <= not(layer1_outputs(8487));
    layer2_outputs(8664) <= layer1_outputs(8123);
    layer2_outputs(8665) <= not(layer1_outputs(1473));
    layer2_outputs(8666) <= not((layer1_outputs(7495)) or (layer1_outputs(677)));
    layer2_outputs(8667) <= not(layer1_outputs(3771));
    layer2_outputs(8668) <= (layer1_outputs(4245)) xor (layer1_outputs(9988));
    layer2_outputs(8669) <= not(layer1_outputs(10082));
    layer2_outputs(8670) <= not((layer1_outputs(1695)) xor (layer1_outputs(8321)));
    layer2_outputs(8671) <= not((layer1_outputs(1451)) or (layer1_outputs(9406)));
    layer2_outputs(8672) <= not(layer1_outputs(6927));
    layer2_outputs(8673) <= not(layer1_outputs(403));
    layer2_outputs(8674) <= (layer1_outputs(77)) xor (layer1_outputs(9736));
    layer2_outputs(8675) <= (layer1_outputs(1398)) and not (layer1_outputs(7045));
    layer2_outputs(8676) <= not(layer1_outputs(9010)) or (layer1_outputs(1425));
    layer2_outputs(8677) <= not(layer1_outputs(7641));
    layer2_outputs(8678) <= layer1_outputs(6110);
    layer2_outputs(8679) <= not(layer1_outputs(5444));
    layer2_outputs(8680) <= not(layer1_outputs(5465));
    layer2_outputs(8681) <= not((layer1_outputs(8686)) xor (layer1_outputs(783)));
    layer2_outputs(8682) <= not(layer1_outputs(2362)) or (layer1_outputs(7856));
    layer2_outputs(8683) <= (layer1_outputs(3233)) and (layer1_outputs(7157));
    layer2_outputs(8684) <= (layer1_outputs(5690)) or (layer1_outputs(9548));
    layer2_outputs(8685) <= '1';
    layer2_outputs(8686) <= '0';
    layer2_outputs(8687) <= '0';
    layer2_outputs(8688) <= not((layer1_outputs(5363)) or (layer1_outputs(2561)));
    layer2_outputs(8689) <= layer1_outputs(6580);
    layer2_outputs(8690) <= layer1_outputs(4139);
    layer2_outputs(8691) <= not((layer1_outputs(3525)) and (layer1_outputs(655)));
    layer2_outputs(8692) <= not((layer1_outputs(5)) and (layer1_outputs(8118)));
    layer2_outputs(8693) <= (layer1_outputs(4032)) xor (layer1_outputs(3718));
    layer2_outputs(8694) <= (layer1_outputs(1837)) or (layer1_outputs(7218));
    layer2_outputs(8695) <= layer1_outputs(4255);
    layer2_outputs(8696) <= layer1_outputs(2751);
    layer2_outputs(8697) <= (layer1_outputs(3438)) and not (layer1_outputs(8162));
    layer2_outputs(8698) <= layer1_outputs(8983);
    layer2_outputs(8699) <= not(layer1_outputs(8719));
    layer2_outputs(8700) <= not(layer1_outputs(147));
    layer2_outputs(8701) <= not(layer1_outputs(6869)) or (layer1_outputs(9533));
    layer2_outputs(8702) <= not(layer1_outputs(10210)) or (layer1_outputs(4073));
    layer2_outputs(8703) <= not((layer1_outputs(8985)) xor (layer1_outputs(2320)));
    layer2_outputs(8704) <= layer1_outputs(2491);
    layer2_outputs(8705) <= layer1_outputs(7526);
    layer2_outputs(8706) <= not(layer1_outputs(2897));
    layer2_outputs(8707) <= not(layer1_outputs(9551));
    layer2_outputs(8708) <= (layer1_outputs(9641)) and not (layer1_outputs(5015));
    layer2_outputs(8709) <= layer1_outputs(10169);
    layer2_outputs(8710) <= not(layer1_outputs(3581)) or (layer1_outputs(9125));
    layer2_outputs(8711) <= not(layer1_outputs(5680)) or (layer1_outputs(5919));
    layer2_outputs(8712) <= layer1_outputs(9787);
    layer2_outputs(8713) <= (layer1_outputs(7659)) and (layer1_outputs(5318));
    layer2_outputs(8714) <= not(layer1_outputs(4194));
    layer2_outputs(8715) <= not(layer1_outputs(2914));
    layer2_outputs(8716) <= layer1_outputs(4629);
    layer2_outputs(8717) <= not((layer1_outputs(5217)) and (layer1_outputs(477)));
    layer2_outputs(8718) <= '0';
    layer2_outputs(8719) <= not(layer1_outputs(8674));
    layer2_outputs(8720) <= not(layer1_outputs(3225));
    layer2_outputs(8721) <= layer1_outputs(6881);
    layer2_outputs(8722) <= not(layer1_outputs(5096));
    layer2_outputs(8723) <= layer1_outputs(8070);
    layer2_outputs(8724) <= layer1_outputs(7562);
    layer2_outputs(8725) <= (layer1_outputs(9070)) and (layer1_outputs(4627));
    layer2_outputs(8726) <= layer1_outputs(3329);
    layer2_outputs(8727) <= not((layer1_outputs(1665)) or (layer1_outputs(10198)));
    layer2_outputs(8728) <= (layer1_outputs(4908)) and (layer1_outputs(7912));
    layer2_outputs(8729) <= not(layer1_outputs(101));
    layer2_outputs(8730) <= not(layer1_outputs(5682));
    layer2_outputs(8731) <= layer1_outputs(1821);
    layer2_outputs(8732) <= layer1_outputs(589);
    layer2_outputs(8733) <= not(layer1_outputs(3257)) or (layer1_outputs(828));
    layer2_outputs(8734) <= not(layer1_outputs(3839));
    layer2_outputs(8735) <= layer1_outputs(3188);
    layer2_outputs(8736) <= (layer1_outputs(9240)) and (layer1_outputs(7446));
    layer2_outputs(8737) <= not(layer1_outputs(9124));
    layer2_outputs(8738) <= not(layer1_outputs(8411)) or (layer1_outputs(6182));
    layer2_outputs(8739) <= (layer1_outputs(9551)) and not (layer1_outputs(7251));
    layer2_outputs(8740) <= (layer1_outputs(4836)) and (layer1_outputs(2722));
    layer2_outputs(8741) <= not(layer1_outputs(3294)) or (layer1_outputs(2518));
    layer2_outputs(8742) <= (layer1_outputs(8968)) and not (layer1_outputs(4731));
    layer2_outputs(8743) <= not(layer1_outputs(3297));
    layer2_outputs(8744) <= '0';
    layer2_outputs(8745) <= (layer1_outputs(851)) or (layer1_outputs(3765));
    layer2_outputs(8746) <= layer1_outputs(4573);
    layer2_outputs(8747) <= not(layer1_outputs(7474));
    layer2_outputs(8748) <= layer1_outputs(7457);
    layer2_outputs(8749) <= (layer1_outputs(9256)) and not (layer1_outputs(3592));
    layer2_outputs(8750) <= (layer1_outputs(7335)) and not (layer1_outputs(8679));
    layer2_outputs(8751) <= not(layer1_outputs(5450));
    layer2_outputs(8752) <= not(layer1_outputs(869)) or (layer1_outputs(6409));
    layer2_outputs(8753) <= layer1_outputs(4026);
    layer2_outputs(8754) <= not(layer1_outputs(3837));
    layer2_outputs(8755) <= layer1_outputs(7004);
    layer2_outputs(8756) <= not(layer1_outputs(2517)) or (layer1_outputs(623));
    layer2_outputs(8757) <= layer1_outputs(5985);
    layer2_outputs(8758) <= layer1_outputs(9991);
    layer2_outputs(8759) <= layer1_outputs(3967);
    layer2_outputs(8760) <= not((layer1_outputs(842)) or (layer1_outputs(9228)));
    layer2_outputs(8761) <= not((layer1_outputs(1091)) xor (layer1_outputs(5689)));
    layer2_outputs(8762) <= (layer1_outputs(6481)) and (layer1_outputs(3069));
    layer2_outputs(8763) <= layer1_outputs(4711);
    layer2_outputs(8764) <= layer1_outputs(8619);
    layer2_outputs(8765) <= (layer1_outputs(5699)) and not (layer1_outputs(6614));
    layer2_outputs(8766) <= layer1_outputs(7296);
    layer2_outputs(8767) <= not(layer1_outputs(5007));
    layer2_outputs(8768) <= not(layer1_outputs(3384));
    layer2_outputs(8769) <= not(layer1_outputs(92));
    layer2_outputs(8770) <= layer1_outputs(5378);
    layer2_outputs(8771) <= (layer1_outputs(160)) and not (layer1_outputs(5639));
    layer2_outputs(8772) <= (layer1_outputs(9038)) and not (layer1_outputs(1300));
    layer2_outputs(8773) <= not((layer1_outputs(197)) xor (layer1_outputs(10076)));
    layer2_outputs(8774) <= not(layer1_outputs(2777));
    layer2_outputs(8775) <= (layer1_outputs(4816)) xor (layer1_outputs(3003));
    layer2_outputs(8776) <= not(layer1_outputs(561));
    layer2_outputs(8777) <= not(layer1_outputs(1409));
    layer2_outputs(8778) <= (layer1_outputs(2032)) xor (layer1_outputs(6134));
    layer2_outputs(8779) <= layer1_outputs(7622);
    layer2_outputs(8780) <= not((layer1_outputs(3313)) xor (layer1_outputs(9665)));
    layer2_outputs(8781) <= not(layer1_outputs(1663));
    layer2_outputs(8782) <= (layer1_outputs(2527)) or (layer1_outputs(9893));
    layer2_outputs(8783) <= layer1_outputs(7348);
    layer2_outputs(8784) <= layer1_outputs(9780);
    layer2_outputs(8785) <= not(layer1_outputs(4596)) or (layer1_outputs(7947));
    layer2_outputs(8786) <= not(layer1_outputs(6957));
    layer2_outputs(8787) <= not(layer1_outputs(9789));
    layer2_outputs(8788) <= '0';
    layer2_outputs(8789) <= (layer1_outputs(4276)) and not (layer1_outputs(4754));
    layer2_outputs(8790) <= (layer1_outputs(638)) and (layer1_outputs(4975));
    layer2_outputs(8791) <= not((layer1_outputs(4483)) xor (layer1_outputs(7857)));
    layer2_outputs(8792) <= not((layer1_outputs(5230)) xor (layer1_outputs(9269)));
    layer2_outputs(8793) <= '1';
    layer2_outputs(8794) <= not(layer1_outputs(9929));
    layer2_outputs(8795) <= layer1_outputs(7023);
    layer2_outputs(8796) <= layer1_outputs(3487);
    layer2_outputs(8797) <= not(layer1_outputs(8705));
    layer2_outputs(8798) <= layer1_outputs(2212);
    layer2_outputs(8799) <= not(layer1_outputs(7657)) or (layer1_outputs(9098));
    layer2_outputs(8800) <= not(layer1_outputs(8386));
    layer2_outputs(8801) <= not(layer1_outputs(4638));
    layer2_outputs(8802) <= (layer1_outputs(8950)) xor (layer1_outputs(3969));
    layer2_outputs(8803) <= (layer1_outputs(7731)) and not (layer1_outputs(2688));
    layer2_outputs(8804) <= not(layer1_outputs(1279));
    layer2_outputs(8805) <= (layer1_outputs(5910)) and not (layer1_outputs(2466));
    layer2_outputs(8806) <= (layer1_outputs(2140)) and (layer1_outputs(3611));
    layer2_outputs(8807) <= layer1_outputs(3544);
    layer2_outputs(8808) <= (layer1_outputs(2150)) and (layer1_outputs(9791));
    layer2_outputs(8809) <= not(layer1_outputs(2675)) or (layer1_outputs(1079));
    layer2_outputs(8810) <= not((layer1_outputs(968)) or (layer1_outputs(10044)));
    layer2_outputs(8811) <= layer1_outputs(778);
    layer2_outputs(8812) <= not((layer1_outputs(3390)) xor (layer1_outputs(5252)));
    layer2_outputs(8813) <= layer1_outputs(6632);
    layer2_outputs(8814) <= not(layer1_outputs(8494)) or (layer1_outputs(339));
    layer2_outputs(8815) <= layer1_outputs(2079);
    layer2_outputs(8816) <= not((layer1_outputs(785)) and (layer1_outputs(6154)));
    layer2_outputs(8817) <= layer1_outputs(1161);
    layer2_outputs(8818) <= (layer1_outputs(4215)) or (layer1_outputs(8355));
    layer2_outputs(8819) <= not(layer1_outputs(4172));
    layer2_outputs(8820) <= (layer1_outputs(8500)) and not (layer1_outputs(6989));
    layer2_outputs(8821) <= not(layer1_outputs(6731));
    layer2_outputs(8822) <= not(layer1_outputs(8612));
    layer2_outputs(8823) <= layer1_outputs(8981);
    layer2_outputs(8824) <= not(layer1_outputs(3396));
    layer2_outputs(8825) <= layer1_outputs(733);
    layer2_outputs(8826) <= not(layer1_outputs(9610));
    layer2_outputs(8827) <= (layer1_outputs(5865)) xor (layer1_outputs(2862));
    layer2_outputs(8828) <= not((layer1_outputs(2766)) or (layer1_outputs(2101)));
    layer2_outputs(8829) <= layer1_outputs(619);
    layer2_outputs(8830) <= not((layer1_outputs(8268)) xor (layer1_outputs(3425)));
    layer2_outputs(8831) <= layer1_outputs(8174);
    layer2_outputs(8832) <= not(layer1_outputs(9363));
    layer2_outputs(8833) <= not((layer1_outputs(6126)) and (layer1_outputs(6943)));
    layer2_outputs(8834) <= (layer1_outputs(8243)) or (layer1_outputs(3377));
    layer2_outputs(8835) <= (layer1_outputs(4021)) and (layer1_outputs(4683));
    layer2_outputs(8836) <= not(layer1_outputs(8202)) or (layer1_outputs(2530));
    layer2_outputs(8837) <= (layer1_outputs(6792)) and not (layer1_outputs(5327));
    layer2_outputs(8838) <= (layer1_outputs(5651)) and not (layer1_outputs(797));
    layer2_outputs(8839) <= not(layer1_outputs(9927)) or (layer1_outputs(9917));
    layer2_outputs(8840) <= not(layer1_outputs(10088));
    layer2_outputs(8841) <= not(layer1_outputs(9328));
    layer2_outputs(8842) <= not(layer1_outputs(3417));
    layer2_outputs(8843) <= layer1_outputs(1335);
    layer2_outputs(8844) <= (layer1_outputs(8839)) and (layer1_outputs(1560));
    layer2_outputs(8845) <= not(layer1_outputs(8033));
    layer2_outputs(8846) <= layer1_outputs(693);
    layer2_outputs(8847) <= (layer1_outputs(8472)) or (layer1_outputs(7485));
    layer2_outputs(8848) <= not(layer1_outputs(7804));
    layer2_outputs(8849) <= layer1_outputs(856);
    layer2_outputs(8850) <= layer1_outputs(9309);
    layer2_outputs(8851) <= layer1_outputs(6896);
    layer2_outputs(8852) <= not((layer1_outputs(8225)) xor (layer1_outputs(7039)));
    layer2_outputs(8853) <= not(layer1_outputs(6395));
    layer2_outputs(8854) <= not(layer1_outputs(7997));
    layer2_outputs(8855) <= (layer1_outputs(1634)) xor (layer1_outputs(5843));
    layer2_outputs(8856) <= layer1_outputs(7981);
    layer2_outputs(8857) <= layer1_outputs(1533);
    layer2_outputs(8858) <= layer1_outputs(4383);
    layer2_outputs(8859) <= not(layer1_outputs(6865));
    layer2_outputs(8860) <= layer1_outputs(5030);
    layer2_outputs(8861) <= (layer1_outputs(7947)) or (layer1_outputs(1570));
    layer2_outputs(8862) <= not((layer1_outputs(7514)) xor (layer1_outputs(5006)));
    layer2_outputs(8863) <= layer1_outputs(3012);
    layer2_outputs(8864) <= not((layer1_outputs(1789)) or (layer1_outputs(9815)));
    layer2_outputs(8865) <= not(layer1_outputs(7989));
    layer2_outputs(8866) <= (layer1_outputs(3693)) and (layer1_outputs(6779));
    layer2_outputs(8867) <= not((layer1_outputs(1060)) xor (layer1_outputs(284)));
    layer2_outputs(8868) <= not((layer1_outputs(2863)) or (layer1_outputs(3922)));
    layer2_outputs(8869) <= (layer1_outputs(1276)) and not (layer1_outputs(3030));
    layer2_outputs(8870) <= not(layer1_outputs(6013));
    layer2_outputs(8871) <= (layer1_outputs(5002)) and not (layer1_outputs(4612));
    layer2_outputs(8872) <= not(layer1_outputs(4089));
    layer2_outputs(8873) <= not(layer1_outputs(5758));
    layer2_outputs(8874) <= layer1_outputs(9137);
    layer2_outputs(8875) <= (layer1_outputs(1750)) or (layer1_outputs(5607));
    layer2_outputs(8876) <= not(layer1_outputs(4856)) or (layer1_outputs(2030));
    layer2_outputs(8877) <= (layer1_outputs(7847)) or (layer1_outputs(8));
    layer2_outputs(8878) <= not((layer1_outputs(3004)) xor (layer1_outputs(2202)));
    layer2_outputs(8879) <= not(layer1_outputs(170)) or (layer1_outputs(8872));
    layer2_outputs(8880) <= (layer1_outputs(4512)) xor (layer1_outputs(9836));
    layer2_outputs(8881) <= (layer1_outputs(4962)) xor (layer1_outputs(7136));
    layer2_outputs(8882) <= (layer1_outputs(206)) xor (layer1_outputs(980));
    layer2_outputs(8883) <= not(layer1_outputs(8481));
    layer2_outputs(8884) <= (layer1_outputs(680)) xor (layer1_outputs(5990));
    layer2_outputs(8885) <= not(layer1_outputs(867));
    layer2_outputs(8886) <= not(layer1_outputs(6295));
    layer2_outputs(8887) <= (layer1_outputs(1271)) xor (layer1_outputs(5980));
    layer2_outputs(8888) <= layer1_outputs(88);
    layer2_outputs(8889) <= layer1_outputs(7841);
    layer2_outputs(8890) <= (layer1_outputs(5904)) and not (layer1_outputs(8532));
    layer2_outputs(8891) <= not(layer1_outputs(4132));
    layer2_outputs(8892) <= (layer1_outputs(7696)) and not (layer1_outputs(5626));
    layer2_outputs(8893) <= not((layer1_outputs(4223)) and (layer1_outputs(1924)));
    layer2_outputs(8894) <= layer1_outputs(7191);
    layer2_outputs(8895) <= layer1_outputs(8485);
    layer2_outputs(8896) <= (layer1_outputs(7521)) and not (layer1_outputs(1698));
    layer2_outputs(8897) <= layer1_outputs(9950);
    layer2_outputs(8898) <= (layer1_outputs(5976)) and (layer1_outputs(3717));
    layer2_outputs(8899) <= layer1_outputs(5342);
    layer2_outputs(8900) <= not((layer1_outputs(1748)) xor (layer1_outputs(6323)));
    layer2_outputs(8901) <= not((layer1_outputs(4441)) or (layer1_outputs(8464)));
    layer2_outputs(8902) <= not(layer1_outputs(857));
    layer2_outputs(8903) <= layer1_outputs(2833);
    layer2_outputs(8904) <= layer1_outputs(5382);
    layer2_outputs(8905) <= (layer1_outputs(3672)) and not (layer1_outputs(4398));
    layer2_outputs(8906) <= layer1_outputs(2100);
    layer2_outputs(8907) <= layer1_outputs(5504);
    layer2_outputs(8908) <= not(layer1_outputs(225)) or (layer1_outputs(5949));
    layer2_outputs(8909) <= layer1_outputs(2904);
    layer2_outputs(8910) <= layer1_outputs(2262);
    layer2_outputs(8911) <= not(layer1_outputs(9253));
    layer2_outputs(8912) <= layer1_outputs(9243);
    layer2_outputs(8913) <= not((layer1_outputs(4657)) and (layer1_outputs(8835)));
    layer2_outputs(8914) <= not((layer1_outputs(6502)) and (layer1_outputs(2441)));
    layer2_outputs(8915) <= not(layer1_outputs(7167));
    layer2_outputs(8916) <= not(layer1_outputs(6482));
    layer2_outputs(8917) <= layer1_outputs(6062);
    layer2_outputs(8918) <= (layer1_outputs(5424)) or (layer1_outputs(7178));
    layer2_outputs(8919) <= layer1_outputs(9103);
    layer2_outputs(8920) <= (layer1_outputs(5550)) and not (layer1_outputs(9858));
    layer2_outputs(8921) <= not(layer1_outputs(8472));
    layer2_outputs(8922) <= not(layer1_outputs(9486));
    layer2_outputs(8923) <= not(layer1_outputs(8250));
    layer2_outputs(8924) <= (layer1_outputs(1735)) and not (layer1_outputs(5666));
    layer2_outputs(8925) <= '1';
    layer2_outputs(8926) <= (layer1_outputs(1009)) or (layer1_outputs(148));
    layer2_outputs(8927) <= not((layer1_outputs(5851)) xor (layer1_outputs(2093)));
    layer2_outputs(8928) <= (layer1_outputs(7121)) and (layer1_outputs(450));
    layer2_outputs(8929) <= not(layer1_outputs(3074));
    layer2_outputs(8930) <= not(layer1_outputs(6877));
    layer2_outputs(8931) <= not(layer1_outputs(4049));
    layer2_outputs(8932) <= not(layer1_outputs(5820)) or (layer1_outputs(8967));
    layer2_outputs(8933) <= layer1_outputs(7184);
    layer2_outputs(8934) <= not(layer1_outputs(7993)) or (layer1_outputs(8014));
    layer2_outputs(8935) <= layer1_outputs(515);
    layer2_outputs(8936) <= not(layer1_outputs(841));
    layer2_outputs(8937) <= not(layer1_outputs(6915));
    layer2_outputs(8938) <= layer1_outputs(3104);
    layer2_outputs(8939) <= not(layer1_outputs(6856)) or (layer1_outputs(4477));
    layer2_outputs(8940) <= not((layer1_outputs(6159)) and (layer1_outputs(7812)));
    layer2_outputs(8941) <= not(layer1_outputs(6332));
    layer2_outputs(8942) <= not(layer1_outputs(9415));
    layer2_outputs(8943) <= not(layer1_outputs(8896)) or (layer1_outputs(7286));
    layer2_outputs(8944) <= layer1_outputs(2727);
    layer2_outputs(8945) <= not(layer1_outputs(2582));
    layer2_outputs(8946) <= not((layer1_outputs(9706)) and (layer1_outputs(7200)));
    layer2_outputs(8947) <= layer1_outputs(1923);
    layer2_outputs(8948) <= (layer1_outputs(4301)) or (layer1_outputs(7285));
    layer2_outputs(8949) <= layer1_outputs(4672);
    layer2_outputs(8950) <= not(layer1_outputs(6626));
    layer2_outputs(8951) <= layer1_outputs(1790);
    layer2_outputs(8952) <= not(layer1_outputs(5882)) or (layer1_outputs(2226));
    layer2_outputs(8953) <= not(layer1_outputs(992));
    layer2_outputs(8954) <= layer1_outputs(3896);
    layer2_outputs(8955) <= layer1_outputs(1415);
    layer2_outputs(8956) <= not(layer1_outputs(1261));
    layer2_outputs(8957) <= (layer1_outputs(2640)) and not (layer1_outputs(5944));
    layer2_outputs(8958) <= layer1_outputs(5368);
    layer2_outputs(8959) <= not((layer1_outputs(2016)) xor (layer1_outputs(6404)));
    layer2_outputs(8960) <= not(layer1_outputs(2302));
    layer2_outputs(8961) <= not(layer1_outputs(1253)) or (layer1_outputs(2683));
    layer2_outputs(8962) <= layer1_outputs(9825);
    layer2_outputs(8963) <= (layer1_outputs(1454)) xor (layer1_outputs(4803));
    layer2_outputs(8964) <= not(layer1_outputs(39));
    layer2_outputs(8965) <= not(layer1_outputs(426));
    layer2_outputs(8966) <= not(layer1_outputs(9055)) or (layer1_outputs(6377));
    layer2_outputs(8967) <= not(layer1_outputs(2108));
    layer2_outputs(8968) <= not(layer1_outputs(953));
    layer2_outputs(8969) <= layer1_outputs(8461);
    layer2_outputs(8970) <= (layer1_outputs(116)) or (layer1_outputs(6271));
    layer2_outputs(8971) <= (layer1_outputs(8130)) or (layer1_outputs(1174));
    layer2_outputs(8972) <= (layer1_outputs(7183)) and not (layer1_outputs(8797));
    layer2_outputs(8973) <= not(layer1_outputs(6755));
    layer2_outputs(8974) <= not(layer1_outputs(5687));
    layer2_outputs(8975) <= not(layer1_outputs(7533)) or (layer1_outputs(6346));
    layer2_outputs(8976) <= not(layer1_outputs(6885)) or (layer1_outputs(499));
    layer2_outputs(8977) <= '1';
    layer2_outputs(8978) <= (layer1_outputs(8037)) and (layer1_outputs(184));
    layer2_outputs(8979) <= layer1_outputs(6984);
    layer2_outputs(8980) <= layer1_outputs(6467);
    layer2_outputs(8981) <= not(layer1_outputs(7694)) or (layer1_outputs(7650));
    layer2_outputs(8982) <= (layer1_outputs(4990)) xor (layer1_outputs(9474));
    layer2_outputs(8983) <= layer1_outputs(3408);
    layer2_outputs(8984) <= layer1_outputs(757);
    layer2_outputs(8985) <= layer1_outputs(1806);
    layer2_outputs(8986) <= (layer1_outputs(8423)) and (layer1_outputs(9102));
    layer2_outputs(8987) <= not(layer1_outputs(4614)) or (layer1_outputs(9929));
    layer2_outputs(8988) <= (layer1_outputs(9699)) xor (layer1_outputs(3702));
    layer2_outputs(8989) <= not((layer1_outputs(7943)) or (layer1_outputs(7725)));
    layer2_outputs(8990) <= '0';
    layer2_outputs(8991) <= layer1_outputs(2960);
    layer2_outputs(8992) <= layer1_outputs(4443);
    layer2_outputs(8993) <= not((layer1_outputs(3327)) xor (layer1_outputs(4562)));
    layer2_outputs(8994) <= (layer1_outputs(7365)) and (layer1_outputs(1455));
    layer2_outputs(8995) <= (layer1_outputs(7370)) and not (layer1_outputs(991));
    layer2_outputs(8996) <= (layer1_outputs(7995)) xor (layer1_outputs(7858));
    layer2_outputs(8997) <= layer1_outputs(5934);
    layer2_outputs(8998) <= not(layer1_outputs(6588)) or (layer1_outputs(8632));
    layer2_outputs(8999) <= not(layer1_outputs(1508));
    layer2_outputs(9000) <= not(layer1_outputs(723));
    layer2_outputs(9001) <= layer1_outputs(3416);
    layer2_outputs(9002) <= layer1_outputs(7201);
    layer2_outputs(9003) <= not((layer1_outputs(4844)) xor (layer1_outputs(9371)));
    layer2_outputs(9004) <= not((layer1_outputs(7727)) and (layer1_outputs(9407)));
    layer2_outputs(9005) <= not(layer1_outputs(1775));
    layer2_outputs(9006) <= '1';
    layer2_outputs(9007) <= not(layer1_outputs(1283));
    layer2_outputs(9008) <= not(layer1_outputs(3904));
    layer2_outputs(9009) <= layer1_outputs(4275);
    layer2_outputs(9010) <= (layer1_outputs(5134)) and (layer1_outputs(2793));
    layer2_outputs(9011) <= not(layer1_outputs(4325));
    layer2_outputs(9012) <= not((layer1_outputs(6177)) or (layer1_outputs(8195)));
    layer2_outputs(9013) <= not(layer1_outputs(9943));
    layer2_outputs(9014) <= not(layer1_outputs(1470));
    layer2_outputs(9015) <= (layer1_outputs(908)) and not (layer1_outputs(1969));
    layer2_outputs(9016) <= (layer1_outputs(7581)) and not (layer1_outputs(6287));
    layer2_outputs(9017) <= layer1_outputs(4864);
    layer2_outputs(9018) <= not((layer1_outputs(1443)) and (layer1_outputs(9739)));
    layer2_outputs(9019) <= not((layer1_outputs(1402)) xor (layer1_outputs(9970)));
    layer2_outputs(9020) <= not((layer1_outputs(754)) xor (layer1_outputs(1239)));
    layer2_outputs(9021) <= layer1_outputs(1589);
    layer2_outputs(9022) <= layer1_outputs(10195);
    layer2_outputs(9023) <= (layer1_outputs(4130)) xor (layer1_outputs(4342));
    layer2_outputs(9024) <= (layer1_outputs(3777)) and (layer1_outputs(6549));
    layer2_outputs(9025) <= not(layer1_outputs(6928));
    layer2_outputs(9026) <= not(layer1_outputs(2037));
    layer2_outputs(9027) <= layer1_outputs(1199);
    layer2_outputs(9028) <= (layer1_outputs(1503)) and not (layer1_outputs(80));
    layer2_outputs(9029) <= not(layer1_outputs(175));
    layer2_outputs(9030) <= not(layer1_outputs(2931));
    layer2_outputs(9031) <= not(layer1_outputs(7745)) or (layer1_outputs(4310));
    layer2_outputs(9032) <= not(layer1_outputs(1421));
    layer2_outputs(9033) <= not(layer1_outputs(4185));
    layer2_outputs(9034) <= not(layer1_outputs(4468)) or (layer1_outputs(7465));
    layer2_outputs(9035) <= not(layer1_outputs(9034)) or (layer1_outputs(4904));
    layer2_outputs(9036) <= (layer1_outputs(2659)) xor (layer1_outputs(7297));
    layer2_outputs(9037) <= not(layer1_outputs(7723));
    layer2_outputs(9038) <= layer1_outputs(2694);
    layer2_outputs(9039) <= layer1_outputs(577);
    layer2_outputs(9040) <= (layer1_outputs(1271)) or (layer1_outputs(5714));
    layer2_outputs(9041) <= (layer1_outputs(8336)) and (layer1_outputs(9242));
    layer2_outputs(9042) <= not((layer1_outputs(497)) xor (layer1_outputs(6219)));
    layer2_outputs(9043) <= layer1_outputs(1994);
    layer2_outputs(9044) <= not(layer1_outputs(2186));
    layer2_outputs(9045) <= not(layer1_outputs(497));
    layer2_outputs(9046) <= layer1_outputs(3241);
    layer2_outputs(9047) <= layer1_outputs(210);
    layer2_outputs(9048) <= (layer1_outputs(4028)) and (layer1_outputs(9478));
    layer2_outputs(9049) <= not(layer1_outputs(4721));
    layer2_outputs(9050) <= not(layer1_outputs(2473)) or (layer1_outputs(4034));
    layer2_outputs(9051) <= not(layer1_outputs(622));
    layer2_outputs(9052) <= layer1_outputs(2841);
    layer2_outputs(9053) <= layer1_outputs(2275);
    layer2_outputs(9054) <= (layer1_outputs(5505)) and not (layer1_outputs(69));
    layer2_outputs(9055) <= not(layer1_outputs(9436));
    layer2_outputs(9056) <= layer1_outputs(2977);
    layer2_outputs(9057) <= (layer1_outputs(6847)) and not (layer1_outputs(8225));
    layer2_outputs(9058) <= layer1_outputs(2770);
    layer2_outputs(9059) <= (layer1_outputs(9491)) and not (layer1_outputs(4967));
    layer2_outputs(9060) <= (layer1_outputs(6285)) and (layer1_outputs(5566));
    layer2_outputs(9061) <= (layer1_outputs(2792)) or (layer1_outputs(2046));
    layer2_outputs(9062) <= layer1_outputs(8977);
    layer2_outputs(9063) <= layer1_outputs(8658);
    layer2_outputs(9064) <= not(layer1_outputs(6049)) or (layer1_outputs(10018));
    layer2_outputs(9065) <= not(layer1_outputs(6894));
    layer2_outputs(9066) <= (layer1_outputs(10032)) or (layer1_outputs(4366));
    layer2_outputs(9067) <= not(layer1_outputs(5630));
    layer2_outputs(9068) <= (layer1_outputs(6606)) or (layer1_outputs(1363));
    layer2_outputs(9069) <= (layer1_outputs(3509)) and not (layer1_outputs(3863));
    layer2_outputs(9070) <= layer1_outputs(7847);
    layer2_outputs(9071) <= layer1_outputs(5249);
    layer2_outputs(9072) <= layer1_outputs(3541);
    layer2_outputs(9073) <= not(layer1_outputs(2049));
    layer2_outputs(9074) <= (layer1_outputs(5038)) and not (layer1_outputs(2332));
    layer2_outputs(9075) <= not((layer1_outputs(9436)) and (layer1_outputs(4098)));
    layer2_outputs(9076) <= layer1_outputs(367);
    layer2_outputs(9077) <= layer1_outputs(3057);
    layer2_outputs(9078) <= not(layer1_outputs(6471));
    layer2_outputs(9079) <= (layer1_outputs(3255)) and (layer1_outputs(9529));
    layer2_outputs(9080) <= not(layer1_outputs(7649));
    layer2_outputs(9081) <= not((layer1_outputs(32)) and (layer1_outputs(3937)));
    layer2_outputs(9082) <= layer1_outputs(4330);
    layer2_outputs(9083) <= (layer1_outputs(286)) and not (layer1_outputs(5324));
    layer2_outputs(9084) <= not(layer1_outputs(1435));
    layer2_outputs(9085) <= layer1_outputs(7093);
    layer2_outputs(9086) <= layer1_outputs(4052);
    layer2_outputs(9087) <= layer1_outputs(3448);
    layer2_outputs(9088) <= not(layer1_outputs(1992));
    layer2_outputs(9089) <= (layer1_outputs(6299)) and not (layer1_outputs(9177));
    layer2_outputs(9090) <= layer1_outputs(7032);
    layer2_outputs(9091) <= not(layer1_outputs(837));
    layer2_outputs(9092) <= not(layer1_outputs(9675)) or (layer1_outputs(7537));
    layer2_outputs(9093) <= not(layer1_outputs(4710));
    layer2_outputs(9094) <= layer1_outputs(5712);
    layer2_outputs(9095) <= (layer1_outputs(6231)) and not (layer1_outputs(8733));
    layer2_outputs(9096) <= not(layer1_outputs(526));
    layer2_outputs(9097) <= not(layer1_outputs(2497));
    layer2_outputs(9098) <= layer1_outputs(1318);
    layer2_outputs(9099) <= not((layer1_outputs(9761)) and (layer1_outputs(4709)));
    layer2_outputs(9100) <= (layer1_outputs(4212)) and not (layer1_outputs(9467));
    layer2_outputs(9101) <= layer1_outputs(7045);
    layer2_outputs(9102) <= layer1_outputs(5694);
    layer2_outputs(9103) <= layer1_outputs(4390);
    layer2_outputs(9104) <= not((layer1_outputs(10162)) or (layer1_outputs(9181)));
    layer2_outputs(9105) <= layer1_outputs(1775);
    layer2_outputs(9106) <= not(layer1_outputs(5192));
    layer2_outputs(9107) <= not(layer1_outputs(5526));
    layer2_outputs(9108) <= layer1_outputs(5482);
    layer2_outputs(9109) <= (layer1_outputs(9153)) or (layer1_outputs(3324));
    layer2_outputs(9110) <= not((layer1_outputs(3763)) xor (layer1_outputs(8863)));
    layer2_outputs(9111) <= '0';
    layer2_outputs(9112) <= not(layer1_outputs(6621));
    layer2_outputs(9113) <= not(layer1_outputs(1915));
    layer2_outputs(9114) <= not(layer1_outputs(8155));
    layer2_outputs(9115) <= not(layer1_outputs(5059));
    layer2_outputs(9116) <= layer1_outputs(6615);
    layer2_outputs(9117) <= layer1_outputs(7067);
    layer2_outputs(9118) <= not(layer1_outputs(893));
    layer2_outputs(9119) <= (layer1_outputs(4621)) and (layer1_outputs(1317));
    layer2_outputs(9120) <= (layer1_outputs(2462)) or (layer1_outputs(8752));
    layer2_outputs(9121) <= not((layer1_outputs(525)) xor (layer1_outputs(7783)));
    layer2_outputs(9122) <= not(layer1_outputs(2740));
    layer2_outputs(9123) <= not(layer1_outputs(4236));
    layer2_outputs(9124) <= not((layer1_outputs(4780)) and (layer1_outputs(2164)));
    layer2_outputs(9125) <= not(layer1_outputs(1382));
    layer2_outputs(9126) <= (layer1_outputs(4501)) xor (layer1_outputs(475));
    layer2_outputs(9127) <= not(layer1_outputs(1567));
    layer2_outputs(9128) <= not(layer1_outputs(6957));
    layer2_outputs(9129) <= not(layer1_outputs(1149));
    layer2_outputs(9130) <= (layer1_outputs(5248)) and not (layer1_outputs(2625));
    layer2_outputs(9131) <= layer1_outputs(8430);
    layer2_outputs(9132) <= not(layer1_outputs(1999));
    layer2_outputs(9133) <= not(layer1_outputs(1485));
    layer2_outputs(9134) <= not(layer1_outputs(4401)) or (layer1_outputs(8107));
    layer2_outputs(9135) <= not((layer1_outputs(8138)) xor (layer1_outputs(10048)));
    layer2_outputs(9136) <= layer1_outputs(3796);
    layer2_outputs(9137) <= not((layer1_outputs(4446)) or (layer1_outputs(3352)));
    layer2_outputs(9138) <= layer1_outputs(8953);
    layer2_outputs(9139) <= not((layer1_outputs(8517)) xor (layer1_outputs(7446)));
    layer2_outputs(9140) <= layer1_outputs(6247);
    layer2_outputs(9141) <= not(layer1_outputs(9711));
    layer2_outputs(9142) <= not(layer1_outputs(6713)) or (layer1_outputs(9862));
    layer2_outputs(9143) <= (layer1_outputs(4128)) and not (layer1_outputs(931));
    layer2_outputs(9144) <= (layer1_outputs(5656)) and (layer1_outputs(797));
    layer2_outputs(9145) <= (layer1_outputs(1881)) and not (layer1_outputs(2332));
    layer2_outputs(9146) <= not(layer1_outputs(2258));
    layer2_outputs(9147) <= layer1_outputs(8941);
    layer2_outputs(9148) <= not(layer1_outputs(3985)) or (layer1_outputs(6416));
    layer2_outputs(9149) <= not(layer1_outputs(3974));
    layer2_outputs(9150) <= not(layer1_outputs(4851));
    layer2_outputs(9151) <= (layer1_outputs(9843)) and not (layer1_outputs(2613));
    layer2_outputs(9152) <= layer1_outputs(1174);
    layer2_outputs(9153) <= layer1_outputs(5015);
    layer2_outputs(9154) <= not(layer1_outputs(5900));
    layer2_outputs(9155) <= (layer1_outputs(1010)) xor (layer1_outputs(2763));
    layer2_outputs(9156) <= (layer1_outputs(1760)) xor (layer1_outputs(3157));
    layer2_outputs(9157) <= layer1_outputs(5159);
    layer2_outputs(9158) <= not((layer1_outputs(8184)) or (layer1_outputs(2264)));
    layer2_outputs(9159) <= layer1_outputs(6303);
    layer2_outputs(9160) <= not(layer1_outputs(154));
    layer2_outputs(9161) <= layer1_outputs(9767);
    layer2_outputs(9162) <= not(layer1_outputs(8176));
    layer2_outputs(9163) <= (layer1_outputs(1054)) or (layer1_outputs(7229));
    layer2_outputs(9164) <= (layer1_outputs(4673)) xor (layer1_outputs(7782));
    layer2_outputs(9165) <= layer1_outputs(5129);
    layer2_outputs(9166) <= (layer1_outputs(1331)) and not (layer1_outputs(5535));
    layer2_outputs(9167) <= (layer1_outputs(3956)) and not (layer1_outputs(1022));
    layer2_outputs(9168) <= not(layer1_outputs(4986)) or (layer1_outputs(8237));
    layer2_outputs(9169) <= not(layer1_outputs(9646));
    layer2_outputs(9170) <= layer1_outputs(6660);
    layer2_outputs(9171) <= '1';
    layer2_outputs(9172) <= not(layer1_outputs(2016));
    layer2_outputs(9173) <= not(layer1_outputs(9884));
    layer2_outputs(9174) <= not(layer1_outputs(1403));
    layer2_outputs(9175) <= (layer1_outputs(379)) xor (layer1_outputs(9715));
    layer2_outputs(9176) <= not(layer1_outputs(7355));
    layer2_outputs(9177) <= layer1_outputs(4479);
    layer2_outputs(9178) <= not(layer1_outputs(8264));
    layer2_outputs(9179) <= layer1_outputs(2878);
    layer2_outputs(9180) <= not(layer1_outputs(1067));
    layer2_outputs(9181) <= not(layer1_outputs(8232));
    layer2_outputs(9182) <= layer1_outputs(3559);
    layer2_outputs(9183) <= layer1_outputs(1557);
    layer2_outputs(9184) <= not(layer1_outputs(2789));
    layer2_outputs(9185) <= (layer1_outputs(3500)) and not (layer1_outputs(1998));
    layer2_outputs(9186) <= (layer1_outputs(4313)) and not (layer1_outputs(9919));
    layer2_outputs(9187) <= (layer1_outputs(2118)) xor (layer1_outputs(9698));
    layer2_outputs(9188) <= (layer1_outputs(4430)) and (layer1_outputs(6188));
    layer2_outputs(9189) <= (layer1_outputs(3867)) and (layer1_outputs(5604));
    layer2_outputs(9190) <= (layer1_outputs(3354)) and not (layer1_outputs(3850));
    layer2_outputs(9191) <= not(layer1_outputs(3512)) or (layer1_outputs(5075));
    layer2_outputs(9192) <= not((layer1_outputs(8714)) or (layer1_outputs(8300)));
    layer2_outputs(9193) <= not(layer1_outputs(10126));
    layer2_outputs(9194) <= not(layer1_outputs(7068));
    layer2_outputs(9195) <= not(layer1_outputs(337));
    layer2_outputs(9196) <= layer1_outputs(7403);
    layer2_outputs(9197) <= not(layer1_outputs(6790));
    layer2_outputs(9198) <= layer1_outputs(4393);
    layer2_outputs(9199) <= not(layer1_outputs(2785));
    layer2_outputs(9200) <= layer1_outputs(8658);
    layer2_outputs(9201) <= not(layer1_outputs(2936));
    layer2_outputs(9202) <= layer1_outputs(9100);
    layer2_outputs(9203) <= (layer1_outputs(7487)) and not (layer1_outputs(9426));
    layer2_outputs(9204) <= (layer1_outputs(4256)) xor (layer1_outputs(5502));
    layer2_outputs(9205) <= not(layer1_outputs(4793));
    layer2_outputs(9206) <= (layer1_outputs(7396)) and (layer1_outputs(8837));
    layer2_outputs(9207) <= (layer1_outputs(1006)) and not (layer1_outputs(1315));
    layer2_outputs(9208) <= (layer1_outputs(9383)) xor (layer1_outputs(300));
    layer2_outputs(9209) <= not(layer1_outputs(4751));
    layer2_outputs(9210) <= (layer1_outputs(9385)) and not (layer1_outputs(6875));
    layer2_outputs(9211) <= layer1_outputs(2799);
    layer2_outputs(9212) <= (layer1_outputs(3803)) or (layer1_outputs(7447));
    layer2_outputs(9213) <= layer1_outputs(5627);
    layer2_outputs(9214) <= not((layer1_outputs(5870)) xor (layer1_outputs(7189)));
    layer2_outputs(9215) <= not(layer1_outputs(8086));
    layer2_outputs(9216) <= layer1_outputs(6221);
    layer2_outputs(9217) <= not(layer1_outputs(817));
    layer2_outputs(9218) <= layer1_outputs(2093);
    layer2_outputs(9219) <= not(layer1_outputs(5573));
    layer2_outputs(9220) <= layer1_outputs(8861);
    layer2_outputs(9221) <= not((layer1_outputs(6393)) xor (layer1_outputs(7807)));
    layer2_outputs(9222) <= (layer1_outputs(5583)) and (layer1_outputs(7637));
    layer2_outputs(9223) <= layer1_outputs(4344);
    layer2_outputs(9224) <= layer1_outputs(9558);
    layer2_outputs(9225) <= not(layer1_outputs(7852));
    layer2_outputs(9226) <= layer1_outputs(8935);
    layer2_outputs(9227) <= layer1_outputs(6603);
    layer2_outputs(9228) <= layer1_outputs(6666);
    layer2_outputs(9229) <= layer1_outputs(5322);
    layer2_outputs(9230) <= not((layer1_outputs(1867)) and (layer1_outputs(7507)));
    layer2_outputs(9231) <= not(layer1_outputs(8723));
    layer2_outputs(9232) <= layer1_outputs(670);
    layer2_outputs(9233) <= layer1_outputs(5060);
    layer2_outputs(9234) <= layer1_outputs(4319);
    layer2_outputs(9235) <= not(layer1_outputs(3254)) or (layer1_outputs(792));
    layer2_outputs(9236) <= (layer1_outputs(6527)) and (layer1_outputs(376));
    layer2_outputs(9237) <= not(layer1_outputs(6902));
    layer2_outputs(9238) <= layer1_outputs(9967);
    layer2_outputs(9239) <= (layer1_outputs(4439)) and not (layer1_outputs(3131));
    layer2_outputs(9240) <= not(layer1_outputs(5290));
    layer2_outputs(9241) <= layer1_outputs(1424);
    layer2_outputs(9242) <= not(layer1_outputs(9913));
    layer2_outputs(9243) <= not(layer1_outputs(3033));
    layer2_outputs(9244) <= (layer1_outputs(9809)) xor (layer1_outputs(3520));
    layer2_outputs(9245) <= (layer1_outputs(9301)) xor (layer1_outputs(9803));
    layer2_outputs(9246) <= not(layer1_outputs(5273)) or (layer1_outputs(8368));
    layer2_outputs(9247) <= (layer1_outputs(961)) xor (layer1_outputs(140));
    layer2_outputs(9248) <= not((layer1_outputs(8113)) xor (layer1_outputs(3240)));
    layer2_outputs(9249) <= layer1_outputs(1188);
    layer2_outputs(9250) <= layer1_outputs(9526);
    layer2_outputs(9251) <= not((layer1_outputs(7143)) or (layer1_outputs(10197)));
    layer2_outputs(9252) <= not(layer1_outputs(8691));
    layer2_outputs(9253) <= not((layer1_outputs(1591)) xor (layer1_outputs(6837)));
    layer2_outputs(9254) <= layer1_outputs(4806);
    layer2_outputs(9255) <= layer1_outputs(86);
    layer2_outputs(9256) <= layer1_outputs(1771);
    layer2_outputs(9257) <= not(layer1_outputs(4944)) or (layer1_outputs(9120));
    layer2_outputs(9258) <= layer1_outputs(6886);
    layer2_outputs(9259) <= not(layer1_outputs(6312));
    layer2_outputs(9260) <= (layer1_outputs(442)) or (layer1_outputs(3681));
    layer2_outputs(9261) <= layer1_outputs(4349);
    layer2_outputs(9262) <= (layer1_outputs(2627)) or (layer1_outputs(4705));
    layer2_outputs(9263) <= not(layer1_outputs(2120));
    layer2_outputs(9264) <= (layer1_outputs(9235)) and not (layer1_outputs(9651));
    layer2_outputs(9265) <= layer1_outputs(6473);
    layer2_outputs(9266) <= not((layer1_outputs(5936)) xor (layer1_outputs(5679)));
    layer2_outputs(9267) <= layer1_outputs(2113);
    layer2_outputs(9268) <= not((layer1_outputs(3326)) or (layer1_outputs(9432)));
    layer2_outputs(9269) <= not((layer1_outputs(1344)) or (layer1_outputs(272)));
    layer2_outputs(9270) <= (layer1_outputs(2117)) and (layer1_outputs(9019));
    layer2_outputs(9271) <= layer1_outputs(3284);
    layer2_outputs(9272) <= layer1_outputs(1694);
    layer2_outputs(9273) <= '1';
    layer2_outputs(9274) <= layer1_outputs(7702);
    layer2_outputs(9275) <= not(layer1_outputs(8585));
    layer2_outputs(9276) <= not(layer1_outputs(5640));
    layer2_outputs(9277) <= layer1_outputs(2159);
    layer2_outputs(9278) <= layer1_outputs(4384);
    layer2_outputs(9279) <= not(layer1_outputs(8349));
    layer2_outputs(9280) <= not(layer1_outputs(9534));
    layer2_outputs(9281) <= not((layer1_outputs(925)) and (layer1_outputs(8904)));
    layer2_outputs(9282) <= not((layer1_outputs(1791)) xor (layer1_outputs(9702)));
    layer2_outputs(9283) <= (layer1_outputs(4457)) and not (layer1_outputs(256));
    layer2_outputs(9284) <= (layer1_outputs(4069)) and (layer1_outputs(3424));
    layer2_outputs(9285) <= layer1_outputs(5428);
    layer2_outputs(9286) <= not(layer1_outputs(1234));
    layer2_outputs(9287) <= not((layer1_outputs(4954)) or (layer1_outputs(2034)));
    layer2_outputs(9288) <= not(layer1_outputs(9172));
    layer2_outputs(9289) <= not((layer1_outputs(8442)) and (layer1_outputs(7724)));
    layer2_outputs(9290) <= (layer1_outputs(9020)) and not (layer1_outputs(3122));
    layer2_outputs(9291) <= not(layer1_outputs(5429));
    layer2_outputs(9292) <= layer1_outputs(8940);
    layer2_outputs(9293) <= not(layer1_outputs(6805));
    layer2_outputs(9294) <= not(layer1_outputs(691));
    layer2_outputs(9295) <= (layer1_outputs(3322)) and (layer1_outputs(1098));
    layer2_outputs(9296) <= not((layer1_outputs(5266)) and (layer1_outputs(5573)));
    layer2_outputs(9297) <= layer1_outputs(8974);
    layer2_outputs(9298) <= not(layer1_outputs(1861));
    layer2_outputs(9299) <= layer1_outputs(2461);
    layer2_outputs(9300) <= not(layer1_outputs(3817));
    layer2_outputs(9301) <= (layer1_outputs(2101)) and not (layer1_outputs(394));
    layer2_outputs(9302) <= not((layer1_outputs(7716)) xor (layer1_outputs(7343)));
    layer2_outputs(9303) <= not(layer1_outputs(9220));
    layer2_outputs(9304) <= layer1_outputs(9768);
    layer2_outputs(9305) <= layer1_outputs(7682);
    layer2_outputs(9306) <= layer1_outputs(7182);
    layer2_outputs(9307) <= layer1_outputs(4772);
    layer2_outputs(9308) <= (layer1_outputs(129)) and (layer1_outputs(9682));
    layer2_outputs(9309) <= not(layer1_outputs(3440));
    layer2_outputs(9310) <= not(layer1_outputs(4145));
    layer2_outputs(9311) <= not(layer1_outputs(6164)) or (layer1_outputs(6370));
    layer2_outputs(9312) <= not(layer1_outputs(1946));
    layer2_outputs(9313) <= layer1_outputs(5329);
    layer2_outputs(9314) <= (layer1_outputs(9983)) xor (layer1_outputs(606));
    layer2_outputs(9315) <= not(layer1_outputs(3355));
    layer2_outputs(9316) <= not(layer1_outputs(5911));
    layer2_outputs(9317) <= layer1_outputs(8139);
    layer2_outputs(9318) <= layer1_outputs(1926);
    layer2_outputs(9319) <= layer1_outputs(2015);
    layer2_outputs(9320) <= not((layer1_outputs(7085)) xor (layer1_outputs(4438)));
    layer2_outputs(9321) <= layer1_outputs(9626);
    layer2_outputs(9322) <= not(layer1_outputs(1612));
    layer2_outputs(9323) <= layer1_outputs(6040);
    layer2_outputs(9324) <= '1';
    layer2_outputs(9325) <= not(layer1_outputs(9109));
    layer2_outputs(9326) <= not(layer1_outputs(1555));
    layer2_outputs(9327) <= layer1_outputs(7419);
    layer2_outputs(9328) <= not(layer1_outputs(1610));
    layer2_outputs(9329) <= layer1_outputs(7113);
    layer2_outputs(9330) <= not(layer1_outputs(3119)) or (layer1_outputs(2121));
    layer2_outputs(9331) <= layer1_outputs(10110);
    layer2_outputs(9332) <= layer1_outputs(6270);
    layer2_outputs(9333) <= layer1_outputs(1553);
    layer2_outputs(9334) <= not(layer1_outputs(1911)) or (layer1_outputs(7866));
    layer2_outputs(9335) <= not(layer1_outputs(8884));
    layer2_outputs(9336) <= not(layer1_outputs(8922));
    layer2_outputs(9337) <= layer1_outputs(1413);
    layer2_outputs(9338) <= not(layer1_outputs(7122));
    layer2_outputs(9339) <= '1';
    layer2_outputs(9340) <= layer1_outputs(550);
    layer2_outputs(9341) <= layer1_outputs(5989);
    layer2_outputs(9342) <= not(layer1_outputs(8213));
    layer2_outputs(9343) <= (layer1_outputs(3547)) xor (layer1_outputs(10042));
    layer2_outputs(9344) <= (layer1_outputs(4138)) or (layer1_outputs(2204));
    layer2_outputs(9345) <= layer1_outputs(4298);
    layer2_outputs(9346) <= not(layer1_outputs(6328));
    layer2_outputs(9347) <= not(layer1_outputs(3397));
    layer2_outputs(9348) <= (layer1_outputs(7686)) xor (layer1_outputs(9066));
    layer2_outputs(9349) <= (layer1_outputs(4159)) xor (layer1_outputs(735));
    layer2_outputs(9350) <= (layer1_outputs(2124)) xor (layer1_outputs(5788));
    layer2_outputs(9351) <= not(layer1_outputs(7096));
    layer2_outputs(9352) <= not(layer1_outputs(6939));
    layer2_outputs(9353) <= (layer1_outputs(1880)) and (layer1_outputs(7666));
    layer2_outputs(9354) <= not(layer1_outputs(4388)) or (layer1_outputs(7330));
    layer2_outputs(9355) <= not(layer1_outputs(2322));
    layer2_outputs(9356) <= layer1_outputs(9243);
    layer2_outputs(9357) <= not(layer1_outputs(1743));
    layer2_outputs(9358) <= not((layer1_outputs(4308)) xor (layer1_outputs(9493)));
    layer2_outputs(9359) <= not(layer1_outputs(55));
    layer2_outputs(9360) <= layer1_outputs(963);
    layer2_outputs(9361) <= layer1_outputs(9060);
    layer2_outputs(9362) <= not((layer1_outputs(1357)) xor (layer1_outputs(6138)));
    layer2_outputs(9363) <= not(layer1_outputs(6100));
    layer2_outputs(9364) <= layer1_outputs(4686);
    layer2_outputs(9365) <= (layer1_outputs(763)) and not (layer1_outputs(7300));
    layer2_outputs(9366) <= not(layer1_outputs(1705));
    layer2_outputs(9367) <= not(layer1_outputs(5762));
    layer2_outputs(9368) <= (layer1_outputs(1148)) and not (layer1_outputs(9573));
    layer2_outputs(9369) <= layer1_outputs(1243);
    layer2_outputs(9370) <= not(layer1_outputs(2354));
    layer2_outputs(9371) <= not(layer1_outputs(9131));
    layer2_outputs(9372) <= not(layer1_outputs(3965));
    layer2_outputs(9373) <= not(layer1_outputs(6333));
    layer2_outputs(9374) <= not((layer1_outputs(7020)) and (layer1_outputs(924)));
    layer2_outputs(9375) <= layer1_outputs(345);
    layer2_outputs(9376) <= not((layer1_outputs(7360)) and (layer1_outputs(5331)));
    layer2_outputs(9377) <= (layer1_outputs(9882)) or (layer1_outputs(5984));
    layer2_outputs(9378) <= not(layer1_outputs(1733));
    layer2_outputs(9379) <= layer1_outputs(8643);
    layer2_outputs(9380) <= not(layer1_outputs(6744));
    layer2_outputs(9381) <= (layer1_outputs(9195)) and not (layer1_outputs(5715));
    layer2_outputs(9382) <= (layer1_outputs(7792)) xor (layer1_outputs(3431));
    layer2_outputs(9383) <= layer1_outputs(6737);
    layer2_outputs(9384) <= '1';
    layer2_outputs(9385) <= not(layer1_outputs(5062)) or (layer1_outputs(7769));
    layer2_outputs(9386) <= not((layer1_outputs(9693)) and (layer1_outputs(9979)));
    layer2_outputs(9387) <= layer1_outputs(5700);
    layer2_outputs(9388) <= not(layer1_outputs(6210));
    layer2_outputs(9389) <= layer1_outputs(6440);
    layer2_outputs(9390) <= (layer1_outputs(1227)) and (layer1_outputs(5712));
    layer2_outputs(9391) <= layer1_outputs(5940);
    layer2_outputs(9392) <= layer1_outputs(1352);
    layer2_outputs(9393) <= (layer1_outputs(9388)) and not (layer1_outputs(723));
    layer2_outputs(9394) <= not(layer1_outputs(4605)) or (layer1_outputs(401));
    layer2_outputs(9395) <= not(layer1_outputs(8341));
    layer2_outputs(9396) <= layer1_outputs(3515);
    layer2_outputs(9397) <= (layer1_outputs(796)) and not (layer1_outputs(702));
    layer2_outputs(9398) <= (layer1_outputs(8796)) xor (layer1_outputs(8913));
    layer2_outputs(9399) <= not((layer1_outputs(9623)) xor (layer1_outputs(6507)));
    layer2_outputs(9400) <= (layer1_outputs(2802)) xor (layer1_outputs(4062));
    layer2_outputs(9401) <= not(layer1_outputs(6257));
    layer2_outputs(9402) <= not(layer1_outputs(5418));
    layer2_outputs(9403) <= layer1_outputs(8701);
    layer2_outputs(9404) <= layer1_outputs(8293);
    layer2_outputs(9405) <= not(layer1_outputs(4181));
    layer2_outputs(9406) <= not(layer1_outputs(4096));
    layer2_outputs(9407) <= (layer1_outputs(9258)) and not (layer1_outputs(9607));
    layer2_outputs(9408) <= not(layer1_outputs(5877));
    layer2_outputs(9409) <= layer1_outputs(1486);
    layer2_outputs(9410) <= not(layer1_outputs(1357));
    layer2_outputs(9411) <= not(layer1_outputs(968));
    layer2_outputs(9412) <= (layer1_outputs(8059)) and not (layer1_outputs(665));
    layer2_outputs(9413) <= layer1_outputs(2476);
    layer2_outputs(9414) <= '1';
    layer2_outputs(9415) <= (layer1_outputs(3805)) xor (layer1_outputs(3268));
    layer2_outputs(9416) <= not(layer1_outputs(2314));
    layer2_outputs(9417) <= layer1_outputs(4956);
    layer2_outputs(9418) <= not(layer1_outputs(4679));
    layer2_outputs(9419) <= not(layer1_outputs(4815));
    layer2_outputs(9420) <= not(layer1_outputs(205));
    layer2_outputs(9421) <= (layer1_outputs(287)) xor (layer1_outputs(2652));
    layer2_outputs(9422) <= not((layer1_outputs(1450)) and (layer1_outputs(8165)));
    layer2_outputs(9423) <= layer1_outputs(775);
    layer2_outputs(9424) <= not((layer1_outputs(7532)) xor (layer1_outputs(6093)));
    layer2_outputs(9425) <= (layer1_outputs(2619)) xor (layer1_outputs(5885));
    layer2_outputs(9426) <= (layer1_outputs(6911)) xor (layer1_outputs(1157));
    layer2_outputs(9427) <= layer1_outputs(9568);
    layer2_outputs(9428) <= layer1_outputs(6940);
    layer2_outputs(9429) <= (layer1_outputs(10189)) xor (layer1_outputs(6880));
    layer2_outputs(9430) <= not(layer1_outputs(2451)) or (layer1_outputs(4991));
    layer2_outputs(9431) <= not(layer1_outputs(2694)) or (layer1_outputs(223));
    layer2_outputs(9432) <= layer1_outputs(3604);
    layer2_outputs(9433) <= layer1_outputs(8455);
    layer2_outputs(9434) <= layer1_outputs(4416);
    layer2_outputs(9435) <= (layer1_outputs(7859)) xor (layer1_outputs(1228));
    layer2_outputs(9436) <= (layer1_outputs(9770)) and (layer1_outputs(9295));
    layer2_outputs(9437) <= not(layer1_outputs(8071));
    layer2_outputs(9438) <= layer1_outputs(1316);
    layer2_outputs(9439) <= layer1_outputs(7504);
    layer2_outputs(9440) <= layer1_outputs(518);
    layer2_outputs(9441) <= not(layer1_outputs(2709));
    layer2_outputs(9442) <= (layer1_outputs(7221)) or (layer1_outputs(2427));
    layer2_outputs(9443) <= layer1_outputs(5118);
    layer2_outputs(9444) <= not(layer1_outputs(8219));
    layer2_outputs(9445) <= layer1_outputs(5253);
    layer2_outputs(9446) <= not(layer1_outputs(2630)) or (layer1_outputs(7918));
    layer2_outputs(9447) <= (layer1_outputs(9832)) and not (layer1_outputs(8707));
    layer2_outputs(9448) <= layer1_outputs(770);
    layer2_outputs(9449) <= (layer1_outputs(6027)) xor (layer1_outputs(3150));
    layer2_outputs(9450) <= (layer1_outputs(7463)) and not (layer1_outputs(5411));
    layer2_outputs(9451) <= layer1_outputs(983);
    layer2_outputs(9452) <= (layer1_outputs(480)) and (layer1_outputs(4839));
    layer2_outputs(9453) <= (layer1_outputs(748)) and not (layer1_outputs(4400));
    layer2_outputs(9454) <= not(layer1_outputs(7688));
    layer2_outputs(9455) <= layer1_outputs(2890);
    layer2_outputs(9456) <= not(layer1_outputs(8762));
    layer2_outputs(9457) <= layer1_outputs(7441);
    layer2_outputs(9458) <= not(layer1_outputs(8987)) or (layer1_outputs(4537));
    layer2_outputs(9459) <= not(layer1_outputs(1330));
    layer2_outputs(9460) <= not(layer1_outputs(2338)) or (layer1_outputs(9378));
    layer2_outputs(9461) <= layer1_outputs(8289);
    layer2_outputs(9462) <= layer1_outputs(11);
    layer2_outputs(9463) <= not(layer1_outputs(8035));
    layer2_outputs(9464) <= not(layer1_outputs(5235)) or (layer1_outputs(8912));
    layer2_outputs(9465) <= (layer1_outputs(1853)) and not (layer1_outputs(9470));
    layer2_outputs(9466) <= not(layer1_outputs(4606));
    layer2_outputs(9467) <= not(layer1_outputs(3844));
    layer2_outputs(9468) <= layer1_outputs(3523);
    layer2_outputs(9469) <= layer1_outputs(8324);
    layer2_outputs(9470) <= not(layer1_outputs(9214)) or (layer1_outputs(5887));
    layer2_outputs(9471) <= not((layer1_outputs(3034)) or (layer1_outputs(2235)));
    layer2_outputs(9472) <= layer1_outputs(3764);
    layer2_outputs(9473) <= not(layer1_outputs(3833)) or (layer1_outputs(3698));
    layer2_outputs(9474) <= (layer1_outputs(5533)) xor (layer1_outputs(6633));
    layer2_outputs(9475) <= (layer1_outputs(8751)) or (layer1_outputs(4589));
    layer2_outputs(9476) <= not((layer1_outputs(9262)) and (layer1_outputs(548)));
    layer2_outputs(9477) <= not((layer1_outputs(4747)) and (layer1_outputs(5943)));
    layer2_outputs(9478) <= not(layer1_outputs(8251));
    layer2_outputs(9479) <= not(layer1_outputs(8332));
    layer2_outputs(9480) <= not(layer1_outputs(7180));
    layer2_outputs(9481) <= not((layer1_outputs(9889)) and (layer1_outputs(5249)));
    layer2_outputs(9482) <= layer1_outputs(121);
    layer2_outputs(9483) <= not(layer1_outputs(6127)) or (layer1_outputs(5641));
    layer2_outputs(9484) <= not(layer1_outputs(2880));
    layer2_outputs(9485) <= (layer1_outputs(6037)) or (layer1_outputs(1774));
    layer2_outputs(9486) <= not((layer1_outputs(3934)) or (layer1_outputs(10231)));
    layer2_outputs(9487) <= not(layer1_outputs(1441));
    layer2_outputs(9488) <= not(layer1_outputs(4048));
    layer2_outputs(9489) <= (layer1_outputs(4354)) xor (layer1_outputs(1930));
    layer2_outputs(9490) <= layer1_outputs(4789);
    layer2_outputs(9491) <= not(layer1_outputs(4771));
    layer2_outputs(9492) <= layer1_outputs(768);
    layer2_outputs(9493) <= layer1_outputs(3026);
    layer2_outputs(9494) <= not(layer1_outputs(10059));
    layer2_outputs(9495) <= (layer1_outputs(4738)) or (layer1_outputs(9176));
    layer2_outputs(9496) <= not((layer1_outputs(737)) or (layer1_outputs(5679)));
    layer2_outputs(9497) <= not(layer1_outputs(5083));
    layer2_outputs(9498) <= not(layer1_outputs(6864));
    layer2_outputs(9499) <= not(layer1_outputs(10136));
    layer2_outputs(9500) <= not(layer1_outputs(579)) or (layer1_outputs(653));
    layer2_outputs(9501) <= layer1_outputs(2600);
    layer2_outputs(9502) <= not(layer1_outputs(4321));
    layer2_outputs(9503) <= not((layer1_outputs(8579)) xor (layer1_outputs(5300)));
    layer2_outputs(9504) <= (layer1_outputs(3257)) xor (layer1_outputs(1862));
    layer2_outputs(9505) <= (layer1_outputs(5876)) xor (layer1_outputs(7829));
    layer2_outputs(9506) <= layer1_outputs(6671);
    layer2_outputs(9507) <= not((layer1_outputs(3535)) and (layer1_outputs(890)));
    layer2_outputs(9508) <= layer1_outputs(4783);
    layer2_outputs(9509) <= layer1_outputs(9329);
    layer2_outputs(9510) <= not(layer1_outputs(888)) or (layer1_outputs(1145));
    layer2_outputs(9511) <= layer1_outputs(6060);
    layer2_outputs(9512) <= not(layer1_outputs(5359));
    layer2_outputs(9513) <= not(layer1_outputs(6685));
    layer2_outputs(9514) <= (layer1_outputs(7840)) and not (layer1_outputs(5926));
    layer2_outputs(9515) <= layer1_outputs(10160);
    layer2_outputs(9516) <= not((layer1_outputs(8019)) xor (layer1_outputs(7172)));
    layer2_outputs(9517) <= layer1_outputs(2811);
    layer2_outputs(9518) <= layer1_outputs(818);
    layer2_outputs(9519) <= not((layer1_outputs(1934)) xor (layer1_outputs(7995)));
    layer2_outputs(9520) <= not(layer1_outputs(1949));
    layer2_outputs(9521) <= not(layer1_outputs(971));
    layer2_outputs(9522) <= layer1_outputs(5575);
    layer2_outputs(9523) <= not((layer1_outputs(7544)) xor (layer1_outputs(2846)));
    layer2_outputs(9524) <= not(layer1_outputs(9278));
    layer2_outputs(9525) <= not(layer1_outputs(9676)) or (layer1_outputs(4855));
    layer2_outputs(9526) <= (layer1_outputs(3282)) or (layer1_outputs(7588));
    layer2_outputs(9527) <= layer1_outputs(7530);
    layer2_outputs(9528) <= not(layer1_outputs(1351));
    layer2_outputs(9529) <= not((layer1_outputs(7693)) or (layer1_outputs(8866)));
    layer2_outputs(9530) <= (layer1_outputs(3624)) xor (layer1_outputs(2861));
    layer2_outputs(9531) <= layer1_outputs(5511);
    layer2_outputs(9532) <= layer1_outputs(5931);
    layer2_outputs(9533) <= (layer1_outputs(8006)) and not (layer1_outputs(2650));
    layer2_outputs(9534) <= not(layer1_outputs(7752));
    layer2_outputs(9535) <= layer1_outputs(5661);
    layer2_outputs(9536) <= not(layer1_outputs(4053));
    layer2_outputs(9537) <= not(layer1_outputs(9381));
    layer2_outputs(9538) <= not((layer1_outputs(8335)) xor (layer1_outputs(6761)));
    layer2_outputs(9539) <= layer1_outputs(2533);
    layer2_outputs(9540) <= not(layer1_outputs(8993));
    layer2_outputs(9541) <= layer1_outputs(2811);
    layer2_outputs(9542) <= not(layer1_outputs(1121));
    layer2_outputs(9543) <= not(layer1_outputs(5656));
    layer2_outputs(9544) <= not(layer1_outputs(2353)) or (layer1_outputs(5792));
    layer2_outputs(9545) <= layer1_outputs(9590);
    layer2_outputs(9546) <= (layer1_outputs(1326)) and (layer1_outputs(4131));
    layer2_outputs(9547) <= not(layer1_outputs(10016));
    layer2_outputs(9548) <= (layer1_outputs(1163)) or (layer1_outputs(5784));
    layer2_outputs(9549) <= not(layer1_outputs(9237));
    layer2_outputs(9550) <= not(layer1_outputs(1259));
    layer2_outputs(9551) <= layer1_outputs(4789);
    layer2_outputs(9552) <= layer1_outputs(5567);
    layer2_outputs(9553) <= layer1_outputs(8835);
    layer2_outputs(9554) <= layer1_outputs(9765);
    layer2_outputs(9555) <= not(layer1_outputs(2876));
    layer2_outputs(9556) <= (layer1_outputs(6506)) and not (layer1_outputs(1339));
    layer2_outputs(9557) <= not(layer1_outputs(2774));
    layer2_outputs(9558) <= (layer1_outputs(9553)) xor (layer1_outputs(3246));
    layer2_outputs(9559) <= not(layer1_outputs(7486));
    layer2_outputs(9560) <= not((layer1_outputs(7971)) or (layer1_outputs(9541)));
    layer2_outputs(9561) <= (layer1_outputs(8850)) xor (layer1_outputs(180));
    layer2_outputs(9562) <= not(layer1_outputs(5316));
    layer2_outputs(9563) <= layer1_outputs(2635);
    layer2_outputs(9564) <= not(layer1_outputs(4544));
    layer2_outputs(9565) <= layer1_outputs(7241);
    layer2_outputs(9566) <= not(layer1_outputs(4023));
    layer2_outputs(9567) <= (layer1_outputs(6062)) and (layer1_outputs(5625));
    layer2_outputs(9568) <= (layer1_outputs(1948)) and not (layer1_outputs(9806));
    layer2_outputs(9569) <= (layer1_outputs(949)) xor (layer1_outputs(1436));
    layer2_outputs(9570) <= not(layer1_outputs(7862));
    layer2_outputs(9571) <= layer1_outputs(2363);
    layer2_outputs(9572) <= layer1_outputs(3552);
    layer2_outputs(9573) <= not(layer1_outputs(8039));
    layer2_outputs(9574) <= '0';
    layer2_outputs(9575) <= layer1_outputs(5567);
    layer2_outputs(9576) <= layer1_outputs(8721);
    layer2_outputs(9577) <= (layer1_outputs(4201)) xor (layer1_outputs(3482));
    layer2_outputs(9578) <= not(layer1_outputs(5962));
    layer2_outputs(9579) <= layer1_outputs(1602);
    layer2_outputs(9580) <= layer1_outputs(3388);
    layer2_outputs(9581) <= not(layer1_outputs(8562));
    layer2_outputs(9582) <= not(layer1_outputs(149)) or (layer1_outputs(3579));
    layer2_outputs(9583) <= not(layer1_outputs(1502));
    layer2_outputs(9584) <= not(layer1_outputs(112)) or (layer1_outputs(6757));
    layer2_outputs(9585) <= (layer1_outputs(6437)) xor (layer1_outputs(2497));
    layer2_outputs(9586) <= '0';
    layer2_outputs(9587) <= not((layer1_outputs(2073)) and (layer1_outputs(786)));
    layer2_outputs(9588) <= layer1_outputs(3932);
    layer2_outputs(9589) <= not(layer1_outputs(6511));
    layer2_outputs(9590) <= layer1_outputs(7358);
    layer2_outputs(9591) <= (layer1_outputs(9476)) and not (layer1_outputs(5806));
    layer2_outputs(9592) <= not(layer1_outputs(10039)) or (layer1_outputs(9230));
    layer2_outputs(9593) <= not(layer1_outputs(4165));
    layer2_outputs(9594) <= not(layer1_outputs(8611)) or (layer1_outputs(2384));
    layer2_outputs(9595) <= not((layer1_outputs(7302)) xor (layer1_outputs(9455)));
    layer2_outputs(9596) <= (layer1_outputs(1628)) or (layer1_outputs(5108));
    layer2_outputs(9597) <= not(layer1_outputs(1424));
    layer2_outputs(9598) <= not(layer1_outputs(1539)) or (layer1_outputs(10060));
    layer2_outputs(9599) <= layer1_outputs(9051);
    layer2_outputs(9600) <= layer1_outputs(4217);
    layer2_outputs(9601) <= layer1_outputs(8349);
    layer2_outputs(9602) <= not((layer1_outputs(3960)) xor (layer1_outputs(6720)));
    layer2_outputs(9603) <= not(layer1_outputs(8419));
    layer2_outputs(9604) <= layer1_outputs(2372);
    layer2_outputs(9605) <= (layer1_outputs(519)) or (layer1_outputs(1644));
    layer2_outputs(9606) <= not(layer1_outputs(1292));
    layer2_outputs(9607) <= not(layer1_outputs(7217));
    layer2_outputs(9608) <= layer1_outputs(3069);
    layer2_outputs(9609) <= (layer1_outputs(5493)) or (layer1_outputs(4449));
    layer2_outputs(9610) <= not(layer1_outputs(6143));
    layer2_outputs(9611) <= not((layer1_outputs(2813)) or (layer1_outputs(4452)));
    layer2_outputs(9612) <= (layer1_outputs(8753)) xor (layer1_outputs(3207));
    layer2_outputs(9613) <= not(layer1_outputs(5789));
    layer2_outputs(9614) <= layer1_outputs(5574);
    layer2_outputs(9615) <= (layer1_outputs(1831)) or (layer1_outputs(4704));
    layer2_outputs(9616) <= not(layer1_outputs(2641));
    layer2_outputs(9617) <= not(layer1_outputs(5863));
    layer2_outputs(9618) <= not(layer1_outputs(7013));
    layer2_outputs(9619) <= '0';
    layer2_outputs(9620) <= (layer1_outputs(3990)) or (layer1_outputs(5405));
    layer2_outputs(9621) <= not(layer1_outputs(5874));
    layer2_outputs(9622) <= (layer1_outputs(9265)) and (layer1_outputs(8441));
    layer2_outputs(9623) <= not(layer1_outputs(1118));
    layer2_outputs(9624) <= layer1_outputs(8647);
    layer2_outputs(9625) <= not((layer1_outputs(5454)) and (layer1_outputs(1720)));
    layer2_outputs(9626) <= not((layer1_outputs(1073)) and (layer1_outputs(10207)));
    layer2_outputs(9627) <= not((layer1_outputs(8770)) xor (layer1_outputs(5551)));
    layer2_outputs(9628) <= not(layer1_outputs(7171)) or (layer1_outputs(5270));
    layer2_outputs(9629) <= not((layer1_outputs(9223)) or (layer1_outputs(5571)));
    layer2_outputs(9630) <= not(layer1_outputs(2024));
    layer2_outputs(9631) <= layer1_outputs(2255);
    layer2_outputs(9632) <= layer1_outputs(5472);
    layer2_outputs(9633) <= layer1_outputs(3432);
    layer2_outputs(9634) <= not((layer1_outputs(1749)) and (layer1_outputs(413)));
    layer2_outputs(9635) <= not(layer1_outputs(720));
    layer2_outputs(9636) <= (layer1_outputs(6112)) and (layer1_outputs(6022));
    layer2_outputs(9637) <= not(layer1_outputs(810));
    layer2_outputs(9638) <= not(layer1_outputs(157));
    layer2_outputs(9639) <= not((layer1_outputs(5774)) or (layer1_outputs(2739)));
    layer2_outputs(9640) <= layer1_outputs(1864);
    layer2_outputs(9641) <= (layer1_outputs(7910)) and not (layer1_outputs(6536));
    layer2_outputs(9642) <= not(layer1_outputs(2864));
    layer2_outputs(9643) <= (layer1_outputs(1512)) or (layer1_outputs(2773));
    layer2_outputs(9644) <= (layer1_outputs(5708)) xor (layer1_outputs(7926));
    layer2_outputs(9645) <= layer1_outputs(8080);
    layer2_outputs(9646) <= not(layer1_outputs(9998));
    layer2_outputs(9647) <= not(layer1_outputs(3699));
    layer2_outputs(9648) <= not(layer1_outputs(4617));
    layer2_outputs(9649) <= not(layer1_outputs(9902));
    layer2_outputs(9650) <= not(layer1_outputs(9528));
    layer2_outputs(9651) <= layer1_outputs(1878);
    layer2_outputs(9652) <= layer1_outputs(8072);
    layer2_outputs(9653) <= not((layer1_outputs(1197)) xor (layer1_outputs(8829)));
    layer2_outputs(9654) <= (layer1_outputs(6111)) xor (layer1_outputs(7869));
    layer2_outputs(9655) <= (layer1_outputs(3582)) and (layer1_outputs(4939));
    layer2_outputs(9656) <= not((layer1_outputs(1616)) and (layer1_outputs(6840)));
    layer2_outputs(9657) <= not(layer1_outputs(2365));
    layer2_outputs(9658) <= layer1_outputs(7009);
    layer2_outputs(9659) <= not(layer1_outputs(1908));
    layer2_outputs(9660) <= layer1_outputs(8556);
    layer2_outputs(9661) <= not(layer1_outputs(8717));
    layer2_outputs(9662) <= not(layer1_outputs(4111));
    layer2_outputs(9663) <= not(layer1_outputs(6728));
    layer2_outputs(9664) <= not(layer1_outputs(4204));
    layer2_outputs(9665) <= (layer1_outputs(346)) or (layer1_outputs(2336));
    layer2_outputs(9666) <= not(layer1_outputs(7978));
    layer2_outputs(9667) <= layer1_outputs(6421);
    layer2_outputs(9668) <= not(layer1_outputs(8045));
    layer2_outputs(9669) <= not((layer1_outputs(4928)) xor (layer1_outputs(7038)));
    layer2_outputs(9670) <= not(layer1_outputs(3191));
    layer2_outputs(9671) <= not(layer1_outputs(4207));
    layer2_outputs(9672) <= layer1_outputs(10079);
    layer2_outputs(9673) <= (layer1_outputs(8223)) xor (layer1_outputs(6121));
    layer2_outputs(9674) <= layer1_outputs(6735);
    layer2_outputs(9675) <= not(layer1_outputs(5351));
    layer2_outputs(9676) <= not(layer1_outputs(5303)) or (layer1_outputs(1599));
    layer2_outputs(9677) <= layer1_outputs(3662);
    layer2_outputs(9678) <= (layer1_outputs(6893)) and not (layer1_outputs(7289));
    layer2_outputs(9679) <= not((layer1_outputs(8754)) xor (layer1_outputs(9075)));
    layer2_outputs(9680) <= layer1_outputs(9814);
    layer2_outputs(9681) <= not(layer1_outputs(2304));
    layer2_outputs(9682) <= not((layer1_outputs(8235)) or (layer1_outputs(3159)));
    layer2_outputs(9683) <= (layer1_outputs(3199)) and (layer1_outputs(7386));
    layer2_outputs(9684) <= layer1_outputs(5394);
    layer2_outputs(9685) <= '1';
    layer2_outputs(9686) <= not(layer1_outputs(8480));
    layer2_outputs(9687) <= layer1_outputs(861);
    layer2_outputs(9688) <= layer1_outputs(6166);
    layer2_outputs(9689) <= (layer1_outputs(8674)) and (layer1_outputs(1598));
    layer2_outputs(9690) <= layer1_outputs(1607);
    layer2_outputs(9691) <= layer1_outputs(9680);
    layer2_outputs(9692) <= layer1_outputs(34);
    layer2_outputs(9693) <= not(layer1_outputs(3020));
    layer2_outputs(9694) <= not(layer1_outputs(4764));
    layer2_outputs(9695) <= (layer1_outputs(595)) and (layer1_outputs(8731));
    layer2_outputs(9696) <= not((layer1_outputs(3178)) or (layer1_outputs(1866)));
    layer2_outputs(9697) <= layer1_outputs(10012);
    layer2_outputs(9698) <= not((layer1_outputs(7627)) and (layer1_outputs(3271)));
    layer2_outputs(9699) <= layer1_outputs(2211);
    layer2_outputs(9700) <= layer1_outputs(2110);
    layer2_outputs(9701) <= (layer1_outputs(9315)) or (layer1_outputs(1863));
    layer2_outputs(9702) <= (layer1_outputs(7508)) and not (layer1_outputs(9058));
    layer2_outputs(9703) <= layer1_outputs(3023);
    layer2_outputs(9704) <= layer1_outputs(3404);
    layer2_outputs(9705) <= not(layer1_outputs(8224));
    layer2_outputs(9706) <= (layer1_outputs(3121)) and (layer1_outputs(2730));
    layer2_outputs(9707) <= not(layer1_outputs(5109));
    layer2_outputs(9708) <= layer1_outputs(6854);
    layer2_outputs(9709) <= not(layer1_outputs(6117));
    layer2_outputs(9710) <= not((layer1_outputs(3439)) xor (layer1_outputs(4012)));
    layer2_outputs(9711) <= not(layer1_outputs(9640));
    layer2_outputs(9712) <= layer1_outputs(6662);
    layer2_outputs(9713) <= not(layer1_outputs(6091)) or (layer1_outputs(5269));
    layer2_outputs(9714) <= not((layer1_outputs(6099)) and (layer1_outputs(7439)));
    layer2_outputs(9715) <= not(layer1_outputs(8236));
    layer2_outputs(9716) <= not((layer1_outputs(9304)) and (layer1_outputs(690)));
    layer2_outputs(9717) <= not(layer1_outputs(2612));
    layer2_outputs(9718) <= not(layer1_outputs(6236));
    layer2_outputs(9719) <= (layer1_outputs(2076)) and (layer1_outputs(4029));
    layer2_outputs(9720) <= (layer1_outputs(6417)) and not (layer1_outputs(8199));
    layer2_outputs(9721) <= layer1_outputs(9718);
    layer2_outputs(9722) <= layer1_outputs(4088);
    layer2_outputs(9723) <= not(layer1_outputs(311));
    layer2_outputs(9724) <= not((layer1_outputs(9884)) xor (layer1_outputs(2704)));
    layer2_outputs(9725) <= layer1_outputs(9013);
    layer2_outputs(9726) <= layer1_outputs(877);
    layer2_outputs(9727) <= not(layer1_outputs(5009)) or (layer1_outputs(4374));
    layer2_outputs(9728) <= not(layer1_outputs(5275));
    layer2_outputs(9729) <= not(layer1_outputs(6110));
    layer2_outputs(9730) <= layer1_outputs(125);
    layer2_outputs(9731) <= not((layer1_outputs(872)) or (layer1_outputs(6294)));
    layer2_outputs(9732) <= layer1_outputs(2454);
    layer2_outputs(9733) <= not(layer1_outputs(8451));
    layer2_outputs(9734) <= not((layer1_outputs(736)) xor (layer1_outputs(4327)));
    layer2_outputs(9735) <= (layer1_outputs(2027)) and not (layer1_outputs(7827));
    layer2_outputs(9736) <= layer1_outputs(7408);
    layer2_outputs(9737) <= not((layer1_outputs(8141)) xor (layer1_outputs(9800)));
    layer2_outputs(9738) <= layer1_outputs(1703);
    layer2_outputs(9739) <= (layer1_outputs(997)) and not (layer1_outputs(8659));
    layer2_outputs(9740) <= layer1_outputs(9303);
    layer2_outputs(9741) <= not(layer1_outputs(4644));
    layer2_outputs(9742) <= not(layer1_outputs(5978));
    layer2_outputs(9743) <= layer1_outputs(4515);
    layer2_outputs(9744) <= not(layer1_outputs(2095));
    layer2_outputs(9745) <= not(layer1_outputs(5276));
    layer2_outputs(9746) <= not((layer1_outputs(7488)) xor (layer1_outputs(6057)));
    layer2_outputs(9747) <= not((layer1_outputs(4706)) xor (layer1_outputs(3430)));
    layer2_outputs(9748) <= not(layer1_outputs(1175)) or (layer1_outputs(7683));
    layer2_outputs(9749) <= not(layer1_outputs(2705));
    layer2_outputs(9750) <= (layer1_outputs(8568)) or (layer1_outputs(1702));
    layer2_outputs(9751) <= not(layer1_outputs(5906));
    layer2_outputs(9752) <= '1';
    layer2_outputs(9753) <= not(layer1_outputs(1936));
    layer2_outputs(9754) <= layer1_outputs(6334);
    layer2_outputs(9755) <= not(layer1_outputs(2114));
    layer2_outputs(9756) <= (layer1_outputs(8878)) xor (layer1_outputs(2064));
    layer2_outputs(9757) <= (layer1_outputs(8934)) or (layer1_outputs(1905));
    layer2_outputs(9758) <= layer1_outputs(3959);
    layer2_outputs(9759) <= not((layer1_outputs(9827)) or (layer1_outputs(1229)));
    layer2_outputs(9760) <= (layer1_outputs(74)) and not (layer1_outputs(8964));
    layer2_outputs(9761) <= layer1_outputs(2829);
    layer2_outputs(9762) <= not(layer1_outputs(240));
    layer2_outputs(9763) <= (layer1_outputs(7670)) and not (layer1_outputs(9673));
    layer2_outputs(9764) <= not(layer1_outputs(6512));
    layer2_outputs(9765) <= layer1_outputs(1805);
    layer2_outputs(9766) <= not((layer1_outputs(4078)) xor (layer1_outputs(2775)));
    layer2_outputs(9767) <= not(layer1_outputs(18)) or (layer1_outputs(7586));
    layer2_outputs(9768) <= layer1_outputs(2969);
    layer2_outputs(9769) <= layer1_outputs(993);
    layer2_outputs(9770) <= not(layer1_outputs(2374));
    layer2_outputs(9771) <= not(layer1_outputs(8229));
    layer2_outputs(9772) <= layer1_outputs(1434);
    layer2_outputs(9773) <= (layer1_outputs(8168)) and not (layer1_outputs(4799));
    layer2_outputs(9774) <= not(layer1_outputs(8366));
    layer2_outputs(9775) <= layer1_outputs(10052);
    layer2_outputs(9776) <= (layer1_outputs(859)) and not (layer1_outputs(8261));
    layer2_outputs(9777) <= (layer1_outputs(5228)) and (layer1_outputs(903));
    layer2_outputs(9778) <= not((layer1_outputs(9921)) and (layer1_outputs(286)));
    layer2_outputs(9779) <= not((layer1_outputs(5462)) and (layer1_outputs(4548)));
    layer2_outputs(9780) <= not(layer1_outputs(2222));
    layer2_outputs(9781) <= not(layer1_outputs(5914));
    layer2_outputs(9782) <= (layer1_outputs(4338)) and not (layer1_outputs(2315));
    layer2_outputs(9783) <= (layer1_outputs(1208)) and not (layer1_outputs(3066));
    layer2_outputs(9784) <= layer1_outputs(4914);
    layer2_outputs(9785) <= layer1_outputs(10125);
    layer2_outputs(9786) <= not(layer1_outputs(7700)) or (layer1_outputs(8126));
    layer2_outputs(9787) <= not(layer1_outputs(4653));
    layer2_outputs(9788) <= layer1_outputs(6255);
    layer2_outputs(9789) <= (layer1_outputs(9006)) and not (layer1_outputs(275));
    layer2_outputs(9790) <= not((layer1_outputs(7422)) xor (layer1_outputs(261)));
    layer2_outputs(9791) <= (layer1_outputs(4234)) or (layer1_outputs(3619));
    layer2_outputs(9792) <= layer1_outputs(1668);
    layer2_outputs(9793) <= not((layer1_outputs(1887)) xor (layer1_outputs(4328)));
    layer2_outputs(9794) <= not((layer1_outputs(4193)) xor (layer1_outputs(5880)));
    layer2_outputs(9795) <= not(layer1_outputs(2119)) or (layer1_outputs(7242));
    layer2_outputs(9796) <= not(layer1_outputs(7843));
    layer2_outputs(9797) <= layer1_outputs(5350);
    layer2_outputs(9798) <= not(layer1_outputs(2225));
    layer2_outputs(9799) <= layer1_outputs(1605);
    layer2_outputs(9800) <= '0';
    layer2_outputs(9801) <= '1';
    layer2_outputs(9802) <= not(layer1_outputs(2033));
    layer2_outputs(9803) <= not(layer1_outputs(4687));
    layer2_outputs(9804) <= not((layer1_outputs(7174)) xor (layer1_outputs(9539)));
    layer2_outputs(9805) <= not(layer1_outputs(7583)) or (layer1_outputs(5906));
    layer2_outputs(9806) <= layer1_outputs(1464);
    layer2_outputs(9807) <= not(layer1_outputs(9027));
    layer2_outputs(9808) <= layer1_outputs(6616);
    layer2_outputs(9809) <= layer1_outputs(4411);
    layer2_outputs(9810) <= not((layer1_outputs(1504)) xor (layer1_outputs(7965)));
    layer2_outputs(9811) <= not(layer1_outputs(7571)) or (layer1_outputs(5945));
    layer2_outputs(9812) <= layer1_outputs(7758);
    layer2_outputs(9813) <= not((layer1_outputs(8701)) or (layer1_outputs(8775)));
    layer2_outputs(9814) <= not(layer1_outputs(9470));
    layer2_outputs(9815) <= not(layer1_outputs(485));
    layer2_outputs(9816) <= not(layer1_outputs(2490));
    layer2_outputs(9817) <= not(layer1_outputs(8296));
    layer2_outputs(9818) <= not(layer1_outputs(6539)) or (layer1_outputs(8697));
    layer2_outputs(9819) <= not(layer1_outputs(7426)) or (layer1_outputs(2019));
    layer2_outputs(9820) <= not((layer1_outputs(6436)) and (layer1_outputs(4937)));
    layer2_outputs(9821) <= layer1_outputs(4263);
    layer2_outputs(9822) <= (layer1_outputs(19)) and (layer1_outputs(3275));
    layer2_outputs(9823) <= layer1_outputs(1013);
    layer2_outputs(9824) <= not(layer1_outputs(3388));
    layer2_outputs(9825) <= layer1_outputs(4222);
    layer2_outputs(9826) <= layer1_outputs(1439);
    layer2_outputs(9827) <= layer1_outputs(1914);
    layer2_outputs(9828) <= not(layer1_outputs(319)) or (layer1_outputs(5928));
    layer2_outputs(9829) <= not(layer1_outputs(3889));
    layer2_outputs(9830) <= not(layer1_outputs(8604));
    layer2_outputs(9831) <= not(layer1_outputs(4175));
    layer2_outputs(9832) <= (layer1_outputs(9157)) and not (layer1_outputs(2220));
    layer2_outputs(9833) <= layer1_outputs(5373);
    layer2_outputs(9834) <= not(layer1_outputs(4521));
    layer2_outputs(9835) <= layer1_outputs(8915);
    layer2_outputs(9836) <= (layer1_outputs(191)) or (layer1_outputs(5883));
    layer2_outputs(9837) <= not(layer1_outputs(6162));
    layer2_outputs(9838) <= not(layer1_outputs(6552)) or (layer1_outputs(2837));
    layer2_outputs(9839) <= not(layer1_outputs(5470));
    layer2_outputs(9840) <= (layer1_outputs(1136)) and not (layer1_outputs(1493));
    layer2_outputs(9841) <= not((layer1_outputs(3531)) xor (layer1_outputs(9653)));
    layer2_outputs(9842) <= not(layer1_outputs(6307));
    layer2_outputs(9843) <= layer1_outputs(7528);
    layer2_outputs(9844) <= not(layer1_outputs(7529));
    layer2_outputs(9845) <= not((layer1_outputs(9819)) xor (layer1_outputs(5459)));
    layer2_outputs(9846) <= layer1_outputs(6380);
    layer2_outputs(9847) <= (layer1_outputs(6493)) and not (layer1_outputs(2855));
    layer2_outputs(9848) <= (layer1_outputs(8253)) and not (layer1_outputs(647));
    layer2_outputs(9849) <= not(layer1_outputs(1814));
    layer2_outputs(9850) <= layer1_outputs(2983);
    layer2_outputs(9851) <= (layer1_outputs(2885)) or (layer1_outputs(4240));
    layer2_outputs(9852) <= not((layer1_outputs(10188)) xor (layer1_outputs(2850)));
    layer2_outputs(9853) <= (layer1_outputs(2527)) and not (layer1_outputs(6946));
    layer2_outputs(9854) <= (layer1_outputs(9586)) and not (layer1_outputs(4630));
    layer2_outputs(9855) <= layer1_outputs(6216);
    layer2_outputs(9856) <= (layer1_outputs(5817)) and not (layer1_outputs(3819));
    layer2_outputs(9857) <= not(layer1_outputs(3277));
    layer2_outputs(9858) <= not(layer1_outputs(5608));
    layer2_outputs(9859) <= layer1_outputs(4608);
    layer2_outputs(9860) <= layer1_outputs(5155);
    layer2_outputs(9861) <= (layer1_outputs(6858)) or (layer1_outputs(1728));
    layer2_outputs(9862) <= not(layer1_outputs(3610));
    layer2_outputs(9863) <= (layer1_outputs(8826)) xor (layer1_outputs(3680));
    layer2_outputs(9864) <= not((layer1_outputs(5199)) and (layer1_outputs(4843)));
    layer2_outputs(9865) <= not(layer1_outputs(8590)) or (layer1_outputs(214));
    layer2_outputs(9866) <= layer1_outputs(7129);
    layer2_outputs(9867) <= layer1_outputs(1746);
    layer2_outputs(9868) <= not(layer1_outputs(1541)) or (layer1_outputs(10134));
    layer2_outputs(9869) <= layer1_outputs(9875);
    layer2_outputs(9870) <= not((layer1_outputs(4339)) xor (layer1_outputs(5696)));
    layer2_outputs(9871) <= not((layer1_outputs(9608)) or (layer1_outputs(4320)));
    layer2_outputs(9872) <= not(layer1_outputs(8447));
    layer2_outputs(9873) <= not(layer1_outputs(8852));
    layer2_outputs(9874) <= '1';
    layer2_outputs(9875) <= not(layer1_outputs(6673)) or (layer1_outputs(8671));
    layer2_outputs(9876) <= layer1_outputs(6825);
    layer2_outputs(9877) <= (layer1_outputs(3492)) and not (layer1_outputs(9223));
    layer2_outputs(9878) <= not((layer1_outputs(5434)) xor (layer1_outputs(9655)));
    layer2_outputs(9879) <= not(layer1_outputs(4294));
    layer2_outputs(9880) <= not(layer1_outputs(8625));
    layer2_outputs(9881) <= layer1_outputs(893);
    layer2_outputs(9882) <= not((layer1_outputs(8497)) xor (layer1_outputs(6454)));
    layer2_outputs(9883) <= (layer1_outputs(9024)) and not (layer1_outputs(8943));
    layer2_outputs(9884) <= not(layer1_outputs(9847));
    layer2_outputs(9885) <= layer1_outputs(2699);
    layer2_outputs(9886) <= not((layer1_outputs(6437)) xor (layer1_outputs(5390)));
    layer2_outputs(9887) <= (layer1_outputs(6362)) and (layer1_outputs(1912));
    layer2_outputs(9888) <= (layer1_outputs(128)) and not (layer1_outputs(8187));
    layer2_outputs(9889) <= layer1_outputs(847);
    layer2_outputs(9890) <= layer1_outputs(6610);
    layer2_outputs(9891) <= '0';
    layer2_outputs(9892) <= layer1_outputs(8163);
    layer2_outputs(9893) <= (layer1_outputs(9249)) or (layer1_outputs(2865));
    layer2_outputs(9894) <= not(layer1_outputs(5338));
    layer2_outputs(9895) <= not(layer1_outputs(2303));
    layer2_outputs(9896) <= (layer1_outputs(3454)) and (layer1_outputs(5286));
    layer2_outputs(9897) <= not(layer1_outputs(1084));
    layer2_outputs(9898) <= not(layer1_outputs(3594));
    layer2_outputs(9899) <= '1';
    layer2_outputs(9900) <= not((layer1_outputs(9224)) and (layer1_outputs(3001)));
    layer2_outputs(9901) <= (layer1_outputs(7845)) xor (layer1_outputs(9074));
    layer2_outputs(9902) <= not(layer1_outputs(5327));
    layer2_outputs(9903) <= layer1_outputs(5738);
    layer2_outputs(9904) <= not(layer1_outputs(3110));
    layer2_outputs(9905) <= not(layer1_outputs(8887));
    layer2_outputs(9906) <= not(layer1_outputs(2022));
    layer2_outputs(9907) <= not(layer1_outputs(9578));
    layer2_outputs(9908) <= not((layer1_outputs(918)) or (layer1_outputs(2401)));
    layer2_outputs(9909) <= not(layer1_outputs(7592));
    layer2_outputs(9910) <= layer1_outputs(8359);
    layer2_outputs(9911) <= not(layer1_outputs(5725));
    layer2_outputs(9912) <= layer1_outputs(6742);
    layer2_outputs(9913) <= not((layer1_outputs(1127)) and (layer1_outputs(8015)));
    layer2_outputs(9914) <= not(layer1_outputs(4336)) or (layer1_outputs(2882));
    layer2_outputs(9915) <= layer1_outputs(1210);
    layer2_outputs(9916) <= not(layer1_outputs(7678));
    layer2_outputs(9917) <= layer1_outputs(9316);
    layer2_outputs(9918) <= (layer1_outputs(3471)) and (layer1_outputs(7393));
    layer2_outputs(9919) <= layer1_outputs(10150);
    layer2_outputs(9920) <= '1';
    layer2_outputs(9921) <= layer1_outputs(1574);
    layer2_outputs(9922) <= not((layer1_outputs(1052)) xor (layer1_outputs(8006)));
    layer2_outputs(9923) <= not((layer1_outputs(6573)) and (layer1_outputs(5126)));
    layer2_outputs(9924) <= layer1_outputs(5706);
    layer2_outputs(9925) <= not(layer1_outputs(7813));
    layer2_outputs(9926) <= not((layer1_outputs(454)) or (layer1_outputs(8324)));
    layer2_outputs(9927) <= (layer1_outputs(4093)) and not (layer1_outputs(1819));
    layer2_outputs(9928) <= (layer1_outputs(505)) or (layer1_outputs(549));
    layer2_outputs(9929) <= (layer1_outputs(2883)) and not (layer1_outputs(2421));
    layer2_outputs(9930) <= layer1_outputs(9790);
    layer2_outputs(9931) <= not(layer1_outputs(4703));
    layer2_outputs(9932) <= layer1_outputs(6111);
    layer2_outputs(9933) <= not(layer1_outputs(2663));
    layer2_outputs(9934) <= (layer1_outputs(8036)) xor (layer1_outputs(1884));
    layer2_outputs(9935) <= layer1_outputs(784);
    layer2_outputs(9936) <= not(layer1_outputs(6391));
    layer2_outputs(9937) <= (layer1_outputs(4927)) and not (layer1_outputs(2245));
    layer2_outputs(9938) <= (layer1_outputs(10185)) xor (layer1_outputs(9241));
    layer2_outputs(9939) <= layer1_outputs(3452);
    layer2_outputs(9940) <= layer1_outputs(766);
    layer2_outputs(9941) <= layer1_outputs(1706);
    layer2_outputs(9942) <= not(layer1_outputs(3629));
    layer2_outputs(9943) <= not(layer1_outputs(3507));
    layer2_outputs(9944) <= (layer1_outputs(1189)) xor (layer1_outputs(7510));
    layer2_outputs(9945) <= (layer1_outputs(7006)) and not (layer1_outputs(264));
    layer2_outputs(9946) <= not(layer1_outputs(8523));
    layer2_outputs(9947) <= not(layer1_outputs(3303));
    layer2_outputs(9948) <= layer1_outputs(7238);
    layer2_outputs(9949) <= (layer1_outputs(5000)) and not (layer1_outputs(4738));
    layer2_outputs(9950) <= (layer1_outputs(9047)) and (layer1_outputs(7438));
    layer2_outputs(9951) <= layer1_outputs(9785);
    layer2_outputs(9952) <= not(layer1_outputs(4129));
    layer2_outputs(9953) <= not(layer1_outputs(4737)) or (layer1_outputs(9368));
    layer2_outputs(9954) <= layer1_outputs(7948);
    layer2_outputs(9955) <= not((layer1_outputs(9480)) and (layer1_outputs(8679)));
    layer2_outputs(9956) <= not(layer1_outputs(6818));
    layer2_outputs(9957) <= not((layer1_outputs(5453)) xor (layer1_outputs(1372)));
    layer2_outputs(9958) <= (layer1_outputs(9227)) or (layer1_outputs(2053));
    layer2_outputs(9959) <= not(layer1_outputs(6567));
    layer2_outputs(9960) <= (layer1_outputs(7882)) xor (layer1_outputs(894));
    layer2_outputs(9961) <= not((layer1_outputs(6370)) xor (layer1_outputs(9601)));
    layer2_outputs(9962) <= layer1_outputs(1245);
    layer2_outputs(9963) <= not(layer1_outputs(2116));
    layer2_outputs(9964) <= (layer1_outputs(7424)) and not (layer1_outputs(357));
    layer2_outputs(9965) <= layer1_outputs(9012);
    layer2_outputs(9966) <= not(layer1_outputs(7586));
    layer2_outputs(9967) <= not(layer1_outputs(9432));
    layer2_outputs(9968) <= not(layer1_outputs(8460));
    layer2_outputs(9969) <= layer1_outputs(6309);
    layer2_outputs(9970) <= not((layer1_outputs(10215)) xor (layer1_outputs(9042)));
    layer2_outputs(9971) <= (layer1_outputs(7538)) xor (layer1_outputs(2840));
    layer2_outputs(9972) <= not(layer1_outputs(6357));
    layer2_outputs(9973) <= not((layer1_outputs(13)) xor (layer1_outputs(9162)));
    layer2_outputs(9974) <= not(layer1_outputs(654));
    layer2_outputs(9975) <= (layer1_outputs(3468)) and (layer1_outputs(3339));
    layer2_outputs(9976) <= (layer1_outputs(10015)) and not (layer1_outputs(1072));
    layer2_outputs(9977) <= (layer1_outputs(5487)) and not (layer1_outputs(8733));
    layer2_outputs(9978) <= (layer1_outputs(10022)) or (layer1_outputs(3063));
    layer2_outputs(9979) <= not((layer1_outputs(6939)) and (layer1_outputs(7591)));
    layer2_outputs(9980) <= not(layer1_outputs(6144));
    layer2_outputs(9981) <= layer1_outputs(4541);
    layer2_outputs(9982) <= not(layer1_outputs(9679));
    layer2_outputs(9983) <= (layer1_outputs(8664)) and (layer1_outputs(5947));
    layer2_outputs(9984) <= '1';
    layer2_outputs(9985) <= layer1_outputs(4825);
    layer2_outputs(9986) <= (layer1_outputs(5648)) and not (layer1_outputs(9627));
    layer2_outputs(9987) <= not(layer1_outputs(368));
    layer2_outputs(9988) <= (layer1_outputs(1441)) and not (layer1_outputs(8767));
    layer2_outputs(9989) <= not(layer1_outputs(798));
    layer2_outputs(9990) <= not(layer1_outputs(7853)) or (layer1_outputs(6153));
    layer2_outputs(9991) <= (layer1_outputs(579)) xor (layer1_outputs(395));
    layer2_outputs(9992) <= not(layer1_outputs(8354));
    layer2_outputs(9993) <= layer1_outputs(1216);
    layer2_outputs(9994) <= not(layer1_outputs(10210));
    layer2_outputs(9995) <= not(layer1_outputs(4215));
    layer2_outputs(9996) <= layer1_outputs(5965);
    layer2_outputs(9997) <= layer1_outputs(1923);
    layer2_outputs(9998) <= layer1_outputs(5026);
    layer2_outputs(9999) <= not(layer1_outputs(9357));
    layer2_outputs(10000) <= not(layer1_outputs(8221)) or (layer1_outputs(3609));
    layer2_outputs(10001) <= not(layer1_outputs(4454));
    layer2_outputs(10002) <= layer1_outputs(312);
    layer2_outputs(10003) <= (layer1_outputs(886)) and (layer1_outputs(7292));
    layer2_outputs(10004) <= layer1_outputs(530);
    layer2_outputs(10005) <= (layer1_outputs(1825)) and not (layer1_outputs(1440));
    layer2_outputs(10006) <= layer1_outputs(3759);
    layer2_outputs(10007) <= layer1_outputs(4355);
    layer2_outputs(10008) <= layer1_outputs(6690);
    layer2_outputs(10009) <= not(layer1_outputs(8454));
    layer2_outputs(10010) <= layer1_outputs(10196);
    layer2_outputs(10011) <= not(layer1_outputs(3335));
    layer2_outputs(10012) <= not(layer1_outputs(3395)) or (layer1_outputs(6450));
    layer2_outputs(10013) <= not(layer1_outputs(9345));
    layer2_outputs(10014) <= not(layer1_outputs(6042));
    layer2_outputs(10015) <= not((layer1_outputs(5054)) or (layer1_outputs(8010)));
    layer2_outputs(10016) <= not((layer1_outputs(1818)) xor (layer1_outputs(5178)));
    layer2_outputs(10017) <= (layer1_outputs(3349)) and (layer1_outputs(994));
    layer2_outputs(10018) <= not(layer1_outputs(4702));
    layer2_outputs(10019) <= not(layer1_outputs(6959));
    layer2_outputs(10020) <= (layer1_outputs(6339)) and not (layer1_outputs(1398));
    layer2_outputs(10021) <= not(layer1_outputs(1988)) or (layer1_outputs(3241));
    layer2_outputs(10022) <= not(layer1_outputs(9475));
    layer2_outputs(10023) <= layer1_outputs(2018);
    layer2_outputs(10024) <= (layer1_outputs(4784)) xor (layer1_outputs(8786));
    layer2_outputs(10025) <= (layer1_outputs(3970)) and (layer1_outputs(3601));
    layer2_outputs(10026) <= layer1_outputs(2637);
    layer2_outputs(10027) <= not((layer1_outputs(1679)) and (layer1_outputs(3566)));
    layer2_outputs(10028) <= not(layer1_outputs(3079));
    layer2_outputs(10029) <= not(layer1_outputs(4437));
    layer2_outputs(10030) <= not(layer1_outputs(7543));
    layer2_outputs(10031) <= not(layer1_outputs(898));
    layer2_outputs(10032) <= layer1_outputs(5874);
    layer2_outputs(10033) <= (layer1_outputs(1448)) and (layer1_outputs(757));
    layer2_outputs(10034) <= not(layer1_outputs(9352));
    layer2_outputs(10035) <= layer1_outputs(1928);
    layer2_outputs(10036) <= (layer1_outputs(6349)) xor (layer1_outputs(2373));
    layer2_outputs(10037) <= not((layer1_outputs(795)) xor (layer1_outputs(3110)));
    layer2_outputs(10038) <= not(layer1_outputs(1110));
    layer2_outputs(10039) <= not(layer1_outputs(3006)) or (layer1_outputs(9380));
    layer2_outputs(10040) <= not(layer1_outputs(8846));
    layer2_outputs(10041) <= (layer1_outputs(925)) and (layer1_outputs(6948));
    layer2_outputs(10042) <= layer1_outputs(1144);
    layer2_outputs(10043) <= not(layer1_outputs(7971));
    layer2_outputs(10044) <= layer1_outputs(776);
    layer2_outputs(10045) <= layer1_outputs(6556);
    layer2_outputs(10046) <= not((layer1_outputs(7830)) and (layer1_outputs(7291)));
    layer2_outputs(10047) <= not(layer1_outputs(7246)) or (layer1_outputs(3909));
    layer2_outputs(10048) <= not((layer1_outputs(5031)) or (layer1_outputs(1445)));
    layer2_outputs(10049) <= layer1_outputs(5772);
    layer2_outputs(10050) <= not((layer1_outputs(5366)) or (layer1_outputs(2223)));
    layer2_outputs(10051) <= layer1_outputs(3118);
    layer2_outputs(10052) <= not(layer1_outputs(1900));
    layer2_outputs(10053) <= (layer1_outputs(3366)) and not (layer1_outputs(1625));
    layer2_outputs(10054) <= not(layer1_outputs(6381));
    layer2_outputs(10055) <= not((layer1_outputs(8682)) xor (layer1_outputs(611)));
    layer2_outputs(10056) <= not((layer1_outputs(4838)) xor (layer1_outputs(2590)));
    layer2_outputs(10057) <= layer1_outputs(5202);
    layer2_outputs(10058) <= layer1_outputs(7426);
    layer2_outputs(10059) <= (layer1_outputs(8805)) and (layer1_outputs(97));
    layer2_outputs(10060) <= not(layer1_outputs(7848));
    layer2_outputs(10061) <= not((layer1_outputs(6638)) xor (layer1_outputs(9096)));
    layer2_outputs(10062) <= layer1_outputs(4744);
    layer2_outputs(10063) <= not(layer1_outputs(2226));
    layer2_outputs(10064) <= layer1_outputs(6871);
    layer2_outputs(10065) <= not(layer1_outputs(7589));
    layer2_outputs(10066) <= (layer1_outputs(978)) xor (layer1_outputs(1658));
    layer2_outputs(10067) <= layer1_outputs(149);
    layer2_outputs(10068) <= layer1_outputs(2412);
    layer2_outputs(10069) <= not(layer1_outputs(9776));
    layer2_outputs(10070) <= not((layer1_outputs(4549)) or (layer1_outputs(9142)));
    layer2_outputs(10071) <= not(layer1_outputs(6804)) or (layer1_outputs(2689));
    layer2_outputs(10072) <= (layer1_outputs(9969)) and (layer1_outputs(2127));
    layer2_outputs(10073) <= (layer1_outputs(109)) and not (layer1_outputs(4569));
    layer2_outputs(10074) <= (layer1_outputs(3467)) xor (layer1_outputs(7726));
    layer2_outputs(10075) <= not(layer1_outputs(9090)) or (layer1_outputs(5913));
    layer2_outputs(10076) <= not((layer1_outputs(9138)) xor (layer1_outputs(9771)));
    layer2_outputs(10077) <= (layer1_outputs(2437)) and not (layer1_outputs(8018));
    layer2_outputs(10078) <= not(layer1_outputs(8862));
    layer2_outputs(10079) <= not((layer1_outputs(8007)) xor (layer1_outputs(8311)));
    layer2_outputs(10080) <= (layer1_outputs(4046)) and (layer1_outputs(6990));
    layer2_outputs(10081) <= layer1_outputs(2457);
    layer2_outputs(10082) <= layer1_outputs(6958);
    layer2_outputs(10083) <= (layer1_outputs(3770)) xor (layer1_outputs(907));
    layer2_outputs(10084) <= not((layer1_outputs(8471)) xor (layer1_outputs(9246)));
    layer2_outputs(10085) <= layer1_outputs(5609);
    layer2_outputs(10086) <= layer1_outputs(1240);
    layer2_outputs(10087) <= (layer1_outputs(1097)) and not (layer1_outputs(3870));
    layer2_outputs(10088) <= not(layer1_outputs(4691));
    layer2_outputs(10089) <= (layer1_outputs(2037)) or (layer1_outputs(1977));
    layer2_outputs(10090) <= not(layer1_outputs(546)) or (layer1_outputs(6218));
    layer2_outputs(10091) <= not(layer1_outputs(5719));
    layer2_outputs(10092) <= layer1_outputs(1897);
    layer2_outputs(10093) <= not(layer1_outputs(7660));
    layer2_outputs(10094) <= not(layer1_outputs(5151));
    layer2_outputs(10095) <= not(layer1_outputs(688)) or (layer1_outputs(3926));
    layer2_outputs(10096) <= not(layer1_outputs(6757));
    layer2_outputs(10097) <= not(layer1_outputs(2203));
    layer2_outputs(10098) <= (layer1_outputs(156)) and not (layer1_outputs(10180));
    layer2_outputs(10099) <= (layer1_outputs(8222)) and (layer1_outputs(3502));
    layer2_outputs(10100) <= not(layer1_outputs(849));
    layer2_outputs(10101) <= not(layer1_outputs(8663));
    layer2_outputs(10102) <= not(layer1_outputs(3141));
    layer2_outputs(10103) <= layer1_outputs(4241);
    layer2_outputs(10104) <= not((layer1_outputs(9783)) or (layer1_outputs(318)));
    layer2_outputs(10105) <= not((layer1_outputs(5546)) or (layer1_outputs(5122)));
    layer2_outputs(10106) <= (layer1_outputs(9431)) and not (layer1_outputs(7541));
    layer2_outputs(10107) <= (layer1_outputs(5821)) and not (layer1_outputs(7595));
    layer2_outputs(10108) <= not((layer1_outputs(9076)) xor (layer1_outputs(3373)));
    layer2_outputs(10109) <= layer1_outputs(1244);
    layer2_outputs(10110) <= not((layer1_outputs(1023)) and (layer1_outputs(5671)));
    layer2_outputs(10111) <= not(layer1_outputs(7177));
    layer2_outputs(10112) <= not((layer1_outputs(10212)) xor (layer1_outputs(8314)));
    layer2_outputs(10113) <= not(layer1_outputs(9334));
    layer2_outputs(10114) <= not((layer1_outputs(6048)) xor (layer1_outputs(7434)));
    layer2_outputs(10115) <= layer1_outputs(1667);
    layer2_outputs(10116) <= not(layer1_outputs(1543)) or (layer1_outputs(3710));
    layer2_outputs(10117) <= not((layer1_outputs(40)) xor (layer1_outputs(6172)));
    layer2_outputs(10118) <= not(layer1_outputs(5645));
    layer2_outputs(10119) <= layer1_outputs(6400);
    layer2_outputs(10120) <= not(layer1_outputs(6329));
    layer2_outputs(10121) <= layer1_outputs(1940);
    layer2_outputs(10122) <= not((layer1_outputs(6548)) or (layer1_outputs(8021)));
    layer2_outputs(10123) <= layer1_outputs(5278);
    layer2_outputs(10124) <= not(layer1_outputs(6154));
    layer2_outputs(10125) <= (layer1_outputs(7727)) and not (layer1_outputs(3332));
    layer2_outputs(10126) <= not(layer1_outputs(3993));
    layer2_outputs(10127) <= not((layer1_outputs(1171)) or (layer1_outputs(7235)));
    layer2_outputs(10128) <= not(layer1_outputs(10041));
    layer2_outputs(10129) <= not((layer1_outputs(4535)) or (layer1_outputs(9737)));
    layer2_outputs(10130) <= (layer1_outputs(3196)) xor (layer1_outputs(2409));
    layer2_outputs(10131) <= (layer1_outputs(1781)) or (layer1_outputs(236));
    layer2_outputs(10132) <= (layer1_outputs(7030)) xor (layer1_outputs(387));
    layer2_outputs(10133) <= '0';
    layer2_outputs(10134) <= layer1_outputs(3478);
    layer2_outputs(10135) <= (layer1_outputs(4140)) or (layer1_outputs(9887));
    layer2_outputs(10136) <= not(layer1_outputs(8105)) or (layer1_outputs(4530));
    layer2_outputs(10137) <= layer1_outputs(1085);
    layer2_outputs(10138) <= '0';
    layer2_outputs(10139) <= layer1_outputs(3664);
    layer2_outputs(10140) <= layer1_outputs(183);
    layer2_outputs(10141) <= (layer1_outputs(1378)) and not (layer1_outputs(5178));
    layer2_outputs(10142) <= not(layer1_outputs(4288));
    layer2_outputs(10143) <= not((layer1_outputs(9129)) or (layer1_outputs(8841)));
    layer2_outputs(10144) <= not(layer1_outputs(2910)) or (layer1_outputs(156));
    layer2_outputs(10145) <= layer1_outputs(5028);
    layer2_outputs(10146) <= layer1_outputs(9252);
    layer2_outputs(10147) <= layer1_outputs(10106);
    layer2_outputs(10148) <= (layer1_outputs(2272)) and not (layer1_outputs(500));
    layer2_outputs(10149) <= not(layer1_outputs(1159));
    layer2_outputs(10150) <= not(layer1_outputs(9286));
    layer2_outputs(10151) <= not(layer1_outputs(3606)) or (layer1_outputs(4892));
    layer2_outputs(10152) <= layer1_outputs(4255);
    layer2_outputs(10153) <= (layer1_outputs(2301)) and not (layer1_outputs(7337));
    layer2_outputs(10154) <= layer1_outputs(1178);
    layer2_outputs(10155) <= layer1_outputs(8247);
    layer2_outputs(10156) <= not(layer1_outputs(7279)) or (layer1_outputs(4091));
    layer2_outputs(10157) <= (layer1_outputs(9092)) and (layer1_outputs(513));
    layer2_outputs(10158) <= not(layer1_outputs(1594)) or (layer1_outputs(4675));
    layer2_outputs(10159) <= not(layer1_outputs(9778));
    layer2_outputs(10160) <= (layer1_outputs(6391)) and (layer1_outputs(5391));
    layer2_outputs(10161) <= layer1_outputs(6137);
    layer2_outputs(10162) <= layer1_outputs(9620);
    layer2_outputs(10163) <= (layer1_outputs(5681)) or (layer1_outputs(9393));
    layer2_outputs(10164) <= not(layer1_outputs(4427));
    layer2_outputs(10165) <= not(layer1_outputs(1188));
    layer2_outputs(10166) <= layer1_outputs(8867);
    layer2_outputs(10167) <= not(layer1_outputs(8986)) or (layer1_outputs(10120));
    layer2_outputs(10168) <= (layer1_outputs(2178)) and (layer1_outputs(2194));
    layer2_outputs(10169) <= layer1_outputs(2913);
    layer2_outputs(10170) <= not((layer1_outputs(9577)) xor (layer1_outputs(7734)));
    layer2_outputs(10171) <= layer1_outputs(8011);
    layer2_outputs(10172) <= (layer1_outputs(4321)) and (layer1_outputs(639));
    layer2_outputs(10173) <= (layer1_outputs(2106)) and not (layer1_outputs(822));
    layer2_outputs(10174) <= not((layer1_outputs(3305)) xor (layer1_outputs(2345)));
    layer2_outputs(10175) <= not(layer1_outputs(315));
    layer2_outputs(10176) <= (layer1_outputs(6147)) xor (layer1_outputs(6808));
    layer2_outputs(10177) <= not(layer1_outputs(5011));
    layer2_outputs(10178) <= not(layer1_outputs(6313));
    layer2_outputs(10179) <= not(layer1_outputs(2215));
    layer2_outputs(10180) <= layer1_outputs(6149);
    layer2_outputs(10181) <= not(layer1_outputs(80));
    layer2_outputs(10182) <= layer1_outputs(7432);
    layer2_outputs(10183) <= layer1_outputs(6067);
    layer2_outputs(10184) <= (layer1_outputs(4564)) xor (layer1_outputs(9440));
    layer2_outputs(10185) <= (layer1_outputs(4901)) or (layer1_outputs(81));
    layer2_outputs(10186) <= (layer1_outputs(9489)) xor (layer1_outputs(275));
    layer2_outputs(10187) <= not((layer1_outputs(1294)) or (layer1_outputs(1090)));
    layer2_outputs(10188) <= (layer1_outputs(8823)) and (layer1_outputs(3724));
    layer2_outputs(10189) <= layer1_outputs(5683);
    layer2_outputs(10190) <= layer1_outputs(4951);
    layer2_outputs(10191) <= not(layer1_outputs(1132));
    layer2_outputs(10192) <= layer1_outputs(8288);
    layer2_outputs(10193) <= (layer1_outputs(5149)) and not (layer1_outputs(3028));
    layer2_outputs(10194) <= layer1_outputs(4728);
    layer2_outputs(10195) <= layer1_outputs(4988);
    layer2_outputs(10196) <= not(layer1_outputs(7260));
    layer2_outputs(10197) <= not(layer1_outputs(2239));
    layer2_outputs(10198) <= (layer1_outputs(1033)) and not (layer1_outputs(982));
    layer2_outputs(10199) <= (layer1_outputs(89)) or (layer1_outputs(627));
    layer2_outputs(10200) <= not((layer1_outputs(6767)) or (layer1_outputs(2750)));
    layer2_outputs(10201) <= not((layer1_outputs(2997)) or (layer1_outputs(6978)));
    layer2_outputs(10202) <= (layer1_outputs(6630)) and not (layer1_outputs(7194));
    layer2_outputs(10203) <= (layer1_outputs(2111)) xor (layer1_outputs(4926));
    layer2_outputs(10204) <= (layer1_outputs(597)) or (layer1_outputs(6912));
    layer2_outputs(10205) <= (layer1_outputs(6651)) and not (layer1_outputs(8713));
    layer2_outputs(10206) <= (layer1_outputs(1620)) xor (layer1_outputs(6923));
    layer2_outputs(10207) <= layer1_outputs(5584);
    layer2_outputs(10208) <= layer1_outputs(3981);
    layer2_outputs(10209) <= layer1_outputs(3504);
    layer2_outputs(10210) <= not((layer1_outputs(2109)) or (layer1_outputs(10163)));
    layer2_outputs(10211) <= not((layer1_outputs(557)) and (layer1_outputs(6751)));
    layer2_outputs(10212) <= (layer1_outputs(7204)) xor (layer1_outputs(9473));
    layer2_outputs(10213) <= layer1_outputs(5599);
    layer2_outputs(10214) <= not(layer1_outputs(977));
    layer2_outputs(10215) <= (layer1_outputs(8357)) and not (layer1_outputs(210));
    layer2_outputs(10216) <= not((layer1_outputs(8382)) xor (layer1_outputs(7554)));
    layer2_outputs(10217) <= layer1_outputs(9679);
    layer2_outputs(10218) <= layer1_outputs(2836);
    layer2_outputs(10219) <= layer1_outputs(4883);
    layer2_outputs(10220) <= layer1_outputs(735);
    layer2_outputs(10221) <= not((layer1_outputs(7707)) or (layer1_outputs(6336)));
    layer2_outputs(10222) <= not((layer1_outputs(6203)) and (layer1_outputs(4625)));
    layer2_outputs(10223) <= not(layer1_outputs(2310)) or (layer1_outputs(9734));
    layer2_outputs(10224) <= not(layer1_outputs(5787));
    layer2_outputs(10225) <= not((layer1_outputs(449)) or (layer1_outputs(708)));
    layer2_outputs(10226) <= layer1_outputs(6834);
    layer2_outputs(10227) <= not((layer1_outputs(8238)) and (layer1_outputs(7429)));
    layer2_outputs(10228) <= layer1_outputs(5476);
    layer2_outputs(10229) <= layer1_outputs(428);
    layer2_outputs(10230) <= (layer1_outputs(1718)) xor (layer1_outputs(8993));
    layer2_outputs(10231) <= not(layer1_outputs(7687));
    layer2_outputs(10232) <= layer1_outputs(9270);
    layer2_outputs(10233) <= (layer1_outputs(4457)) and not (layer1_outputs(4284));
    layer2_outputs(10234) <= not(layer1_outputs(8235)) or (layer1_outputs(9595));
    layer2_outputs(10235) <= not((layer1_outputs(725)) and (layer1_outputs(5703)));
    layer2_outputs(10236) <= (layer1_outputs(8789)) xor (layer1_outputs(4611));
    layer2_outputs(10237) <= not(layer1_outputs(9979));
    layer2_outputs(10238) <= not(layer1_outputs(8942));
    layer2_outputs(10239) <= (layer1_outputs(4947)) and not (layer1_outputs(7359));
    outputs(0) <= (layer2_outputs(1662)) xor (layer2_outputs(7339));
    outputs(1) <= (layer2_outputs(3597)) and (layer2_outputs(538));
    outputs(2) <= not(layer2_outputs(2397));
    outputs(3) <= not(layer2_outputs(3560)) or (layer2_outputs(1977));
    outputs(4) <= not(layer2_outputs(9731));
    outputs(5) <= (layer2_outputs(1645)) and not (layer2_outputs(677));
    outputs(6) <= (layer2_outputs(3657)) or (layer2_outputs(8514));
    outputs(7) <= layer2_outputs(7);
    outputs(8) <= layer2_outputs(4740);
    outputs(9) <= not(layer2_outputs(6575));
    outputs(10) <= not((layer2_outputs(7916)) xor (layer2_outputs(5614)));
    outputs(11) <= layer2_outputs(9210);
    outputs(12) <= (layer2_outputs(8947)) and not (layer2_outputs(491));
    outputs(13) <= not((layer2_outputs(6418)) and (layer2_outputs(4148)));
    outputs(14) <= not(layer2_outputs(8715)) or (layer2_outputs(9688));
    outputs(15) <= layer2_outputs(2266);
    outputs(16) <= layer2_outputs(908);
    outputs(17) <= not((layer2_outputs(3614)) xor (layer2_outputs(9929)));
    outputs(18) <= not((layer2_outputs(3885)) and (layer2_outputs(371)));
    outputs(19) <= (layer2_outputs(6099)) xor (layer2_outputs(1733));
    outputs(20) <= not(layer2_outputs(5500));
    outputs(21) <= not((layer2_outputs(7325)) xor (layer2_outputs(10156)));
    outputs(22) <= not(layer2_outputs(7981)) or (layer2_outputs(9281));
    outputs(23) <= not(layer2_outputs(1939));
    outputs(24) <= not(layer2_outputs(988)) or (layer2_outputs(1694));
    outputs(25) <= layer2_outputs(7372);
    outputs(26) <= layer2_outputs(4095);
    outputs(27) <= not((layer2_outputs(5906)) and (layer2_outputs(3129)));
    outputs(28) <= layer2_outputs(1188);
    outputs(29) <= not(layer2_outputs(3338));
    outputs(30) <= not(layer2_outputs(3521)) or (layer2_outputs(6797));
    outputs(31) <= layer2_outputs(9113);
    outputs(32) <= not(layer2_outputs(1705));
    outputs(33) <= not(layer2_outputs(1473));
    outputs(34) <= layer2_outputs(6962);
    outputs(35) <= not(layer2_outputs(6768));
    outputs(36) <= not(layer2_outputs(8430));
    outputs(37) <= layer2_outputs(9677);
    outputs(38) <= layer2_outputs(8610);
    outputs(39) <= (layer2_outputs(6503)) xor (layer2_outputs(1));
    outputs(40) <= not(layer2_outputs(8714)) or (layer2_outputs(7469));
    outputs(41) <= (layer2_outputs(2155)) or (layer2_outputs(4159));
    outputs(42) <= not(layer2_outputs(444));
    outputs(43) <= (layer2_outputs(5184)) or (layer2_outputs(4475));
    outputs(44) <= layer2_outputs(8176);
    outputs(45) <= (layer2_outputs(5296)) and (layer2_outputs(8311));
    outputs(46) <= not(layer2_outputs(1757));
    outputs(47) <= not(layer2_outputs(3965));
    outputs(48) <= not(layer2_outputs(3454));
    outputs(49) <= layer2_outputs(1045);
    outputs(50) <= layer2_outputs(195);
    outputs(51) <= not((layer2_outputs(4438)) or (layer2_outputs(6149)));
    outputs(52) <= not(layer2_outputs(834));
    outputs(53) <= not(layer2_outputs(1613));
    outputs(54) <= not(layer2_outputs(7050));
    outputs(55) <= (layer2_outputs(4533)) xor (layer2_outputs(5103));
    outputs(56) <= layer2_outputs(9840);
    outputs(57) <= not(layer2_outputs(1623));
    outputs(58) <= not(layer2_outputs(7137));
    outputs(59) <= not(layer2_outputs(360));
    outputs(60) <= (layer2_outputs(6263)) and not (layer2_outputs(3457));
    outputs(61) <= not(layer2_outputs(5859));
    outputs(62) <= layer2_outputs(279);
    outputs(63) <= (layer2_outputs(5996)) and not (layer2_outputs(9449));
    outputs(64) <= layer2_outputs(6074);
    outputs(65) <= not(layer2_outputs(2010));
    outputs(66) <= (layer2_outputs(10131)) or (layer2_outputs(4773));
    outputs(67) <= (layer2_outputs(2888)) and not (layer2_outputs(1656));
    outputs(68) <= not(layer2_outputs(6643));
    outputs(69) <= not(layer2_outputs(9524));
    outputs(70) <= not(layer2_outputs(6694));
    outputs(71) <= layer2_outputs(9796);
    outputs(72) <= layer2_outputs(1192);
    outputs(73) <= not(layer2_outputs(8919));
    outputs(74) <= (layer2_outputs(7510)) xor (layer2_outputs(5877));
    outputs(75) <= (layer2_outputs(9413)) and not (layer2_outputs(2433));
    outputs(76) <= not(layer2_outputs(3485));
    outputs(77) <= not((layer2_outputs(3073)) xor (layer2_outputs(10130)));
    outputs(78) <= not(layer2_outputs(6902));
    outputs(79) <= layer2_outputs(7329);
    outputs(80) <= (layer2_outputs(6607)) xor (layer2_outputs(8894));
    outputs(81) <= not(layer2_outputs(2997));
    outputs(82) <= not(layer2_outputs(137));
    outputs(83) <= not(layer2_outputs(7489));
    outputs(84) <= not(layer2_outputs(2662));
    outputs(85) <= not(layer2_outputs(2369));
    outputs(86) <= layer2_outputs(3573);
    outputs(87) <= (layer2_outputs(4693)) xor (layer2_outputs(8368));
    outputs(88) <= not(layer2_outputs(1513));
    outputs(89) <= not((layer2_outputs(7925)) and (layer2_outputs(3526)));
    outputs(90) <= not(layer2_outputs(8903));
    outputs(91) <= layer2_outputs(4943);
    outputs(92) <= not(layer2_outputs(10098));
    outputs(93) <= not(layer2_outputs(9177));
    outputs(94) <= not(layer2_outputs(82));
    outputs(95) <= not(layer2_outputs(2349));
    outputs(96) <= (layer2_outputs(5344)) or (layer2_outputs(4323));
    outputs(97) <= (layer2_outputs(4244)) and not (layer2_outputs(4866));
    outputs(98) <= (layer2_outputs(3363)) xor (layer2_outputs(7514));
    outputs(99) <= (layer2_outputs(1981)) or (layer2_outputs(7068));
    outputs(100) <= not(layer2_outputs(6821));
    outputs(101) <= layer2_outputs(9189);
    outputs(102) <= (layer2_outputs(4953)) xor (layer2_outputs(808));
    outputs(103) <= not(layer2_outputs(7987));
    outputs(104) <= not((layer2_outputs(8700)) and (layer2_outputs(4794)));
    outputs(105) <= (layer2_outputs(2746)) or (layer2_outputs(6737));
    outputs(106) <= not(layer2_outputs(4125));
    outputs(107) <= layer2_outputs(5674);
    outputs(108) <= (layer2_outputs(6561)) and not (layer2_outputs(587));
    outputs(109) <= not(layer2_outputs(1498)) or (layer2_outputs(9664));
    outputs(110) <= not(layer2_outputs(5058)) or (layer2_outputs(1682));
    outputs(111) <= layer2_outputs(870);
    outputs(112) <= layer2_outputs(1669);
    outputs(113) <= not(layer2_outputs(5806));
    outputs(114) <= not((layer2_outputs(1148)) or (layer2_outputs(8131)));
    outputs(115) <= not(layer2_outputs(3543));
    outputs(116) <= not(layer2_outputs(1771));
    outputs(117) <= (layer2_outputs(9635)) and not (layer2_outputs(5992));
    outputs(118) <= not(layer2_outputs(9781));
    outputs(119) <= (layer2_outputs(9027)) and (layer2_outputs(9470));
    outputs(120) <= not(layer2_outputs(6933));
    outputs(121) <= not(layer2_outputs(5720));
    outputs(122) <= not((layer2_outputs(56)) xor (layer2_outputs(269)));
    outputs(123) <= layer2_outputs(787);
    outputs(124) <= (layer2_outputs(4514)) xor (layer2_outputs(7622));
    outputs(125) <= (layer2_outputs(6599)) and (layer2_outputs(7291));
    outputs(126) <= not((layer2_outputs(633)) xor (layer2_outputs(1856)));
    outputs(127) <= not(layer2_outputs(803));
    outputs(128) <= not(layer2_outputs(387));
    outputs(129) <= layer2_outputs(4907);
    outputs(130) <= not((layer2_outputs(3272)) xor (layer2_outputs(2020)));
    outputs(131) <= layer2_outputs(9417);
    outputs(132) <= layer2_outputs(4071);
    outputs(133) <= not(layer2_outputs(8103));
    outputs(134) <= (layer2_outputs(7930)) and (layer2_outputs(5831));
    outputs(135) <= (layer2_outputs(3265)) and not (layer2_outputs(5954));
    outputs(136) <= layer2_outputs(6632);
    outputs(137) <= (layer2_outputs(3917)) and not (layer2_outputs(6140));
    outputs(138) <= not(layer2_outputs(1794)) or (layer2_outputs(8446));
    outputs(139) <= layer2_outputs(4085);
    outputs(140) <= layer2_outputs(2684);
    outputs(141) <= layer2_outputs(7484);
    outputs(142) <= layer2_outputs(7337);
    outputs(143) <= layer2_outputs(8078);
    outputs(144) <= layer2_outputs(9629);
    outputs(145) <= not(layer2_outputs(9577));
    outputs(146) <= layer2_outputs(8260);
    outputs(147) <= not(layer2_outputs(4393));
    outputs(148) <= not(layer2_outputs(9888)) or (layer2_outputs(8589));
    outputs(149) <= not(layer2_outputs(1871));
    outputs(150) <= layer2_outputs(1208);
    outputs(151) <= (layer2_outputs(2999)) xor (layer2_outputs(744));
    outputs(152) <= not(layer2_outputs(314));
    outputs(153) <= layer2_outputs(4359);
    outputs(154) <= not((layer2_outputs(1128)) or (layer2_outputs(5452)));
    outputs(155) <= layer2_outputs(8833);
    outputs(156) <= layer2_outputs(1033);
    outputs(157) <= layer2_outputs(3666);
    outputs(158) <= layer2_outputs(3290);
    outputs(159) <= not((layer2_outputs(7841)) xor (layer2_outputs(9014)));
    outputs(160) <= not(layer2_outputs(2558));
    outputs(161) <= not(layer2_outputs(5770));
    outputs(162) <= layer2_outputs(8101);
    outputs(163) <= (layer2_outputs(9662)) and not (layer2_outputs(7050));
    outputs(164) <= not(layer2_outputs(9049));
    outputs(165) <= layer2_outputs(1499);
    outputs(166) <= (layer2_outputs(6709)) xor (layer2_outputs(4701));
    outputs(167) <= layer2_outputs(5413);
    outputs(168) <= (layer2_outputs(1416)) and (layer2_outputs(6885));
    outputs(169) <= not(layer2_outputs(8181));
    outputs(170) <= not(layer2_outputs(597));
    outputs(171) <= (layer2_outputs(5626)) and not (layer2_outputs(8056));
    outputs(172) <= not(layer2_outputs(3233));
    outputs(173) <= layer2_outputs(4804);
    outputs(174) <= (layer2_outputs(9898)) xor (layer2_outputs(5980));
    outputs(175) <= not(layer2_outputs(2984));
    outputs(176) <= layer2_outputs(6454);
    outputs(177) <= not((layer2_outputs(4165)) xor (layer2_outputs(4819)));
    outputs(178) <= (layer2_outputs(2088)) xor (layer2_outputs(7978));
    outputs(179) <= (layer2_outputs(9957)) xor (layer2_outputs(6638));
    outputs(180) <= not(layer2_outputs(2573));
    outputs(181) <= (layer2_outputs(924)) and not (layer2_outputs(4889));
    outputs(182) <= not(layer2_outputs(276));
    outputs(183) <= not(layer2_outputs(6643));
    outputs(184) <= not(layer2_outputs(6941));
    outputs(185) <= layer2_outputs(3306);
    outputs(186) <= layer2_outputs(8984);
    outputs(187) <= (layer2_outputs(9557)) and (layer2_outputs(10009));
    outputs(188) <= not(layer2_outputs(440));
    outputs(189) <= layer2_outputs(2975);
    outputs(190) <= layer2_outputs(9832);
    outputs(191) <= layer2_outputs(9563);
    outputs(192) <= layer2_outputs(2641);
    outputs(193) <= not((layer2_outputs(6881)) and (layer2_outputs(6723)));
    outputs(194) <= layer2_outputs(6997);
    outputs(195) <= not(layer2_outputs(5723));
    outputs(196) <= (layer2_outputs(5838)) xor (layer2_outputs(9141));
    outputs(197) <= not((layer2_outputs(6667)) and (layer2_outputs(9718)));
    outputs(198) <= not(layer2_outputs(9873));
    outputs(199) <= not((layer2_outputs(2234)) and (layer2_outputs(8363)));
    outputs(200) <= layer2_outputs(4289);
    outputs(201) <= not(layer2_outputs(2973));
    outputs(202) <= layer2_outputs(1834);
    outputs(203) <= layer2_outputs(6700);
    outputs(204) <= not(layer2_outputs(1060));
    outputs(205) <= (layer2_outputs(912)) and not (layer2_outputs(9671));
    outputs(206) <= (layer2_outputs(8566)) xor (layer2_outputs(5547));
    outputs(207) <= (layer2_outputs(4053)) and not (layer2_outputs(3608));
    outputs(208) <= layer2_outputs(6100);
    outputs(209) <= layer2_outputs(6028);
    outputs(210) <= layer2_outputs(1467);
    outputs(211) <= layer2_outputs(5807);
    outputs(212) <= (layer2_outputs(6676)) and not (layer2_outputs(3512));
    outputs(213) <= not(layer2_outputs(3547));
    outputs(214) <= not(layer2_outputs(1870));
    outputs(215) <= not(layer2_outputs(8358));
    outputs(216) <= layer2_outputs(5096);
    outputs(217) <= layer2_outputs(1088);
    outputs(218) <= layer2_outputs(6817);
    outputs(219) <= layer2_outputs(8819);
    outputs(220) <= (layer2_outputs(2298)) and not (layer2_outputs(1836));
    outputs(221) <= layer2_outputs(589);
    outputs(222) <= not(layer2_outputs(6442)) or (layer2_outputs(1157));
    outputs(223) <= layer2_outputs(415);
    outputs(224) <= not(layer2_outputs(9642));
    outputs(225) <= (layer2_outputs(637)) xor (layer2_outputs(4200));
    outputs(226) <= not(layer2_outputs(7516));
    outputs(227) <= not(layer2_outputs(6277));
    outputs(228) <= not(layer2_outputs(1949));
    outputs(229) <= not(layer2_outputs(4226));
    outputs(230) <= not(layer2_outputs(1623));
    outputs(231) <= not(layer2_outputs(5679));
    outputs(232) <= (layer2_outputs(9735)) and (layer2_outputs(7499));
    outputs(233) <= layer2_outputs(977);
    outputs(234) <= layer2_outputs(3641);
    outputs(235) <= not(layer2_outputs(5991)) or (layer2_outputs(421));
    outputs(236) <= not(layer2_outputs(8234));
    outputs(237) <= layer2_outputs(535);
    outputs(238) <= (layer2_outputs(7244)) and (layer2_outputs(5107));
    outputs(239) <= not(layer2_outputs(7179));
    outputs(240) <= (layer2_outputs(2219)) and not (layer2_outputs(3871));
    outputs(241) <= not((layer2_outputs(8626)) and (layer2_outputs(6655)));
    outputs(242) <= not(layer2_outputs(2454));
    outputs(243) <= layer2_outputs(7295);
    outputs(244) <= not((layer2_outputs(9295)) xor (layer2_outputs(9517)));
    outputs(245) <= layer2_outputs(5757);
    outputs(246) <= not(layer2_outputs(5476));
    outputs(247) <= layer2_outputs(7511);
    outputs(248) <= (layer2_outputs(2326)) xor (layer2_outputs(4776));
    outputs(249) <= (layer2_outputs(6038)) and not (layer2_outputs(7932));
    outputs(250) <= not(layer2_outputs(762));
    outputs(251) <= layer2_outputs(9933);
    outputs(252) <= layer2_outputs(1335);
    outputs(253) <= layer2_outputs(8161);
    outputs(254) <= not((layer2_outputs(9046)) or (layer2_outputs(3474)));
    outputs(255) <= layer2_outputs(1348);
    outputs(256) <= (layer2_outputs(5192)) xor (layer2_outputs(8877));
    outputs(257) <= layer2_outputs(3362);
    outputs(258) <= layer2_outputs(4869);
    outputs(259) <= not((layer2_outputs(7496)) xor (layer2_outputs(2154)));
    outputs(260) <= not(layer2_outputs(9437));
    outputs(261) <= not(layer2_outputs(1097));
    outputs(262) <= not(layer2_outputs(2064));
    outputs(263) <= not(layer2_outputs(2363));
    outputs(264) <= not(layer2_outputs(2037));
    outputs(265) <= layer2_outputs(4846);
    outputs(266) <= layer2_outputs(9397);
    outputs(267) <= (layer2_outputs(8282)) and not (layer2_outputs(2401));
    outputs(268) <= (layer2_outputs(8939)) xor (layer2_outputs(1662));
    outputs(269) <= layer2_outputs(5331);
    outputs(270) <= not((layer2_outputs(3729)) xor (layer2_outputs(880)));
    outputs(271) <= not(layer2_outputs(9944));
    outputs(272) <= not(layer2_outputs(1031));
    outputs(273) <= layer2_outputs(871);
    outputs(274) <= (layer2_outputs(7845)) and not (layer2_outputs(8967));
    outputs(275) <= not((layer2_outputs(8691)) xor (layer2_outputs(6882)));
    outputs(276) <= layer2_outputs(791);
    outputs(277) <= not(layer2_outputs(8701));
    outputs(278) <= not(layer2_outputs(4395));
    outputs(279) <= (layer2_outputs(7075)) xor (layer2_outputs(2494));
    outputs(280) <= (layer2_outputs(8876)) xor (layer2_outputs(6594));
    outputs(281) <= (layer2_outputs(9055)) xor (layer2_outputs(6820));
    outputs(282) <= layer2_outputs(2872);
    outputs(283) <= not(layer2_outputs(9070));
    outputs(284) <= not(layer2_outputs(9994));
    outputs(285) <= not((layer2_outputs(1299)) and (layer2_outputs(6584)));
    outputs(286) <= layer2_outputs(4745);
    outputs(287) <= not(layer2_outputs(1871));
    outputs(288) <= (layer2_outputs(20)) and not (layer2_outputs(234));
    outputs(289) <= not(layer2_outputs(3051));
    outputs(290) <= not(layer2_outputs(4302));
    outputs(291) <= layer2_outputs(5502);
    outputs(292) <= not(layer2_outputs(7251));
    outputs(293) <= layer2_outputs(6621);
    outputs(294) <= (layer2_outputs(9911)) xor (layer2_outputs(4731));
    outputs(295) <= not(layer2_outputs(2743));
    outputs(296) <= not((layer2_outputs(945)) and (layer2_outputs(1342)));
    outputs(297) <= not(layer2_outputs(10124));
    outputs(298) <= not((layer2_outputs(6217)) xor (layer2_outputs(9618)));
    outputs(299) <= not((layer2_outputs(7324)) and (layer2_outputs(6920)));
    outputs(300) <= layer2_outputs(589);
    outputs(301) <= not(layer2_outputs(1096));
    outputs(302) <= (layer2_outputs(5129)) and (layer2_outputs(7903));
    outputs(303) <= not((layer2_outputs(8570)) xor (layer2_outputs(6983)));
    outputs(304) <= (layer2_outputs(668)) and not (layer2_outputs(8411));
    outputs(305) <= not(layer2_outputs(1061));
    outputs(306) <= layer2_outputs(4042);
    outputs(307) <= layer2_outputs(6806);
    outputs(308) <= layer2_outputs(7334);
    outputs(309) <= (layer2_outputs(6714)) xor (layer2_outputs(8775));
    outputs(310) <= not(layer2_outputs(7790));
    outputs(311) <= not(layer2_outputs(9680));
    outputs(312) <= not(layer2_outputs(4339));
    outputs(313) <= not(layer2_outputs(8408));
    outputs(314) <= layer2_outputs(1094);
    outputs(315) <= layer2_outputs(9462);
    outputs(316) <= layer2_outputs(1384);
    outputs(317) <= (layer2_outputs(5325)) and (layer2_outputs(580));
    outputs(318) <= not(layer2_outputs(7839));
    outputs(319) <= layer2_outputs(7611);
    outputs(320) <= not(layer2_outputs(5148));
    outputs(321) <= not(layer2_outputs(1292));
    outputs(322) <= not(layer2_outputs(19));
    outputs(323) <= layer2_outputs(9563);
    outputs(324) <= layer2_outputs(7719);
    outputs(325) <= layer2_outputs(5827);
    outputs(326) <= (layer2_outputs(7819)) and not (layer2_outputs(2838));
    outputs(327) <= not(layer2_outputs(7240));
    outputs(328) <= not((layer2_outputs(5991)) and (layer2_outputs(6145)));
    outputs(329) <= not(layer2_outputs(8861));
    outputs(330) <= (layer2_outputs(5517)) xor (layer2_outputs(2212));
    outputs(331) <= layer2_outputs(7433);
    outputs(332) <= (layer2_outputs(2545)) and not (layer2_outputs(9118));
    outputs(333) <= not(layer2_outputs(2356));
    outputs(334) <= not((layer2_outputs(4971)) and (layer2_outputs(2115)));
    outputs(335) <= (layer2_outputs(3859)) and not (layer2_outputs(2183));
    outputs(336) <= not(layer2_outputs(275)) or (layer2_outputs(8554));
    outputs(337) <= not((layer2_outputs(4625)) or (layer2_outputs(8752)));
    outputs(338) <= layer2_outputs(7959);
    outputs(339) <= not(layer2_outputs(9900));
    outputs(340) <= layer2_outputs(5423);
    outputs(341) <= layer2_outputs(7272);
    outputs(342) <= layer2_outputs(4308);
    outputs(343) <= not((layer2_outputs(489)) or (layer2_outputs(1783)));
    outputs(344) <= not((layer2_outputs(1000)) xor (layer2_outputs(2446)));
    outputs(345) <= layer2_outputs(2934);
    outputs(346) <= (layer2_outputs(4734)) and not (layer2_outputs(6857));
    outputs(347) <= (layer2_outputs(1834)) and not (layer2_outputs(3054));
    outputs(348) <= not((layer2_outputs(2641)) xor (layer2_outputs(8793)));
    outputs(349) <= not(layer2_outputs(5780));
    outputs(350) <= layer2_outputs(941);
    outputs(351) <= not((layer2_outputs(6415)) xor (layer2_outputs(7379)));
    outputs(352) <= not(layer2_outputs(2407));
    outputs(353) <= layer2_outputs(5347);
    outputs(354) <= not(layer2_outputs(8264)) or (layer2_outputs(576));
    outputs(355) <= not(layer2_outputs(1540));
    outputs(356) <= layer2_outputs(7710);
    outputs(357) <= layer2_outputs(7344);
    outputs(358) <= not(layer2_outputs(2054));
    outputs(359) <= layer2_outputs(5096);
    outputs(360) <= not(layer2_outputs(8580));
    outputs(361) <= layer2_outputs(7188);
    outputs(362) <= not((layer2_outputs(4135)) or (layer2_outputs(5465)));
    outputs(363) <= not((layer2_outputs(8412)) or (layer2_outputs(8914)));
    outputs(364) <= not(layer2_outputs(7095));
    outputs(365) <= layer2_outputs(8190);
    outputs(366) <= (layer2_outputs(8589)) and not (layer2_outputs(5327));
    outputs(367) <= not((layer2_outputs(2518)) or (layer2_outputs(5936)));
    outputs(368) <= (layer2_outputs(4857)) and (layer2_outputs(2814));
    outputs(369) <= layer2_outputs(3290);
    outputs(370) <= layer2_outputs(6532);
    outputs(371) <= layer2_outputs(7933);
    outputs(372) <= (layer2_outputs(9001)) xor (layer2_outputs(3330));
    outputs(373) <= layer2_outputs(4103);
    outputs(374) <= not(layer2_outputs(5452));
    outputs(375) <= not(layer2_outputs(5707)) or (layer2_outputs(2511));
    outputs(376) <= not(layer2_outputs(4268));
    outputs(377) <= layer2_outputs(9796);
    outputs(378) <= layer2_outputs(2294);
    outputs(379) <= not((layer2_outputs(2524)) xor (layer2_outputs(3395)));
    outputs(380) <= not(layer2_outputs(1167));
    outputs(381) <= not((layer2_outputs(4902)) xor (layer2_outputs(1547)));
    outputs(382) <= not(layer2_outputs(6370));
    outputs(383) <= layer2_outputs(9426);
    outputs(384) <= not(layer2_outputs(443));
    outputs(385) <= layer2_outputs(8898);
    outputs(386) <= not(layer2_outputs(10125));
    outputs(387) <= not((layer2_outputs(10103)) or (layer2_outputs(2910)));
    outputs(388) <= layer2_outputs(3298);
    outputs(389) <= not(layer2_outputs(7491));
    outputs(390) <= not(layer2_outputs(8848));
    outputs(391) <= (layer2_outputs(6960)) and (layer2_outputs(9305));
    outputs(392) <= not(layer2_outputs(3870));
    outputs(393) <= not((layer2_outputs(3846)) xor (layer2_outputs(5791)));
    outputs(394) <= (layer2_outputs(3564)) or (layer2_outputs(1121));
    outputs(395) <= not(layer2_outputs(8553)) or (layer2_outputs(5235));
    outputs(396) <= not((layer2_outputs(7408)) xor (layer2_outputs(3173)));
    outputs(397) <= layer2_outputs(1779);
    outputs(398) <= not(layer2_outputs(9086)) or (layer2_outputs(8555));
    outputs(399) <= (layer2_outputs(7390)) xor (layer2_outputs(3514));
    outputs(400) <= not(layer2_outputs(45));
    outputs(401) <= (layer2_outputs(9714)) and not (layer2_outputs(5450));
    outputs(402) <= not(layer2_outputs(1641));
    outputs(403) <= (layer2_outputs(7188)) and not (layer2_outputs(2397));
    outputs(404) <= not(layer2_outputs(788));
    outputs(405) <= not(layer2_outputs(3373));
    outputs(406) <= (layer2_outputs(8573)) and not (layer2_outputs(2801));
    outputs(407) <= (layer2_outputs(4034)) xor (layer2_outputs(2999));
    outputs(408) <= layer2_outputs(3114);
    outputs(409) <= (layer2_outputs(6249)) or (layer2_outputs(3068));
    outputs(410) <= not((layer2_outputs(494)) xor (layer2_outputs(524)));
    outputs(411) <= not(layer2_outputs(7695));
    outputs(412) <= layer2_outputs(6869);
    outputs(413) <= not((layer2_outputs(5036)) or (layer2_outputs(3570)));
    outputs(414) <= (layer2_outputs(1669)) and not (layer2_outputs(7013));
    outputs(415) <= (layer2_outputs(7856)) or (layer2_outputs(511));
    outputs(416) <= not(layer2_outputs(8415));
    outputs(417) <= not(layer2_outputs(2243));
    outputs(418) <= not(layer2_outputs(4489));
    outputs(419) <= not(layer2_outputs(7193));
    outputs(420) <= (layer2_outputs(6228)) or (layer2_outputs(7411));
    outputs(421) <= (layer2_outputs(7934)) xor (layer2_outputs(8309));
    outputs(422) <= not(layer2_outputs(4301));
    outputs(423) <= not((layer2_outputs(4438)) xor (layer2_outputs(8851)));
    outputs(424) <= not((layer2_outputs(2549)) xor (layer2_outputs(7323)));
    outputs(425) <= not(layer2_outputs(7574));
    outputs(426) <= (layer2_outputs(1464)) xor (layer2_outputs(8813));
    outputs(427) <= not((layer2_outputs(5305)) xor (layer2_outputs(3597)));
    outputs(428) <= not(layer2_outputs(7840));
    outputs(429) <= layer2_outputs(270);
    outputs(430) <= layer2_outputs(2758);
    outputs(431) <= layer2_outputs(6732);
    outputs(432) <= not(layer2_outputs(3344));
    outputs(433) <= not(layer2_outputs(5796)) or (layer2_outputs(4233));
    outputs(434) <= not(layer2_outputs(7449));
    outputs(435) <= layer2_outputs(3565);
    outputs(436) <= layer2_outputs(3896);
    outputs(437) <= (layer2_outputs(5080)) and (layer2_outputs(5793));
    outputs(438) <= (layer2_outputs(8043)) and (layer2_outputs(1728));
    outputs(439) <= not(layer2_outputs(9932));
    outputs(440) <= not(layer2_outputs(309));
    outputs(441) <= not((layer2_outputs(6387)) and (layer2_outputs(4979)));
    outputs(442) <= layer2_outputs(372);
    outputs(443) <= layer2_outputs(2661);
    outputs(444) <= not(layer2_outputs(1890));
    outputs(445) <= not(layer2_outputs(3060));
    outputs(446) <= not(layer2_outputs(5897));
    outputs(447) <= layer2_outputs(823);
    outputs(448) <= layer2_outputs(176);
    outputs(449) <= layer2_outputs(3528);
    outputs(450) <= not(layer2_outputs(1361));
    outputs(451) <= (layer2_outputs(8707)) and not (layer2_outputs(4684));
    outputs(452) <= not(layer2_outputs(8456));
    outputs(453) <= not((layer2_outputs(6472)) xor (layer2_outputs(3343)));
    outputs(454) <= not((layer2_outputs(7451)) and (layer2_outputs(7918)));
    outputs(455) <= layer2_outputs(9249);
    outputs(456) <= not(layer2_outputs(5177));
    outputs(457) <= not(layer2_outputs(6786));
    outputs(458) <= not(layer2_outputs(3646));
    outputs(459) <= (layer2_outputs(1707)) and (layer2_outputs(4451));
    outputs(460) <= layer2_outputs(5890);
    outputs(461) <= layer2_outputs(8322);
    outputs(462) <= (layer2_outputs(322)) and not (layer2_outputs(8837));
    outputs(463) <= not(layer2_outputs(9999));
    outputs(464) <= not((layer2_outputs(5845)) xor (layer2_outputs(7335)));
    outputs(465) <= not(layer2_outputs(5672));
    outputs(466) <= not(layer2_outputs(7529));
    outputs(467) <= not(layer2_outputs(8256));
    outputs(468) <= layer2_outputs(3664);
    outputs(469) <= not(layer2_outputs(4348));
    outputs(470) <= layer2_outputs(8732);
    outputs(471) <= (layer2_outputs(96)) or (layer2_outputs(4520));
    outputs(472) <= not((layer2_outputs(1136)) and (layer2_outputs(1851)));
    outputs(473) <= not(layer2_outputs(5024));
    outputs(474) <= not(layer2_outputs(9059));
    outputs(475) <= layer2_outputs(9367);
    outputs(476) <= not(layer2_outputs(6410));
    outputs(477) <= (layer2_outputs(3231)) and not (layer2_outputs(2794));
    outputs(478) <= layer2_outputs(2325);
    outputs(479) <= not(layer2_outputs(2703));
    outputs(480) <= layer2_outputs(252);
    outputs(481) <= not((layer2_outputs(3431)) xor (layer2_outputs(1130)));
    outputs(482) <= layer2_outputs(8479);
    outputs(483) <= not(layer2_outputs(615));
    outputs(484) <= not(layer2_outputs(5421));
    outputs(485) <= (layer2_outputs(9061)) xor (layer2_outputs(6659));
    outputs(486) <= not(layer2_outputs(1116));
    outputs(487) <= layer2_outputs(33);
    outputs(488) <= (layer2_outputs(1731)) and not (layer2_outputs(3142));
    outputs(489) <= not(layer2_outputs(9968));
    outputs(490) <= not(layer2_outputs(4163));
    outputs(491) <= not((layer2_outputs(1334)) and (layer2_outputs(7614)));
    outputs(492) <= layer2_outputs(1555);
    outputs(493) <= not(layer2_outputs(2283));
    outputs(494) <= (layer2_outputs(5700)) or (layer2_outputs(10018));
    outputs(495) <= not(layer2_outputs(7332));
    outputs(496) <= not(layer2_outputs(7834));
    outputs(497) <= layer2_outputs(2934);
    outputs(498) <= not(layer2_outputs(6681)) or (layer2_outputs(9815));
    outputs(499) <= not(layer2_outputs(7393)) or (layer2_outputs(306));
    outputs(500) <= not(layer2_outputs(10124));
    outputs(501) <= not(layer2_outputs(5472)) or (layer2_outputs(2824));
    outputs(502) <= layer2_outputs(1260);
    outputs(503) <= layer2_outputs(3120);
    outputs(504) <= (layer2_outputs(4492)) and not (layer2_outputs(23));
    outputs(505) <= layer2_outputs(6467);
    outputs(506) <= not(layer2_outputs(10106));
    outputs(507) <= not(layer2_outputs(2717)) or (layer2_outputs(143));
    outputs(508) <= (layer2_outputs(9137)) and not (layer2_outputs(8777));
    outputs(509) <= not(layer2_outputs(9078));
    outputs(510) <= not(layer2_outputs(199));
    outputs(511) <= (layer2_outputs(1387)) xor (layer2_outputs(8913));
    outputs(512) <= not(layer2_outputs(9777));
    outputs(513) <= not(layer2_outputs(3172));
    outputs(514) <= layer2_outputs(4183);
    outputs(515) <= not(layer2_outputs(1847));
    outputs(516) <= (layer2_outputs(7121)) or (layer2_outputs(9706));
    outputs(517) <= layer2_outputs(9444);
    outputs(518) <= layer2_outputs(4973);
    outputs(519) <= not(layer2_outputs(6333));
    outputs(520) <= layer2_outputs(7368);
    outputs(521) <= layer2_outputs(4026);
    outputs(522) <= not(layer2_outputs(5190));
    outputs(523) <= layer2_outputs(60);
    outputs(524) <= not(layer2_outputs(4138));
    outputs(525) <= layer2_outputs(7736);
    outputs(526) <= layer2_outputs(870);
    outputs(527) <= (layer2_outputs(1413)) xor (layer2_outputs(6481));
    outputs(528) <= (layer2_outputs(2685)) and (layer2_outputs(363));
    outputs(529) <= not(layer2_outputs(4406));
    outputs(530) <= not((layer2_outputs(7513)) xor (layer2_outputs(3237)));
    outputs(531) <= not((layer2_outputs(974)) xor (layer2_outputs(2806)));
    outputs(532) <= (layer2_outputs(6516)) xor (layer2_outputs(7687));
    outputs(533) <= not((layer2_outputs(8196)) xor (layer2_outputs(6471)));
    outputs(534) <= not(layer2_outputs(8612));
    outputs(535) <= not(layer2_outputs(1089));
    outputs(536) <= layer2_outputs(9543);
    outputs(537) <= not(layer2_outputs(425)) or (layer2_outputs(7301));
    outputs(538) <= not((layer2_outputs(9862)) or (layer2_outputs(362)));
    outputs(539) <= not(layer2_outputs(2731));
    outputs(540) <= not((layer2_outputs(3273)) xor (layer2_outputs(4907)));
    outputs(541) <= not(layer2_outputs(5836));
    outputs(542) <= not(layer2_outputs(3085));
    outputs(543) <= not((layer2_outputs(8659)) or (layer2_outputs(3570)));
    outputs(544) <= layer2_outputs(6132);
    outputs(545) <= not(layer2_outputs(1533));
    outputs(546) <= not(layer2_outputs(6405));
    outputs(547) <= layer2_outputs(9378);
    outputs(548) <= (layer2_outputs(8261)) and not (layer2_outputs(2112));
    outputs(549) <= not(layer2_outputs(2080));
    outputs(550) <= not((layer2_outputs(5104)) xor (layer2_outputs(4937)));
    outputs(551) <= not((layer2_outputs(965)) xor (layer2_outputs(5114)));
    outputs(552) <= (layer2_outputs(6892)) or (layer2_outputs(5039));
    outputs(553) <= not(layer2_outputs(9483));
    outputs(554) <= not(layer2_outputs(4509));
    outputs(555) <= not(layer2_outputs(10075));
    outputs(556) <= not(layer2_outputs(8546));
    outputs(557) <= not(layer2_outputs(4741));
    outputs(558) <= (layer2_outputs(5394)) or (layer2_outputs(8336));
    outputs(559) <= layer2_outputs(7066);
    outputs(560) <= not(layer2_outputs(5511));
    outputs(561) <= not(layer2_outputs(7506));
    outputs(562) <= layer2_outputs(9631);
    outputs(563) <= not(layer2_outputs(5828));
    outputs(564) <= not(layer2_outputs(1556)) or (layer2_outputs(9342));
    outputs(565) <= not(layer2_outputs(6830));
    outputs(566) <= not((layer2_outputs(2770)) xor (layer2_outputs(1440)));
    outputs(567) <= (layer2_outputs(9697)) xor (layer2_outputs(2866));
    outputs(568) <= layer2_outputs(396);
    outputs(569) <= (layer2_outputs(2570)) xor (layer2_outputs(6671));
    outputs(570) <= not(layer2_outputs(9726));
    outputs(571) <= (layer2_outputs(1081)) and (layer2_outputs(10183));
    outputs(572) <= not(layer2_outputs(7919));
    outputs(573) <= not((layer2_outputs(4850)) or (layer2_outputs(2725)));
    outputs(574) <= (layer2_outputs(2505)) and not (layer2_outputs(7969));
    outputs(575) <= layer2_outputs(7429);
    outputs(576) <= layer2_outputs(169);
    outputs(577) <= (layer2_outputs(5230)) xor (layer2_outputs(4613));
    outputs(578) <= not(layer2_outputs(9932));
    outputs(579) <= not(layer2_outputs(7349));
    outputs(580) <= not((layer2_outputs(2802)) xor (layer2_outputs(8974)));
    outputs(581) <= not(layer2_outputs(1619));
    outputs(582) <= not(layer2_outputs(658));
    outputs(583) <= not(layer2_outputs(254));
    outputs(584) <= not(layer2_outputs(1754));
    outputs(585) <= not(layer2_outputs(9608));
    outputs(586) <= layer2_outputs(2257);
    outputs(587) <= layer2_outputs(5328);
    outputs(588) <= (layer2_outputs(9896)) or (layer2_outputs(8344));
    outputs(589) <= not((layer2_outputs(7431)) and (layer2_outputs(2479)));
    outputs(590) <= layer2_outputs(3508);
    outputs(591) <= not(layer2_outputs(1352));
    outputs(592) <= layer2_outputs(270);
    outputs(593) <= (layer2_outputs(2800)) xor (layer2_outputs(6580));
    outputs(594) <= layer2_outputs(1499);
    outputs(595) <= not(layer2_outputs(2389));
    outputs(596) <= layer2_outputs(7804);
    outputs(597) <= (layer2_outputs(7929)) and not (layer2_outputs(9882));
    outputs(598) <= (layer2_outputs(10235)) xor (layer2_outputs(8493));
    outputs(599) <= not((layer2_outputs(1900)) xor (layer2_outputs(8716)));
    outputs(600) <= (layer2_outputs(3675)) xor (layer2_outputs(3081));
    outputs(601) <= not(layer2_outputs(2163));
    outputs(602) <= (layer2_outputs(2520)) xor (layer2_outputs(4579));
    outputs(603) <= not(layer2_outputs(4648)) or (layer2_outputs(3257));
    outputs(604) <= layer2_outputs(6864);
    outputs(605) <= not(layer2_outputs(2223));
    outputs(606) <= not((layer2_outputs(5791)) xor (layer2_outputs(7901)));
    outputs(607) <= layer2_outputs(6788);
    outputs(608) <= layer2_outputs(4029);
    outputs(609) <= (layer2_outputs(2198)) or (layer2_outputs(2910));
    outputs(610) <= layer2_outputs(6095);
    outputs(611) <= (layer2_outputs(3329)) and not (layer2_outputs(9608));
    outputs(612) <= (layer2_outputs(9374)) and not (layer2_outputs(4591));
    outputs(613) <= not(layer2_outputs(1100));
    outputs(614) <= not(layer2_outputs(3867));
    outputs(615) <= layer2_outputs(7675);
    outputs(616) <= layer2_outputs(3886);
    outputs(617) <= (layer2_outputs(2871)) and not (layer2_outputs(2526));
    outputs(618) <= not(layer2_outputs(3560));
    outputs(619) <= not(layer2_outputs(2115)) or (layer2_outputs(3204));
    outputs(620) <= (layer2_outputs(572)) xor (layer2_outputs(6191));
    outputs(621) <= not(layer2_outputs(6319));
    outputs(622) <= layer2_outputs(5582);
    outputs(623) <= (layer2_outputs(7654)) xor (layer2_outputs(8009));
    outputs(624) <= not(layer2_outputs(7590));
    outputs(625) <= not((layer2_outputs(256)) xor (layer2_outputs(4814)));
    outputs(626) <= layer2_outputs(3154);
    outputs(627) <= not(layer2_outputs(2281));
    outputs(628) <= not(layer2_outputs(7421));
    outputs(629) <= layer2_outputs(6894);
    outputs(630) <= (layer2_outputs(4816)) and not (layer2_outputs(7357));
    outputs(631) <= not(layer2_outputs(353));
    outputs(632) <= (layer2_outputs(4714)) and (layer2_outputs(5399));
    outputs(633) <= not(layer2_outputs(125));
    outputs(634) <= not(layer2_outputs(7975));
    outputs(635) <= layer2_outputs(2101);
    outputs(636) <= not(layer2_outputs(2966));
    outputs(637) <= not((layer2_outputs(7183)) or (layer2_outputs(8734)));
    outputs(638) <= not(layer2_outputs(2183));
    outputs(639) <= not(layer2_outputs(5046));
    outputs(640) <= not(layer2_outputs(7638));
    outputs(641) <= not(layer2_outputs(7516));
    outputs(642) <= layer2_outputs(5922);
    outputs(643) <= not((layer2_outputs(10006)) or (layer2_outputs(2370)));
    outputs(644) <= not(layer2_outputs(3831));
    outputs(645) <= not(layer2_outputs(1757));
    outputs(646) <= layer2_outputs(2099);
    outputs(647) <= (layer2_outputs(9479)) and (layer2_outputs(2368));
    outputs(648) <= not((layer2_outputs(6886)) and (layer2_outputs(1025)));
    outputs(649) <= not(layer2_outputs(2593));
    outputs(650) <= not(layer2_outputs(2998)) or (layer2_outputs(2927));
    outputs(651) <= not((layer2_outputs(4453)) and (layer2_outputs(3083)));
    outputs(652) <= layer2_outputs(9341);
    outputs(653) <= layer2_outputs(166);
    outputs(654) <= layer2_outputs(6650);
    outputs(655) <= not(layer2_outputs(5908));
    outputs(656) <= not((layer2_outputs(8476)) xor (layer2_outputs(2472)));
    outputs(657) <= layer2_outputs(1512);
    outputs(658) <= layer2_outputs(297);
    outputs(659) <= not(layer2_outputs(3776));
    outputs(660) <= layer2_outputs(6289);
    outputs(661) <= not(layer2_outputs(5848));
    outputs(662) <= layer2_outputs(7832);
    outputs(663) <= not(layer2_outputs(483)) or (layer2_outputs(8908));
    outputs(664) <= not(layer2_outputs(6487));
    outputs(665) <= layer2_outputs(2568);
    outputs(666) <= not(layer2_outputs(2856));
    outputs(667) <= not((layer2_outputs(5717)) and (layer2_outputs(3933)));
    outputs(668) <= not(layer2_outputs(1702));
    outputs(669) <= layer2_outputs(8556);
    outputs(670) <= not(layer2_outputs(3226));
    outputs(671) <= not(layer2_outputs(379)) or (layer2_outputs(9130));
    outputs(672) <= not((layer2_outputs(4159)) xor (layer2_outputs(9590)));
    outputs(673) <= not(layer2_outputs(6871));
    outputs(674) <= not(layer2_outputs(8777));
    outputs(675) <= not(layer2_outputs(700));
    outputs(676) <= not(layer2_outputs(8278));
    outputs(677) <= (layer2_outputs(3293)) and not (layer2_outputs(7283));
    outputs(678) <= not(layer2_outputs(3188));
    outputs(679) <= layer2_outputs(1569);
    outputs(680) <= layer2_outputs(9315);
    outputs(681) <= layer2_outputs(9009);
    outputs(682) <= not(layer2_outputs(2660));
    outputs(683) <= (layer2_outputs(8137)) xor (layer2_outputs(4404));
    outputs(684) <= not(layer2_outputs(5803));
    outputs(685) <= (layer2_outputs(2478)) or (layer2_outputs(8007));
    outputs(686) <= (layer2_outputs(1320)) xor (layer2_outputs(5084));
    outputs(687) <= not((layer2_outputs(8617)) and (layer2_outputs(9552)));
    outputs(688) <= layer2_outputs(6788);
    outputs(689) <= layer2_outputs(10039);
    outputs(690) <= (layer2_outputs(8214)) or (layer2_outputs(717));
    outputs(691) <= layer2_outputs(8321);
    outputs(692) <= not((layer2_outputs(3676)) and (layer2_outputs(8445)));
    outputs(693) <= not((layer2_outputs(471)) or (layer2_outputs(7723)));
    outputs(694) <= not(layer2_outputs(328));
    outputs(695) <= not((layer2_outputs(4709)) xor (layer2_outputs(8469)));
    outputs(696) <= layer2_outputs(13);
    outputs(697) <= layer2_outputs(849);
    outputs(698) <= not(layer2_outputs(5549));
    outputs(699) <= not((layer2_outputs(2517)) xor (layer2_outputs(2954)));
    outputs(700) <= not(layer2_outputs(5306));
    outputs(701) <= (layer2_outputs(311)) and (layer2_outputs(9967));
    outputs(702) <= not(layer2_outputs(1139)) or (layer2_outputs(4377));
    outputs(703) <= not(layer2_outputs(5490));
    outputs(704) <= not(layer2_outputs(8711));
    outputs(705) <= not(layer2_outputs(4079));
    outputs(706) <= not((layer2_outputs(9556)) xor (layer2_outputs(1617)));
    outputs(707) <= layer2_outputs(1241);
    outputs(708) <= layer2_outputs(6734);
    outputs(709) <= layer2_outputs(6206);
    outputs(710) <= not(layer2_outputs(8747));
    outputs(711) <= layer2_outputs(30);
    outputs(712) <= not(layer2_outputs(5220));
    outputs(713) <= layer2_outputs(748);
    outputs(714) <= not((layer2_outputs(2776)) xor (layer2_outputs(2968)));
    outputs(715) <= (layer2_outputs(3036)) and not (layer2_outputs(7689));
    outputs(716) <= not((layer2_outputs(6639)) xor (layer2_outputs(7749)));
    outputs(717) <= not(layer2_outputs(8135));
    outputs(718) <= layer2_outputs(3503);
    outputs(719) <= not(layer2_outputs(8115));
    outputs(720) <= not(layer2_outputs(9399));
    outputs(721) <= '0';
    outputs(722) <= not(layer2_outputs(720));
    outputs(723) <= (layer2_outputs(4652)) xor (layer2_outputs(8187));
    outputs(724) <= layer2_outputs(5966);
    outputs(725) <= layer2_outputs(3432);
    outputs(726) <= layer2_outputs(7493);
    outputs(727) <= not((layer2_outputs(7592)) and (layer2_outputs(6922)));
    outputs(728) <= (layer2_outputs(5946)) and not (layer2_outputs(1572));
    outputs(729) <= layer2_outputs(222);
    outputs(730) <= not(layer2_outputs(6633));
    outputs(731) <= (layer2_outputs(910)) and not (layer2_outputs(6320));
    outputs(732) <= (layer2_outputs(3980)) or (layer2_outputs(9281));
    outputs(733) <= not(layer2_outputs(3477));
    outputs(734) <= layer2_outputs(1741);
    outputs(735) <= not(layer2_outputs(1152));
    outputs(736) <= layer2_outputs(7946);
    outputs(737) <= layer2_outputs(4088);
    outputs(738) <= not(layer2_outputs(5112));
    outputs(739) <= layer2_outputs(3536);
    outputs(740) <= (layer2_outputs(2907)) and (layer2_outputs(3917));
    outputs(741) <= layer2_outputs(3947);
    outputs(742) <= not((layer2_outputs(1155)) xor (layer2_outputs(839)));
    outputs(743) <= not(layer2_outputs(2623)) or (layer2_outputs(2003));
    outputs(744) <= not(layer2_outputs(185));
    outputs(745) <= not(layer2_outputs(1766));
    outputs(746) <= not(layer2_outputs(334));
    outputs(747) <= layer2_outputs(2487);
    outputs(748) <= layer2_outputs(8697);
    outputs(749) <= not((layer2_outputs(4955)) or (layer2_outputs(8818)));
    outputs(750) <= not(layer2_outputs(3179));
    outputs(751) <= not(layer2_outputs(5887));
    outputs(752) <= not(layer2_outputs(1321));
    outputs(753) <= not(layer2_outputs(6476));
    outputs(754) <= layer2_outputs(6183);
    outputs(755) <= (layer2_outputs(617)) and not (layer2_outputs(7040));
    outputs(756) <= layer2_outputs(8660);
    outputs(757) <= not(layer2_outputs(531));
    outputs(758) <= layer2_outputs(1023);
    outputs(759) <= not(layer2_outputs(8388));
    outputs(760) <= not(layer2_outputs(3787));
    outputs(761) <= (layer2_outputs(140)) xor (layer2_outputs(5098));
    outputs(762) <= layer2_outputs(97);
    outputs(763) <= not(layer2_outputs(5721));
    outputs(764) <= not(layer2_outputs(3446));
    outputs(765) <= layer2_outputs(4498);
    outputs(766) <= (layer2_outputs(5832)) xor (layer2_outputs(9821));
    outputs(767) <= layer2_outputs(6856);
    outputs(768) <= not(layer2_outputs(5887)) or (layer2_outputs(6705));
    outputs(769) <= not(layer2_outputs(8414));
    outputs(770) <= layer2_outputs(2391);
    outputs(771) <= not(layer2_outputs(1294));
    outputs(772) <= not(layer2_outputs(139));
    outputs(773) <= not((layer2_outputs(4519)) xor (layer2_outputs(6050)));
    outputs(774) <= not(layer2_outputs(1324));
    outputs(775) <= layer2_outputs(9844);
    outputs(776) <= layer2_outputs(3442);
    outputs(777) <= layer2_outputs(3851);
    outputs(778) <= not(layer2_outputs(9979));
    outputs(779) <= layer2_outputs(4384);
    outputs(780) <= (layer2_outputs(5077)) xor (layer2_outputs(8992));
    outputs(781) <= not(layer2_outputs(2571));
    outputs(782) <= (layer2_outputs(4921)) or (layer2_outputs(4877));
    outputs(783) <= layer2_outputs(3649);
    outputs(784) <= layer2_outputs(1345);
    outputs(785) <= not(layer2_outputs(8640)) or (layer2_outputs(825));
    outputs(786) <= layer2_outputs(10118);
    outputs(787) <= layer2_outputs(7559);
    outputs(788) <= layer2_outputs(2384);
    outputs(789) <= not((layer2_outputs(6946)) or (layer2_outputs(8905)));
    outputs(790) <= layer2_outputs(6009);
    outputs(791) <= not(layer2_outputs(1702));
    outputs(792) <= (layer2_outputs(7109)) and not (layer2_outputs(4210));
    outputs(793) <= not(layer2_outputs(8634));
    outputs(794) <= not(layer2_outputs(816)) or (layer2_outputs(7892));
    outputs(795) <= not(layer2_outputs(9792));
    outputs(796) <= layer2_outputs(7123);
    outputs(797) <= layer2_outputs(8503);
    outputs(798) <= layer2_outputs(5819);
    outputs(799) <= (layer2_outputs(5875)) xor (layer2_outputs(109));
    outputs(800) <= not(layer2_outputs(737));
    outputs(801) <= not(layer2_outputs(1097));
    outputs(802) <= (layer2_outputs(793)) xor (layer2_outputs(9705));
    outputs(803) <= layer2_outputs(7546);
    outputs(804) <= not(layer2_outputs(9759));
    outputs(805) <= layer2_outputs(3097);
    outputs(806) <= layer2_outputs(5492);
    outputs(807) <= not(layer2_outputs(1908));
    outputs(808) <= not(layer2_outputs(4778));
    outputs(809) <= not(layer2_outputs(2670));
    outputs(810) <= layer2_outputs(9758);
    outputs(811) <= not(layer2_outputs(8644));
    outputs(812) <= layer2_outputs(5751);
    outputs(813) <= not(layer2_outputs(181));
    outputs(814) <= layer2_outputs(3157);
    outputs(815) <= not(layer2_outputs(5798));
    outputs(816) <= not((layer2_outputs(9235)) and (layer2_outputs(6315)));
    outputs(817) <= not(layer2_outputs(478));
    outputs(818) <= not(layer2_outputs(7662));
    outputs(819) <= not(layer2_outputs(4392));
    outputs(820) <= layer2_outputs(4466);
    outputs(821) <= not(layer2_outputs(3194));
    outputs(822) <= (layer2_outputs(1241)) and not (layer2_outputs(2825));
    outputs(823) <= layer2_outputs(7759);
    outputs(824) <= not((layer2_outputs(4718)) xor (layer2_outputs(3952)));
    outputs(825) <= layer2_outputs(4318);
    outputs(826) <= not(layer2_outputs(3617));
    outputs(827) <= layer2_outputs(7822);
    outputs(828) <= (layer2_outputs(143)) xor (layer2_outputs(5402));
    outputs(829) <= not(layer2_outputs(8415));
    outputs(830) <= layer2_outputs(8770);
    outputs(831) <= not((layer2_outputs(6680)) xor (layer2_outputs(6344)));
    outputs(832) <= not(layer2_outputs(8637));
    outputs(833) <= not(layer2_outputs(6223));
    outputs(834) <= (layer2_outputs(6651)) or (layer2_outputs(4091));
    outputs(835) <= not((layer2_outputs(2490)) or (layer2_outputs(8036)));
    outputs(836) <= layer2_outputs(8049);
    outputs(837) <= not((layer2_outputs(8937)) or (layer2_outputs(334)));
    outputs(838) <= layer2_outputs(3546);
    outputs(839) <= layer2_outputs(6379);
    outputs(840) <= not((layer2_outputs(10141)) xor (layer2_outputs(7991)));
    outputs(841) <= layer2_outputs(3019);
    outputs(842) <= layer2_outputs(6539);
    outputs(843) <= not(layer2_outputs(4859));
    outputs(844) <= layer2_outputs(5109);
    outputs(845) <= not((layer2_outputs(6719)) or (layer2_outputs(7201)));
    outputs(846) <= (layer2_outputs(1744)) and (layer2_outputs(1420));
    outputs(847) <= not(layer2_outputs(9876)) or (layer2_outputs(1390));
    outputs(848) <= not(layer2_outputs(6634));
    outputs(849) <= not(layer2_outputs(9396));
    outputs(850) <= layer2_outputs(3258);
    outputs(851) <= layer2_outputs(574);
    outputs(852) <= layer2_outputs(6591);
    outputs(853) <= (layer2_outputs(9594)) and not (layer2_outputs(10049));
    outputs(854) <= (layer2_outputs(4434)) xor (layer2_outputs(4822));
    outputs(855) <= not(layer2_outputs(4455));
    outputs(856) <= (layer2_outputs(10103)) xor (layer2_outputs(8590));
    outputs(857) <= (layer2_outputs(4917)) xor (layer2_outputs(6559));
    outputs(858) <= (layer2_outputs(959)) and not (layer2_outputs(1098));
    outputs(859) <= layer2_outputs(3705);
    outputs(860) <= layer2_outputs(7359);
    outputs(861) <= not((layer2_outputs(6372)) xor (layer2_outputs(6688)));
    outputs(862) <= not((layer2_outputs(4717)) or (layer2_outputs(5118)));
    outputs(863) <= not((layer2_outputs(7973)) xor (layer2_outputs(8597)));
    outputs(864) <= not(layer2_outputs(3541));
    outputs(865) <= layer2_outputs(7080);
    outputs(866) <= layer2_outputs(8829);
    outputs(867) <= (layer2_outputs(9715)) and (layer2_outputs(9507));
    outputs(868) <= not(layer2_outputs(2485));
    outputs(869) <= not((layer2_outputs(7036)) xor (layer2_outputs(6863)));
    outputs(870) <= not(layer2_outputs(710)) or (layer2_outputs(7239));
    outputs(871) <= (layer2_outputs(6424)) xor (layer2_outputs(7417));
    outputs(872) <= not(layer2_outputs(788));
    outputs(873) <= not(layer2_outputs(2538));
    outputs(874) <= layer2_outputs(9122);
    outputs(875) <= not(layer2_outputs(997));
    outputs(876) <= layer2_outputs(621);
    outputs(877) <= not((layer2_outputs(4162)) xor (layer2_outputs(526)));
    outputs(878) <= not(layer2_outputs(9660));
    outputs(879) <= not(layer2_outputs(9642));
    outputs(880) <= (layer2_outputs(3915)) and (layer2_outputs(2200));
    outputs(881) <= not(layer2_outputs(7826));
    outputs(882) <= not(layer2_outputs(9102));
    outputs(883) <= not(layer2_outputs(2885));
    outputs(884) <= layer2_outputs(8005);
    outputs(885) <= not(layer2_outputs(3698));
    outputs(886) <= not(layer2_outputs(6280));
    outputs(887) <= (layer2_outputs(135)) xor (layer2_outputs(2601));
    outputs(888) <= not((layer2_outputs(9741)) xor (layer2_outputs(3113)));
    outputs(889) <= layer2_outputs(5676);
    outputs(890) <= layer2_outputs(214);
    outputs(891) <= layer2_outputs(6282);
    outputs(892) <= not(layer2_outputs(9704));
    outputs(893) <= not((layer2_outputs(4772)) or (layer2_outputs(7177)));
    outputs(894) <= (layer2_outputs(4910)) xor (layer2_outputs(3195));
    outputs(895) <= (layer2_outputs(355)) xor (layer2_outputs(2745));
    outputs(896) <= (layer2_outputs(3371)) and not (layer2_outputs(9239));
    outputs(897) <= (layer2_outputs(3121)) and (layer2_outputs(4793));
    outputs(898) <= layer2_outputs(1451);
    outputs(899) <= (layer2_outputs(1416)) xor (layer2_outputs(7020));
    outputs(900) <= not(layer2_outputs(2593));
    outputs(901) <= not(layer2_outputs(9440));
    outputs(902) <= not(layer2_outputs(613));
    outputs(903) <= layer2_outputs(5222);
    outputs(904) <= (layer2_outputs(322)) xor (layer2_outputs(9184));
    outputs(905) <= layer2_outputs(7520);
    outputs(906) <= not(layer2_outputs(1806));
    outputs(907) <= (layer2_outputs(1396)) and not (layer2_outputs(8124));
    outputs(908) <= not(layer2_outputs(8612));
    outputs(909) <= layer2_outputs(4527);
    outputs(910) <= not(layer2_outputs(2349));
    outputs(911) <= (layer2_outputs(4688)) and (layer2_outputs(5906));
    outputs(912) <= (layer2_outputs(7059)) xor (layer2_outputs(5621));
    outputs(913) <= layer2_outputs(575);
    outputs(914) <= not(layer2_outputs(6151));
    outputs(915) <= not(layer2_outputs(2596));
    outputs(916) <= (layer2_outputs(7732)) and not (layer2_outputs(7781));
    outputs(917) <= not(layer2_outputs(7106));
    outputs(918) <= (layer2_outputs(2273)) xor (layer2_outputs(1937));
    outputs(919) <= layer2_outputs(5590);
    outputs(920) <= not((layer2_outputs(6342)) or (layer2_outputs(4301)));
    outputs(921) <= not(layer2_outputs(8901));
    outputs(922) <= layer2_outputs(6591);
    outputs(923) <= (layer2_outputs(8893)) xor (layer2_outputs(6780));
    outputs(924) <= (layer2_outputs(6976)) and (layer2_outputs(2260));
    outputs(925) <= layer2_outputs(7460);
    outputs(926) <= not(layer2_outputs(6349));
    outputs(927) <= layer2_outputs(1594);
    outputs(928) <= (layer2_outputs(8300)) xor (layer2_outputs(1804));
    outputs(929) <= layer2_outputs(8632);
    outputs(930) <= layer2_outputs(1486);
    outputs(931) <= layer2_outputs(9342);
    outputs(932) <= layer2_outputs(8401);
    outputs(933) <= not(layer2_outputs(368));
    outputs(934) <= not(layer2_outputs(6176));
    outputs(935) <= not(layer2_outputs(164));
    outputs(936) <= (layer2_outputs(1037)) and not (layer2_outputs(3829));
    outputs(937) <= (layer2_outputs(9857)) and not (layer2_outputs(5969));
    outputs(938) <= (layer2_outputs(4060)) or (layer2_outputs(1082));
    outputs(939) <= not(layer2_outputs(6426)) or (layer2_outputs(4347));
    outputs(940) <= not((layer2_outputs(7472)) and (layer2_outputs(3444)));
    outputs(941) <= not(layer2_outputs(4883));
    outputs(942) <= not((layer2_outputs(3044)) and (layer2_outputs(5724)));
    outputs(943) <= not(layer2_outputs(7166));
    outputs(944) <= not((layer2_outputs(8018)) xor (layer2_outputs(1887)));
    outputs(945) <= layer2_outputs(7475);
    outputs(946) <= not((layer2_outputs(8361)) or (layer2_outputs(8762)));
    outputs(947) <= not(layer2_outputs(10172));
    outputs(948) <= layer2_outputs(2843);
    outputs(949) <= not(layer2_outputs(7275));
    outputs(950) <= not((layer2_outputs(7407)) xor (layer2_outputs(8959)));
    outputs(951) <= layer2_outputs(6368);
    outputs(952) <= (layer2_outputs(8726)) xor (layer2_outputs(3180));
    outputs(953) <= not(layer2_outputs(262));
    outputs(954) <= (layer2_outputs(7352)) or (layer2_outputs(8972));
    outputs(955) <= layer2_outputs(2697);
    outputs(956) <= (layer2_outputs(6036)) and not (layer2_outputs(94));
    outputs(957) <= layer2_outputs(5817);
    outputs(958) <= (layer2_outputs(7037)) and not (layer2_outputs(8316));
    outputs(959) <= not(layer2_outputs(2718));
    outputs(960) <= layer2_outputs(4694);
    outputs(961) <= not((layer2_outputs(3849)) and (layer2_outputs(2342)));
    outputs(962) <= (layer2_outputs(7928)) xor (layer2_outputs(1811));
    outputs(963) <= layer2_outputs(890);
    outputs(964) <= not((layer2_outputs(3695)) xor (layer2_outputs(7928)));
    outputs(965) <= not((layer2_outputs(7768)) xor (layer2_outputs(7597)));
    outputs(966) <= not(layer2_outputs(8663));
    outputs(967) <= (layer2_outputs(9357)) xor (layer2_outputs(5758));
    outputs(968) <= not(layer2_outputs(2243));
    outputs(969) <= not(layer2_outputs(9299));
    outputs(970) <= layer2_outputs(776);
    outputs(971) <= not(layer2_outputs(1334));
    outputs(972) <= layer2_outputs(7793);
    outputs(973) <= not(layer2_outputs(8031));
    outputs(974) <= layer2_outputs(4906);
    outputs(975) <= layer2_outputs(9139);
    outputs(976) <= layer2_outputs(10116);
    outputs(977) <= layer2_outputs(7404);
    outputs(978) <= (layer2_outputs(3315)) and not (layer2_outputs(9658));
    outputs(979) <= layer2_outputs(4703);
    outputs(980) <= layer2_outputs(55);
    outputs(981) <= layer2_outputs(4667);
    outputs(982) <= not((layer2_outputs(4454)) xor (layer2_outputs(1599)));
    outputs(983) <= not(layer2_outputs(2));
    outputs(984) <= not(layer2_outputs(10077));
    outputs(985) <= not(layer2_outputs(5032));
    outputs(986) <= (layer2_outputs(1923)) xor (layer2_outputs(477));
    outputs(987) <= layer2_outputs(3435);
    outputs(988) <= (layer2_outputs(8349)) xor (layer2_outputs(5911));
    outputs(989) <= not(layer2_outputs(4927));
    outputs(990) <= layer2_outputs(963);
    outputs(991) <= layer2_outputs(5419);
    outputs(992) <= (layer2_outputs(6001)) xor (layer2_outputs(5198));
    outputs(993) <= (layer2_outputs(4031)) and not (layer2_outputs(5629));
    outputs(994) <= layer2_outputs(10086);
    outputs(995) <= layer2_outputs(5555);
    outputs(996) <= not(layer2_outputs(7821));
    outputs(997) <= layer2_outputs(1545);
    outputs(998) <= not(layer2_outputs(9439));
    outputs(999) <= layer2_outputs(1830);
    outputs(1000) <= not(layer2_outputs(4372));
    outputs(1001) <= not(layer2_outputs(2079)) or (layer2_outputs(8969));
    outputs(1002) <= layer2_outputs(5686);
    outputs(1003) <= layer2_outputs(9904);
    outputs(1004) <= not(layer2_outputs(6207));
    outputs(1005) <= layer2_outputs(6841);
    outputs(1006) <= layer2_outputs(2881);
    outputs(1007) <= not(layer2_outputs(1272));
    outputs(1008) <= layer2_outputs(5081);
    outputs(1009) <= not(layer2_outputs(4366));
    outputs(1010) <= not((layer2_outputs(6546)) and (layer2_outputs(133)));
    outputs(1011) <= not(layer2_outputs(1216));
    outputs(1012) <= not((layer2_outputs(8647)) xor (layer2_outputs(3952)));
    outputs(1013) <= (layer2_outputs(9037)) and not (layer2_outputs(2766));
    outputs(1014) <= (layer2_outputs(5127)) xor (layer2_outputs(2158));
    outputs(1015) <= not(layer2_outputs(3981));
    outputs(1016) <= not(layer2_outputs(544));
    outputs(1017) <= not(layer2_outputs(8760));
    outputs(1018) <= (layer2_outputs(10170)) xor (layer2_outputs(4252));
    outputs(1019) <= not(layer2_outputs(7693));
    outputs(1020) <= not(layer2_outputs(731)) or (layer2_outputs(5935));
    outputs(1021) <= not(layer2_outputs(8880));
    outputs(1022) <= not((layer2_outputs(9894)) xor (layer2_outputs(6618)));
    outputs(1023) <= layer2_outputs(2697);
    outputs(1024) <= layer2_outputs(2217);
    outputs(1025) <= not(layer2_outputs(2052));
    outputs(1026) <= layer2_outputs(772);
    outputs(1027) <= (layer2_outputs(2779)) and (layer2_outputs(1777));
    outputs(1028) <= not(layer2_outputs(4952));
    outputs(1029) <= not(layer2_outputs(1321)) or (layer2_outputs(1795));
    outputs(1030) <= layer2_outputs(5125);
    outputs(1031) <= (layer2_outputs(5365)) xor (layer2_outputs(9797));
    outputs(1032) <= layer2_outputs(9096);
    outputs(1033) <= not(layer2_outputs(8277));
    outputs(1034) <= (layer2_outputs(1980)) and not (layer2_outputs(2500));
    outputs(1035) <= not((layer2_outputs(4349)) xor (layer2_outputs(8647)));
    outputs(1036) <= not(layer2_outputs(3394));
    outputs(1037) <= (layer2_outputs(3383)) and (layer2_outputs(5681));
    outputs(1038) <= (layer2_outputs(9370)) and not (layer2_outputs(7823));
    outputs(1039) <= (layer2_outputs(2289)) and (layer2_outputs(6022));
    outputs(1040) <= (layer2_outputs(2655)) xor (layer2_outputs(2403));
    outputs(1041) <= not((layer2_outputs(10036)) or (layer2_outputs(4063)));
    outputs(1042) <= layer2_outputs(8230);
    outputs(1043) <= not(layer2_outputs(4572));
    outputs(1044) <= layer2_outputs(4790);
    outputs(1045) <= (layer2_outputs(9556)) or (layer2_outputs(908));
    outputs(1046) <= not(layer2_outputs(4096));
    outputs(1047) <= not((layer2_outputs(2505)) xor (layer2_outputs(9600)));
    outputs(1048) <= not((layer2_outputs(706)) xor (layer2_outputs(1671)));
    outputs(1049) <= layer2_outputs(130);
    outputs(1050) <= not((layer2_outputs(7777)) or (layer2_outputs(393)));
    outputs(1051) <= not((layer2_outputs(8403)) xor (layer2_outputs(4203)));
    outputs(1052) <= (layer2_outputs(7300)) and not (layer2_outputs(6146));
    outputs(1053) <= not((layer2_outputs(1837)) or (layer2_outputs(10185)));
    outputs(1054) <= not(layer2_outputs(7829));
    outputs(1055) <= not(layer2_outputs(7729));
    outputs(1056) <= (layer2_outputs(6041)) and not (layer2_outputs(9345));
    outputs(1057) <= (layer2_outputs(6761)) xor (layer2_outputs(5528));
    outputs(1058) <= layer2_outputs(1193);
    outputs(1059) <= (layer2_outputs(224)) xor (layer2_outputs(6757));
    outputs(1060) <= not(layer2_outputs(10177));
    outputs(1061) <= not((layer2_outputs(6785)) or (layer2_outputs(9913)));
    outputs(1062) <= not(layer2_outputs(8346));
    outputs(1063) <= not(layer2_outputs(2959));
    outputs(1064) <= (layer2_outputs(2154)) and not (layer2_outputs(5763));
    outputs(1065) <= not(layer2_outputs(10039));
    outputs(1066) <= (layer2_outputs(7289)) and (layer2_outputs(2523));
    outputs(1067) <= not((layer2_outputs(655)) xor (layer2_outputs(2240)));
    outputs(1068) <= not(layer2_outputs(2322));
    outputs(1069) <= (layer2_outputs(2903)) xor (layer2_outputs(9106));
    outputs(1070) <= not((layer2_outputs(6279)) xor (layer2_outputs(2329)));
    outputs(1071) <= not((layer2_outputs(9034)) xor (layer2_outputs(7776)));
    outputs(1072) <= (layer2_outputs(8360)) and (layer2_outputs(5714));
    outputs(1073) <= (layer2_outputs(3613)) and not (layer2_outputs(9935));
    outputs(1074) <= not(layer2_outputs(2002));
    outputs(1075) <= (layer2_outputs(352)) xor (layer2_outputs(5057));
    outputs(1076) <= layer2_outputs(9917);
    outputs(1077) <= not(layer2_outputs(781));
    outputs(1078) <= layer2_outputs(3356);
    outputs(1079) <= (layer2_outputs(721)) and (layer2_outputs(4789));
    outputs(1080) <= (layer2_outputs(1502)) and not (layer2_outputs(3552));
    outputs(1081) <= layer2_outputs(2457);
    outputs(1082) <= not(layer2_outputs(7774));
    outputs(1083) <= '0';
    outputs(1084) <= layer2_outputs(1258);
    outputs(1085) <= not(layer2_outputs(7504));
    outputs(1086) <= layer2_outputs(157);
    outputs(1087) <= layer2_outputs(9484);
    outputs(1088) <= layer2_outputs(7802);
    outputs(1089) <= not((layer2_outputs(9754)) or (layer2_outputs(2057)));
    outputs(1090) <= not((layer2_outputs(3665)) xor (layer2_outputs(7404)));
    outputs(1091) <= not(layer2_outputs(4903));
    outputs(1092) <= not(layer2_outputs(2385));
    outputs(1093) <= layer2_outputs(1108);
    outputs(1094) <= (layer2_outputs(618)) xor (layer2_outputs(3174));
    outputs(1095) <= not(layer2_outputs(652));
    outputs(1096) <= (layer2_outputs(6781)) xor (layer2_outputs(5841));
    outputs(1097) <= not(layer2_outputs(4530));
    outputs(1098) <= not((layer2_outputs(8505)) xor (layer2_outputs(2100)));
    outputs(1099) <= layer2_outputs(7623);
    outputs(1100) <= (layer2_outputs(5942)) xor (layer2_outputs(9757));
    outputs(1101) <= (layer2_outputs(1397)) and not (layer2_outputs(9242));
    outputs(1102) <= not((layer2_outputs(4053)) or (layer2_outputs(3551)));
    outputs(1103) <= not(layer2_outputs(1610));
    outputs(1104) <= not(layer2_outputs(6849));
    outputs(1105) <= (layer2_outputs(5473)) and not (layer2_outputs(3991));
    outputs(1106) <= layer2_outputs(7576);
    outputs(1107) <= layer2_outputs(8285);
    outputs(1108) <= not(layer2_outputs(1467));
    outputs(1109) <= (layer2_outputs(2602)) xor (layer2_outputs(5414));
    outputs(1110) <= not(layer2_outputs(9606));
    outputs(1111) <= not(layer2_outputs(946));
    outputs(1112) <= not(layer2_outputs(9756));
    outputs(1113) <= not(layer2_outputs(847)) or (layer2_outputs(7073));
    outputs(1114) <= (layer2_outputs(8069)) and (layer2_outputs(4654));
    outputs(1115) <= not(layer2_outputs(10143));
    outputs(1116) <= not((layer2_outputs(7542)) xor (layer2_outputs(1214)));
    outputs(1117) <= not(layer2_outputs(5380));
    outputs(1118) <= (layer2_outputs(6502)) and not (layer2_outputs(7208));
    outputs(1119) <= layer2_outputs(5749);
    outputs(1120) <= layer2_outputs(3697);
    outputs(1121) <= (layer2_outputs(6810)) and (layer2_outputs(2282));
    outputs(1122) <= not((layer2_outputs(1196)) xor (layer2_outputs(3672)));
    outputs(1123) <= not(layer2_outputs(246));
    outputs(1124) <= not(layer2_outputs(6021));
    outputs(1125) <= not(layer2_outputs(4810));
    outputs(1126) <= not(layer2_outputs(8536));
    outputs(1127) <= (layer2_outputs(6611)) and not (layer2_outputs(9603));
    outputs(1128) <= (layer2_outputs(1951)) and not (layer2_outputs(1024));
    outputs(1129) <= not(layer2_outputs(1849));
    outputs(1130) <= not(layer2_outputs(937)) or (layer2_outputs(4741));
    outputs(1131) <= not(layer2_outputs(7906));
    outputs(1132) <= (layer2_outputs(2167)) and not (layer2_outputs(3805));
    outputs(1133) <= layer2_outputs(7698);
    outputs(1134) <= (layer2_outputs(10187)) xor (layer2_outputs(9276));
    outputs(1135) <= not(layer2_outputs(3176));
    outputs(1136) <= layer2_outputs(6425);
    outputs(1137) <= not(layer2_outputs(5918));
    outputs(1138) <= not(layer2_outputs(9026));
    outputs(1139) <= layer2_outputs(7592);
    outputs(1140) <= (layer2_outputs(9691)) xor (layer2_outputs(6928));
    outputs(1141) <= (layer2_outputs(4762)) and not (layer2_outputs(10107));
    outputs(1142) <= layer2_outputs(3723);
    outputs(1143) <= not(layer2_outputs(9820));
    outputs(1144) <= not((layer2_outputs(1053)) or (layer2_outputs(7778)));
    outputs(1145) <= layer2_outputs(3703);
    outputs(1146) <= (layer2_outputs(4950)) and not (layer2_outputs(2161));
    outputs(1147) <= not(layer2_outputs(6420));
    outputs(1148) <= layer2_outputs(5734);
    outputs(1149) <= (layer2_outputs(4681)) and not (layer2_outputs(2828));
    outputs(1150) <= layer2_outputs(707);
    outputs(1151) <= not((layer2_outputs(7480)) xor (layer2_outputs(9798)));
    outputs(1152) <= (layer2_outputs(1456)) and (layer2_outputs(2689));
    outputs(1153) <= not(layer2_outputs(6552));
    outputs(1154) <= not(layer2_outputs(7097));
    outputs(1155) <= not((layer2_outputs(9779)) or (layer2_outputs(5126)));
    outputs(1156) <= layer2_outputs(5716);
    outputs(1157) <= not(layer2_outputs(4938));
    outputs(1158) <= not(layer2_outputs(8140));
    outputs(1159) <= (layer2_outputs(3930)) xor (layer2_outputs(103));
    outputs(1160) <= not((layer2_outputs(8599)) xor (layer2_outputs(8131)));
    outputs(1161) <= (layer2_outputs(7173)) xor (layer2_outputs(9595));
    outputs(1162) <= (layer2_outputs(9405)) and not (layer2_outputs(7426));
    outputs(1163) <= layer2_outputs(8362);
    outputs(1164) <= layer2_outputs(86);
    outputs(1165) <= layer2_outputs(3741);
    outputs(1166) <= layer2_outputs(8670);
    outputs(1167) <= not((layer2_outputs(4769)) xor (layer2_outputs(10127)));
    outputs(1168) <= layer2_outputs(10200);
    outputs(1169) <= not(layer2_outputs(8855));
    outputs(1170) <= (layer2_outputs(674)) and not (layer2_outputs(5520));
    outputs(1171) <= not(layer2_outputs(9477));
    outputs(1172) <= layer2_outputs(10029);
    outputs(1173) <= layer2_outputs(9761);
    outputs(1174) <= (layer2_outputs(1147)) xor (layer2_outputs(4341));
    outputs(1175) <= not((layer2_outputs(8221)) or (layer2_outputs(3274)));
    outputs(1176) <= (layer2_outputs(9415)) xor (layer2_outputs(4525));
    outputs(1177) <= (layer2_outputs(10064)) xor (layer2_outputs(1014));
    outputs(1178) <= layer2_outputs(10003);
    outputs(1179) <= layer2_outputs(9176);
    outputs(1180) <= not(layer2_outputs(227));
    outputs(1181) <= (layer2_outputs(4005)) xor (layer2_outputs(8626));
    outputs(1182) <= (layer2_outputs(1766)) and not (layer2_outputs(6159));
    outputs(1183) <= not(layer2_outputs(1990));
    outputs(1184) <= (layer2_outputs(5079)) and (layer2_outputs(3403));
    outputs(1185) <= layer2_outputs(9860);
    outputs(1186) <= layer2_outputs(6958);
    outputs(1187) <= (layer2_outputs(7129)) and not (layer2_outputs(1012));
    outputs(1188) <= layer2_outputs(5762);
    outputs(1189) <= (layer2_outputs(10132)) and not (layer2_outputs(8060));
    outputs(1190) <= layer2_outputs(9953);
    outputs(1191) <= not(layer2_outputs(4692));
    outputs(1192) <= (layer2_outputs(1280)) and (layer2_outputs(2579));
    outputs(1193) <= not(layer2_outputs(2234));
    outputs(1194) <= layer2_outputs(8053);
    outputs(1195) <= (layer2_outputs(5318)) and (layer2_outputs(5756));
    outputs(1196) <= layer2_outputs(8611);
    outputs(1197) <= not(layer2_outputs(859));
    outputs(1198) <= not((layer2_outputs(6397)) xor (layer2_outputs(4328)));
    outputs(1199) <= layer2_outputs(6609);
    outputs(1200) <= (layer2_outputs(10001)) and (layer2_outputs(7308));
    outputs(1201) <= (layer2_outputs(9990)) and (layer2_outputs(9912));
    outputs(1202) <= layer2_outputs(50);
    outputs(1203) <= not(layer2_outputs(4560));
    outputs(1204) <= (layer2_outputs(6944)) and not (layer2_outputs(9740));
    outputs(1205) <= (layer2_outputs(9959)) and not (layer2_outputs(2424));
    outputs(1206) <= layer2_outputs(1429);
    outputs(1207) <= not(layer2_outputs(2987));
    outputs(1208) <= layer2_outputs(9994);
    outputs(1209) <= (layer2_outputs(5129)) or (layer2_outputs(6484));
    outputs(1210) <= not((layer2_outputs(9071)) or (layer2_outputs(6102)));
    outputs(1211) <= layer2_outputs(692);
    outputs(1212) <= not(layer2_outputs(4583));
    outputs(1213) <= not(layer2_outputs(9753));
    outputs(1214) <= layer2_outputs(1932);
    outputs(1215) <= layer2_outputs(2937);
    outputs(1216) <= layer2_outputs(1915);
    outputs(1217) <= not((layer2_outputs(445)) xor (layer2_outputs(1819)));
    outputs(1218) <= not(layer2_outputs(10169));
    outputs(1219) <= layer2_outputs(9193);
    outputs(1220) <= (layer2_outputs(7391)) and (layer2_outputs(9842));
    outputs(1221) <= not((layer2_outputs(8842)) xor (layer2_outputs(8073)));
    outputs(1222) <= (layer2_outputs(5865)) xor (layer2_outputs(1411));
    outputs(1223) <= layer2_outputs(5234);
    outputs(1224) <= not(layer2_outputs(1340));
    outputs(1225) <= (layer2_outputs(6298)) xor (layer2_outputs(4048));
    outputs(1226) <= not((layer2_outputs(8847)) or (layer2_outputs(6720)));
    outputs(1227) <= layer2_outputs(1113);
    outputs(1228) <= layer2_outputs(7199);
    outputs(1229) <= (layer2_outputs(3517)) xor (layer2_outputs(976));
    outputs(1230) <= (layer2_outputs(4932)) and not (layer2_outputs(3942));
    outputs(1231) <= layer2_outputs(5247);
    outputs(1232) <= (layer2_outputs(6361)) or (layer2_outputs(2648));
    outputs(1233) <= not(layer2_outputs(315));
    outputs(1234) <= not((layer2_outputs(7774)) xor (layer2_outputs(5969)));
    outputs(1235) <= not((layer2_outputs(6698)) or (layer2_outputs(7363)));
    outputs(1236) <= layer2_outputs(8050);
    outputs(1237) <= (layer2_outputs(4842)) and not (layer2_outputs(3967));
    outputs(1238) <= (layer2_outputs(6820)) and not (layer2_outputs(7647));
    outputs(1239) <= (layer2_outputs(6549)) and not (layer2_outputs(2832));
    outputs(1240) <= not(layer2_outputs(4282));
    outputs(1241) <= not((layer2_outputs(2189)) xor (layer2_outputs(7235)));
    outputs(1242) <= (layer2_outputs(2979)) and not (layer2_outputs(9472));
    outputs(1243) <= not((layer2_outputs(7887)) xor (layer2_outputs(9553)));
    outputs(1244) <= not((layer2_outputs(7536)) or (layer2_outputs(9294)));
    outputs(1245) <= (layer2_outputs(5228)) xor (layer2_outputs(3651));
    outputs(1246) <= (layer2_outputs(2476)) and (layer2_outputs(7557));
    outputs(1247) <= (layer2_outputs(8215)) xor (layer2_outputs(216));
    outputs(1248) <= layer2_outputs(1906);
    outputs(1249) <= (layer2_outputs(4860)) and not (layer2_outputs(659));
    outputs(1250) <= not(layer2_outputs(9027));
    outputs(1251) <= not(layer2_outputs(4670)) or (layer2_outputs(5104));
    outputs(1252) <= not(layer2_outputs(7564));
    outputs(1253) <= layer2_outputs(8198);
    outputs(1254) <= not((layer2_outputs(4378)) xor (layer2_outputs(2966)));
    outputs(1255) <= not((layer2_outputs(7539)) or (layer2_outputs(781)));
    outputs(1256) <= not(layer2_outputs(4583));
    outputs(1257) <= not(layer2_outputs(8819));
    outputs(1258) <= (layer2_outputs(9049)) xor (layer2_outputs(9649));
    outputs(1259) <= (layer2_outputs(8812)) xor (layer2_outputs(4941));
    outputs(1260) <= (layer2_outputs(559)) and not (layer2_outputs(9666));
    outputs(1261) <= not((layer2_outputs(1586)) or (layer2_outputs(681)));
    outputs(1262) <= (layer2_outputs(2799)) and (layer2_outputs(1344));
    outputs(1263) <= (layer2_outputs(4306)) and not (layer2_outputs(2239));
    outputs(1264) <= (layer2_outputs(9566)) xor (layer2_outputs(3529));
    outputs(1265) <= not(layer2_outputs(8462));
    outputs(1266) <= layer2_outputs(1461);
    outputs(1267) <= layer2_outputs(6027);
    outputs(1268) <= not((layer2_outputs(5547)) xor (layer2_outputs(1596)));
    outputs(1269) <= (layer2_outputs(3215)) and not (layer2_outputs(1419));
    outputs(1270) <= (layer2_outputs(9713)) xor (layer2_outputs(8924));
    outputs(1271) <= not(layer2_outputs(2362));
    outputs(1272) <= (layer2_outputs(8876)) and not (layer2_outputs(5211));
    outputs(1273) <= (layer2_outputs(7167)) and not (layer2_outputs(705));
    outputs(1274) <= not(layer2_outputs(2673));
    outputs(1275) <= not((layer2_outputs(7687)) or (layer2_outputs(9233)));
    outputs(1276) <= not((layer2_outputs(1269)) xor (layer2_outputs(4603)));
    outputs(1277) <= (layer2_outputs(2242)) and (layer2_outputs(4018));
    outputs(1278) <= not((layer2_outputs(686)) xor (layer2_outputs(7573)));
    outputs(1279) <= (layer2_outputs(8657)) xor (layer2_outputs(8084));
    outputs(1280) <= (layer2_outputs(7440)) and not (layer2_outputs(3099));
    outputs(1281) <= not((layer2_outputs(4315)) or (layer2_outputs(5000)));
    outputs(1282) <= not((layer2_outputs(5554)) or (layer2_outputs(2640)));
    outputs(1283) <= (layer2_outputs(5152)) xor (layer2_outputs(1128));
    outputs(1284) <= (layer2_outputs(7937)) and (layer2_outputs(7939));
    outputs(1285) <= not(layer2_outputs(6136));
    outputs(1286) <= not((layer2_outputs(6079)) or (layer2_outputs(6563)));
    outputs(1287) <= not(layer2_outputs(1500));
    outputs(1288) <= not(layer2_outputs(4812));
    outputs(1289) <= layer2_outputs(3717);
    outputs(1290) <= not((layer2_outputs(5072)) or (layer2_outputs(2757)));
    outputs(1291) <= not((layer2_outputs(1045)) or (layer2_outputs(259)));
    outputs(1292) <= (layer2_outputs(10213)) xor (layer2_outputs(10185));
    outputs(1293) <= layer2_outputs(9665);
    outputs(1294) <= (layer2_outputs(4925)) and (layer2_outputs(735));
    outputs(1295) <= (layer2_outputs(1132)) xor (layer2_outputs(8402));
    outputs(1296) <= layer2_outputs(2304);
    outputs(1297) <= layer2_outputs(7171);
    outputs(1298) <= not(layer2_outputs(5446));
    outputs(1299) <= (layer2_outputs(4500)) and not (layer2_outputs(8651));
    outputs(1300) <= not(layer2_outputs(9195));
    outputs(1301) <= not((layer2_outputs(5152)) xor (layer2_outputs(3708)));
    outputs(1302) <= not(layer2_outputs(3239));
    outputs(1303) <= not(layer2_outputs(8202));
    outputs(1304) <= layer2_outputs(10159);
    outputs(1305) <= not((layer2_outputs(1843)) or (layer2_outputs(1261)));
    outputs(1306) <= not((layer2_outputs(9115)) or (layer2_outputs(9330)));
    outputs(1307) <= (layer2_outputs(193)) xor (layer2_outputs(9935));
    outputs(1308) <= layer2_outputs(858);
    outputs(1309) <= not(layer2_outputs(9786));
    outputs(1310) <= (layer2_outputs(556)) and not (layer2_outputs(664));
    outputs(1311) <= not(layer2_outputs(10197));
    outputs(1312) <= not((layer2_outputs(8347)) or (layer2_outputs(2715)));
    outputs(1313) <= layer2_outputs(3240);
    outputs(1314) <= layer2_outputs(3742);
    outputs(1315) <= (layer2_outputs(5054)) and not (layer2_outputs(6729));
    outputs(1316) <= (layer2_outputs(7135)) xor (layer2_outputs(7233));
    outputs(1317) <= (layer2_outputs(9076)) xor (layer2_outputs(4851));
    outputs(1318) <= (layer2_outputs(4319)) and not (layer2_outputs(3590));
    outputs(1319) <= layer2_outputs(3057);
    outputs(1320) <= (layer2_outputs(7631)) and not (layer2_outputs(3027));
    outputs(1321) <= not((layer2_outputs(6253)) xor (layer2_outputs(965)));
    outputs(1322) <= (layer2_outputs(1013)) and not (layer2_outputs(4284));
    outputs(1323) <= (layer2_outputs(7089)) and not (layer2_outputs(8950));
    outputs(1324) <= not((layer2_outputs(2953)) or (layer2_outputs(3792)));
    outputs(1325) <= (layer2_outputs(4258)) and not (layer2_outputs(10147));
    outputs(1326) <= not(layer2_outputs(4661));
    outputs(1327) <= layer2_outputs(497);
    outputs(1328) <= (layer2_outputs(6603)) and not (layer2_outputs(8315));
    outputs(1329) <= not((layer2_outputs(6104)) or (layer2_outputs(9689)));
    outputs(1330) <= (layer2_outputs(6931)) and (layer2_outputs(8502));
    outputs(1331) <= layer2_outputs(502);
    outputs(1332) <= not(layer2_outputs(8382));
    outputs(1333) <= (layer2_outputs(9671)) and (layer2_outputs(1968));
    outputs(1334) <= layer2_outputs(8412);
    outputs(1335) <= (layer2_outputs(3335)) and (layer2_outputs(9926));
    outputs(1336) <= not(layer2_outputs(2271));
    outputs(1337) <= (layer2_outputs(4233)) xor (layer2_outputs(6787));
    outputs(1338) <= (layer2_outputs(35)) xor (layer2_outputs(2477));
    outputs(1339) <= (layer2_outputs(8226)) xor (layer2_outputs(2345));
    outputs(1340) <= not(layer2_outputs(7444));
    outputs(1341) <= (layer2_outputs(6800)) xor (layer2_outputs(3203));
    outputs(1342) <= (layer2_outputs(1453)) xor (layer2_outputs(1781));
    outputs(1343) <= not((layer2_outputs(8294)) or (layer2_outputs(6172)));
    outputs(1344) <= (layer2_outputs(4435)) and not (layer2_outputs(5578));
    outputs(1345) <= not(layer2_outputs(6135));
    outputs(1346) <= not(layer2_outputs(4710));
    outputs(1347) <= (layer2_outputs(4835)) xor (layer2_outputs(6145));
    outputs(1348) <= (layer2_outputs(7499)) xor (layer2_outputs(6596));
    outputs(1349) <= not(layer2_outputs(7252));
    outputs(1350) <= not((layer2_outputs(3345)) xor (layer2_outputs(6341)));
    outputs(1351) <= (layer2_outputs(7658)) and not (layer2_outputs(7799));
    outputs(1352) <= (layer2_outputs(6595)) and (layer2_outputs(7746));
    outputs(1353) <= not((layer2_outputs(8024)) xor (layer2_outputs(3430)));
    outputs(1354) <= not(layer2_outputs(7311));
    outputs(1355) <= not(layer2_outputs(9500));
    outputs(1356) <= not(layer2_outputs(4788));
    outputs(1357) <= '0';
    outputs(1358) <= not((layer2_outputs(7022)) or (layer2_outputs(3731)));
    outputs(1359) <= not(layer2_outputs(542));
    outputs(1360) <= not(layer2_outputs(3062));
    outputs(1361) <= layer2_outputs(6381);
    outputs(1362) <= layer2_outputs(3871);
    outputs(1363) <= (layer2_outputs(2368)) xor (layer2_outputs(3883));
    outputs(1364) <= (layer2_outputs(7155)) xor (layer2_outputs(4490));
    outputs(1365) <= (layer2_outputs(2000)) xor (layer2_outputs(9475));
    outputs(1366) <= '0';
    outputs(1367) <= (layer2_outputs(5473)) and (layer2_outputs(3198));
    outputs(1368) <= layer2_outputs(3723);
    outputs(1369) <= not(layer2_outputs(6894));
    outputs(1370) <= layer2_outputs(6272);
    outputs(1371) <= layer2_outputs(3862);
    outputs(1372) <= not((layer2_outputs(5600)) xor (layer2_outputs(8489)));
    outputs(1373) <= not(layer2_outputs(5286));
    outputs(1374) <= (layer2_outputs(2274)) and not (layer2_outputs(4150));
    outputs(1375) <= (layer2_outputs(2125)) and (layer2_outputs(7661));
    outputs(1376) <= (layer2_outputs(5259)) and not (layer2_outputs(3674));
    outputs(1377) <= (layer2_outputs(287)) and (layer2_outputs(5396));
    outputs(1378) <= not(layer2_outputs(3801));
    outputs(1379) <= (layer2_outputs(4962)) and (layer2_outputs(8857));
    outputs(1380) <= (layer2_outputs(3612)) and not (layer2_outputs(6650));
    outputs(1381) <= not((layer2_outputs(8223)) xor (layer2_outputs(9459)));
    outputs(1382) <= (layer2_outputs(7100)) and not (layer2_outputs(8070));
    outputs(1383) <= (layer2_outputs(8000)) and (layer2_outputs(5301));
    outputs(1384) <= not((layer2_outputs(205)) or (layer2_outputs(4942)));
    outputs(1385) <= not((layer2_outputs(1105)) or (layer2_outputs(991)));
    outputs(1386) <= layer2_outputs(7373);
    outputs(1387) <= (layer2_outputs(8262)) xor (layer2_outputs(3490));
    outputs(1388) <= not((layer2_outputs(8504)) xor (layer2_outputs(3701)));
    outputs(1389) <= layer2_outputs(4101);
    outputs(1390) <= layer2_outputs(7846);
    outputs(1391) <= not((layer2_outputs(2841)) or (layer2_outputs(3751)));
    outputs(1392) <= (layer2_outputs(5724)) and not (layer2_outputs(8756));
    outputs(1393) <= not(layer2_outputs(6242));
    outputs(1394) <= not(layer2_outputs(243));
    outputs(1395) <= not(layer2_outputs(1253));
    outputs(1396) <= not(layer2_outputs(7625));
    outputs(1397) <= (layer2_outputs(9643)) and not (layer2_outputs(5108));
    outputs(1398) <= (layer2_outputs(1052)) and (layer2_outputs(9011));
    outputs(1399) <= layer2_outputs(7750);
    outputs(1400) <= layer2_outputs(9505);
    outputs(1401) <= layer2_outputs(9335);
    outputs(1402) <= not((layer2_outputs(405)) or (layer2_outputs(6513)));
    outputs(1403) <= layer2_outputs(5118);
    outputs(1404) <= (layer2_outputs(1199)) and not (layer2_outputs(5411));
    outputs(1405) <= not(layer2_outputs(2909));
    outputs(1406) <= (layer2_outputs(10005)) and (layer2_outputs(262));
    outputs(1407) <= not(layer2_outputs(3493));
    outputs(1408) <= not(layer2_outputs(2771)) or (layer2_outputs(1621));
    outputs(1409) <= not((layer2_outputs(9742)) xor (layer2_outputs(2545)));
    outputs(1410) <= (layer2_outputs(4510)) and not (layer2_outputs(5132));
    outputs(1411) <= layer2_outputs(3137);
    outputs(1412) <= not((layer2_outputs(4567)) or (layer2_outputs(2923)));
    outputs(1413) <= not((layer2_outputs(760)) xor (layer2_outputs(2885)));
    outputs(1414) <= (layer2_outputs(891)) and not (layer2_outputs(1739));
    outputs(1415) <= (layer2_outputs(9983)) and (layer2_outputs(303));
    outputs(1416) <= layer2_outputs(3671);
    outputs(1417) <= not((layer2_outputs(9065)) xor (layer2_outputs(2318)));
    outputs(1418) <= not(layer2_outputs(5492));
    outputs(1419) <= (layer2_outputs(5952)) xor (layer2_outputs(2377));
    outputs(1420) <= not((layer2_outputs(5828)) xor (layer2_outputs(2970)));
    outputs(1421) <= not(layer2_outputs(2119));
    outputs(1422) <= layer2_outputs(4624);
    outputs(1423) <= not(layer2_outputs(9238));
    outputs(1424) <= layer2_outputs(9399);
    outputs(1425) <= not((layer2_outputs(5371)) xor (layer2_outputs(8963)));
    outputs(1426) <= layer2_outputs(3680);
    outputs(1427) <= not(layer2_outputs(9910));
    outputs(1428) <= (layer2_outputs(6990)) and not (layer2_outputs(93));
    outputs(1429) <= not(layer2_outputs(2470));
    outputs(1430) <= layer2_outputs(5464);
    outputs(1431) <= layer2_outputs(7082);
    outputs(1432) <= not((layer2_outputs(7285)) xor (layer2_outputs(8719)));
    outputs(1433) <= not(layer2_outputs(7906));
    outputs(1434) <= (layer2_outputs(9018)) and not (layer2_outputs(407));
    outputs(1435) <= (layer2_outputs(3269)) and (layer2_outputs(4));
    outputs(1436) <= (layer2_outputs(2233)) or (layer2_outputs(2409));
    outputs(1437) <= not(layer2_outputs(6238));
    outputs(1438) <= (layer2_outputs(284)) and not (layer2_outputs(8588));
    outputs(1439) <= layer2_outputs(1984);
    outputs(1440) <= not(layer2_outputs(5593));
    outputs(1441) <= (layer2_outputs(9267)) and not (layer2_outputs(1026));
    outputs(1442) <= not(layer2_outputs(462));
    outputs(1443) <= layer2_outputs(10210);
    outputs(1444) <= (layer2_outputs(4883)) and not (layer2_outputs(9177));
    outputs(1445) <= layer2_outputs(4316);
    outputs(1446) <= (layer2_outputs(1377)) xor (layer2_outputs(7882));
    outputs(1447) <= not((layer2_outputs(4292)) xor (layer2_outputs(1194)));
    outputs(1448) <= (layer2_outputs(5173)) xor (layer2_outputs(206));
    outputs(1449) <= not((layer2_outputs(2708)) and (layer2_outputs(3764)));
    outputs(1450) <= (layer2_outputs(1243)) and (layer2_outputs(3907));
    outputs(1451) <= (layer2_outputs(4340)) and not (layer2_outputs(8707));
    outputs(1452) <= not(layer2_outputs(8485));
    outputs(1453) <= not(layer2_outputs(5769));
    outputs(1454) <= not((layer2_outputs(9057)) or (layer2_outputs(9488)));
    outputs(1455) <= not(layer2_outputs(7963));
    outputs(1456) <= (layer2_outputs(8242)) xor (layer2_outputs(660));
    outputs(1457) <= (layer2_outputs(137)) or (layer2_outputs(3968));
    outputs(1458) <= not(layer2_outputs(1824));
    outputs(1459) <= layer2_outputs(2532);
    outputs(1460) <= (layer2_outputs(8758)) xor (layer2_outputs(8298));
    outputs(1461) <= (layer2_outputs(583)) and not (layer2_outputs(7479));
    outputs(1462) <= not((layer2_outputs(10007)) xor (layer2_outputs(6032)));
    outputs(1463) <= not(layer2_outputs(3375));
    outputs(1464) <= (layer2_outputs(611)) xor (layer2_outputs(1033));
    outputs(1465) <= not(layer2_outputs(1899));
    outputs(1466) <= (layer2_outputs(9285)) and not (layer2_outputs(8868));
    outputs(1467) <= (layer2_outputs(7686)) xor (layer2_outputs(1083));
    outputs(1468) <= (layer2_outputs(7011)) and (layer2_outputs(4695));
    outputs(1469) <= not(layer2_outputs(2219));
    outputs(1470) <= not(layer2_outputs(2435));
    outputs(1471) <= not(layer2_outputs(4945));
    outputs(1472) <= not((layer2_outputs(3516)) xor (layer2_outputs(868)));
    outputs(1473) <= not((layer2_outputs(2308)) xor (layer2_outputs(4192)));
    outputs(1474) <= layer2_outputs(7529);
    outputs(1475) <= layer2_outputs(3626);
    outputs(1476) <= (layer2_outputs(9119)) and not (layer2_outputs(7213));
    outputs(1477) <= not(layer2_outputs(1610));
    outputs(1478) <= not(layer2_outputs(9795));
    outputs(1479) <= layer2_outputs(6603);
    outputs(1480) <= not(layer2_outputs(2216));
    outputs(1481) <= not(layer2_outputs(2123)) or (layer2_outputs(3683));
    outputs(1482) <= (layer2_outputs(8022)) xor (layer2_outputs(9416));
    outputs(1483) <= (layer2_outputs(4185)) or (layer2_outputs(3494));
    outputs(1484) <= not(layer2_outputs(1022));
    outputs(1485) <= layer2_outputs(5666);
    outputs(1486) <= (layer2_outputs(6805)) and not (layer2_outputs(9847));
    outputs(1487) <= (layer2_outputs(4871)) xor (layer2_outputs(3653));
    outputs(1488) <= not(layer2_outputs(2963));
    outputs(1489) <= not((layer2_outputs(3216)) xor (layer2_outputs(7752)));
    outputs(1490) <= not(layer2_outputs(6920));
    outputs(1491) <= not(layer2_outputs(1257));
    outputs(1492) <= (layer2_outputs(4922)) and not (layer2_outputs(9266));
    outputs(1493) <= not((layer2_outputs(4686)) or (layer2_outputs(8143)));
    outputs(1494) <= layer2_outputs(9151);
    outputs(1495) <= not(layer2_outputs(2086));
    outputs(1496) <= not(layer2_outputs(5292));
    outputs(1497) <= (layer2_outputs(5818)) xor (layer2_outputs(6340));
    outputs(1498) <= not(layer2_outputs(4636));
    outputs(1499) <= (layer2_outputs(10216)) and (layer2_outputs(7234));
    outputs(1500) <= not((layer2_outputs(636)) or (layer2_outputs(2070)));
    outputs(1501) <= not(layer2_outputs(9006));
    outputs(1502) <= (layer2_outputs(9560)) or (layer2_outputs(1795));
    outputs(1503) <= (layer2_outputs(5599)) and (layer2_outputs(3368));
    outputs(1504) <= not((layer2_outputs(7598)) xor (layer2_outputs(8939)));
    outputs(1505) <= layer2_outputs(6982);
    outputs(1506) <= not(layer2_outputs(7599));
    outputs(1507) <= layer2_outputs(2997);
    outputs(1508) <= (layer2_outputs(2376)) xor (layer2_outputs(4482));
    outputs(1509) <= (layer2_outputs(6371)) and not (layer2_outputs(2983));
    outputs(1510) <= (layer2_outputs(5424)) and not (layer2_outputs(1008));
    outputs(1511) <= (layer2_outputs(2892)) xor (layer2_outputs(8162));
    outputs(1512) <= not((layer2_outputs(9427)) or (layer2_outputs(6339)));
    outputs(1513) <= (layer2_outputs(7446)) xor (layer2_outputs(6568));
    outputs(1514) <= layer2_outputs(4589);
    outputs(1515) <= not((layer2_outputs(6880)) or (layer2_outputs(6988)));
    outputs(1516) <= (layer2_outputs(7813)) and not (layer2_outputs(10052));
    outputs(1517) <= layer2_outputs(7082);
    outputs(1518) <= not((layer2_outputs(7983)) xor (layer2_outputs(5779)));
    outputs(1519) <= layer2_outputs(1937);
    outputs(1520) <= not((layer2_outputs(6722)) xor (layer2_outputs(9760)));
    outputs(1521) <= not(layer2_outputs(4682));
    outputs(1522) <= not(layer2_outputs(5141));
    outputs(1523) <= layer2_outputs(3313);
    outputs(1524) <= not(layer2_outputs(7752));
    outputs(1525) <= layer2_outputs(3227);
    outputs(1526) <= (layer2_outputs(2543)) xor (layer2_outputs(2629));
    outputs(1527) <= not((layer2_outputs(3513)) xor (layer2_outputs(2024)));
    outputs(1528) <= (layer2_outputs(6722)) xor (layer2_outputs(4778));
    outputs(1529) <= (layer2_outputs(4350)) and not (layer2_outputs(6715));
    outputs(1530) <= layer2_outputs(6405);
    outputs(1531) <= layer2_outputs(4295);
    outputs(1532) <= not(layer2_outputs(345));
    outputs(1533) <= not(layer2_outputs(2851));
    outputs(1534) <= not(layer2_outputs(42));
    outputs(1535) <= not(layer2_outputs(9795));
    outputs(1536) <= (layer2_outputs(8713)) xor (layer2_outputs(323));
    outputs(1537) <= layer2_outputs(2481);
    outputs(1538) <= not((layer2_outputs(9349)) xor (layer2_outputs(675)));
    outputs(1539) <= layer2_outputs(9237);
    outputs(1540) <= layer2_outputs(5200);
    outputs(1541) <= (layer2_outputs(3767)) xor (layer2_outputs(6635));
    outputs(1542) <= not(layer2_outputs(5226));
    outputs(1543) <= (layer2_outputs(5056)) and (layer2_outputs(10062));
    outputs(1544) <= layer2_outputs(5577);
    outputs(1545) <= not((layer2_outputs(56)) xor (layer2_outputs(8438)));
    outputs(1546) <= not((layer2_outputs(4298)) xor (layer2_outputs(1106)));
    outputs(1547) <= not(layer2_outputs(5031));
    outputs(1548) <= (layer2_outputs(936)) and not (layer2_outputs(8713));
    outputs(1549) <= (layer2_outputs(8454)) and not (layer2_outputs(6264));
    outputs(1550) <= not(layer2_outputs(9508));
    outputs(1551) <= layer2_outputs(8118);
    outputs(1552) <= (layer2_outputs(4293)) and (layer2_outputs(6114));
    outputs(1553) <= layer2_outputs(10133);
    outputs(1554) <= not(layer2_outputs(4174));
    outputs(1555) <= not((layer2_outputs(1789)) or (layer2_outputs(9296)));
    outputs(1556) <= (layer2_outputs(5474)) and (layer2_outputs(8814));
    outputs(1557) <= not(layer2_outputs(3128));
    outputs(1558) <= (layer2_outputs(8349)) xor (layer2_outputs(9222));
    outputs(1559) <= not(layer2_outputs(1989));
    outputs(1560) <= (layer2_outputs(1131)) and not (layer2_outputs(10195));
    outputs(1561) <= (layer2_outputs(76)) xor (layer2_outputs(2708));
    outputs(1562) <= (layer2_outputs(6068)) and not (layer2_outputs(8065));
    outputs(1563) <= layer2_outputs(10057);
    outputs(1564) <= not((layer2_outputs(5321)) xor (layer2_outputs(1517)));
    outputs(1565) <= not(layer2_outputs(6907));
    outputs(1566) <= (layer2_outputs(4602)) xor (layer2_outputs(7945));
    outputs(1567) <= not(layer2_outputs(833));
    outputs(1568) <= (layer2_outputs(4340)) xor (layer2_outputs(4643));
    outputs(1569) <= (layer2_outputs(6467)) and not (layer2_outputs(10180));
    outputs(1570) <= (layer2_outputs(7186)) and not (layer2_outputs(1568));
    outputs(1571) <= not((layer2_outputs(6226)) xor (layer2_outputs(60)));
    outputs(1572) <= not((layer2_outputs(3010)) xor (layer2_outputs(7080)));
    outputs(1573) <= (layer2_outputs(6538)) and (layer2_outputs(6568));
    outputs(1574) <= layer2_outputs(9505);
    outputs(1575) <= not((layer2_outputs(9976)) or (layer2_outputs(734)));
    outputs(1576) <= layer2_outputs(388);
    outputs(1577) <= not(layer2_outputs(3647));
    outputs(1578) <= (layer2_outputs(6255)) or (layer2_outputs(7515));
    outputs(1579) <= (layer2_outputs(9900)) xor (layer2_outputs(4415));
    outputs(1580) <= not(layer2_outputs(4432));
    outputs(1581) <= layer2_outputs(186);
    outputs(1582) <= not((layer2_outputs(4536)) or (layer2_outputs(8422)));
    outputs(1583) <= layer2_outputs(9663);
    outputs(1584) <= not(layer2_outputs(7530));
    outputs(1585) <= not(layer2_outputs(6283));
    outputs(1586) <= (layer2_outputs(6814)) and not (layer2_outputs(8120));
    outputs(1587) <= not(layer2_outputs(1022));
    outputs(1588) <= (layer2_outputs(1745)) xor (layer2_outputs(9656));
    outputs(1589) <= not((layer2_outputs(5218)) or (layer2_outputs(8536)));
    outputs(1590) <= (layer2_outputs(1605)) and not (layer2_outputs(6055));
    outputs(1591) <= layer2_outputs(8855);
    outputs(1592) <= not((layer2_outputs(1024)) xor (layer2_outputs(8265)));
    outputs(1593) <= not(layer2_outputs(6705));
    outputs(1594) <= not((layer2_outputs(9908)) xor (layer2_outputs(8709)));
    outputs(1595) <= layer2_outputs(9021);
    outputs(1596) <= not(layer2_outputs(5346));
    outputs(1597) <= (layer2_outputs(4932)) and (layer2_outputs(8477));
    outputs(1598) <= not((layer2_outputs(9486)) xor (layer2_outputs(3718)));
    outputs(1599) <= not((layer2_outputs(4886)) xor (layer2_outputs(5729)));
    outputs(1600) <= (layer2_outputs(2425)) xor (layer2_outputs(1587));
    outputs(1601) <= layer2_outputs(2690);
    outputs(1602) <= not(layer2_outputs(7640));
    outputs(1603) <= not((layer2_outputs(3063)) or (layer2_outputs(6111)));
    outputs(1604) <= (layer2_outputs(4798)) and not (layer2_outputs(7791));
    outputs(1605) <= (layer2_outputs(3601)) and not (layer2_outputs(9028));
    outputs(1606) <= layer2_outputs(3255);
    outputs(1607) <= not((layer2_outputs(7507)) or (layer2_outputs(294)));
    outputs(1608) <= (layer2_outputs(6649)) and (layer2_outputs(2504));
    outputs(1609) <= (layer2_outputs(6050)) and not (layer2_outputs(7075));
    outputs(1610) <= not((layer2_outputs(4384)) or (layer2_outputs(6775)));
    outputs(1611) <= (layer2_outputs(4707)) and not (layer2_outputs(5294));
    outputs(1612) <= not(layer2_outputs(6588));
    outputs(1613) <= not((layer2_outputs(7960)) or (layer2_outputs(8544)));
    outputs(1614) <= not((layer2_outputs(3364)) xor (layer2_outputs(692)));
    outputs(1615) <= not((layer2_outputs(8248)) xor (layer2_outputs(4891)));
    outputs(1616) <= layer2_outputs(6147);
    outputs(1617) <= (layer2_outputs(9626)) and (layer2_outputs(1515));
    outputs(1618) <= not(layer2_outputs(4646));
    outputs(1619) <= not(layer2_outputs(5617));
    outputs(1620) <= not(layer2_outputs(1023));
    outputs(1621) <= not(layer2_outputs(3308));
    outputs(1622) <= (layer2_outputs(8702)) xor (layer2_outputs(4082));
    outputs(1623) <= not(layer2_outputs(3647));
    outputs(1624) <= layer2_outputs(488);
    outputs(1625) <= not(layer2_outputs(3588));
    outputs(1626) <= (layer2_outputs(9546)) xor (layer2_outputs(650));
    outputs(1627) <= (layer2_outputs(6397)) or (layer2_outputs(9763));
    outputs(1628) <= (layer2_outputs(819)) xor (layer2_outputs(3082));
    outputs(1629) <= not(layer2_outputs(9154));
    outputs(1630) <= not(layer2_outputs(3993));
    outputs(1631) <= not(layer2_outputs(6091));
    outputs(1632) <= not(layer2_outputs(1415));
    outputs(1633) <= not(layer2_outputs(6875));
    outputs(1634) <= not(layer2_outputs(5380));
    outputs(1635) <= not((layer2_outputs(2331)) or (layer2_outputs(1354)));
    outputs(1636) <= not(layer2_outputs(8956));
    outputs(1637) <= not((layer2_outputs(5930)) xor (layer2_outputs(10136)));
    outputs(1638) <= layer2_outputs(5880);
    outputs(1639) <= not(layer2_outputs(9097));
    outputs(1640) <= not(layer2_outputs(4992));
    outputs(1641) <= (layer2_outputs(621)) xor (layer2_outputs(1259));
    outputs(1642) <= not((layer2_outputs(2118)) and (layer2_outputs(4706)));
    outputs(1643) <= layer2_outputs(820);
    outputs(1644) <= not(layer2_outputs(6555));
    outputs(1645) <= not(layer2_outputs(196));
    outputs(1646) <= (layer2_outputs(6867)) and (layer2_outputs(7943));
    outputs(1647) <= (layer2_outputs(5025)) and not (layer2_outputs(727));
    outputs(1648) <= layer2_outputs(9352);
    outputs(1649) <= layer2_outputs(1199);
    outputs(1650) <= layer2_outputs(1066);
    outputs(1651) <= (layer2_outputs(3842)) xor (layer2_outputs(9905));
    outputs(1652) <= not((layer2_outputs(4752)) or (layer2_outputs(4131)));
    outputs(1653) <= layer2_outputs(8212);
    outputs(1654) <= not((layer2_outputs(1764)) or (layer2_outputs(7422)));
    outputs(1655) <= not((layer2_outputs(8318)) or (layer2_outputs(4170)));
    outputs(1656) <= not(layer2_outputs(5457)) or (layer2_outputs(459));
    outputs(1657) <= not(layer2_outputs(3876));
    outputs(1658) <= layer2_outputs(4586);
    outputs(1659) <= (layer2_outputs(6489)) and (layer2_outputs(8765));
    outputs(1660) <= not(layer2_outputs(1493));
    outputs(1661) <= not(layer2_outputs(8142));
    outputs(1662) <= not(layer2_outputs(8564));
    outputs(1663) <= layer2_outputs(2779);
    outputs(1664) <= not(layer2_outputs(1102));
    outputs(1665) <= (layer2_outputs(8916)) and (layer2_outputs(5570));
    outputs(1666) <= not(layer2_outputs(3946));
    outputs(1667) <= layer2_outputs(2126);
    outputs(1668) <= not(layer2_outputs(7873));
    outputs(1669) <= (layer2_outputs(1270)) and not (layer2_outputs(7187));
    outputs(1670) <= not((layer2_outputs(3064)) xor (layer2_outputs(9551)));
    outputs(1671) <= layer2_outputs(8334);
    outputs(1672) <= not((layer2_outputs(7242)) xor (layer2_outputs(407)));
    outputs(1673) <= layer2_outputs(148);
    outputs(1674) <= layer2_outputs(7138);
    outputs(1675) <= not(layer2_outputs(7387));
    outputs(1676) <= not(layer2_outputs(9527));
    outputs(1677) <= '0';
    outputs(1678) <= not(layer2_outputs(3690));
    outputs(1679) <= not(layer2_outputs(3898));
    outputs(1680) <= (layer2_outputs(4678)) and not (layer2_outputs(9301));
    outputs(1681) <= not((layer2_outputs(593)) xor (layer2_outputs(6554)));
    outputs(1682) <= not((layer2_outputs(3730)) or (layer2_outputs(759)));
    outputs(1683) <= (layer2_outputs(3009)) and (layer2_outputs(7333));
    outputs(1684) <= layer2_outputs(4518);
    outputs(1685) <= not(layer2_outputs(7817)) or (layer2_outputs(5774));
    outputs(1686) <= not((layer2_outputs(1856)) xor (layer2_outputs(2387)));
    outputs(1687) <= not((layer2_outputs(7412)) xor (layer2_outputs(5772)));
    outputs(1688) <= layer2_outputs(5899);
    outputs(1689) <= layer2_outputs(3448);
    outputs(1690) <= not(layer2_outputs(1053));
    outputs(1691) <= (layer2_outputs(9000)) and (layer2_outputs(5314));
    outputs(1692) <= not((layer2_outputs(8378)) or (layer2_outputs(7301)));
    outputs(1693) <= not(layer2_outputs(1319)) or (layer2_outputs(2696));
    outputs(1694) <= layer2_outputs(5441);
    outputs(1695) <= not(layer2_outputs(4188));
    outputs(1696) <= (layer2_outputs(2913)) xor (layer2_outputs(4280));
    outputs(1697) <= not(layer2_outputs(2305));
    outputs(1698) <= not((layer2_outputs(3111)) xor (layer2_outputs(3713)));
    outputs(1699) <= (layer2_outputs(7735)) xor (layer2_outputs(8345));
    outputs(1700) <= layer2_outputs(127);
    outputs(1701) <= (layer2_outputs(2868)) and not (layer2_outputs(39));
    outputs(1702) <= (layer2_outputs(6312)) and (layer2_outputs(7935));
    outputs(1703) <= not((layer2_outputs(8335)) xor (layer2_outputs(2942)));
    outputs(1704) <= not((layer2_outputs(2585)) xor (layer2_outputs(3507)));
    outputs(1705) <= layer2_outputs(5592);
    outputs(1706) <= not(layer2_outputs(887));
    outputs(1707) <= not(layer2_outputs(8217));
    outputs(1708) <= layer2_outputs(9098);
    outputs(1709) <= layer2_outputs(9370);
    outputs(1710) <= not(layer2_outputs(8322));
    outputs(1711) <= not(layer2_outputs(1137));
    outputs(1712) <= (layer2_outputs(5948)) or (layer2_outputs(7745));
    outputs(1713) <= not((layer2_outputs(64)) xor (layer2_outputs(8085)));
    outputs(1714) <= not((layer2_outputs(149)) or (layer2_outputs(7982)));
    outputs(1715) <= not((layer2_outputs(8786)) xor (layer2_outputs(8286)));
    outputs(1716) <= not(layer2_outputs(4230));
    outputs(1717) <= (layer2_outputs(4203)) and not (layer2_outputs(3046));
    outputs(1718) <= (layer2_outputs(7954)) xor (layer2_outputs(2569));
    outputs(1719) <= not((layer2_outputs(9717)) xor (layer2_outputs(3417)));
    outputs(1720) <= not(layer2_outputs(8609));
    outputs(1721) <= layer2_outputs(7381);
    outputs(1722) <= not(layer2_outputs(9115));
    outputs(1723) <= not(layer2_outputs(9830));
    outputs(1724) <= not(layer2_outputs(9433));
    outputs(1725) <= not(layer2_outputs(7116));
    outputs(1726) <= not(layer2_outputs(782));
    outputs(1727) <= not((layer2_outputs(630)) or (layer2_outputs(1745)));
    outputs(1728) <= layer2_outputs(9201);
    outputs(1729) <= layer2_outputs(2229);
    outputs(1730) <= not((layer2_outputs(239)) or (layer2_outputs(9991)));
    outputs(1731) <= layer2_outputs(5026);
    outputs(1732) <= not(layer2_outputs(625));
    outputs(1733) <= not(layer2_outputs(293)) or (layer2_outputs(8532));
    outputs(1734) <= not(layer2_outputs(9165));
    outputs(1735) <= not(layer2_outputs(8435));
    outputs(1736) <= not(layer2_outputs(341));
    outputs(1737) <= not(layer2_outputs(68));
    outputs(1738) <= (layer2_outputs(8211)) and not (layer2_outputs(7838));
    outputs(1739) <= not(layer2_outputs(9320));
    outputs(1740) <= layer2_outputs(1974);
    outputs(1741) <= (layer2_outputs(10156)) and not (layer2_outputs(5086));
    outputs(1742) <= layer2_outputs(6437);
    outputs(1743) <= (layer2_outputs(2287)) xor (layer2_outputs(3357));
    outputs(1744) <= not(layer2_outputs(6582)) or (layer2_outputs(1495));
    outputs(1745) <= not(layer2_outputs(3355));
    outputs(1746) <= not(layer2_outputs(8544));
    outputs(1747) <= not(layer2_outputs(3138));
    outputs(1748) <= not(layer2_outputs(8759));
    outputs(1749) <= layer2_outputs(2381);
    outputs(1750) <= layer2_outputs(3535);
    outputs(1751) <= layer2_outputs(3679);
    outputs(1752) <= (layer2_outputs(7382)) xor (layer2_outputs(1262));
    outputs(1753) <= not(layer2_outputs(4982));
    outputs(1754) <= not(layer2_outputs(7108));
    outputs(1755) <= not(layer2_outputs(2870)) or (layer2_outputs(3361));
    outputs(1756) <= not(layer2_outputs(2210));
    outputs(1757) <= (layer2_outputs(2941)) and not (layer2_outputs(1458));
    outputs(1758) <= (layer2_outputs(4696)) and not (layer2_outputs(4426));
    outputs(1759) <= (layer2_outputs(78)) and not (layer2_outputs(7054));
    outputs(1760) <= layer2_outputs(3628);
    outputs(1761) <= (layer2_outputs(1312)) and not (layer2_outputs(2327));
    outputs(1762) <= layer2_outputs(6845);
    outputs(1763) <= layer2_outputs(4374);
    outputs(1764) <= (layer2_outputs(2075)) xor (layer2_outputs(9202));
    outputs(1765) <= not(layer2_outputs(3806));
    outputs(1766) <= (layer2_outputs(10165)) and (layer2_outputs(1984));
    outputs(1767) <= not(layer2_outputs(2537));
    outputs(1768) <= layer2_outputs(4722);
    outputs(1769) <= (layer2_outputs(10164)) and not (layer2_outputs(2462));
    outputs(1770) <= (layer2_outputs(6211)) xor (layer2_outputs(3899));
    outputs(1771) <= not(layer2_outputs(5617));
    outputs(1772) <= not((layer2_outputs(3726)) or (layer2_outputs(1819)));
    outputs(1773) <= not((layer2_outputs(3696)) xor (layer2_outputs(6787)));
    outputs(1774) <= not((layer2_outputs(4206)) xor (layer2_outputs(2259)));
    outputs(1775) <= layer2_outputs(1710);
    outputs(1776) <= (layer2_outputs(3933)) and not (layer2_outputs(1163));
    outputs(1777) <= layer2_outputs(7122);
    outputs(1778) <= layer2_outputs(5692);
    outputs(1779) <= not(layer2_outputs(9516));
    outputs(1780) <= layer2_outputs(7505);
    outputs(1781) <= layer2_outputs(7063);
    outputs(1782) <= layer2_outputs(8067);
    outputs(1783) <= not((layer2_outputs(7302)) xor (layer2_outputs(10101)));
    outputs(1784) <= not((layer2_outputs(3025)) xor (layer2_outputs(3721)));
    outputs(1785) <= not((layer2_outputs(2149)) xor (layer2_outputs(7485)));
    outputs(1786) <= layer2_outputs(2904);
    outputs(1787) <= not((layer2_outputs(3222)) or (layer2_outputs(9840)));
    outputs(1788) <= (layer2_outputs(8035)) and not (layer2_outputs(3911));
    outputs(1789) <= layer2_outputs(4687);
    outputs(1790) <= not(layer2_outputs(1441));
    outputs(1791) <= not((layer2_outputs(4836)) xor (layer2_outputs(4831)));
    outputs(1792) <= not((layer2_outputs(2231)) xor (layer2_outputs(3771)));
    outputs(1793) <= not(layer2_outputs(9183));
    outputs(1794) <= layer2_outputs(7895);
    outputs(1795) <= layer2_outputs(5482);
    outputs(1796) <= not(layer2_outputs(3481));
    outputs(1797) <= not(layer2_outputs(9008));
    outputs(1798) <= not((layer2_outputs(899)) or (layer2_outputs(3640)));
    outputs(1799) <= not(layer2_outputs(8395));
    outputs(1800) <= not(layer2_outputs(3872));
    outputs(1801) <= layer2_outputs(7795);
    outputs(1802) <= not(layer2_outputs(1409));
    outputs(1803) <= (layer2_outputs(3082)) xor (layer2_outputs(1643));
    outputs(1804) <= (layer2_outputs(6275)) and not (layer2_outputs(6734));
    outputs(1805) <= not(layer2_outputs(404));
    outputs(1806) <= not(layer2_outputs(5253));
    outputs(1807) <= not(layer2_outputs(2412));
    outputs(1808) <= (layer2_outputs(9218)) and not (layer2_outputs(926));
    outputs(1809) <= not(layer2_outputs(2380));
    outputs(1810) <= not((layer2_outputs(3288)) xor (layer2_outputs(6946)));
    outputs(1811) <= layer2_outputs(4054);
    outputs(1812) <= (layer2_outputs(4484)) xor (layer2_outputs(9613));
    outputs(1813) <= not(layer2_outputs(4665));
    outputs(1814) <= (layer2_outputs(1399)) and (layer2_outputs(5862));
    outputs(1815) <= layer2_outputs(902);
    outputs(1816) <= layer2_outputs(9100);
    outputs(1817) <= not(layer2_outputs(3365));
    outputs(1818) <= layer2_outputs(1465);
    outputs(1819) <= layer2_outputs(7636);
    outputs(1820) <= not((layer2_outputs(6018)) xor (layer2_outputs(2125)));
    outputs(1821) <= layer2_outputs(9853);
    outputs(1822) <= (layer2_outputs(6772)) and (layer2_outputs(1167));
    outputs(1823) <= not(layer2_outputs(8434));
    outputs(1824) <= (layer2_outputs(9360)) and not (layer2_outputs(8774));
    outputs(1825) <= not(layer2_outputs(1765));
    outputs(1826) <= not(layer2_outputs(4450));
    outputs(1827) <= (layer2_outputs(3193)) xor (layer2_outputs(3596));
    outputs(1828) <= not(layer2_outputs(9738));
    outputs(1829) <= layer2_outputs(3422);
    outputs(1830) <= (layer2_outputs(2996)) xor (layer2_outputs(1277));
    outputs(1831) <= not(layer2_outputs(3852));
    outputs(1832) <= layer2_outputs(6460);
    outputs(1833) <= not((layer2_outputs(8040)) xor (layer2_outputs(308)));
    outputs(1834) <= layer2_outputs(6620);
    outputs(1835) <= not(layer2_outputs(5348));
    outputs(1836) <= not(layer2_outputs(7216));
    outputs(1837) <= not((layer2_outputs(5895)) xor (layer2_outputs(8016)));
    outputs(1838) <= not(layer2_outputs(4281));
    outputs(1839) <= not(layer2_outputs(7398));
    outputs(1840) <= layer2_outputs(9873);
    outputs(1841) <= layer2_outputs(4749);
    outputs(1842) <= '0';
    outputs(1843) <= (layer2_outputs(4828)) and (layer2_outputs(3612));
    outputs(1844) <= (layer2_outputs(4959)) and not (layer2_outputs(4644));
    outputs(1845) <= (layer2_outputs(3187)) and not (layer2_outputs(5712));
    outputs(1846) <= not(layer2_outputs(4161));
    outputs(1847) <= layer2_outputs(4139);
    outputs(1848) <= (layer2_outputs(3308)) xor (layer2_outputs(6940));
    outputs(1849) <= (layer2_outputs(9452)) and not (layer2_outputs(8627));
    outputs(1850) <= (layer2_outputs(9454)) and (layer2_outputs(3215));
    outputs(1851) <= not((layer2_outputs(6294)) or (layer2_outputs(6868)));
    outputs(1852) <= layer2_outputs(2580);
    outputs(1853) <= not((layer2_outputs(3883)) xor (layer2_outputs(6071)));
    outputs(1854) <= (layer2_outputs(6438)) xor (layer2_outputs(6711));
    outputs(1855) <= (layer2_outputs(1067)) and not (layer2_outputs(1796));
    outputs(1856) <= not(layer2_outputs(5831));
    outputs(1857) <= layer2_outputs(8077);
    outputs(1858) <= not(layer2_outputs(494));
    outputs(1859) <= (layer2_outputs(5438)) xor (layer2_outputs(2178));
    outputs(1860) <= (layer2_outputs(9408)) and (layer2_outputs(6122));
    outputs(1861) <= (layer2_outputs(7821)) and not (layer2_outputs(7459));
    outputs(1862) <= not(layer2_outputs(1287));
    outputs(1863) <= not(layer2_outputs(7533));
    outputs(1864) <= layer2_outputs(3791);
    outputs(1865) <= not((layer2_outputs(5331)) xor (layer2_outputs(4373)));
    outputs(1866) <= layer2_outputs(3893);
    outputs(1867) <= layer2_outputs(7807);
    outputs(1868) <= not((layer2_outputs(3762)) or (layer2_outputs(4494)));
    outputs(1869) <= layer2_outputs(9837);
    outputs(1870) <= layer2_outputs(638);
    outputs(1871) <= layer2_outputs(7858);
    outputs(1872) <= layer2_outputs(6353);
    outputs(1873) <= not(layer2_outputs(8005));
    outputs(1874) <= (layer2_outputs(5115)) xor (layer2_outputs(3058));
    outputs(1875) <= not((layer2_outputs(6039)) or (layer2_outputs(8996)));
    outputs(1876) <= not(layer2_outputs(2647));
    outputs(1877) <= not((layer2_outputs(3364)) xor (layer2_outputs(4166)));
    outputs(1878) <= layer2_outputs(3779);
    outputs(1879) <= layer2_outputs(10114);
    outputs(1880) <= (layer2_outputs(2004)) and not (layer2_outputs(8346));
    outputs(1881) <= (layer2_outputs(3104)) and not (layer2_outputs(8292));
    outputs(1882) <= (layer2_outputs(338)) xor (layer2_outputs(2309));
    outputs(1883) <= not((layer2_outputs(9226)) xor (layer2_outputs(3059)));
    outputs(1884) <= (layer2_outputs(6678)) and not (layer2_outputs(5874));
    outputs(1885) <= not((layer2_outputs(3267)) or (layer2_outputs(3152)));
    outputs(1886) <= layer2_outputs(1450);
    outputs(1887) <= layer2_outputs(8437);
    outputs(1888) <= not(layer2_outputs(6320));
    outputs(1889) <= (layer2_outputs(2752)) and (layer2_outputs(649));
    outputs(1890) <= not((layer2_outputs(9170)) xor (layer2_outputs(1210)));
    outputs(1891) <= layer2_outputs(1425);
    outputs(1892) <= not((layer2_outputs(6447)) or (layer2_outputs(3936)));
    outputs(1893) <= layer2_outputs(7506);
    outputs(1894) <= not((layer2_outputs(2765)) or (layer2_outputs(3416)));
    outputs(1895) <= (layer2_outputs(451)) and (layer2_outputs(9382));
    outputs(1896) <= layer2_outputs(5790);
    outputs(1897) <= layer2_outputs(6268);
    outputs(1898) <= (layer2_outputs(2498)) and (layer2_outputs(761));
    outputs(1899) <= (layer2_outputs(7437)) and not (layer2_outputs(6837));
    outputs(1900) <= not(layer2_outputs(2026));
    outputs(1901) <= not(layer2_outputs(8242));
    outputs(1902) <= not(layer2_outputs(4296));
    outputs(1903) <= '0';
    outputs(1904) <= not(layer2_outputs(3028));
    outputs(1905) <= layer2_outputs(9544);
    outputs(1906) <= (layer2_outputs(4036)) and not (layer2_outputs(6688));
    outputs(1907) <= (layer2_outputs(4944)) or (layer2_outputs(2682));
    outputs(1908) <= layer2_outputs(7225);
    outputs(1909) <= (layer2_outputs(7779)) xor (layer2_outputs(4381));
    outputs(1910) <= (layer2_outputs(438)) xor (layer2_outputs(4621));
    outputs(1911) <= layer2_outputs(7652);
    outputs(1912) <= layer2_outputs(9287);
    outputs(1913) <= (layer2_outputs(4506)) and (layer2_outputs(9083));
    outputs(1914) <= not(layer2_outputs(8015));
    outputs(1915) <= not(layer2_outputs(1958));
    outputs(1916) <= (layer2_outputs(9525)) and not (layer2_outputs(4193));
    outputs(1917) <= not((layer2_outputs(7377)) xor (layer2_outputs(3465)));
    outputs(1918) <= not(layer2_outputs(6136));
    outputs(1919) <= (layer2_outputs(9628)) xor (layer2_outputs(935));
    outputs(1920) <= (layer2_outputs(6723)) and (layer2_outputs(9856));
    outputs(1921) <= layer2_outputs(9483);
    outputs(1922) <= not((layer2_outputs(6637)) xor (layer2_outputs(6653)));
    outputs(1923) <= (layer2_outputs(7038)) xor (layer2_outputs(1086));
    outputs(1924) <= (layer2_outputs(7052)) and (layer2_outputs(3965));
    outputs(1925) <= not((layer2_outputs(6638)) xor (layer2_outputs(7207)));
    outputs(1926) <= layer2_outputs(3910);
    outputs(1927) <= layer2_outputs(4240);
    outputs(1928) <= (layer2_outputs(5559)) and not (layer2_outputs(6371));
    outputs(1929) <= layer2_outputs(7704);
    outputs(1930) <= (layer2_outputs(337)) or (layer2_outputs(1767));
    outputs(1931) <= not((layer2_outputs(3108)) or (layer2_outputs(2395)));
    outputs(1932) <= layer2_outputs(5333);
    outputs(1933) <= not(layer2_outputs(5294));
    outputs(1934) <= not(layer2_outputs(9991));
    outputs(1935) <= not(layer2_outputs(4807));
    outputs(1936) <= (layer2_outputs(4516)) and not (layer2_outputs(7297));
    outputs(1937) <= (layer2_outputs(8748)) and not (layer2_outputs(3610));
    outputs(1938) <= (layer2_outputs(549)) or (layer2_outputs(1145));
    outputs(1939) <= (layer2_outputs(6485)) and not (layer2_outputs(1127));
    outputs(1940) <= (layer2_outputs(6252)) and (layer2_outputs(6108));
    outputs(1941) <= (layer2_outputs(4632)) xor (layer2_outputs(345));
    outputs(1942) <= not(layer2_outputs(8983));
    outputs(1943) <= not(layer2_outputs(183));
    outputs(1944) <= (layer2_outputs(9669)) and (layer2_outputs(8954));
    outputs(1945) <= not(layer2_outputs(198));
    outputs(1946) <= not(layer2_outputs(3231));
    outputs(1947) <= (layer2_outputs(6013)) and not (layer2_outputs(2608));
    outputs(1948) <= not(layer2_outputs(1140));
    outputs(1949) <= (layer2_outputs(8054)) xor (layer2_outputs(6482));
    outputs(1950) <= layer2_outputs(7087);
    outputs(1951) <= not(layer2_outputs(6885));
    outputs(1952) <= not(layer2_outputs(850));
    outputs(1953) <= layer2_outputs(8134);
    outputs(1954) <= not(layer2_outputs(2554));
    outputs(1955) <= not(layer2_outputs(8948));
    outputs(1956) <= layer2_outputs(8189);
    outputs(1957) <= not((layer2_outputs(1617)) or (layer2_outputs(1082)));
    outputs(1958) <= (layer2_outputs(9768)) and not (layer2_outputs(6286));
    outputs(1959) <= not((layer2_outputs(47)) and (layer2_outputs(6402)));
    outputs(1960) <= not((layer2_outputs(4008)) xor (layer2_outputs(9634)));
    outputs(1961) <= (layer2_outputs(4160)) xor (layer2_outputs(7884));
    outputs(1962) <= (layer2_outputs(5915)) or (layer2_outputs(682));
    outputs(1963) <= (layer2_outputs(3530)) and not (layer2_outputs(6360));
    outputs(1964) <= not((layer2_outputs(8468)) or (layer2_outputs(3785)));
    outputs(1965) <= not(layer2_outputs(3548));
    outputs(1966) <= not(layer2_outputs(3987));
    outputs(1967) <= layer2_outputs(5266);
    outputs(1968) <= (layer2_outputs(4398)) and not (layer2_outputs(416));
    outputs(1969) <= not(layer2_outputs(1150));
    outputs(1970) <= layer2_outputs(1625);
    outputs(1971) <= layer2_outputs(3616);
    outputs(1972) <= (layer2_outputs(5737)) and not (layer2_outputs(5041));
    outputs(1973) <= not((layer2_outputs(1201)) xor (layer2_outputs(8835)));
    outputs(1974) <= layer2_outputs(3031);
    outputs(1975) <= not(layer2_outputs(5415));
    outputs(1976) <= not(layer2_outputs(8232));
    outputs(1977) <= not(layer2_outputs(6198));
    outputs(1978) <= not(layer2_outputs(2171));
    outputs(1979) <= '0';
    outputs(1980) <= layer2_outputs(3556);
    outputs(1981) <= not(layer2_outputs(1689));
    outputs(1982) <= not((layer2_outputs(6251)) or (layer2_outputs(2032)));
    outputs(1983) <= (layer2_outputs(6497)) and not (layer2_outputs(8439));
    outputs(1984) <= not(layer2_outputs(7611));
    outputs(1985) <= not((layer2_outputs(2144)) or (layer2_outputs(195)));
    outputs(1986) <= not(layer2_outputs(6019));
    outputs(1987) <= layer2_outputs(9240);
    outputs(1988) <= layer2_outputs(5532);
    outputs(1989) <= not((layer2_outputs(7273)) xor (layer2_outputs(8811)));
    outputs(1990) <= layer2_outputs(6271);
    outputs(1991) <= not(layer2_outputs(4505));
    outputs(1992) <= not(layer2_outputs(1177));
    outputs(1993) <= layer2_outputs(7765);
    outputs(1994) <= not((layer2_outputs(1927)) or (layer2_outputs(7331)));
    outputs(1995) <= (layer2_outputs(1988)) xor (layer2_outputs(8018));
    outputs(1996) <= not(layer2_outputs(5923));
    outputs(1997) <= (layer2_outputs(3132)) xor (layer2_outputs(2335));
    outputs(1998) <= not((layer2_outputs(2566)) or (layer2_outputs(6834)));
    outputs(1999) <= (layer2_outputs(8528)) and not (layer2_outputs(4387));
    outputs(2000) <= not(layer2_outputs(7964));
    outputs(2001) <= not(layer2_outputs(1616));
    outputs(2002) <= layer2_outputs(3537);
    outputs(2003) <= layer2_outputs(338);
    outputs(2004) <= (layer2_outputs(6004)) xor (layer2_outputs(5891));
    outputs(2005) <= (layer2_outputs(2930)) and not (layer2_outputs(6553));
    outputs(2006) <= layer2_outputs(3619);
    outputs(2007) <= (layer2_outputs(3444)) and not (layer2_outputs(8114));
    outputs(2008) <= (layer2_outputs(986)) and (layer2_outputs(1440));
    outputs(2009) <= (layer2_outputs(1882)) and (layer2_outputs(7918));
    outputs(2010) <= not(layer2_outputs(2530));
    outputs(2011) <= (layer2_outputs(6503)) and (layer2_outputs(8957));
    outputs(2012) <= (layer2_outputs(4398)) and (layer2_outputs(1077));
    outputs(2013) <= layer2_outputs(2358);
    outputs(2014) <= not((layer2_outputs(483)) xor (layer2_outputs(8690)));
    outputs(2015) <= layer2_outputs(3772);
    outputs(2016) <= not((layer2_outputs(6446)) xor (layer2_outputs(604)));
    outputs(2017) <= not(layer2_outputs(8424));
    outputs(2018) <= not(layer2_outputs(749));
    outputs(2019) <= not((layer2_outputs(1570)) xor (layer2_outputs(2064)));
    outputs(2020) <= (layer2_outputs(9523)) and (layer2_outputs(1025));
    outputs(2021) <= not(layer2_outputs(1278));
    outputs(2022) <= layer2_outputs(7583);
    outputs(2023) <= not(layer2_outputs(3868));
    outputs(2024) <= (layer2_outputs(8907)) xor (layer2_outputs(9305));
    outputs(2025) <= not(layer2_outputs(8113));
    outputs(2026) <= (layer2_outputs(4547)) and not (layer2_outputs(1805));
    outputs(2027) <= not(layer2_outputs(2216));
    outputs(2028) <= (layer2_outputs(530)) and not (layer2_outputs(109));
    outputs(2029) <= not(layer2_outputs(6325));
    outputs(2030) <= (layer2_outputs(8840)) and not (layer2_outputs(2950));
    outputs(2031) <= not((layer2_outputs(1969)) or (layer2_outputs(767)));
    outputs(2032) <= not(layer2_outputs(7725));
    outputs(2033) <= layer2_outputs(9410);
    outputs(2034) <= (layer2_outputs(10164)) and not (layer2_outputs(8466));
    outputs(2035) <= layer2_outputs(1122);
    outputs(2036) <= (layer2_outputs(9348)) and not (layer2_outputs(10066));
    outputs(2037) <= layer2_outputs(5025);
    outputs(2038) <= layer2_outputs(7226);
    outputs(2039) <= not(layer2_outputs(922));
    outputs(2040) <= not(layer2_outputs(1521));
    outputs(2041) <= (layer2_outputs(2159)) and not (layer2_outputs(9053));
    outputs(2042) <= not(layer2_outputs(7853));
    outputs(2043) <= layer2_outputs(7277);
    outputs(2044) <= not(layer2_outputs(4351));
    outputs(2045) <= layer2_outputs(527);
    outputs(2046) <= (layer2_outputs(9830)) xor (layer2_outputs(1488));
    outputs(2047) <= (layer2_outputs(237)) and not (layer2_outputs(8270));
    outputs(2048) <= layer2_outputs(4855);
    outputs(2049) <= layer2_outputs(1066);
    outputs(2050) <= (layer2_outputs(4873)) and not (layer2_outputs(4234));
    outputs(2051) <= layer2_outputs(5673);
    outputs(2052) <= (layer2_outputs(859)) xor (layer2_outputs(889));
    outputs(2053) <= layer2_outputs(5197);
    outputs(2054) <= not(layer2_outputs(5137));
    outputs(2055) <= not(layer2_outputs(9113));
    outputs(2056) <= not((layer2_outputs(9209)) and (layer2_outputs(8226)));
    outputs(2057) <= not(layer2_outputs(6304));
    outputs(2058) <= layer2_outputs(8133);
    outputs(2059) <= layer2_outputs(4326);
    outputs(2060) <= layer2_outputs(6762);
    outputs(2061) <= layer2_outputs(3861);
    outputs(2062) <= not((layer2_outputs(1919)) and (layer2_outputs(6567)));
    outputs(2063) <= not(layer2_outputs(9215));
    outputs(2064) <= layer2_outputs(4033);
    outputs(2065) <= layer2_outputs(4575);
    outputs(2066) <= layer2_outputs(900);
    outputs(2067) <= not(layer2_outputs(3995));
    outputs(2068) <= not((layer2_outputs(5608)) xor (layer2_outputs(7243)));
    outputs(2069) <= not(layer2_outputs(6303));
    outputs(2070) <= not(layer2_outputs(9253));
    outputs(2071) <= not(layer2_outputs(3502));
    outputs(2072) <= not(layer2_outputs(1515)) or (layer2_outputs(1497));
    outputs(2073) <= (layer2_outputs(6573)) xor (layer2_outputs(708));
    outputs(2074) <= (layer2_outputs(6711)) and (layer2_outputs(4698));
    outputs(2075) <= not(layer2_outputs(5442));
    outputs(2076) <= not((layer2_outputs(6141)) xor (layer2_outputs(6378)));
    outputs(2077) <= not(layer2_outputs(4086));
    outputs(2078) <= layer2_outputs(1780);
    outputs(2079) <= layer2_outputs(9454);
    outputs(2080) <= not(layer2_outputs(598));
    outputs(2081) <= layer2_outputs(1903);
    outputs(2082) <= not((layer2_outputs(9903)) xor (layer2_outputs(7749)));
    outputs(2083) <= not(layer2_outputs(3630));
    outputs(2084) <= layer2_outputs(9000);
    outputs(2085) <= not((layer2_outputs(9467)) xor (layer2_outputs(7796)));
    outputs(2086) <= (layer2_outputs(9702)) and (layer2_outputs(1196));
    outputs(2087) <= (layer2_outputs(5010)) and not (layer2_outputs(9879));
    outputs(2088) <= not(layer2_outputs(4275));
    outputs(2089) <= not(layer2_outputs(7696));
    outputs(2090) <= (layer2_outputs(5335)) xor (layer2_outputs(9519));
    outputs(2091) <= (layer2_outputs(1987)) or (layer2_outputs(5805));
    outputs(2092) <= not(layer2_outputs(4824));
    outputs(2093) <= not((layer2_outputs(3356)) and (layer2_outputs(3214)));
    outputs(2094) <= not(layer2_outputs(7236));
    outputs(2095) <= layer2_outputs(8342);
    outputs(2096) <= layer2_outputs(3409);
    outputs(2097) <= layer2_outputs(1306);
    outputs(2098) <= not(layer2_outputs(3567));
    outputs(2099) <= not((layer2_outputs(2736)) or (layer2_outputs(5103)));
    outputs(2100) <= layer2_outputs(8413);
    outputs(2101) <= not(layer2_outputs(9250));
    outputs(2102) <= not(layer2_outputs(9593));
    outputs(2103) <= layer2_outputs(5181);
    outputs(2104) <= not((layer2_outputs(461)) or (layer2_outputs(4984)));
    outputs(2105) <= layer2_outputs(1524);
    outputs(2106) <= (layer2_outputs(2288)) xor (layer2_outputs(9478));
    outputs(2107) <= not(layer2_outputs(1603));
    outputs(2108) <= layer2_outputs(2623);
    outputs(2109) <= not(layer2_outputs(7357));
    outputs(2110) <= not(layer2_outputs(1909));
    outputs(2111) <= not(layer2_outputs(9317));
    outputs(2112) <= layer2_outputs(2678);
    outputs(2113) <= not((layer2_outputs(4997)) and (layer2_outputs(7868)));
    outputs(2114) <= layer2_outputs(3476);
    outputs(2115) <= layer2_outputs(4175);
    outputs(2116) <= layer2_outputs(952);
    outputs(2117) <= not(layer2_outputs(3456));
    outputs(2118) <= not(layer2_outputs(1918));
    outputs(2119) <= not((layer2_outputs(8993)) and (layer2_outputs(1193)));
    outputs(2120) <= not((layer2_outputs(6660)) xor (layer2_outputs(3084)));
    outputs(2121) <= not(layer2_outputs(1031));
    outputs(2122) <= layer2_outputs(2177);
    outputs(2123) <= not((layer2_outputs(8320)) or (layer2_outputs(7241)));
    outputs(2124) <= not(layer2_outputs(6563)) or (layer2_outputs(1480));
    outputs(2125) <= not(layer2_outputs(29));
    outputs(2126) <= layer2_outputs(4180);
    outputs(2127) <= layer2_outputs(9790);
    outputs(2128) <= layer2_outputs(2178);
    outputs(2129) <= (layer2_outputs(8740)) and not (layer2_outputs(8066));
    outputs(2130) <= not(layer2_outputs(6966));
    outputs(2131) <= not(layer2_outputs(3671));
    outputs(2132) <= layer2_outputs(2742);
    outputs(2133) <= not(layer2_outputs(5506));
    outputs(2134) <= layer2_outputs(305);
    outputs(2135) <= (layer2_outputs(3012)) and not (layer2_outputs(3853));
    outputs(2136) <= (layer2_outputs(8769)) and (layer2_outputs(5463));
    outputs(2137) <= layer2_outputs(1315);
    outputs(2138) <= layer2_outputs(565);
    outputs(2139) <= layer2_outputs(170);
    outputs(2140) <= not(layer2_outputs(2357));
    outputs(2141) <= layer2_outputs(4892);
    outputs(2142) <= not(layer2_outputs(1633));
    outputs(2143) <= not((layer2_outputs(9751)) and (layer2_outputs(8523)));
    outputs(2144) <= not((layer2_outputs(7311)) xor (layer2_outputs(4739)));
    outputs(2145) <= not((layer2_outputs(3963)) or (layer2_outputs(6840)));
    outputs(2146) <= layer2_outputs(9398);
    outputs(2147) <= layer2_outputs(6358);
    outputs(2148) <= not(layer2_outputs(4969));
    outputs(2149) <= not(layer2_outputs(3855));
    outputs(2150) <= not((layer2_outputs(2556)) and (layer2_outputs(2212)));
    outputs(2151) <= layer2_outputs(205);
    outputs(2152) <= not(layer2_outputs(2624));
    outputs(2153) <= layer2_outputs(1225);
    outputs(2154) <= not(layer2_outputs(3821));
    outputs(2155) <= (layer2_outputs(6415)) and not (layer2_outputs(6478));
    outputs(2156) <= layer2_outputs(8831);
    outputs(2157) <= layer2_outputs(9735);
    outputs(2158) <= (layer2_outputs(8181)) and (layer2_outputs(7276));
    outputs(2159) <= layer2_outputs(775);
    outputs(2160) <= not(layer2_outputs(9624));
    outputs(2161) <= layer2_outputs(3110);
    outputs(2162) <= not(layer2_outputs(2217));
    outputs(2163) <= layer2_outputs(927);
    outputs(2164) <= layer2_outputs(6927);
    outputs(2165) <= layer2_outputs(696);
    outputs(2166) <= layer2_outputs(6103);
    outputs(2167) <= (layer2_outputs(321)) and (layer2_outputs(1462));
    outputs(2168) <= layer2_outputs(7232);
    outputs(2169) <= not((layer2_outputs(4367)) and (layer2_outputs(413)));
    outputs(2170) <= not((layer2_outputs(244)) and (layer2_outputs(9847)));
    outputs(2171) <= not(layer2_outputs(2205));
    outputs(2172) <= layer2_outputs(4866);
    outputs(2173) <= not(layer2_outputs(5873));
    outputs(2174) <= layer2_outputs(8983);
    outputs(2175) <= layer2_outputs(7844);
    outputs(2176) <= layer2_outputs(4995);
    outputs(2177) <= not((layer2_outputs(7109)) or (layer2_outputs(2689)));
    outputs(2178) <= layer2_outputs(1624);
    outputs(2179) <= not(layer2_outputs(7536));
    outputs(2180) <= layer2_outputs(6388);
    outputs(2181) <= not((layer2_outputs(9252)) xor (layer2_outputs(9463)));
    outputs(2182) <= (layer2_outputs(3861)) and not (layer2_outputs(576));
    outputs(2183) <= not((layer2_outputs(4303)) or (layer2_outputs(383)));
    outputs(2184) <= not((layer2_outputs(8860)) xor (layer2_outputs(2527)));
    outputs(2185) <= not(layer2_outputs(1021));
    outputs(2186) <= not(layer2_outputs(9401));
    outputs(2187) <= layer2_outputs(1885);
    outputs(2188) <= (layer2_outputs(9380)) or (layer2_outputs(9308));
    outputs(2189) <= not((layer2_outputs(4328)) and (layer2_outputs(4191)));
    outputs(2190) <= layer2_outputs(5576);
    outputs(2191) <= layer2_outputs(5758);
    outputs(2192) <= not((layer2_outputs(9482)) xor (layer2_outputs(10090)));
    outputs(2193) <= not(layer2_outputs(3470));
    outputs(2194) <= not((layer2_outputs(7985)) and (layer2_outputs(6784)));
    outputs(2195) <= layer2_outputs(2928);
    outputs(2196) <= (layer2_outputs(7391)) and not (layer2_outputs(4432));
    outputs(2197) <= not(layer2_outputs(8500));
    outputs(2198) <= not((layer2_outputs(1229)) or (layer2_outputs(5597)));
    outputs(2199) <= layer2_outputs(7042);
    outputs(2200) <= layer2_outputs(558);
    outputs(2201) <= not(layer2_outputs(517));
    outputs(2202) <= layer2_outputs(8258);
    outputs(2203) <= layer2_outputs(1833);
    outputs(2204) <= layer2_outputs(2742);
    outputs(2205) <= layer2_outputs(6298);
    outputs(2206) <= not(layer2_outputs(330)) or (layer2_outputs(8722));
    outputs(2207) <= not(layer2_outputs(7405));
    outputs(2208) <= not((layer2_outputs(4560)) xor (layer2_outputs(8724)));
    outputs(2209) <= not((layer2_outputs(3398)) xor (layer2_outputs(6987)));
    outputs(2210) <= not((layer2_outputs(3335)) or (layer2_outputs(8706)));
    outputs(2211) <= layer2_outputs(9266);
    outputs(2212) <= (layer2_outputs(6528)) or (layer2_outputs(2829));
    outputs(2213) <= not(layer2_outputs(4442));
    outputs(2214) <= not(layer2_outputs(2270));
    outputs(2215) <= (layer2_outputs(5761)) xor (layer2_outputs(7623));
    outputs(2216) <= layer2_outputs(1237);
    outputs(2217) <= not(layer2_outputs(9447));
    outputs(2218) <= not(layer2_outputs(2996));
    outputs(2219) <= not(layer2_outputs(5461));
    outputs(2220) <= layer2_outputs(5984);
    outputs(2221) <= layer2_outputs(4091);
    outputs(2222) <= layer2_outputs(8889);
    outputs(2223) <= (layer2_outputs(1501)) and not (layer2_outputs(3380));
    outputs(2224) <= layer2_outputs(4865);
    outputs(2225) <= not(layer2_outputs(3351));
    outputs(2226) <= not(layer2_outputs(8879));
    outputs(2227) <= layer2_outputs(1190);
    outputs(2228) <= not(layer2_outputs(8984));
    outputs(2229) <= layer2_outputs(5440);
    outputs(2230) <= not(layer2_outputs(7371));
    outputs(2231) <= not(layer2_outputs(10047)) or (layer2_outputs(7500));
    outputs(2232) <= not((layer2_outputs(9167)) and (layer2_outputs(3720)));
    outputs(2233) <= not(layer2_outputs(8129));
    outputs(2234) <= not(layer2_outputs(2392)) or (layer2_outputs(6065));
    outputs(2235) <= (layer2_outputs(3178)) and (layer2_outputs(9196));
    outputs(2236) <= not(layer2_outputs(1701));
    outputs(2237) <= not(layer2_outputs(3253)) or (layer2_outputs(8127));
    outputs(2238) <= not(layer2_outputs(8170)) or (layer2_outputs(3154));
    outputs(2239) <= not(layer2_outputs(7720));
    outputs(2240) <= not(layer2_outputs(8273));
    outputs(2241) <= not((layer2_outputs(2922)) xor (layer2_outputs(1556)));
    outputs(2242) <= layer2_outputs(3177);
    outputs(2243) <= (layer2_outputs(3522)) xor (layer2_outputs(10024));
    outputs(2244) <= not(layer2_outputs(8669)) or (layer2_outputs(1373));
    outputs(2245) <= not(layer2_outputs(8306));
    outputs(2246) <= not(layer2_outputs(8587)) or (layer2_outputs(9052));
    outputs(2247) <= not(layer2_outputs(7476));
    outputs(2248) <= not((layer2_outputs(6157)) and (layer2_outputs(433)));
    outputs(2249) <= layer2_outputs(5598);
    outputs(2250) <= (layer2_outputs(8466)) or (layer2_outputs(8792));
    outputs(2251) <= not((layer2_outputs(6295)) xor (layer2_outputs(6192)));
    outputs(2252) <= not(layer2_outputs(6426));
    outputs(2253) <= not(layer2_outputs(8337)) or (layer2_outputs(3576));
    outputs(2254) <= not((layer2_outputs(3848)) xor (layer2_outputs(3272)));
    outputs(2255) <= (layer2_outputs(9037)) xor (layer2_outputs(6783));
    outputs(2256) <= not(layer2_outputs(8138));
    outputs(2257) <= not((layer2_outputs(8252)) xor (layer2_outputs(8341)));
    outputs(2258) <= not(layer2_outputs(5309)) or (layer2_outputs(1780));
    outputs(2259) <= not((layer2_outputs(1192)) and (layer2_outputs(4763)));
    outputs(2260) <= not(layer2_outputs(215));
    outputs(2261) <= not(layer2_outputs(2740));
    outputs(2262) <= layer2_outputs(4374);
    outputs(2263) <= not((layer2_outputs(1408)) or (layer2_outputs(2587)));
    outputs(2264) <= not(layer2_outputs(5027)) or (layer2_outputs(9451));
    outputs(2265) <= layer2_outputs(1484);
    outputs(2266) <= not(layer2_outputs(5050));
    outputs(2267) <= not(layer2_outputs(1228));
    outputs(2268) <= not((layer2_outputs(2297)) xor (layer2_outputs(2194)));
    outputs(2269) <= (layer2_outputs(5154)) xor (layer2_outputs(5709));
    outputs(2270) <= (layer2_outputs(5782)) and not (layer2_outputs(6249));
    outputs(2271) <= layer2_outputs(9162);
    outputs(2272) <= layer2_outputs(4735);
    outputs(2273) <= layer2_outputs(10019);
    outputs(2274) <= not(layer2_outputs(6975));
    outputs(2275) <= (layer2_outputs(2455)) or (layer2_outputs(1839));
    outputs(2276) <= layer2_outputs(4905);
    outputs(2277) <= layer2_outputs(8689);
    outputs(2278) <= (layer2_outputs(5174)) or (layer2_outputs(333));
    outputs(2279) <= layer2_outputs(10073);
    outputs(2280) <= not(layer2_outputs(4024));
    outputs(2281) <= (layer2_outputs(2439)) xor (layer2_outputs(2139));
    outputs(2282) <= layer2_outputs(2393);
    outputs(2283) <= (layer2_outputs(6040)) and not (layer2_outputs(4849));
    outputs(2284) <= layer2_outputs(5037);
    outputs(2285) <= not((layer2_outputs(8728)) and (layer2_outputs(3392)));
    outputs(2286) <= layer2_outputs(144);
    outputs(2287) <= not(layer2_outputs(8704)) or (layer2_outputs(7179));
    outputs(2288) <= layer2_outputs(1252);
    outputs(2289) <= not((layer2_outputs(4007)) and (layer2_outputs(10042)));
    outputs(2290) <= layer2_outputs(4608);
    outputs(2291) <= layer2_outputs(1968);
    outputs(2292) <= layer2_outputs(9846);
    outputs(2293) <= not((layer2_outputs(2702)) xor (layer2_outputs(3781)));
    outputs(2294) <= (layer2_outputs(2671)) and not (layer2_outputs(4729));
    outputs(2295) <= not((layer2_outputs(7579)) and (layer2_outputs(4953)));
    outputs(2296) <= not(layer2_outputs(1433)) or (layer2_outputs(8259));
    outputs(2297) <= layer2_outputs(2122);
    outputs(2298) <= not(layer2_outputs(7677));
    outputs(2299) <= not(layer2_outputs(2468));
    outputs(2300) <= not(layer2_outputs(6391));
    outputs(2301) <= (layer2_outputs(5640)) and not (layer2_outputs(610));
    outputs(2302) <= not(layer2_outputs(2926));
    outputs(2303) <= layer2_outputs(160);
    outputs(2304) <= not(layer2_outputs(7365)) or (layer2_outputs(2511));
    outputs(2305) <= not(layer2_outputs(8797));
    outputs(2306) <= layer2_outputs(8751);
    outputs(2307) <= (layer2_outputs(4813)) xor (layer2_outputs(5631));
    outputs(2308) <= layer2_outputs(6758);
    outputs(2309) <= not(layer2_outputs(7244));
    outputs(2310) <= layer2_outputs(6034);
    outputs(2311) <= not((layer2_outputs(1468)) xor (layer2_outputs(5949)));
    outputs(2312) <= not(layer2_outputs(5810));
    outputs(2313) <= layer2_outputs(3274);
    outputs(2314) <= (layer2_outputs(2146)) and not (layer2_outputs(6202));
    outputs(2315) <= layer2_outputs(2420);
    outputs(2316) <= not(layer2_outputs(7965));
    outputs(2317) <= (layer2_outputs(2611)) or (layer2_outputs(3568));
    outputs(2318) <= not((layer2_outputs(4954)) xor (layer2_outputs(38)));
    outputs(2319) <= not((layer2_outputs(5486)) xor (layer2_outputs(6674)));
    outputs(2320) <= (layer2_outputs(2916)) or (layer2_outputs(2191));
    outputs(2321) <= layer2_outputs(493);
    outputs(2322) <= not(layer2_outputs(3692)) or (layer2_outputs(6825));
    outputs(2323) <= (layer2_outputs(1881)) and (layer2_outputs(7001));
    outputs(2324) <= layer2_outputs(918);
    outputs(2325) <= (layer2_outputs(2280)) or (layer2_outputs(9779));
    outputs(2326) <= (layer2_outputs(1152)) xor (layer2_outputs(9254));
    outputs(2327) <= (layer2_outputs(5015)) or (layer2_outputs(592));
    outputs(2328) <= (layer2_outputs(9259)) xor (layer2_outputs(6466));
    outputs(2329) <= (layer2_outputs(4464)) or (layer2_outputs(8672));
    outputs(2330) <= (layer2_outputs(61)) and not (layer2_outputs(1814));
    outputs(2331) <= layer2_outputs(8784);
    outputs(2332) <= not((layer2_outputs(9978)) xor (layer2_outputs(10163)));
    outputs(2333) <= not(layer2_outputs(7931)) or (layer2_outputs(5662));
    outputs(2334) <= layer2_outputs(9223);
    outputs(2335) <= not(layer2_outputs(5436));
    outputs(2336) <= not((layer2_outputs(2824)) or (layer2_outputs(4102)));
    outputs(2337) <= (layer2_outputs(5978)) and not (layer2_outputs(9889));
    outputs(2338) <= (layer2_outputs(6448)) xor (layer2_outputs(9698));
    outputs(2339) <= layer2_outputs(478);
    outputs(2340) <= (layer2_outputs(7128)) and not (layer2_outputs(5049));
    outputs(2341) <= not((layer2_outputs(9135)) and (layer2_outputs(9967)));
    outputs(2342) <= not(layer2_outputs(2089));
    outputs(2343) <= not(layer2_outputs(3582));
    outputs(2344) <= not(layer2_outputs(4397));
    outputs(2345) <= not(layer2_outputs(8679));
    outputs(2346) <= not(layer2_outputs(2373)) or (layer2_outputs(967));
    outputs(2347) <= not((layer2_outputs(1960)) xor (layer2_outputs(410)));
    outputs(2348) <= not((layer2_outputs(9774)) xor (layer2_outputs(6458)));
    outputs(2349) <= layer2_outputs(8328);
    outputs(2350) <= (layer2_outputs(3729)) and not (layer2_outputs(4424));
    outputs(2351) <= not(layer2_outputs(4485)) or (layer2_outputs(1494));
    outputs(2352) <= not(layer2_outputs(437));
    outputs(2353) <= not(layer2_outputs(8444));
    outputs(2354) <= not(layer2_outputs(3712));
    outputs(2355) <= not(layer2_outputs(2384));
    outputs(2356) <= not((layer2_outputs(4786)) or (layer2_outputs(2645)));
    outputs(2357) <= not((layer2_outputs(2899)) xor (layer2_outputs(8160)));
    outputs(2358) <= not(layer2_outputs(809));
    outputs(2359) <= not(layer2_outputs(8311));
    outputs(2360) <= layer2_outputs(4368);
    outputs(2361) <= not(layer2_outputs(2933));
    outputs(2362) <= not(layer2_outputs(9911));
    outputs(2363) <= layer2_outputs(8946);
    outputs(2364) <= not(layer2_outputs(8136)) or (layer2_outputs(4081));
    outputs(2365) <= layer2_outputs(3324);
    outputs(2366) <= layer2_outputs(2274);
    outputs(2367) <= (layer2_outputs(5045)) and not (layer2_outputs(3427));
    outputs(2368) <= layer2_outputs(915);
    outputs(2369) <= not((layer2_outputs(5076)) xor (layer2_outputs(901)));
    outputs(2370) <= not(layer2_outputs(2456));
    outputs(2371) <= layer2_outputs(4723);
    outputs(2372) <= layer2_outputs(308);
    outputs(2373) <= not(layer2_outputs(4842));
    outputs(2374) <= not(layer2_outputs(344));
    outputs(2375) <= layer2_outputs(9364);
    outputs(2376) <= not(layer2_outputs(3439)) or (layer2_outputs(429));
    outputs(2377) <= layer2_outputs(4552);
    outputs(2378) <= layer2_outputs(1161);
    outputs(2379) <= not(layer2_outputs(2009));
    outputs(2380) <= not(layer2_outputs(10045));
    outputs(2381) <= (layer2_outputs(2005)) or (layer2_outputs(8464));
    outputs(2382) <= not(layer2_outputs(9676));
    outputs(2383) <= not(layer2_outputs(5678));
    outputs(2384) <= layer2_outputs(5299);
    outputs(2385) <= (layer2_outputs(6767)) and not (layer2_outputs(4577));
    outputs(2386) <= layer2_outputs(2226);
    outputs(2387) <= layer2_outputs(9841);
    outputs(2388) <= not(layer2_outputs(3139));
    outputs(2389) <= not((layer2_outputs(2247)) xor (layer2_outputs(8149)));
    outputs(2390) <= not((layer2_outputs(1347)) and (layer2_outputs(9512)));
    outputs(2391) <= layer2_outputs(5187);
    outputs(2392) <= not((layer2_outputs(6109)) and (layer2_outputs(4638)));
    outputs(2393) <= not((layer2_outputs(5956)) xor (layer2_outputs(8935)));
    outputs(2394) <= not((layer2_outputs(7174)) xor (layer2_outputs(1723)));
    outputs(2395) <= not(layer2_outputs(647));
    outputs(2396) <= (layer2_outputs(7324)) and not (layer2_outputs(3380));
    outputs(2397) <= not((layer2_outputs(1493)) xor (layer2_outputs(7191)));
    outputs(2398) <= layer2_outputs(9736);
    outputs(2399) <= (layer2_outputs(5082)) xor (layer2_outputs(1431));
    outputs(2400) <= (layer2_outputs(6801)) xor (layer2_outputs(6047));
    outputs(2401) <= not(layer2_outputs(1771));
    outputs(2402) <= layer2_outputs(1223);
    outputs(2403) <= not(layer2_outputs(8917));
    outputs(2404) <= not(layer2_outputs(9031));
    outputs(2405) <= not(layer2_outputs(3101));
    outputs(2406) <= (layer2_outputs(5088)) or (layer2_outputs(9132));
    outputs(2407) <= not(layer2_outputs(666));
    outputs(2408) <= not(layer2_outputs(2782));
    outputs(2409) <= layer2_outputs(6281);
    outputs(2410) <= not(layer2_outputs(8546));
    outputs(2411) <= layer2_outputs(2398);
    outputs(2412) <= not((layer2_outputs(1026)) xor (layer2_outputs(4773)));
    outputs(2413) <= layer2_outputs(5272);
    outputs(2414) <= layer2_outputs(1225);
    outputs(2415) <= not(layer2_outputs(4421));
    outputs(2416) <= layer2_outputs(2471);
    outputs(2417) <= layer2_outputs(2981);
    outputs(2418) <= not((layer2_outputs(4056)) or (layer2_outputs(7017)));
    outputs(2419) <= not(layer2_outputs(8177));
    outputs(2420) <= (layer2_outputs(7003)) xor (layer2_outputs(8820));
    outputs(2421) <= not((layer2_outputs(8081)) xor (layer2_outputs(3052)));
    outputs(2422) <= not(layer2_outputs(5725));
    outputs(2423) <= (layer2_outputs(5649)) or (layer2_outputs(6153));
    outputs(2424) <= not(layer2_outputs(9511));
    outputs(2425) <= not(layer2_outputs(3606));
    outputs(2426) <= not(layer2_outputs(8432)) or (layer2_outputs(1700));
    outputs(2427) <= not(layer2_outputs(5811));
    outputs(2428) <= (layer2_outputs(6208)) xor (layer2_outputs(1422));
    outputs(2429) <= (layer2_outputs(221)) xor (layer2_outputs(2012));
    outputs(2430) <= not(layer2_outputs(9204));
    outputs(2431) <= not(layer2_outputs(951));
    outputs(2432) <= layer2_outputs(6092);
    outputs(2433) <= not(layer2_outputs(1542));
    outputs(2434) <= not(layer2_outputs(1982));
    outputs(2435) <= not(layer2_outputs(847));
    outputs(2436) <= layer2_outputs(2291);
    outputs(2437) <= not(layer2_outputs(4675));
    outputs(2438) <= layer2_outputs(5765);
    outputs(2439) <= not((layer2_outputs(509)) xor (layer2_outputs(7852)));
    outputs(2440) <= layer2_outputs(4523);
    outputs(2441) <= layer2_outputs(5628);
    outputs(2442) <= not((layer2_outputs(3263)) xor (layer2_outputs(8560)));
    outputs(2443) <= not(layer2_outputs(2621)) or (layer2_outputs(3378));
    outputs(2444) <= (layer2_outputs(9435)) xor (layer2_outputs(982));
    outputs(2445) <= not(layer2_outputs(1295));
    outputs(2446) <= not(layer2_outputs(9784)) or (layer2_outputs(2218));
    outputs(2447) <= layer2_outputs(8650);
    outputs(2448) <= (layer2_outputs(1931)) xor (layer2_outputs(8533));
    outputs(2449) <= not(layer2_outputs(9815));
    outputs(2450) <= not((layer2_outputs(9924)) and (layer2_outputs(6815)));
    outputs(2451) <= not((layer2_outputs(9172)) xor (layer2_outputs(3880)));
    outputs(2452) <= not(layer2_outputs(4310));
    outputs(2453) <= not(layer2_outputs(7130));
    outputs(2454) <= layer2_outputs(257);
    outputs(2455) <= not((layer2_outputs(6080)) and (layer2_outputs(7772)));
    outputs(2456) <= layer2_outputs(227);
    outputs(2457) <= layer2_outputs(6943);
    outputs(2458) <= not(layer2_outputs(1867));
    outputs(2459) <= layer2_outputs(465);
    outputs(2460) <= (layer2_outputs(340)) xor (layer2_outputs(6083));
    outputs(2461) <= not(layer2_outputs(6012));
    outputs(2462) <= (layer2_outputs(4115)) and not (layer2_outputs(7920));
    outputs(2463) <= layer2_outputs(7572);
    outputs(2464) <= not(layer2_outputs(738));
    outputs(2465) <= not((layer2_outputs(2888)) and (layer2_outputs(7261)));
    outputs(2466) <= not(layer2_outputs(9249));
    outputs(2467) <= not(layer2_outputs(5760));
    outputs(2468) <= layer2_outputs(2390);
    outputs(2469) <= layer2_outputs(7480);
    outputs(2470) <= layer2_outputs(7967);
    outputs(2471) <= layer2_outputs(4235);
    outputs(2472) <= layer2_outputs(1751);
    outputs(2473) <= layer2_outputs(1155);
    outputs(2474) <= layer2_outputs(6035);
    outputs(2475) <= (layer2_outputs(8088)) xor (layer2_outputs(146));
    outputs(2476) <= not(layer2_outputs(5785));
    outputs(2477) <= layer2_outputs(2344);
    outputs(2478) <= layer2_outputs(7883);
    outputs(2479) <= (layer2_outputs(6033)) xor (layer2_outputs(6395));
    outputs(2480) <= not(layer2_outputs(7067));
    outputs(2481) <= not(layer2_outputs(7055)) or (layer2_outputs(7589));
    outputs(2482) <= (layer2_outputs(3798)) xor (layer2_outputs(3117));
    outputs(2483) <= layer2_outputs(7777);
    outputs(2484) <= layer2_outputs(9846);
    outputs(2485) <= layer2_outputs(3576);
    outputs(2486) <= (layer2_outputs(4067)) xor (layer2_outputs(998));
    outputs(2487) <= layer2_outputs(6495);
    outputs(2488) <= not(layer2_outputs(3431)) or (layer2_outputs(1955));
    outputs(2489) <= not(layer2_outputs(6081));
    outputs(2490) <= not(layer2_outputs(5074));
    outputs(2491) <= not(layer2_outputs(6517));
    outputs(2492) <= layer2_outputs(2169);
    outputs(2493) <= not((layer2_outputs(1374)) and (layer2_outputs(10223)));
    outputs(2494) <= layer2_outputs(2195);
    outputs(2495) <= (layer2_outputs(10204)) and not (layer2_outputs(5851));
    outputs(2496) <= not(layer2_outputs(9129));
    outputs(2497) <= layer2_outputs(6943);
    outputs(2498) <= layer2_outputs(196);
    outputs(2499) <= layer2_outputs(8015);
    outputs(2500) <= layer2_outputs(6870);
    outputs(2501) <= not(layer2_outputs(7145));
    outputs(2502) <= not(layer2_outputs(4291));
    outputs(2503) <= (layer2_outputs(7728)) xor (layer2_outputs(1307));
    outputs(2504) <= not(layer2_outputs(496)) or (layer2_outputs(8013));
    outputs(2505) <= (layer2_outputs(577)) xor (layer2_outputs(4289));
    outputs(2506) <= layer2_outputs(7989);
    outputs(2507) <= (layer2_outputs(8207)) xor (layer2_outputs(428));
    outputs(2508) <= not((layer2_outputs(5059)) or (layer2_outputs(5557)));
    outputs(2509) <= not((layer2_outputs(1774)) xor (layer2_outputs(5310)));
    outputs(2510) <= (layer2_outputs(1421)) and not (layer2_outputs(9759));
    outputs(2511) <= layer2_outputs(6716);
    outputs(2512) <= layer2_outputs(5060);
    outputs(2513) <= not((layer2_outputs(6352)) or (layer2_outputs(3487)));
    outputs(2514) <= (layer2_outputs(6433)) and (layer2_outputs(5889));
    outputs(2515) <= not((layer2_outputs(4861)) and (layer2_outputs(8461)));
    outputs(2516) <= not((layer2_outputs(3441)) xor (layer2_outputs(9)));
    outputs(2517) <= (layer2_outputs(9190)) or (layer2_outputs(5789));
    outputs(2518) <= layer2_outputs(6764);
    outputs(2519) <= not((layer2_outputs(1496)) and (layer2_outputs(9171)));
    outputs(2520) <= not(layer2_outputs(2878));
    outputs(2521) <= not(layer2_outputs(9958)) or (layer2_outputs(2311));
    outputs(2522) <= not(layer2_outputs(3712)) or (layer2_outputs(9443));
    outputs(2523) <= (layer2_outputs(1779)) and not (layer2_outputs(3367));
    outputs(2524) <= layer2_outputs(5149);
    outputs(2525) <= not(layer2_outputs(2114));
    outputs(2526) <= not((layer2_outputs(6800)) xor (layer2_outputs(6833)));
    outputs(2527) <= (layer2_outputs(8152)) xor (layer2_outputs(10063));
    outputs(2528) <= not((layer2_outputs(9774)) xor (layer2_outputs(393)));
    outputs(2529) <= not(layer2_outputs(2367));
    outputs(2530) <= not(layer2_outputs(7646));
    outputs(2531) <= not(layer2_outputs(7902));
    outputs(2532) <= not((layer2_outputs(8192)) and (layer2_outputs(9004)));
    outputs(2533) <= not((layer2_outputs(8473)) or (layer2_outputs(3381)));
    outputs(2534) <= (layer2_outputs(9688)) xor (layer2_outputs(9196));
    outputs(2535) <= not((layer2_outputs(4367)) xor (layer2_outputs(8023)));
    outputs(2536) <= not(layer2_outputs(5723));
    outputs(2537) <= not(layer2_outputs(5847));
    outputs(2538) <= not(layer2_outputs(812));
    outputs(2539) <= not((layer2_outputs(2085)) xor (layer2_outputs(9931)));
    outputs(2540) <= layer2_outputs(6243);
    outputs(2541) <= not(layer2_outputs(6416)) or (layer2_outputs(8190));
    outputs(2542) <= layer2_outputs(7089);
    outputs(2543) <= not(layer2_outputs(5690));
    outputs(2544) <= not(layer2_outputs(4273));
    outputs(2545) <= not(layer2_outputs(7817));
    outputs(2546) <= not(layer2_outputs(1011));
    outputs(2547) <= layer2_outputs(9869);
    outputs(2548) <= (layer2_outputs(8042)) and not (layer2_outputs(4574));
    outputs(2549) <= (layer2_outputs(8976)) and (layer2_outputs(1290));
    outputs(2550) <= not((layer2_outputs(8614)) or (layer2_outputs(6779)));
    outputs(2551) <= (layer2_outputs(6047)) xor (layer2_outputs(543));
    outputs(2552) <= layer2_outputs(2812);
    outputs(2553) <= layer2_outputs(2483);
    outputs(2554) <= not(layer2_outputs(7875));
    outputs(2555) <= layer2_outputs(2157);
    outputs(2556) <= layer2_outputs(1143);
    outputs(2557) <= layer2_outputs(10205);
    outputs(2558) <= layer2_outputs(7479);
    outputs(2559) <= (layer2_outputs(8089)) and not (layer2_outputs(6950));
    outputs(2560) <= not(layer2_outputs(1391));
    outputs(2561) <= layer2_outputs(9965);
    outputs(2562) <= (layer2_outputs(9387)) xor (layer2_outputs(6878));
    outputs(2563) <= layer2_outputs(4074);
    outputs(2564) <= layer2_outputs(4791);
    outputs(2565) <= not(layer2_outputs(6529));
    outputs(2566) <= (layer2_outputs(3702)) xor (layer2_outputs(9227));
    outputs(2567) <= not(layer2_outputs(7019));
    outputs(2568) <= (layer2_outputs(8771)) xor (layer2_outputs(5962));
    outputs(2569) <= layer2_outputs(1997);
    outputs(2570) <= (layer2_outputs(3814)) or (layer2_outputs(3724));
    outputs(2571) <= layer2_outputs(4401);
    outputs(2572) <= not(layer2_outputs(4060));
    outputs(2573) <= layer2_outputs(6481);
    outputs(2574) <= not((layer2_outputs(9181)) and (layer2_outputs(2100)));
    outputs(2575) <= not(layer2_outputs(6502));
    outputs(2576) <= layer2_outputs(4330);
    outputs(2577) <= not(layer2_outputs(499));
    outputs(2578) <= not(layer2_outputs(885));
    outputs(2579) <= (layer2_outputs(8628)) and not (layer2_outputs(4920));
    outputs(2580) <= not(layer2_outputs(4688));
    outputs(2581) <= not(layer2_outputs(3507));
    outputs(2582) <= not(layer2_outputs(266));
    outputs(2583) <= (layer2_outputs(7326)) or (layer2_outputs(5938));
    outputs(2584) <= not((layer2_outputs(8480)) xor (layer2_outputs(7940)));
    outputs(2585) <= layer2_outputs(5874);
    outputs(2586) <= (layer2_outputs(5321)) xor (layer2_outputs(10235));
    outputs(2587) <= not(layer2_outputs(10095));
    outputs(2588) <= not(layer2_outputs(6241)) or (layer2_outputs(802));
    outputs(2589) <= not(layer2_outputs(5668));
    outputs(2590) <= (layer2_outputs(6754)) and (layer2_outputs(4184));
    outputs(2591) <= not(layer2_outputs(6139)) or (layer2_outputs(2074));
    outputs(2592) <= layer2_outputs(3240);
    outputs(2593) <= not(layer2_outputs(5740));
    outputs(2594) <= layer2_outputs(6335);
    outputs(2595) <= not(layer2_outputs(320));
    outputs(2596) <= layer2_outputs(7052);
    outputs(2597) <= layer2_outputs(863);
    outputs(2598) <= (layer2_outputs(4426)) and (layer2_outputs(3323));
    outputs(2599) <= not(layer2_outputs(2706));
    outputs(2600) <= layer2_outputs(7663);
    outputs(2601) <= layer2_outputs(618);
    outputs(2602) <= not(layer2_outputs(8450));
    outputs(2603) <= not(layer2_outputs(5002)) or (layer2_outputs(9441));
    outputs(2604) <= not(layer2_outputs(6081));
    outputs(2605) <= (layer2_outputs(2661)) and (layer2_outputs(2177));
    outputs(2606) <= layer2_outputs(858);
    outputs(2607) <= layer2_outputs(9265);
    outputs(2608) <= not(layer2_outputs(1434));
    outputs(2609) <= not(layer2_outputs(4390));
    outputs(2610) <= layer2_outputs(5518);
    outputs(2611) <= layer2_outputs(8521);
    outputs(2612) <= not(layer2_outputs(8635));
    outputs(2613) <= layer2_outputs(2911);
    outputs(2614) <= layer2_outputs(5918);
    outputs(2615) <= layer2_outputs(1826);
    outputs(2616) <= layer2_outputs(9379);
    outputs(2617) <= layer2_outputs(4483);
    outputs(2618) <= not(layer2_outputs(6763));
    outputs(2619) <= layer2_outputs(2754);
    outputs(2620) <= (layer2_outputs(4498)) and not (layer2_outputs(3050));
    outputs(2621) <= not(layer2_outputs(2241)) or (layer2_outputs(5533));
    outputs(2622) <= not(layer2_outputs(7342));
    outputs(2623) <= not(layer2_outputs(6780));
    outputs(2624) <= not(layer2_outputs(940));
    outputs(2625) <= (layer2_outputs(9288)) and (layer2_outputs(5173));
    outputs(2626) <= (layer2_outputs(8293)) xor (layer2_outputs(5124));
    outputs(2627) <= (layer2_outputs(6270)) xor (layer2_outputs(9369));
    outputs(2628) <= not(layer2_outputs(435));
    outputs(2629) <= layer2_outputs(6307);
    outputs(2630) <= layer2_outputs(5217);
    outputs(2631) <= (layer2_outputs(5469)) and (layer2_outputs(3691));
    outputs(2632) <= not(layer2_outputs(6938));
    outputs(2633) <= not((layer2_outputs(8953)) or (layer2_outputs(9809)));
    outputs(2634) <= not(layer2_outputs(277));
    outputs(2635) <= not(layer2_outputs(2038));
    outputs(2636) <= (layer2_outputs(10204)) and not (layer2_outputs(2066));
    outputs(2637) <= (layer2_outputs(6317)) or (layer2_outputs(8826));
    outputs(2638) <= not(layer2_outputs(5919));
    outputs(2639) <= not(layer2_outputs(9557));
    outputs(2640) <= not((layer2_outputs(6647)) xor (layer2_outputs(9106)));
    outputs(2641) <= not(layer2_outputs(2933));
    outputs(2642) <= not(layer2_outputs(9693)) or (layer2_outputs(9095));
    outputs(2643) <= not((layer2_outputs(978)) xor (layer2_outputs(2586)));
    outputs(2644) <= not(layer2_outputs(8450));
    outputs(2645) <= not(layer2_outputs(7097));
    outputs(2646) <= not(layer2_outputs(2730));
    outputs(2647) <= not(layer2_outputs(4286));
    outputs(2648) <= not((layer2_outputs(5429)) xor (layer2_outputs(1983)));
    outputs(2649) <= not(layer2_outputs(7105)) or (layer2_outputs(7615));
    outputs(2650) <= not((layer2_outputs(6978)) and (layer2_outputs(3573)));
    outputs(2651) <= not(layer2_outputs(9448));
    outputs(2652) <= layer2_outputs(9198);
    outputs(2653) <= layer2_outputs(8133);
    outputs(2654) <= (layer2_outputs(1140)) or (layer2_outputs(7403));
    outputs(2655) <= (layer2_outputs(3916)) and not (layer2_outputs(1249));
    outputs(2656) <= layer2_outputs(8325);
    outputs(2657) <= not(layer2_outputs(7299));
    outputs(2658) <= not(layer2_outputs(7986));
    outputs(2659) <= not((layer2_outputs(8418)) xor (layer2_outputs(1844)));
    outputs(2660) <= not(layer2_outputs(4120));
    outputs(2661) <= not(layer2_outputs(5623));
    outputs(2662) <= not(layer2_outputs(4798));
    outputs(2663) <= not((layer2_outputs(5087)) and (layer2_outputs(5784)));
    outputs(2664) <= not(layer2_outputs(5574));
    outputs(2665) <= not(layer2_outputs(5282));
    outputs(2666) <= layer2_outputs(863);
    outputs(2667) <= layer2_outputs(458);
    outputs(2668) <= not(layer2_outputs(5229));
    outputs(2669) <= (layer2_outputs(4755)) and (layer2_outputs(7724));
    outputs(2670) <= not((layer2_outputs(9730)) or (layer2_outputs(3716)));
    outputs(2671) <= layer2_outputs(3070);
    outputs(2672) <= layer2_outputs(7276);
    outputs(2673) <= not(layer2_outputs(9025));
    outputs(2674) <= layer2_outputs(7057);
    outputs(2675) <= (layer2_outputs(546)) xor (layer2_outputs(2819));
    outputs(2676) <= (layer2_outputs(9191)) xor (layer2_outputs(522));
    outputs(2677) <= not(layer2_outputs(1124));
    outputs(2678) <= layer2_outputs(5560);
    outputs(2679) <= (layer2_outputs(2900)) xor (layer2_outputs(1532));
    outputs(2680) <= not(layer2_outputs(1776)) or (layer2_outputs(290));
    outputs(2681) <= not(layer2_outputs(5863)) or (layer2_outputs(6306));
    outputs(2682) <= layer2_outputs(4309);
    outputs(2683) <= layer2_outputs(280);
    outputs(2684) <= not(layer2_outputs(8671));
    outputs(2685) <= not(layer2_outputs(7198));
    outputs(2686) <= layer2_outputs(3845);
    outputs(2687) <= (layer2_outputs(314)) xor (layer2_outputs(6253));
    outputs(2688) <= not(layer2_outputs(8197));
    outputs(2689) <= not(layer2_outputs(2132));
    outputs(2690) <= not(layer2_outputs(6));
    outputs(2691) <= (layer2_outputs(4873)) or (layer2_outputs(2846));
    outputs(2692) <= layer2_outputs(1337);
    outputs(2693) <= not(layer2_outputs(733));
    outputs(2694) <= not(layer2_outputs(1548));
    outputs(2695) <= not(layer2_outputs(8962));
    outputs(2696) <= (layer2_outputs(3268)) xor (layer2_outputs(8093));
    outputs(2697) <= layer2_outputs(7239);
    outputs(2698) <= layer2_outputs(4317);
    outputs(2699) <= layer2_outputs(5819);
    outputs(2700) <= layer2_outputs(3545);
    outputs(2701) <= not(layer2_outputs(8255));
    outputs(2702) <= layer2_outputs(3619);
    outputs(2703) <= not((layer2_outputs(8)) and (layer2_outputs(7086)));
    outputs(2704) <= layer2_outputs(3639);
    outputs(2705) <= not(layer2_outputs(2263)) or (layer2_outputs(2369));
    outputs(2706) <= not((layer2_outputs(4521)) xor (layer2_outputs(8827)));
    outputs(2707) <= not(layer2_outputs(241));
    outputs(2708) <= layer2_outputs(4924);
    outputs(2709) <= layer2_outputs(5272);
    outputs(2710) <= not((layer2_outputs(6248)) xor (layer2_outputs(1222)));
    outputs(2711) <= not(layer2_outputs(2105));
    outputs(2712) <= not(layer2_outputs(4840));
    outputs(2713) <= not(layer2_outputs(3654));
    outputs(2714) <= layer2_outputs(5338);
    outputs(2715) <= layer2_outputs(450);
    outputs(2716) <= not((layer2_outputs(1744)) xor (layer2_outputs(5974)));
    outputs(2717) <= (layer2_outputs(7638)) and (layer2_outputs(2719));
    outputs(2718) <= not(layer2_outputs(9295));
    outputs(2719) <= layer2_outputs(9528);
    outputs(2720) <= layer2_outputs(7256);
    outputs(2721) <= (layer2_outputs(53)) or (layer2_outputs(2382));
    outputs(2722) <= not(layer2_outputs(4164));
    outputs(2723) <= not(layer2_outputs(4265));
    outputs(2724) <= not(layer2_outputs(9361));
    outputs(2725) <= not(layer2_outputs(2131));
    outputs(2726) <= not(layer2_outputs(8117));
    outputs(2727) <= layer2_outputs(4705);
    outputs(2728) <= not(layer2_outputs(2472));
    outputs(2729) <= not(layer2_outputs(3139));
    outputs(2730) <= (layer2_outputs(9434)) xor (layer2_outputs(8521));
    outputs(2731) <= layer2_outputs(6346);
    outputs(2732) <= not(layer2_outputs(5276));
    outputs(2733) <= not((layer2_outputs(785)) xor (layer2_outputs(1281)));
    outputs(2734) <= (layer2_outputs(1129)) and not (layer2_outputs(7376));
    outputs(2735) <= not(layer2_outputs(7322));
    outputs(2736) <= not((layer2_outputs(8729)) xor (layer2_outputs(6875)));
    outputs(2737) <= layer2_outputs(6146);
    outputs(2738) <= not((layer2_outputs(1750)) xor (layer2_outputs(91)));
    outputs(2739) <= not(layer2_outputs(1243)) or (layer2_outputs(4151));
    outputs(2740) <= (layer2_outputs(9255)) xor (layer2_outputs(9686));
    outputs(2741) <= not(layer2_outputs(8593));
    outputs(2742) <= (layer2_outputs(2528)) xor (layer2_outputs(9499));
    outputs(2743) <= (layer2_outputs(3471)) and not (layer2_outputs(921));
    outputs(2744) <= not(layer2_outputs(2769));
    outputs(2745) <= not(layer2_outputs(5236)) or (layer2_outputs(3124));
    outputs(2746) <= not(layer2_outputs(10173));
    outputs(2747) <= not((layer2_outputs(5315)) xor (layer2_outputs(7800)));
    outputs(2748) <= not((layer2_outputs(6981)) xor (layer2_outputs(5442)));
    outputs(2749) <= layer2_outputs(6150);
    outputs(2750) <= (layer2_outputs(9978)) xor (layer2_outputs(5890));
    outputs(2751) <= not(layer2_outputs(4502)) or (layer2_outputs(7278));
    outputs(2752) <= not(layer2_outputs(8880));
    outputs(2753) <= not(layer2_outputs(7591));
    outputs(2754) <= not(layer2_outputs(2431));
    outputs(2755) <= not(layer2_outputs(5208));
    outputs(2756) <= layer2_outputs(8823);
    outputs(2757) <= (layer2_outputs(3874)) and (layer2_outputs(8121));
    outputs(2758) <= not(layer2_outputs(1005));
    outputs(2759) <= not(layer2_outputs(9390));
    outputs(2760) <= not((layer2_outputs(639)) or (layer2_outputs(4342)));
    outputs(2761) <= (layer2_outputs(6067)) xor (layer2_outputs(3041));
    outputs(2762) <= not(layer2_outputs(482));
    outputs(2763) <= not(layer2_outputs(9524));
    outputs(2764) <= layer2_outputs(4353);
    outputs(2765) <= layer2_outputs(8906);
    outputs(2766) <= not(layer2_outputs(3819));
    outputs(2767) <= not((layer2_outputs(7192)) xor (layer2_outputs(48)));
    outputs(2768) <= not(layer2_outputs(3402));
    outputs(2769) <= not(layer2_outputs(5089));
    outputs(2770) <= layer2_outputs(4845);
    outputs(2771) <= not(layer2_outputs(2038));
    outputs(2772) <= (layer2_outputs(2141)) xor (layer2_outputs(5512));
    outputs(2773) <= not((layer2_outputs(7083)) xor (layer2_outputs(9800)));
    outputs(2774) <= not(layer2_outputs(6597)) or (layer2_outputs(2923));
    outputs(2775) <= layer2_outputs(2037);
    outputs(2776) <= layer2_outputs(3018);
    outputs(2777) <= not((layer2_outputs(6451)) and (layer2_outputs(4260)));
    outputs(2778) <= not((layer2_outputs(2475)) and (layer2_outputs(957)));
    outputs(2779) <= layer2_outputs(10116);
    outputs(2780) <= not((layer2_outputs(2143)) xor (layer2_outputs(5710)));
    outputs(2781) <= (layer2_outputs(8594)) and not (layer2_outputs(2150));
    outputs(2782) <= not(layer2_outputs(7992));
    outputs(2783) <= not(layer2_outputs(6896));
    outputs(2784) <= not(layer2_outputs(1117));
    outputs(2785) <= layer2_outputs(1343);
    outputs(2786) <= not((layer2_outputs(265)) and (layer2_outputs(6948)));
    outputs(2787) <= not((layer2_outputs(4111)) and (layer2_outputs(1159)));
    outputs(2788) <= not(layer2_outputs(4837));
    outputs(2789) <= not((layer2_outputs(648)) or (layer2_outputs(5242)));
    outputs(2790) <= not(layer2_outputs(3175));
    outputs(2791) <= layer2_outputs(7957);
    outputs(2792) <= layer2_outputs(10009);
    outputs(2793) <= layer2_outputs(6427);
    outputs(2794) <= not(layer2_outputs(9655));
    outputs(2795) <= layer2_outputs(4963);
    outputs(2796) <= layer2_outputs(3568);
    outputs(2797) <= not(layer2_outputs(2827));
    outputs(2798) <= layer2_outputs(4611);
    outputs(2799) <= (layer2_outputs(1111)) or (layer2_outputs(1531));
    outputs(2800) <= not((layer2_outputs(8592)) xor (layer2_outputs(3972)));
    outputs(2801) <= not(layer2_outputs(10104));
    outputs(2802) <= layer2_outputs(8040);
    outputs(2803) <= (layer2_outputs(473)) or (layer2_outputs(2186));
    outputs(2804) <= layer2_outputs(7980);
    outputs(2805) <= not(layer2_outputs(5231)) or (layer2_outputs(3954));
    outputs(2806) <= not(layer2_outputs(3682));
    outputs(2807) <= not(layer2_outputs(2224));
    outputs(2808) <= (layer2_outputs(9047)) and not (layer2_outputs(4857));
    outputs(2809) <= layer2_outputs(2041);
    outputs(2810) <= not(layer2_outputs(7289));
    outputs(2811) <= (layer2_outputs(5542)) and not (layer2_outputs(6986));
    outputs(2812) <= layer2_outputs(6340);
    outputs(2813) <= not(layer2_outputs(9179));
    outputs(2814) <= (layer2_outputs(9922)) or (layer2_outputs(9194));
    outputs(2815) <= not(layer2_outputs(586));
    outputs(2816) <= (layer2_outputs(7823)) or (layer2_outputs(7530));
    outputs(2817) <= layer2_outputs(1355);
    outputs(2818) <= not(layer2_outputs(1626));
    outputs(2819) <= layer2_outputs(4949);
    outputs(2820) <= layer2_outputs(4999);
    outputs(2821) <= (layer2_outputs(8910)) xor (layer2_outputs(3590));
    outputs(2822) <= layer2_outputs(9792);
    outputs(2823) <= layer2_outputs(5628);
    outputs(2824) <= (layer2_outputs(8694)) and not (layer2_outputs(4155));
    outputs(2825) <= layer2_outputs(103);
    outputs(2826) <= not(layer2_outputs(7528)) or (layer2_outputs(5450));
    outputs(2827) <= layer2_outputs(9379);
    outputs(2828) <= (layer2_outputs(2972)) or (layer2_outputs(2380));
    outputs(2829) <= not((layer2_outputs(776)) xor (layer2_outputs(7474)));
    outputs(2830) <= layer2_outputs(7141);
    outputs(2831) <= layer2_outputs(8424);
    outputs(2832) <= (layer2_outputs(9703)) xor (layer2_outputs(10097));
    outputs(2833) <= not((layer2_outputs(9193)) and (layer2_outputs(10014)));
    outputs(2834) <= (layer2_outputs(6044)) xor (layer2_outputs(8577));
    outputs(2835) <= layer2_outputs(406);
    outputs(2836) <= layer2_outputs(3217);
    outputs(2837) <= (layer2_outputs(3596)) or (layer2_outputs(9603));
    outputs(2838) <= not(layer2_outputs(5320));
    outputs(2839) <= layer2_outputs(6985);
    outputs(2840) <= not(layer2_outputs(6804));
    outputs(2841) <= not(layer2_outputs(8700)) or (layer2_outputs(5067));
    outputs(2842) <= not(layer2_outputs(4508)) or (layer2_outputs(927));
    outputs(2843) <= layer2_outputs(8681);
    outputs(2844) <= layer2_outputs(3879);
    outputs(2845) <= layer2_outputs(1279);
    outputs(2846) <= not(layer2_outputs(5760));
    outputs(2847) <= layer2_outputs(8806);
    outputs(2848) <= (layer2_outputs(1719)) and (layer2_outputs(2004));
    outputs(2849) <= not(layer2_outputs(4277));
    outputs(2850) <= layer2_outputs(2882);
    outputs(2851) <= '1';
    outputs(2852) <= layer2_outputs(8061);
    outputs(2853) <= layer2_outputs(2793);
    outputs(2854) <= not(layer2_outputs(5426));
    outputs(2855) <= not(layer2_outputs(6109));
    outputs(2856) <= not(layer2_outputs(7402)) or (layer2_outputs(4770));
    outputs(2857) <= (layer2_outputs(2352)) and not (layer2_outputs(2580));
    outputs(2858) <= not(layer2_outputs(2174));
    outputs(2859) <= not(layer2_outputs(8496));
    outputs(2860) <= (layer2_outputs(9304)) xor (layer2_outputs(6736));
    outputs(2861) <= layer2_outputs(9990);
    outputs(2862) <= not(layer2_outputs(6935)) or (layer2_outputs(9816));
    outputs(2863) <= layer2_outputs(3044);
    outputs(2864) <= not(layer2_outputs(8712));
    outputs(2865) <= (layer2_outputs(9220)) xor (layer2_outputs(4501));
    outputs(2866) <= layer2_outputs(6132);
    outputs(2867) <= not(layer2_outputs(1632));
    outputs(2868) <= not(layer2_outputs(5013));
    outputs(2869) <= not((layer2_outputs(9674)) xor (layer2_outputs(8701)));
    outputs(2870) <= layer2_outputs(2238);
    outputs(2871) <= not(layer2_outputs(6614));
    outputs(2872) <= layer2_outputs(1672);
    outputs(2873) <= not((layer2_outputs(3722)) xor (layer2_outputs(6105)));
    outputs(2874) <= not((layer2_outputs(6302)) and (layer2_outputs(3611)));
    outputs(2875) <= not(layer2_outputs(1704));
    outputs(2876) <= (layer2_outputs(7481)) xor (layer2_outputs(2270));
    outputs(2877) <= not(layer2_outputs(7498));
    outputs(2878) <= not(layer2_outputs(4187)) or (layer2_outputs(9475));
    outputs(2879) <= (layer2_outputs(833)) xor (layer2_outputs(7401));
    outputs(2880) <= not((layer2_outputs(3588)) or (layer2_outputs(171)));
    outputs(2881) <= layer2_outputs(688);
    outputs(2882) <= layer2_outputs(9861);
    outputs(2883) <= layer2_outputs(8115);
    outputs(2884) <= layer2_outputs(8504);
    outputs(2885) <= not((layer2_outputs(4386)) and (layer2_outputs(8037)));
    outputs(2886) <= not(layer2_outputs(486));
    outputs(2887) <= not(layer2_outputs(6991));
    outputs(2888) <= not(layer2_outputs(7144));
    outputs(2889) <= not(layer2_outputs(7465));
    outputs(2890) <= not(layer2_outputs(8175));
    outputs(2891) <= not(layer2_outputs(3808));
    outputs(2892) <= not(layer2_outputs(9854));
    outputs(2893) <= layer2_outputs(2165);
    outputs(2894) <= layer2_outputs(8743);
    outputs(2895) <= (layer2_outputs(2744)) xor (layer2_outputs(265));
    outputs(2896) <= layer2_outputs(8501);
    outputs(2897) <= (layer2_outputs(1309)) or (layer2_outputs(4415));
    outputs(2898) <= layer2_outputs(1039);
    outputs(2899) <= not(layer2_outputs(8551));
    outputs(2900) <= (layer2_outputs(8841)) xor (layer2_outputs(6339));
    outputs(2901) <= (layer2_outputs(2033)) and (layer2_outputs(8678));
    outputs(2902) <= layer2_outputs(895);
    outputs(2903) <= not(layer2_outputs(9772));
    outputs(2904) <= layer2_outputs(8413);
    outputs(2905) <= layer2_outputs(4429);
    outputs(2906) <= not(layer2_outputs(8020));
    outputs(2907) <= layer2_outputs(1337);
    outputs(2908) <= layer2_outputs(7890);
    outputs(2909) <= not(layer2_outputs(10050));
    outputs(2910) <= not(layer2_outputs(9232));
    outputs(2911) <= not(layer2_outputs(5153));
    outputs(2912) <= not(layer2_outputs(8080));
    outputs(2913) <= not(layer2_outputs(3112));
    outputs(2914) <= layer2_outputs(7099);
    outputs(2915) <= not(layer2_outputs(504));
    outputs(2916) <= not((layer2_outputs(5212)) xor (layer2_outputs(8379)));
    outputs(2917) <= not(layer2_outputs(897));
    outputs(2918) <= not((layer2_outputs(5059)) xor (layer2_outputs(1963)));
    outputs(2919) <= (layer2_outputs(2194)) and (layer2_outputs(9973));
    outputs(2920) <= not(layer2_outputs(5517));
    outputs(2921) <= (layer2_outputs(4321)) xor (layer2_outputs(7917));
    outputs(2922) <= not((layer2_outputs(8432)) xor (layer2_outputs(9183)));
    outputs(2923) <= not(layer2_outputs(3141));
    outputs(2924) <= (layer2_outputs(5878)) xor (layer2_outputs(9886));
    outputs(2925) <= layer2_outputs(5009);
    outputs(2926) <= not(layer2_outputs(6461)) or (layer2_outputs(8768));
    outputs(2927) <= layer2_outputs(1514);
    outputs(2928) <= layer2_outputs(3833);
    outputs(2929) <= layer2_outputs(2982);
    outputs(2930) <= (layer2_outputs(6654)) xor (layer2_outputs(5761));
    outputs(2931) <= not(layer2_outputs(5810));
    outputs(2932) <= (layer2_outputs(9939)) and not (layer2_outputs(3566));
    outputs(2933) <= (layer2_outputs(3318)) and not (layer2_outputs(1089));
    outputs(2934) <= not(layer2_outputs(1609));
    outputs(2935) <= not(layer2_outputs(9494));
    outputs(2936) <= not(layer2_outputs(5972)) or (layer2_outputs(7983));
    outputs(2937) <= layer2_outputs(2804);
    outputs(2938) <= not(layer2_outputs(3988)) or (layer2_outputs(6596));
    outputs(2939) <= layer2_outputs(2969);
    outputs(2940) <= not((layer2_outputs(5972)) xor (layer2_outputs(6251)));
    outputs(2941) <= not(layer2_outputs(690));
    outputs(2942) <= not((layer2_outputs(1720)) xor (layer2_outputs(7359)));
    outputs(2943) <= not(layer2_outputs(5559));
    outputs(2944) <= not(layer2_outputs(2187));
    outputs(2945) <= not(layer2_outputs(3167));
    outputs(2946) <= layer2_outputs(9246);
    outputs(2947) <= layer2_outputs(7855);
    outputs(2948) <= not(layer2_outputs(7991));
    outputs(2949) <= not(layer2_outputs(9416));
    outputs(2950) <= not(layer2_outputs(7408));
    outputs(2951) <= not((layer2_outputs(3996)) and (layer2_outputs(7603)));
    outputs(2952) <= (layer2_outputs(8110)) and not (layer2_outputs(10069));
    outputs(2953) <= not(layer2_outputs(2174));
    outputs(2954) <= not(layer2_outputs(7783));
    outputs(2955) <= (layer2_outputs(5861)) or (layer2_outputs(9706));
    outputs(2956) <= layer2_outputs(5820);
    outputs(2957) <= not(layer2_outputs(7715));
    outputs(2958) <= layer2_outputs(9067);
    outputs(2959) <= (layer2_outputs(1445)) or (layer2_outputs(9009));
    outputs(2960) <= (layer2_outputs(8459)) and not (layer2_outputs(5052));
    outputs(2961) <= not(layer2_outputs(7873));
    outputs(2962) <= layer2_outputs(3246);
    outputs(2963) <= layer2_outputs(4995);
    outputs(2964) <= not(layer2_outputs(4635));
    outputs(2965) <= not(layer2_outputs(8496));
    outputs(2966) <= layer2_outputs(8583);
    outputs(2967) <= not(layer2_outputs(2878));
    outputs(2968) <= (layer2_outputs(5051)) xor (layer2_outputs(1109));
    outputs(2969) <= not(layer2_outputs(5759));
    outputs(2970) <= layer2_outputs(523);
    outputs(2971) <= layer2_outputs(8806);
    outputs(2972) <= not(layer2_outputs(5919)) or (layer2_outputs(8591));
    outputs(2973) <= layer2_outputs(3232);
    outputs(2974) <= not((layer2_outputs(7473)) and (layer2_outputs(6710)));
    outputs(2975) <= (layer2_outputs(7049)) xor (layer2_outputs(6297));
    outputs(2976) <= layer2_outputs(3146);
    outputs(2977) <= layer2_outputs(1511);
    outputs(2978) <= layer2_outputs(8464);
    outputs(2979) <= layer2_outputs(1703);
    outputs(2980) <= not((layer2_outputs(3563)) xor (layer2_outputs(2280)));
    outputs(2981) <= not((layer2_outputs(5502)) xor (layer2_outputs(1181)));
    outputs(2982) <= not(layer2_outputs(3850));
    outputs(2983) <= not((layer2_outputs(2319)) and (layer2_outputs(9422)));
    outputs(2984) <= not(layer2_outputs(7837));
    outputs(2985) <= (layer2_outputs(9580)) and not (layer2_outputs(6973));
    outputs(2986) <= layer2_outputs(9775);
    outputs(2987) <= not(layer2_outputs(1961));
    outputs(2988) <= not(layer2_outputs(1580));
    outputs(2989) <= not(layer2_outputs(819));
    outputs(2990) <= layer2_outputs(4785);
    outputs(2991) <= (layer2_outputs(7369)) and not (layer2_outputs(5436));
    outputs(2992) <= layer2_outputs(8334);
    outputs(2993) <= layer2_outputs(6217);
    outputs(2994) <= layer2_outputs(6909);
    outputs(2995) <= not(layer2_outputs(3705));
    outputs(2996) <= layer2_outputs(2087);
    outputs(2997) <= layer2_outputs(7042);
    outputs(2998) <= not(layer2_outputs(4594));
    outputs(2999) <= layer2_outputs(8410);
    outputs(3000) <= layer2_outputs(6988);
    outputs(3001) <= not(layer2_outputs(9211));
    outputs(3002) <= layer2_outputs(1027);
    outputs(3003) <= not(layer2_outputs(5313));
    outputs(3004) <= not(layer2_outputs(3370));
    outputs(3005) <= (layer2_outputs(3583)) xor (layer2_outputs(4599));
    outputs(3006) <= not(layer2_outputs(4610)) or (layer2_outputs(7602));
    outputs(3007) <= layer2_outputs(2594);
    outputs(3008) <= layer2_outputs(855);
    outputs(3009) <= layer2_outputs(94);
    outputs(3010) <= not((layer2_outputs(4282)) xor (layer2_outputs(2529)));
    outputs(3011) <= layer2_outputs(4080);
    outputs(3012) <= layer2_outputs(1843);
    outputs(3013) <= layer2_outputs(7842);
    outputs(3014) <= layer2_outputs(1553);
    outputs(3015) <= (layer2_outputs(7923)) or (layer2_outputs(2430));
    outputs(3016) <= layer2_outputs(767);
    outputs(3017) <= not(layer2_outputs(5226));
    outputs(3018) <= not(layer2_outputs(783));
    outputs(3019) <= layer2_outputs(9883);
    outputs(3020) <= not((layer2_outputs(1628)) xor (layer2_outputs(5266)));
    outputs(3021) <= layer2_outputs(5201);
    outputs(3022) <= not((layer2_outputs(6701)) or (layer2_outputs(8564)));
    outputs(3023) <= layer2_outputs(5230);
    outputs(3024) <= layer2_outputs(9469);
    outputs(3025) <= (layer2_outputs(3021)) xor (layer2_outputs(9539));
    outputs(3026) <= not((layer2_outputs(8264)) xor (layer2_outputs(7401)));
    outputs(3027) <= not(layer2_outputs(1591)) or (layer2_outputs(280));
    outputs(3028) <= not(layer2_outputs(6096));
    outputs(3029) <= not(layer2_outputs(2135));
    outputs(3030) <= (layer2_outputs(5843)) and (layer2_outputs(3696));
    outputs(3031) <= (layer2_outputs(8063)) or (layer2_outputs(6053));
    outputs(3032) <= (layer2_outputs(3346)) xor (layer2_outputs(4237));
    outputs(3033) <= layer2_outputs(4592);
    outputs(3034) <= layer2_outputs(6233);
    outputs(3035) <= layer2_outputs(9888);
    outputs(3036) <= (layer2_outputs(1194)) xor (layer2_outputs(135));
    outputs(3037) <= not(layer2_outputs(6304));
    outputs(3038) <= (layer2_outputs(8641)) xor (layer2_outputs(6640));
    outputs(3039) <= not(layer2_outputs(6593)) or (layer2_outputs(2145));
    outputs(3040) <= not(layer2_outputs(1996)) or (layer2_outputs(4425));
    outputs(3041) <= layer2_outputs(2300);
    outputs(3042) <= (layer2_outputs(6652)) and (layer2_outputs(7691));
    outputs(3043) <= layer2_outputs(9951);
    outputs(3044) <= not(layer2_outputs(3141));
    outputs(3045) <= not(layer2_outputs(6665));
    outputs(3046) <= (layer2_outputs(7551)) or (layer2_outputs(3884));
    outputs(3047) <= not(layer2_outputs(4043));
    outputs(3048) <= not(layer2_outputs(2929));
    outputs(3049) <= not(layer2_outputs(1005)) or (layer2_outputs(8672));
    outputs(3050) <= not((layer2_outputs(3752)) or (layer2_outputs(4141)));
    outputs(3051) <= (layer2_outputs(5852)) xor (layer2_outputs(8384));
    outputs(3052) <= not(layer2_outputs(6222)) or (layer2_outputs(6260));
    outputs(3053) <= not(layer2_outputs(3319)) or (layer2_outputs(6309));
    outputs(3054) <= not(layer2_outputs(108));
    outputs(3055) <= layer2_outputs(4457);
    outputs(3056) <= (layer2_outputs(4523)) and not (layer2_outputs(8037));
    outputs(3057) <= not(layer2_outputs(5802)) or (layer2_outputs(9975));
    outputs(3058) <= (layer2_outputs(3368)) and not (layer2_outputs(2153));
    outputs(3059) <= layer2_outputs(8044);
    outputs(3060) <= not(layer2_outputs(7091)) or (layer2_outputs(7648));
    outputs(3061) <= not(layer2_outputs(7140));
    outputs(3062) <= not((layer2_outputs(7044)) xor (layer2_outputs(7941)));
    outputs(3063) <= not(layer2_outputs(6836));
    outputs(3064) <= not(layer2_outputs(4391));
    outputs(3065) <= layer2_outputs(6953);
    outputs(3066) <= not((layer2_outputs(6917)) xor (layer2_outputs(3277)));
    outputs(3067) <= (layer2_outputs(2406)) xor (layer2_outputs(3437));
    outputs(3068) <= not((layer2_outputs(7332)) xor (layer2_outputs(474)));
    outputs(3069) <= not(layer2_outputs(1918));
    outputs(3070) <= not(layer2_outputs(1541));
    outputs(3071) <= not(layer2_outputs(1114));
    outputs(3072) <= not(layer2_outputs(3841));
    outputs(3073) <= layer2_outputs(7701);
    outputs(3074) <= layer2_outputs(4291);
    outputs(3075) <= (layer2_outputs(5876)) and not (layer2_outputs(8633));
    outputs(3076) <= layer2_outputs(4210);
    outputs(3077) <= not(layer2_outputs(6610));
    outputs(3078) <= layer2_outputs(5501);
    outputs(3079) <= (layer2_outputs(7419)) xor (layer2_outputs(7947));
    outputs(3080) <= layer2_outputs(5390);
    outputs(3081) <= not((layer2_outputs(8986)) xor (layer2_outputs(9766)));
    outputs(3082) <= layer2_outputs(1377);
    outputs(3083) <= layer2_outputs(5544);
    outputs(3084) <= not(layer2_outputs(5494));
    outputs(3085) <= (layer2_outputs(624)) xor (layer2_outputs(1971));
    outputs(3086) <= (layer2_outputs(1683)) xor (layer2_outputs(1883));
    outputs(3087) <= layer2_outputs(1248);
    outputs(3088) <= not((layer2_outputs(5768)) xor (layer2_outputs(1019)));
    outputs(3089) <= layer2_outputs(949);
    outputs(3090) <= layer2_outputs(4217);
    outputs(3091) <= not(layer2_outputs(5086));
    outputs(3092) <= layer2_outputs(6521);
    outputs(3093) <= layer2_outputs(4419);
    outputs(3094) <= not(layer2_outputs(4585));
    outputs(3095) <= layer2_outputs(8228);
    outputs(3096) <= not(layer2_outputs(6674));
    outputs(3097) <= not((layer2_outputs(5330)) xor (layer2_outputs(9054)));
    outputs(3098) <= not(layer2_outputs(2857));
    outputs(3099) <= not(layer2_outputs(7426));
    outputs(3100) <= not(layer2_outputs(1395));
    outputs(3101) <= (layer2_outputs(8875)) xor (layer2_outputs(4754));
    outputs(3102) <= not((layer2_outputs(8991)) and (layer2_outputs(5508)));
    outputs(3103) <= layer2_outputs(4918);
    outputs(3104) <= not((layer2_outputs(9594)) xor (layer2_outputs(2658)));
    outputs(3105) <= layer2_outputs(5078);
    outputs(3106) <= layer2_outputs(3436);
    outputs(3107) <= not(layer2_outputs(861));
    outputs(3108) <= not((layer2_outputs(2561)) xor (layer2_outputs(4899)));
    outputs(3109) <= not(layer2_outputs(1646));
    outputs(3110) <= (layer2_outputs(5011)) xor (layer2_outputs(1637));
    outputs(3111) <= not((layer2_outputs(5172)) xor (layer2_outputs(1092)));
    outputs(3112) <= (layer2_outputs(8631)) xor (layer2_outputs(139));
    outputs(3113) <= layer2_outputs(1439);
    outputs(3114) <= layer2_outputs(3863);
    outputs(3115) <= not(layer2_outputs(7694));
    outputs(3116) <= not(layer2_outputs(5860));
    outputs(3117) <= (layer2_outputs(9753)) xor (layer2_outputs(4470));
    outputs(3118) <= not((layer2_outputs(4759)) and (layer2_outputs(7441)));
    outputs(3119) <= layer2_outputs(8918);
    outputs(3120) <= not((layer2_outputs(4651)) xor (layer2_outputs(1736)));
    outputs(3121) <= layer2_outputs(9292);
    outputs(3122) <= (layer2_outputs(3617)) xor (layer2_outputs(5913));
    outputs(3123) <= not(layer2_outputs(1153));
    outputs(3124) <= layer2_outputs(8978);
    outputs(3125) <= (layer2_outputs(910)) and (layer2_outputs(5119));
    outputs(3126) <= not((layer2_outputs(9854)) or (layer2_outputs(7620)));
    outputs(3127) <= layer2_outputs(1828);
    outputs(3128) <= not(layer2_outputs(877));
    outputs(3129) <= not(layer2_outputs(7761));
    outputs(3130) <= not(layer2_outputs(9711));
    outputs(3131) <= not(layer2_outputs(5359));
    outputs(3132) <= not((layer2_outputs(1165)) xor (layer2_outputs(3316)));
    outputs(3133) <= layer2_outputs(897);
    outputs(3134) <= not(layer2_outputs(5503));
    outputs(3135) <= not((layer2_outputs(2528)) xor (layer2_outputs(519)));
    outputs(3136) <= not(layer2_outputs(6645));
    outputs(3137) <= not(layer2_outputs(1974));
    outputs(3138) <= layer2_outputs(2029);
    outputs(3139) <= not(layer2_outputs(6972));
    outputs(3140) <= (layer2_outputs(5706)) xor (layer2_outputs(83));
    outputs(3141) <= layer2_outputs(4922);
    outputs(3142) <= (layer2_outputs(2419)) xor (layer2_outputs(2768));
    outputs(3143) <= not(layer2_outputs(7292));
    outputs(3144) <= layer2_outputs(802);
    outputs(3145) <= layer2_outputs(2508);
    outputs(3146) <= not(layer2_outputs(391));
    outputs(3147) <= not((layer2_outputs(6639)) xor (layer2_outputs(8250)));
    outputs(3148) <= (layer2_outputs(4392)) and not (layer2_outputs(2946));
    outputs(3149) <= layer2_outputs(639);
    outputs(3150) <= layer2_outputs(7697);
    outputs(3151) <= (layer2_outputs(9590)) and not (layer2_outputs(8791));
    outputs(3152) <= layer2_outputs(4624);
    outputs(3153) <= not(layer2_outputs(9131));
    outputs(3154) <= not(layer2_outputs(1582));
    outputs(3155) <= (layer2_outputs(5196)) and not (layer2_outputs(2666));
    outputs(3156) <= layer2_outputs(838);
    outputs(3157) <= not(layer2_outputs(3152));
    outputs(3158) <= layer2_outputs(10218);
    outputs(3159) <= (layer2_outputs(7307)) xor (layer2_outputs(7338));
    outputs(3160) <= not(layer2_outputs(2604));
    outputs(3161) <= layer2_outputs(2313);
    outputs(3162) <= not(layer2_outputs(8117));
    outputs(3163) <= layer2_outputs(6016);
    outputs(3164) <= not(layer2_outputs(4058));
    outputs(3165) <= not(layer2_outputs(8510));
    outputs(3166) <= not(layer2_outputs(3384));
    outputs(3167) <= not(layer2_outputs(4063));
    outputs(3168) <= layer2_outputs(8519);
    outputs(3169) <= not(layer2_outputs(1956));
    outputs(3170) <= layer2_outputs(10064);
    outputs(3171) <= not(layer2_outputs(1651));
    outputs(3172) <= not(layer2_outputs(1831));
    outputs(3173) <= not((layer2_outputs(592)) xor (layer2_outputs(9175)));
    outputs(3174) <= layer2_outputs(10074);
    outputs(3175) <= not(layer2_outputs(5888)) or (layer2_outputs(6162));
    outputs(3176) <= (layer2_outputs(1786)) xor (layer2_outputs(9527));
    outputs(3177) <= not(layer2_outputs(5727));
    outputs(3178) <= layer2_outputs(7926);
    outputs(3179) <= not((layer2_outputs(6271)) xor (layer2_outputs(3260)));
    outputs(3180) <= not((layer2_outputs(4811)) xor (layer2_outputs(377)));
    outputs(3181) <= layer2_outputs(4101);
    outputs(3182) <= (layer2_outputs(5054)) and not (layer2_outputs(9664));
    outputs(3183) <= (layer2_outputs(3377)) xor (layer2_outputs(6331));
    outputs(3184) <= not(layer2_outputs(4201));
    outputs(3185) <= layer2_outputs(177);
    outputs(3186) <= (layer2_outputs(9474)) and (layer2_outputs(7852));
    outputs(3187) <= not((layer2_outputs(3827)) xor (layer2_outputs(9366)));
    outputs(3188) <= not((layer2_outputs(7736)) xor (layer2_outputs(1291)));
    outputs(3189) <= layer2_outputs(4559);
    outputs(3190) <= not(layer2_outputs(7721));
    outputs(3191) <= not((layer2_outputs(5701)) xor (layer2_outputs(2721)));
    outputs(3192) <= layer2_outputs(6973);
    outputs(3193) <= not((layer2_outputs(507)) xor (layer2_outputs(2206)));
    outputs(3194) <= layer2_outputs(7008);
    outputs(3195) <= layer2_outputs(5341);
    outputs(3196) <= layer2_outputs(3116);
    outputs(3197) <= not(layer2_outputs(5721));
    outputs(3198) <= not(layer2_outputs(8688));
    outputs(3199) <= layer2_outputs(5808);
    outputs(3200) <= not(layer2_outputs(9158));
    outputs(3201) <= not(layer2_outputs(9588));
    outputs(3202) <= layer2_outputs(1954);
    outputs(3203) <= not(layer2_outputs(4544));
    outputs(3204) <= (layer2_outputs(2662)) xor (layer2_outputs(2407));
    outputs(3205) <= layer2_outputs(1079);
    outputs(3206) <= not(layer2_outputs(9022));
    outputs(3207) <= not(layer2_outputs(6048));
    outputs(3208) <= not((layer2_outputs(6420)) and (layer2_outputs(1240)));
    outputs(3209) <= not((layer2_outputs(6170)) xor (layer2_outputs(6613)));
    outputs(3210) <= not(layer2_outputs(6911));
    outputs(3211) <= layer2_outputs(7442);
    outputs(3212) <= layer2_outputs(7754);
    outputs(3213) <= not(layer2_outputs(10217));
    outputs(3214) <= layer2_outputs(3076);
    outputs(3215) <= layer2_outputs(3939);
    outputs(3216) <= layer2_outputs(5311);
    outputs(3217) <= not(layer2_outputs(9278));
    outputs(3218) <= layer2_outputs(2042);
    outputs(3219) <= not(layer2_outputs(4311));
    outputs(3220) <= not(layer2_outputs(9786));
    outputs(3221) <= layer2_outputs(9567);
    outputs(3222) <= not(layer2_outputs(7673));
    outputs(3223) <= layer2_outputs(2158);
    outputs(3224) <= not(layer2_outputs(8082));
    outputs(3225) <= (layer2_outputs(6901)) xor (layer2_outputs(10052));
    outputs(3226) <= not((layer2_outputs(7651)) xor (layer2_outputs(3163)));
    outputs(3227) <= layer2_outputs(6974);
    outputs(3228) <= layer2_outputs(3265);
    outputs(3229) <= not((layer2_outputs(1447)) xor (layer2_outputs(1768)));
    outputs(3230) <= layer2_outputs(3860);
    outputs(3231) <= layer2_outputs(5357);
    outputs(3232) <= not(layer2_outputs(5661));
    outputs(3233) <= not(layer2_outputs(7460));
    outputs(3234) <= not(layer2_outputs(2653));
    outputs(3235) <= (layer2_outputs(1233)) or (layer2_outputs(1753));
    outputs(3236) <= not(layer2_outputs(2383));
    outputs(3237) <= layer2_outputs(8611);
    outputs(3238) <= not(layer2_outputs(3823));
    outputs(3239) <= not(layer2_outputs(5704));
    outputs(3240) <= not(layer2_outputs(8952));
    outputs(3241) <= (layer2_outputs(8470)) xor (layer2_outputs(1868));
    outputs(3242) <= not(layer2_outputs(1275));
    outputs(3243) <= not(layer2_outputs(4654));
    outputs(3244) <= (layer2_outputs(7669)) xor (layer2_outputs(2131));
    outputs(3245) <= not(layer2_outputs(8090));
    outputs(3246) <= not(layer2_outputs(9428));
    outputs(3247) <= (layer2_outputs(2388)) xor (layer2_outputs(3270));
    outputs(3248) <= not(layer2_outputs(6630));
    outputs(3249) <= '0';
    outputs(3250) <= not(layer2_outputs(1250));
    outputs(3251) <= not((layer2_outputs(6957)) xor (layer2_outputs(902)));
    outputs(3252) <= not(layer2_outputs(4628));
    outputs(3253) <= layer2_outputs(6753);
    outputs(3254) <= (layer2_outputs(1068)) and (layer2_outputs(5035));
    outputs(3255) <= (layer2_outputs(2515)) xor (layer2_outputs(3765));
    outputs(3256) <= (layer2_outputs(7810)) xor (layer2_outputs(4075));
    outputs(3257) <= (layer2_outputs(418)) or (layer2_outputs(8942));
    outputs(3258) <= not((layer2_outputs(5728)) xor (layer2_outputs(1204)));
    outputs(3259) <= layer2_outputs(6525);
    outputs(3260) <= (layer2_outputs(6053)) xor (layer2_outputs(5841));
    outputs(3261) <= layer2_outputs(7048);
    outputs(3262) <= not(layer2_outputs(8576));
    outputs(3263) <= (layer2_outputs(6038)) and not (layer2_outputs(9348));
    outputs(3264) <= layer2_outputs(6413);
    outputs(3265) <= not(layer2_outputs(5157));
    outputs(3266) <= layer2_outputs(6515);
    outputs(3267) <= (layer2_outputs(5312)) xor (layer2_outputs(9271));
    outputs(3268) <= (layer2_outputs(8374)) xor (layer2_outputs(2325));
    outputs(3269) <= layer2_outputs(753);
    outputs(3270) <= not(layer2_outputs(8951));
    outputs(3271) <= not(layer2_outputs(7602));
    outputs(3272) <= not(layer2_outputs(3454));
    outputs(3273) <= not(layer2_outputs(2351));
    outputs(3274) <= (layer2_outputs(3827)) and not (layer2_outputs(21));
    outputs(3275) <= layer2_outputs(8598);
    outputs(3276) <= (layer2_outputs(1521)) xor (layer2_outputs(7979));
    outputs(3277) <= (layer2_outputs(6399)) or (layer2_outputs(1073));
    outputs(3278) <= not(layer2_outputs(5156));
    outputs(3279) <= not((layer2_outputs(6771)) or (layer2_outputs(6309)));
    outputs(3280) <= not(layer2_outputs(10148));
    outputs(3281) <= layer2_outputs(8600);
    outputs(3282) <= layer2_outputs(5589);
    outputs(3283) <= not(layer2_outputs(8743));
    outputs(3284) <= layer2_outputs(3449);
    outputs(3285) <= not((layer2_outputs(7283)) xor (layer2_outputs(6385)));
    outputs(3286) <= layer2_outputs(4017);
    outputs(3287) <= (layer2_outputs(9863)) xor (layer2_outputs(4894));
    outputs(3288) <= not((layer2_outputs(8304)) or (layer2_outputs(930)));
    outputs(3289) <= (layer2_outputs(5145)) and not (layer2_outputs(4496));
    outputs(3290) <= layer2_outputs(6330);
    outputs(3291) <= not(layer2_outputs(1436));
    outputs(3292) <= (layer2_outputs(7450)) and not (layer2_outputs(3727));
    outputs(3293) <= (layer2_outputs(9377)) and not (layer2_outputs(2354));
    outputs(3294) <= not(layer2_outputs(2702));
    outputs(3295) <= layer2_outputs(7775);
    outputs(3296) <= layer2_outputs(7674);
    outputs(3297) <= layer2_outputs(5140);
    outputs(3298) <= layer2_outputs(7785);
    outputs(3299) <= not(layer2_outputs(2482));
    outputs(3300) <= (layer2_outputs(3381)) or (layer2_outputs(5513));
    outputs(3301) <= not((layer2_outputs(3769)) or (layer2_outputs(8365)));
    outputs(3302) <= (layer2_outputs(9901)) xor (layer2_outputs(5715));
    outputs(3303) <= layer2_outputs(5698);
    outputs(3304) <= not(layer2_outputs(4730));
    outputs(3305) <= not(layer2_outputs(1574));
    outputs(3306) <= not(layer2_outputs(2682));
    outputs(3307) <= not(layer2_outputs(4930));
    outputs(3308) <= layer2_outputs(191);
    outputs(3309) <= not(layer2_outputs(7111));
    outputs(3310) <= (layer2_outputs(1357)) and not (layer2_outputs(1561));
    outputs(3311) <= (layer2_outputs(6753)) xor (layer2_outputs(9898));
    outputs(3312) <= not(layer2_outputs(2956));
    outputs(3313) <= (layer2_outputs(2886)) and not (layer2_outputs(3079));
    outputs(3314) <= layer2_outputs(3209);
    outputs(3315) <= layer2_outputs(6332);
    outputs(3316) <= layer2_outputs(89);
    outputs(3317) <= not(layer2_outputs(953));
    outputs(3318) <= layer2_outputs(1391);
    outputs(3319) <= not((layer2_outputs(5285)) or (layer2_outputs(7568)));
    outputs(3320) <= (layer2_outputs(4936)) and not (layer2_outputs(4566));
    outputs(3321) <= not((layer2_outputs(10199)) xor (layer2_outputs(2050)));
    outputs(3322) <= layer2_outputs(6238);
    outputs(3323) <= not(layer2_outputs(5223));
    outputs(3324) <= layer2_outputs(2224);
    outputs(3325) <= (layer2_outputs(8336)) xor (layer2_outputs(8000));
    outputs(3326) <= layer2_outputs(5149);
    outputs(3327) <= layer2_outputs(422);
    outputs(3328) <= not((layer2_outputs(4930)) xor (layer2_outputs(1134)));
    outputs(3329) <= not(layer2_outputs(1120));
    outputs(3330) <= not(layer2_outputs(3126));
    outputs(3331) <= layer2_outputs(9575);
    outputs(3332) <= layer2_outputs(1077);
    outputs(3333) <= not(layer2_outputs(5146));
    outputs(3334) <= not(layer2_outputs(8585));
    outputs(3335) <= not(layer2_outputs(8490));
    outputs(3336) <= (layer2_outputs(7257)) and not (layer2_outputs(8305));
    outputs(3337) <= layer2_outputs(8245);
    outputs(3338) <= not(layer2_outputs(8763));
    outputs(3339) <= layer2_outputs(3637);
    outputs(3340) <= layer2_outputs(9150);
    outputs(3341) <= not(layer2_outputs(7246));
    outputs(3342) <= not(layer2_outputs(2814)) or (layer2_outputs(9490));
    outputs(3343) <= not(layer2_outputs(5461));
    outputs(3344) <= (layer2_outputs(7070)) and not (layer2_outputs(2017));
    outputs(3345) <= (layer2_outputs(7274)) and not (layer2_outputs(1195));
    outputs(3346) <= not(layer2_outputs(5892));
    outputs(3347) <= not((layer2_outputs(3328)) xor (layer2_outputs(8218)));
    outputs(3348) <= not((layer2_outputs(7827)) and (layer2_outputs(8879)));
    outputs(3349) <= layer2_outputs(1522);
    outputs(3350) <= layer2_outputs(5427);
    outputs(3351) <= not(layer2_outputs(9923));
    outputs(3352) <= not(layer2_outputs(8095));
    outputs(3353) <= not((layer2_outputs(3967)) xor (layer2_outputs(7228)));
    outputs(3354) <= not(layer2_outputs(9048));
    outputs(3355) <= layer2_outputs(1928);
    outputs(3356) <= (layer2_outputs(832)) and not (layer2_outputs(4176));
    outputs(3357) <= (layer2_outputs(4227)) xor (layer2_outputs(1497));
    outputs(3358) <= not(layer2_outputs(392));
    outputs(3359) <= layer2_outputs(327);
    outputs(3360) <= not((layer2_outputs(7084)) and (layer2_outputs(4554)));
    outputs(3361) <= not(layer2_outputs(3088));
    outputs(3362) <= layer2_outputs(3127);
    outputs(3363) <= (layer2_outputs(4059)) xor (layer2_outputs(2635));
    outputs(3364) <= (layer2_outputs(8937)) xor (layer2_outputs(7609));
    outputs(3365) <= not(layer2_outputs(5630));
    outputs(3366) <= not((layer2_outputs(4787)) xor (layer2_outputs(6001)));
    outputs(3367) <= (layer2_outputs(3516)) xor (layer2_outputs(7792));
    outputs(3368) <= layer2_outputs(448);
    outputs(3369) <= (layer2_outputs(3834)) and not (layer2_outputs(2547));
    outputs(3370) <= not(layer2_outputs(6592)) or (layer2_outputs(7558));
    outputs(3371) <= not(layer2_outputs(4595));
    outputs(3372) <= not(layer2_outputs(2655));
    outputs(3373) <= layer2_outputs(4996);
    outputs(3374) <= (layer2_outputs(10237)) xor (layer2_outputs(7660));
    outputs(3375) <= layer2_outputs(1726);
    outputs(3376) <= layer2_outputs(3330);
    outputs(3377) <= layer2_outputs(2795);
    outputs(3378) <= not((layer2_outputs(5742)) and (layer2_outputs(5872)));
    outputs(3379) <= layer2_outputs(1813);
    outputs(3380) <= (layer2_outputs(1587)) xor (layer2_outputs(2129));
    outputs(3381) <= not(layer2_outputs(7467));
    outputs(3382) <= layer2_outputs(1717);
    outputs(3383) <= layer2_outputs(1572);
    outputs(3384) <= layer2_outputs(3073);
    outputs(3385) <= not(layer2_outputs(6614));
    outputs(3386) <= (layer2_outputs(1461)) xor (layer2_outputs(2675));
    outputs(3387) <= not((layer2_outputs(3939)) xor (layer2_outputs(8366)));
    outputs(3388) <= (layer2_outputs(5978)) xor (layer2_outputs(3128));
    outputs(3389) <= not(layer2_outputs(10083));
    outputs(3390) <= layer2_outputs(9647);
    outputs(3391) <= (layer2_outputs(7351)) xor (layer2_outputs(3776));
    outputs(3392) <= (layer2_outputs(9038)) xor (layer2_outputs(8747));
    outputs(3393) <= not((layer2_outputs(4683)) xor (layer2_outputs(8168)));
    outputs(3394) <= not((layer2_outputs(1280)) xor (layer2_outputs(9054)));
    outputs(3395) <= (layer2_outputs(9088)) xor (layer2_outputs(4294));
    outputs(3396) <= layer2_outputs(8869);
    outputs(3397) <= not(layer2_outputs(1866));
    outputs(3398) <= layer2_outputs(3775);
    outputs(3399) <= layer2_outputs(5340);
    outputs(3400) <= not(layer2_outputs(7205));
    outputs(3401) <= layer2_outputs(7538);
    outputs(3402) <= not((layer2_outputs(1917)) xor (layer2_outputs(5181)));
    outputs(3403) <= layer2_outputs(8936);
    outputs(3404) <= layer2_outputs(2895);
    outputs(3405) <= (layer2_outputs(3357)) xor (layer2_outputs(3579));
    outputs(3406) <= not((layer2_outputs(2473)) or (layer2_outputs(9558)));
    outputs(3407) <= layer2_outputs(8097);
    outputs(3408) <= layer2_outputs(7346);
    outputs(3409) <= not((layer2_outputs(7782)) or (layer2_outputs(906)));
    outputs(3410) <= layer2_outputs(6889);
    outputs(3411) <= not(layer2_outputs(6492));
    outputs(3412) <= layer2_outputs(7543);
    outputs(3413) <= (layer2_outputs(7091)) and not (layer2_outputs(4391));
    outputs(3414) <= not(layer2_outputs(1550));
    outputs(3415) <= layer2_outputs(4576);
    outputs(3416) <= layer2_outputs(1677);
    outputs(3417) <= layer2_outputs(5992);
    outputs(3418) <= not((layer2_outputs(9764)) and (layer2_outputs(8774)));
    outputs(3419) <= layer2_outputs(4220);
    outputs(3420) <= not((layer2_outputs(2764)) xor (layer2_outputs(259)));
    outputs(3421) <= not(layer2_outputs(8083));
    outputs(3422) <= not(layer2_outputs(1189));
    outputs(3423) <= not(layer2_outputs(9149));
    outputs(3424) <= layer2_outputs(2877);
    outputs(3425) <= not(layer2_outputs(427));
    outputs(3426) <= layer2_outputs(5976);
    outputs(3427) <= layer2_outputs(9806);
    outputs(3428) <= layer2_outputs(331);
    outputs(3429) <= not(layer2_outputs(7939));
    outputs(3430) <= not(layer2_outputs(3538));
    outputs(3431) <= not(layer2_outputs(6079));
    outputs(3432) <= not(layer2_outputs(7217));
    outputs(3433) <= layer2_outputs(2868);
    outputs(3434) <= (layer2_outputs(9044)) xor (layer2_outputs(619));
    outputs(3435) <= not(layer2_outputs(574));
    outputs(3436) <= layer2_outputs(658);
    outputs(3437) <= layer2_outputs(9184);
    outputs(3438) <= not(layer2_outputs(9312));
    outputs(3439) <= layer2_outputs(4517);
    outputs(3440) <= not(layer2_outputs(2140));
    outputs(3441) <= layer2_outputs(2221);
    outputs(3442) <= not((layer2_outputs(8021)) xor (layer2_outputs(5800)));
    outputs(3443) <= layer2_outputs(5363);
    outputs(3444) <= layer2_outputs(1289);
    outputs(3445) <= not((layer2_outputs(2778)) xor (layer2_outputs(5731)));
    outputs(3446) <= layer2_outputs(9750);
    outputs(3447) <= not(layer2_outputs(7703));
    outputs(3448) <= not(layer2_outputs(5869));
    outputs(3449) <= layer2_outputs(6658);
    outputs(3450) <= not(layer2_outputs(6645));
    outputs(3451) <= not(layer2_outputs(6572)) or (layer2_outputs(1010));
    outputs(3452) <= not((layer2_outputs(8193)) and (layer2_outputs(5826)));
    outputs(3453) <= (layer2_outputs(2912)) xor (layer2_outputs(1481));
    outputs(3454) <= layer2_outputs(4698);
    outputs(3455) <= not((layer2_outputs(6537)) xor (layer2_outputs(8422)));
    outputs(3456) <= not((layer2_outputs(411)) and (layer2_outputs(1123)));
    outputs(3457) <= not(layer2_outputs(6428));
    outputs(3458) <= layer2_outputs(4797);
    outputs(3459) <= (layer2_outputs(8878)) xor (layer2_outputs(623));
    outputs(3460) <= not(layer2_outputs(2058));
    outputs(3461) <= layer2_outputs(8163);
    outputs(3462) <= not(layer2_outputs(304)) or (layer2_outputs(5662));
    outputs(3463) <= layer2_outputs(2508);
    outputs(3464) <= (layer2_outputs(9466)) xor (layer2_outputs(2046));
    outputs(3465) <= (layer2_outputs(763)) xor (layer2_outputs(2938));
    outputs(3466) <= layer2_outputs(5616);
    outputs(3467) <= (layer2_outputs(7367)) and not (layer2_outputs(4585));
    outputs(3468) <= (layer2_outputs(7361)) and not (layer2_outputs(4786));
    outputs(3469) <= not(layer2_outputs(9941)) or (layer2_outputs(5799));
    outputs(3470) <= not(layer2_outputs(2395));
    outputs(3471) <= not(layer2_outputs(463));
    outputs(3472) <= not((layer2_outputs(8330)) xor (layer2_outputs(907)));
    outputs(3473) <= layer2_outputs(6602);
    outputs(3474) <= layer2_outputs(5657);
    outputs(3475) <= not((layer2_outputs(6209)) xor (layer2_outputs(6746)));
    outputs(3476) <= not(layer2_outputs(4345));
    outputs(3477) <= layer2_outputs(7028);
    outputs(3478) <= layer2_outputs(6700);
    outputs(3479) <= not(layer2_outputs(5291));
    outputs(3480) <= layer2_outputs(7081);
    outputs(3481) <= layer2_outputs(9420);
    outputs(3482) <= layer2_outputs(5248);
    outputs(3483) <= layer2_outputs(1355);
    outputs(3484) <= layer2_outputs(4911);
    outputs(3485) <= (layer2_outputs(7994)) or (layer2_outputs(676));
    outputs(3486) <= layer2_outputs(511);
    outputs(3487) <= not((layer2_outputs(9498)) xor (layer2_outputs(6085)));
    outputs(3488) <= not((layer2_outputs(8407)) xor (layer2_outputs(8933)));
    outputs(3489) <= not(layer2_outputs(6150));
    outputs(3490) <= layer2_outputs(6670);
    outputs(3491) <= not((layer2_outputs(3034)) or (layer2_outputs(2790)));
    outputs(3492) <= not((layer2_outputs(5398)) xor (layer2_outputs(6118)));
    outputs(3493) <= layer2_outputs(9621);
    outputs(3494) <= (layer2_outputs(8421)) and not (layer2_outputs(4247));
    outputs(3495) <= not((layer2_outputs(1787)) and (layer2_outputs(5030)));
    outputs(3496) <= layer2_outputs(5009);
    outputs(3497) <= layer2_outputs(2971);
    outputs(3498) <= not((layer2_outputs(8532)) xor (layer2_outputs(4682)));
    outputs(3499) <= not(layer2_outputs(2527));
    outputs(3500) <= not((layer2_outputs(7908)) or (layer2_outputs(4649)));
    outputs(3501) <= not((layer2_outputs(8180)) xor (layer2_outputs(9689)));
    outputs(3502) <= not((layer2_outputs(9949)) or (layer2_outputs(2578)));
    outputs(3503) <= not((layer2_outputs(2117)) xor (layer2_outputs(7025)));
    outputs(3504) <= not(layer2_outputs(8220));
    outputs(3505) <= layer2_outputs(7027);
    outputs(3506) <= not((layer2_outputs(2525)) xor (layer2_outputs(1695)));
    outputs(3507) <= (layer2_outputs(4006)) and (layer2_outputs(165));
    outputs(3508) <= not(layer2_outputs(8656));
    outputs(3509) <= not(layer2_outputs(5957));
    outputs(3510) <= (layer2_outputs(326)) xor (layer2_outputs(7483));
    outputs(3511) <= not((layer2_outputs(1831)) xor (layer2_outputs(5633)));
    outputs(3512) <= layer2_outputs(4543);
    outputs(3513) <= not((layer2_outputs(10149)) xor (layer2_outputs(6468)));
    outputs(3514) <= layer2_outputs(276);
    outputs(3515) <= (layer2_outputs(1691)) xor (layer2_outputs(8351));
    outputs(3516) <= not(layer2_outputs(2045));
    outputs(3517) <= (layer2_outputs(6499)) xor (layer2_outputs(307));
    outputs(3518) <= not(layer2_outputs(88));
    outputs(3519) <= not((layer2_outputs(987)) xor (layer2_outputs(2751)));
    outputs(3520) <= not(layer2_outputs(6996)) or (layer2_outputs(6123));
    outputs(3521) <= layer2_outputs(5744);
    outputs(3522) <= not((layer2_outputs(8348)) xor (layer2_outputs(9950)));
    outputs(3523) <= layer2_outputs(8038);
    outputs(3524) <= layer2_outputs(5475);
    outputs(3525) <= (layer2_outputs(3578)) xor (layer2_outputs(939));
    outputs(3526) <= layer2_outputs(2719);
    outputs(3527) <= (layer2_outputs(6703)) and not (layer2_outputs(2981));
    outputs(3528) <= not(layer2_outputs(8070));
    outputs(3529) <= not(layer2_outputs(875));
    outputs(3530) <= layer2_outputs(9306);
    outputs(3531) <= not(layer2_outputs(7327));
    outputs(3532) <= layer2_outputs(152);
    outputs(3533) <= layer2_outputs(3511);
    outputs(3534) <= not(layer2_outputs(2948));
    outputs(3535) <= layer2_outputs(8822);
    outputs(3536) <= not(layer2_outputs(4335));
    outputs(3537) <= not(layer2_outputs(5829));
    outputs(3538) <= not((layer2_outputs(10140)) xor (layer2_outputs(1687)));
    outputs(3539) <= (layer2_outputs(8804)) xor (layer2_outputs(5097));
    outputs(3540) <= not(layer2_outputs(2700));
    outputs(3541) <= not(layer2_outputs(5273));
    outputs(3542) <= layer2_outputs(730);
    outputs(3543) <= layer2_outputs(7069);
    outputs(3544) <= not(layer2_outputs(9620));
    outputs(3545) <= (layer2_outputs(9793)) xor (layer2_outputs(5064));
    outputs(3546) <= (layer2_outputs(6844)) xor (layer2_outputs(9536));
    outputs(3547) <= not(layer2_outputs(985));
    outputs(3548) <= (layer2_outputs(7345)) xor (layer2_outputs(9359));
    outputs(3549) <= not(layer2_outputs(3971));
    outputs(3550) <= layer2_outputs(7319);
    outputs(3551) <= layer2_outputs(1065);
    outputs(3552) <= not((layer2_outputs(5001)) or (layer2_outputs(10040)));
    outputs(3553) <= not(layer2_outputs(4815));
    outputs(3554) <= layer2_outputs(4495);
    outputs(3555) <= not((layer2_outputs(6374)) xor (layer2_outputs(5767)));
    outputs(3556) <= not((layer2_outputs(7458)) xor (layer2_outputs(5795)));
    outputs(3557) <= layer2_outputs(5645);
    outputs(3558) <= not(layer2_outputs(7723));
    outputs(3559) <= layer2_outputs(4606);
    outputs(3560) <= not(layer2_outputs(8158));
    outputs(3561) <= not(layer2_outputs(497));
    outputs(3562) <= not(layer2_outputs(8142));
    outputs(3563) <= (layer2_outputs(8597)) and not (layer2_outputs(9344));
    outputs(3564) <= not(layer2_outputs(5751));
    outputs(3565) <= not(layer2_outputs(7195)) or (layer2_outputs(4589));
    outputs(3566) <= layer2_outputs(8953);
    outputs(3567) <= layer2_outputs(6811);
    outputs(3568) <= not((layer2_outputs(3935)) xor (layer2_outputs(8603)));
    outputs(3569) <= (layer2_outputs(4746)) xor (layer2_outputs(1536));
    outputs(3570) <= layer2_outputs(10092);
    outputs(3571) <= not(layer2_outputs(1311));
    outputs(3572) <= layer2_outputs(7435);
    outputs(3573) <= (layer2_outputs(2195)) and not (layer2_outputs(6796));
    outputs(3574) <= not(layer2_outputs(1777));
    outputs(3575) <= not(layer2_outputs(10160));
    outputs(3576) <= layer2_outputs(7056);
    outputs(3577) <= not((layer2_outputs(3140)) xor (layer2_outputs(9257)));
    outputs(3578) <= not(layer2_outputs(9974)) or (layer2_outputs(10070));
    outputs(3579) <= layer2_outputs(2032);
    outputs(3580) <= not((layer2_outputs(9024)) xor (layer2_outputs(1640)));
    outputs(3581) <= layer2_outputs(7797);
    outputs(3582) <= layer2_outputs(825);
    outputs(3583) <= (layer2_outputs(7336)) xor (layer2_outputs(5736));
    outputs(3584) <= not(layer2_outputs(8837));
    outputs(3585) <= not(layer2_outputs(738));
    outputs(3586) <= not(layer2_outputs(6137));
    outputs(3587) <= not(layer2_outputs(10178));
    outputs(3588) <= layer2_outputs(4981);
    outputs(3589) <= not((layer2_outputs(9725)) xor (layer2_outputs(3226)));
    outputs(3590) <= not(layer2_outputs(8274));
    outputs(3591) <= layer2_outputs(4493);
    outputs(3592) <= layer2_outputs(6593);
    outputs(3593) <= not((layer2_outputs(5296)) xor (layer2_outputs(6449)));
    outputs(3594) <= layer2_outputs(7440);
    outputs(3595) <= not(layer2_outputs(9400));
    outputs(3596) <= (layer2_outputs(7995)) and not (layer2_outputs(7000));
    outputs(3597) <= (layer2_outputs(8718)) or (layer2_outputs(6123));
    outputs(3598) <= not(layer2_outputs(9609));
    outputs(3599) <= layer2_outputs(9032);
    outputs(3600) <= (layer2_outputs(8697)) or (layer2_outputs(2088));
    outputs(3601) <= not(layer2_outputs(5356));
    outputs(3602) <= not((layer2_outputs(9651)) or (layer2_outputs(9626)));
    outputs(3603) <= not(layer2_outputs(4707));
    outputs(3604) <= not(layer2_outputs(352));
    outputs(3605) <= layer2_outputs(219);
    outputs(3606) <= (layer2_outputs(117)) and not (layer2_outputs(10225));
    outputs(3607) <= not(layer2_outputs(5786));
    outputs(3608) <= not(layer2_outputs(1670));
    outputs(3609) <= not(layer2_outputs(8583));
    outputs(3610) <= not(layer2_outputs(1586));
    outputs(3611) <= not((layer2_outputs(1344)) xor (layer2_outputs(2989)));
    outputs(3612) <= layer2_outputs(9995);
    outputs(3613) <= (layer2_outputs(8128)) xor (layer2_outputs(3831));
    outputs(3614) <= not(layer2_outputs(4146));
    outputs(3615) <= not((layer2_outputs(7455)) xor (layer2_outputs(293)));
    outputs(3616) <= not(layer2_outputs(6991));
    outputs(3617) <= layer2_outputs(769);
    outputs(3618) <= not(layer2_outputs(2512));
    outputs(3619) <= layer2_outputs(4965);
    outputs(3620) <= not(layer2_outputs(7182));
    outputs(3621) <= not(layer2_outputs(10033));
    outputs(3622) <= layer2_outputs(2920);
    outputs(3623) <= not((layer2_outputs(4046)) xor (layer2_outputs(6741)));
    outputs(3624) <= (layer2_outputs(212)) and not (layer2_outputs(10152));
    outputs(3625) <= (layer2_outputs(3064)) xor (layer2_outputs(1798));
    outputs(3626) <= layer2_outputs(6958);
    outputs(3627) <= not((layer2_outputs(8100)) xor (layer2_outputs(6404)));
    outputs(3628) <= layer2_outputs(1636);
    outputs(3629) <= not(layer2_outputs(2334));
    outputs(3630) <= not(layer2_outputs(2893)) or (layer2_outputs(3420));
    outputs(3631) <= layer2_outputs(1);
    outputs(3632) <= not(layer2_outputs(1322));
    outputs(3633) <= not(layer2_outputs(3902));
    outputs(3634) <= layer2_outputs(1751);
    outputs(3635) <= (layer2_outputs(1629)) xor (layer2_outputs(4687));
    outputs(3636) <= not(layer2_outputs(1943));
    outputs(3637) <= (layer2_outputs(6413)) and (layer2_outputs(5297));
    outputs(3638) <= (layer2_outputs(8284)) xor (layer2_outputs(5261));
    outputs(3639) <= not((layer2_outputs(5726)) xor (layer2_outputs(3348)));
    outputs(3640) <= layer2_outputs(3061);
    outputs(3641) <= layer2_outputs(1770);
    outputs(3642) <= not(layer2_outputs(2018));
    outputs(3643) <= layer2_outputs(1668);
    outputs(3644) <= not(layer2_outputs(9338));
    outputs(3645) <= (layer2_outputs(4359)) xor (layer2_outputs(5128));
    outputs(3646) <= not(layer2_outputs(8159));
    outputs(3647) <= not(layer2_outputs(1135));
    outputs(3648) <= not((layer2_outputs(6163)) xor (layer2_outputs(7870)));
    outputs(3649) <= layer2_outputs(6125);
    outputs(3650) <= layer2_outputs(2434);
    outputs(3651) <= not(layer2_outputs(920));
    outputs(3652) <= not(layer2_outputs(9794));
    outputs(3653) <= not(layer2_outputs(3574));
    outputs(3654) <= not(layer2_outputs(7568));
    outputs(3655) <= (layer2_outputs(348)) xor (layer2_outputs(8301));
    outputs(3656) <= layer2_outputs(9444);
    outputs(3657) <= layer2_outputs(794);
    outputs(3658) <= not(layer2_outputs(6064));
    outputs(3659) <= not((layer2_outputs(4116)) xor (layer2_outputs(5263)));
    outputs(3660) <= not(layer2_outputs(4451));
    outputs(3661) <= layer2_outputs(8279);
    outputs(3662) <= layer2_outputs(7014);
    outputs(3663) <= not(layer2_outputs(8985));
    outputs(3664) <= layer2_outputs(444);
    outputs(3665) <= layer2_outputs(3422);
    outputs(3666) <= (layer2_outputs(6193)) and not (layer2_outputs(7120));
    outputs(3667) <= layer2_outputs(6744);
    outputs(3668) <= layer2_outputs(1536);
    outputs(3669) <= not((layer2_outputs(2484)) xor (layer2_outputs(6119)));
    outputs(3670) <= not(layer2_outputs(750));
    outputs(3671) <= not(layer2_outputs(4586));
    outputs(3672) <= layer2_outputs(1380);
    outputs(3673) <= layer2_outputs(3964);
    outputs(3674) <= layer2_outputs(1705);
    outputs(3675) <= not((layer2_outputs(4808)) xor (layer2_outputs(8122)));
    outputs(3676) <= layer2_outputs(4106);
    outputs(3677) <= layer2_outputs(10100);
    outputs(3678) <= layer2_outputs(7373);
    outputs(3679) <= not(layer2_outputs(8499));
    outputs(3680) <= layer2_outputs(6473);
    outputs(3681) <= not(layer2_outputs(1088));
    outputs(3682) <= not((layer2_outputs(4636)) xor (layer2_outputs(9083)));
    outputs(3683) <= not(layer2_outputs(818));
    outputs(3684) <= not(layer2_outputs(569));
    outputs(3685) <= (layer2_outputs(9318)) or (layer2_outputs(1847));
    outputs(3686) <= not(layer2_outputs(1043));
    outputs(3687) <= not(layer2_outputs(10051));
    outputs(3688) <= not(layer2_outputs(5646));
    outputs(3689) <= layer2_outputs(255);
    outputs(3690) <= layer2_outputs(439);
    outputs(3691) <= (layer2_outputs(979)) and not (layer2_outputs(1762));
    outputs(3692) <= not(layer2_outputs(7733)) or (layer2_outputs(6219));
    outputs(3693) <= not(layer2_outputs(4977));
    outputs(3694) <= layer2_outputs(1482);
    outputs(3695) <= not(layer2_outputs(8083));
    outputs(3696) <= layer2_outputs(5616);
    outputs(3697) <= layer2_outputs(4223);
    outputs(3698) <= not(layer2_outputs(667)) or (layer2_outputs(9789));
    outputs(3699) <= not(layer2_outputs(7579));
    outputs(3700) <= layer2_outputs(3341);
    outputs(3701) <= not(layer2_outputs(6507));
    outputs(3702) <= layer2_outputs(6818);
    outputs(3703) <= not(layer2_outputs(7706));
    outputs(3704) <= not(layer2_outputs(8831));
    outputs(3705) <= (layer2_outputs(2152)) xor (layer2_outputs(456));
    outputs(3706) <= (layer2_outputs(8667)) xor (layer2_outputs(8791));
    outputs(3707) <= (layer2_outputs(9373)) xor (layer2_outputs(9569));
    outputs(3708) <= layer2_outputs(8235);
    outputs(3709) <= not(layer2_outputs(5574));
    outputs(3710) <= not(layer2_outputs(3604));
    outputs(3711) <= (layer2_outputs(3479)) xor (layer2_outputs(10084));
    outputs(3712) <= (layer2_outputs(4503)) and not (layer2_outputs(3084));
    outputs(3713) <= (layer2_outputs(1986)) and not (layer2_outputs(2746));
    outputs(3714) <= (layer2_outputs(9502)) xor (layer2_outputs(6013));
    outputs(3715) <= layer2_outputs(4699);
    outputs(3716) <= layer2_outputs(9871);
    outputs(3717) <= not(layer2_outputs(8998)) or (layer2_outputs(4833));
    outputs(3718) <= not(layer2_outputs(4720));
    outputs(3719) <= not(layer2_outputs(3805));
    outputs(3720) <= layer2_outputs(7785);
    outputs(3721) <= not((layer2_outputs(8371)) xor (layer2_outputs(2605)));
    outputs(3722) <= (layer2_outputs(1447)) xor (layer2_outputs(9699));
    outputs(3723) <= not((layer2_outputs(4422)) xor (layer2_outputs(377)));
    outputs(3724) <= layer2_outputs(6473);
    outputs(3725) <= not((layer2_outputs(7385)) xor (layer2_outputs(9852)));
    outputs(3726) <= layer2_outputs(6576);
    outputs(3727) <= not(layer2_outputs(2739)) or (layer2_outputs(2788));
    outputs(3728) <= layer2_outputs(5931);
    outputs(3729) <= not(layer2_outputs(7125));
    outputs(3730) <= not((layer2_outputs(515)) or (layer2_outputs(4844)));
    outputs(3731) <= not((layer2_outputs(4515)) xor (layer2_outputs(732)));
    outputs(3732) <= not((layer2_outputs(4870)) xor (layer2_outputs(6955)));
    outputs(3733) <= not(layer2_outputs(8891));
    outputs(3734) <= not(layer2_outputs(2562));
    outputs(3735) <= layer2_outputs(10208);
    outputs(3736) <= not(layer2_outputs(7126));
    outputs(3737) <= layer2_outputs(3542);
    outputs(3738) <= layer2_outputs(9380);
    outputs(3739) <= layer2_outputs(3416);
    outputs(3740) <= not((layer2_outputs(9849)) xor (layer2_outputs(8123)));
    outputs(3741) <= (layer2_outputs(6106)) and not (layer2_outputs(146));
    outputs(3742) <= not(layer2_outputs(90));
    outputs(3743) <= layer2_outputs(6725);
    outputs(3744) <= layer2_outputs(7394);
    outputs(3745) <= not(layer2_outputs(3815));
    outputs(3746) <= layer2_outputs(43);
    outputs(3747) <= layer2_outputs(2943);
    outputs(3748) <= layer2_outputs(10082);
    outputs(3749) <= not(layer2_outputs(3644));
    outputs(3750) <= not(layer2_outputs(8472));
    outputs(3751) <= layer2_outputs(2312);
    outputs(3752) <= (layer2_outputs(2925)) and (layer2_outputs(8266));
    outputs(3753) <= layer2_outputs(225);
    outputs(3754) <= not(layer2_outputs(4455)) or (layer2_outputs(987));
    outputs(3755) <= layer2_outputs(8856);
    outputs(3756) <= layer2_outputs(248);
    outputs(3757) <= layer2_outputs(5383);
    outputs(3758) <= not(layer2_outputs(9616));
    outputs(3759) <= layer2_outputs(1074);
    outputs(3760) <= not((layer2_outputs(8565)) or (layer2_outputs(5870)));
    outputs(3761) <= not(layer2_outputs(6861));
    outputs(3762) <= layer2_outputs(8625);
    outputs(3763) <= (layer2_outputs(1131)) and not (layer2_outputs(2974));
    outputs(3764) <= not(layer2_outputs(7523));
    outputs(3765) <= not(layer2_outputs(7938));
    outputs(3766) <= not((layer2_outputs(1273)) and (layer2_outputs(8056)));
    outputs(3767) <= (layer2_outputs(5650)) xor (layer2_outputs(3836));
    outputs(3768) <= layer2_outputs(2798);
    outputs(3769) <= not((layer2_outputs(9765)) and (layer2_outputs(3796)));
    outputs(3770) <= not(layer2_outputs(9114));
    outputs(3771) <= not(layer2_outputs(4967));
    outputs(3772) <= not(layer2_outputs(2841));
    outputs(3773) <= (layer2_outputs(2000)) xor (layer2_outputs(6579));
    outputs(3774) <= not((layer2_outputs(4712)) xor (layer2_outputs(9323)));
    outputs(3775) <= layer2_outputs(464);
    outputs(3776) <= not((layer2_outputs(9396)) xor (layer2_outputs(3532)));
    outputs(3777) <= (layer2_outputs(5250)) and (layer2_outputs(8573));
    outputs(3778) <= layer2_outputs(1363);
    outputs(3779) <= not((layer2_outputs(2924)) xor (layer2_outputs(7831)));
    outputs(3780) <= not((layer2_outputs(5644)) or (layer2_outputs(6318)));
    outputs(3781) <= not(layer2_outputs(2517));
    outputs(3782) <= not(layer2_outputs(5019));
    outputs(3783) <= (layer2_outputs(6338)) xor (layer2_outputs(7560));
    outputs(3784) <= (layer2_outputs(6160)) xor (layer2_outputs(4874));
    outputs(3785) <= (layer2_outputs(3311)) xor (layer2_outputs(8890));
    outputs(3786) <= (layer2_outputs(5939)) and not (layer2_outputs(5604));
    outputs(3787) <= not(layer2_outputs(8409));
    outputs(3788) <= not(layer2_outputs(8699));
    outputs(3789) <= layer2_outputs(2889);
    outputs(3790) <= not(layer2_outputs(2168));
    outputs(3791) <= layer2_outputs(8650);
    outputs(3792) <= not(layer2_outputs(10199)) or (layer2_outputs(7350));
    outputs(3793) <= (layer2_outputs(9476)) xor (layer2_outputs(8854));
    outputs(3794) <= layer2_outputs(9039);
    outputs(3795) <= (layer2_outputs(7606)) or (layer2_outputs(8575));
    outputs(3796) <= layer2_outputs(9353);
    outputs(3797) <= not(layer2_outputs(4094));
    outputs(3798) <= not(layer2_outputs(1737));
    outputs(3799) <= not(layer2_outputs(4184));
    outputs(3800) <= (layer2_outputs(9467)) and not (layer2_outputs(3447));
    outputs(3801) <= (layer2_outputs(6825)) and not (layer2_outputs(1684));
    outputs(3802) <= (layer2_outputs(1668)) or (layer2_outputs(2990));
    outputs(3803) <= not(layer2_outputs(1460)) or (layer2_outputs(4753));
    outputs(3804) <= not(layer2_outputs(2872));
    outputs(3805) <= layer2_outputs(2884);
    outputs(3806) <= (layer2_outputs(4271)) and not (layer2_outputs(5979));
    outputs(3807) <= not((layer2_outputs(4146)) xor (layer2_outputs(3490)));
    outputs(3808) <= not(layer2_outputs(1020));
    outputs(3809) <= layer2_outputs(9041);
    outputs(3810) <= (layer2_outputs(5873)) xor (layer2_outputs(690));
    outputs(3811) <= (layer2_outputs(9346)) xor (layer2_outputs(8898));
    outputs(3812) <= not(layer2_outputs(1311));
    outputs(3813) <= layer2_outputs(8988);
    outputs(3814) <= layer2_outputs(3405);
    outputs(3815) <= layer2_outputs(9233);
    outputs(3816) <= not(layer2_outputs(4467));
    outputs(3817) <= not((layer2_outputs(4177)) xor (layer2_outputs(9350)));
    outputs(3818) <= layer2_outputs(54);
    outputs(3819) <= not((layer2_outputs(2400)) xor (layer2_outputs(7764)));
    outputs(3820) <= not(layer2_outputs(9163));
    outputs(3821) <= layer2_outputs(2262);
    outputs(3822) <= layer2_outputs(4576);
    outputs(3823) <= not(layer2_outputs(696));
    outputs(3824) <= not(layer2_outputs(3163));
    outputs(3825) <= layer2_outputs(10048);
    outputs(3826) <= layer2_outputs(4933);
    outputs(3827) <= not(layer2_outputs(9455));
    outputs(3828) <= not(layer2_outputs(4452)) or (layer2_outputs(6696));
    outputs(3829) <= not((layer2_outputs(4122)) xor (layer2_outputs(3892)));
    outputs(3830) <= layer2_outputs(715);
    outputs(3831) <= not((layer2_outputs(8394)) and (layer2_outputs(9897)));
    outputs(3832) <= not(layer2_outputs(9302));
    outputs(3833) <= (layer2_outputs(2597)) and (layer2_outputs(9377));
    outputs(3834) <= not(layer2_outputs(7498));
    outputs(3835) <= layer2_outputs(3557);
    outputs(3836) <= layer2_outputs(5698);
    outputs(3837) <= not(layer2_outputs(5062));
    outputs(3838) <= layer2_outputs(7857);
    outputs(3839) <= not(layer2_outputs(790)) or (layer2_outputs(6494));
    outputs(3840) <= layer2_outputs(3089);
    outputs(3841) <= (layer2_outputs(9893)) xor (layer2_outputs(4604));
    outputs(3842) <= not(layer2_outputs(5921));
    outputs(3843) <= not(layer2_outputs(1697));
    outputs(3844) <= not(layer2_outputs(3646));
    outputs(3845) <= layer2_outputs(3799);
    outputs(3846) <= (layer2_outputs(8195)) and not (layer2_outputs(1090));
    outputs(3847) <= (layer2_outputs(9656)) and not (layer2_outputs(1239));
    outputs(3848) <= not((layer2_outputs(1917)) xor (layer2_outputs(3314)));
    outputs(3849) <= (layer2_outputs(2225)) and (layer2_outputs(5401));
    outputs(3850) <= not(layer2_outputs(5572));
    outputs(3851) <= not(layer2_outputs(6654));
    outputs(3852) <= (layer2_outputs(3891)) and (layer2_outputs(4946));
    outputs(3853) <= layer2_outputs(2875);
    outputs(3854) <= not(layer2_outputs(4997));
    outputs(3855) <= layer2_outputs(3280);
    outputs(3856) <= not(layer2_outputs(9105));
    outputs(3857) <= not(layer2_outputs(3174));
    outputs(3858) <= not((layer2_outputs(9361)) xor (layer2_outputs(5892)));
    outputs(3859) <= layer2_outputs(6627);
    outputs(3860) <= layer2_outputs(9554);
    outputs(3861) <= layer2_outputs(1065);
    outputs(3862) <= not(layer2_outputs(7921));
    outputs(3863) <= layer2_outputs(3540);
    outputs(3864) <= not(layer2_outputs(3125));
    outputs(3865) <= not(layer2_outputs(6996));
    outputs(3866) <= layer2_outputs(9039);
    outputs(3867) <= layer2_outputs(8556);
    outputs(3868) <= (layer2_outputs(7281)) and (layer2_outputs(9858));
    outputs(3869) <= (layer2_outputs(2244)) and (layer2_outputs(3852));
    outputs(3870) <= (layer2_outputs(6937)) and (layer2_outputs(1877));
    outputs(3871) <= not((layer2_outputs(324)) xor (layer2_outputs(5884)));
    outputs(3872) <= layer2_outputs(7696);
    outputs(3873) <= (layer2_outputs(7466)) and not (layer2_outputs(7380));
    outputs(3874) <= layer2_outputs(7163);
    outputs(3875) <= not(layer2_outputs(1103));
    outputs(3876) <= not(layer2_outputs(3906));
    outputs(3877) <= layer2_outputs(4570);
    outputs(3878) <= not(layer2_outputs(9818));
    outputs(3879) <= layer2_outputs(2789);
    outputs(3880) <= not(layer2_outputs(3369));
    outputs(3881) <= (layer2_outputs(2976)) or (layer2_outputs(9162));
    outputs(3882) <= not((layer2_outputs(8175)) or (layer2_outputs(8484)));
    outputs(3883) <= layer2_outputs(152);
    outputs(3884) <= not(layer2_outputs(9163));
    outputs(3885) <= layer2_outputs(5006);
    outputs(3886) <= not(layer2_outputs(5694)) or (layer2_outputs(9945));
    outputs(3887) <= layer2_outputs(7532);
    outputs(3888) <= layer2_outputs(5248);
    outputs(3889) <= layer2_outputs(2215);
    outputs(3890) <= (layer2_outputs(3159)) xor (layer2_outputs(3314));
    outputs(3891) <= not((layer2_outputs(1188)) xor (layer2_outputs(175)));
    outputs(3892) <= layer2_outputs(423);
    outputs(3893) <= layer2_outputs(584);
    outputs(3894) <= not((layer2_outputs(3133)) xor (layer2_outputs(6248)));
    outputs(3895) <= (layer2_outputs(1200)) and not (layer2_outputs(5938));
    outputs(3896) <= layer2_outputs(1577);
    outputs(3897) <= layer2_outputs(5901);
    outputs(3898) <= not((layer2_outputs(1366)) xor (layer2_outputs(9394)));
    outputs(3899) <= not(layer2_outputs(5358));
    outputs(3900) <= not(layer2_outputs(3527));
    outputs(3901) <= layer2_outputs(2137);
    outputs(3902) <= not(layer2_outputs(3704));
    outputs(3903) <= layer2_outputs(9092);
    outputs(3904) <= (layer2_outputs(6741)) xor (layer2_outputs(3749));
    outputs(3905) <= (layer2_outputs(7287)) xor (layer2_outputs(836));
    outputs(3906) <= not(layer2_outputs(4468));
    outputs(3907) <= (layer2_outputs(7243)) and not (layer2_outputs(2067));
    outputs(3908) <= layer2_outputs(9485);
    outputs(3909) <= (layer2_outputs(9747)) and not (layer2_outputs(6470));
    outputs(3910) <= not(layer2_outputs(9667));
    outputs(3911) <= (layer2_outputs(4083)) xor (layer2_outputs(3058));
    outputs(3912) <= not((layer2_outputs(7924)) xor (layer2_outputs(7927)));
    outputs(3913) <= not((layer2_outputs(9654)) xor (layer2_outputs(5437)));
    outputs(3914) <= layer2_outputs(3429);
    outputs(3915) <= not(layer2_outputs(4140)) or (layer2_outputs(605));
    outputs(3916) <= not((layer2_outputs(7740)) xor (layer2_outputs(2651)));
    outputs(3917) <= layer2_outputs(4712);
    outputs(3918) <= layer2_outputs(6666);
    outputs(3919) <= layer2_outputs(5318);
    outputs(3920) <= '0';
    outputs(3921) <= (layer2_outputs(8395)) xor (layer2_outputs(9948));
    outputs(3922) <= not((layer2_outputs(5085)) xor (layer2_outputs(2410)));
    outputs(3923) <= layer2_outputs(1285);
    outputs(3924) <= layer2_outputs(9465);
    outputs(3925) <= layer2_outputs(6914);
    outputs(3926) <= (layer2_outputs(531)) xor (layer2_outputs(868));
    outputs(3927) <= (layer2_outputs(1232)) xor (layer2_outputs(7735));
    outputs(3928) <= layer2_outputs(4218);
    outputs(3929) <= not(layer2_outputs(6293));
    outputs(3930) <= layer2_outputs(3382);
    outputs(3931) <= (layer2_outputs(8398)) and not (layer2_outputs(5814));
    outputs(3932) <= not(layer2_outputs(6779));
    outputs(3933) <= not((layer2_outputs(1737)) and (layer2_outputs(3387)));
    outputs(3934) <= not(layer2_outputs(8453));
    outputs(3935) <= not(layer2_outputs(8782));
    outputs(3936) <= not(layer2_outputs(1106)) or (layer2_outputs(5746));
    outputs(3937) <= not(layer2_outputs(2056));
    outputs(3938) <= not(layer2_outputs(283));
    outputs(3939) <= not((layer2_outputs(6548)) xor (layer2_outputs(2695)));
    outputs(3940) <= layer2_outputs(7564);
    outputs(3941) <= not(layer2_outputs(9084));
    outputs(3942) <= layer2_outputs(8002);
    outputs(3943) <= (layer2_outputs(5138)) or (layer2_outputs(2614));
    outputs(3944) <= not(layer2_outputs(9178));
    outputs(3945) <= not(layer2_outputs(3734));
    outputs(3946) <= not((layer2_outputs(3455)) xor (layer2_outputs(3451)));
    outputs(3947) <= layer2_outputs(4240);
    outputs(3948) <= layer2_outputs(4994);
    outputs(3949) <= layer2_outputs(420);
    outputs(3950) <= not(layer2_outputs(4512));
    outputs(3951) <= (layer2_outputs(2886)) and (layer2_outputs(6615));
    outputs(3952) <= not(layer2_outputs(1424));
    outputs(3953) <= (layer2_outputs(3881)) and not (layer2_outputs(9988));
    outputs(3954) <= (layer2_outputs(3806)) and (layer2_outputs(2711));
    outputs(3955) <= layer2_outputs(975);
    outputs(3956) <= not(layer2_outputs(8447));
    outputs(3957) <= not(layer2_outputs(6321));
    outputs(3958) <= layer2_outputs(631);
    outputs(3959) <= not(layer2_outputs(1036));
    outputs(3960) <= not(layer2_outputs(2724)) or (layer2_outputs(4272));
    outputs(3961) <= layer2_outputs(8379);
    outputs(3962) <= layer2_outputs(1211);
    outputs(3963) <= layer2_outputs(7436);
    outputs(3964) <= not((layer2_outputs(5915)) or (layer2_outputs(2291)));
    outputs(3965) <= not(layer2_outputs(966));
    outputs(3966) <= not((layer2_outputs(2842)) xor (layer2_outputs(4081)));
    outputs(3967) <= layer2_outputs(1132);
    outputs(3968) <= layer2_outputs(5174);
    outputs(3969) <= (layer2_outputs(4834)) xor (layer2_outputs(2010));
    outputs(3970) <= (layer2_outputs(1926)) xor (layer2_outputs(8921));
    outputs(3971) <= layer2_outputs(5364);
    outputs(3972) <= layer2_outputs(7582);
    outputs(3973) <= not(layer2_outputs(2035));
    outputs(3974) <= (layer2_outputs(4540)) xor (layer2_outputs(9432));
    outputs(3975) <= layer2_outputs(8852);
    outputs(3976) <= not((layer2_outputs(7074)) xor (layer2_outputs(3654)));
    outputs(3977) <= not(layer2_outputs(1967));
    outputs(3978) <= not((layer2_outputs(2461)) or (layer2_outputs(9534)));
    outputs(3979) <= (layer2_outputs(591)) or (layer2_outputs(1598));
    outputs(3980) <= not(layer2_outputs(8042)) or (layer2_outputs(7117));
    outputs(3981) <= layer2_outputs(537);
    outputs(3982) <= not(layer2_outputs(7366));
    outputs(3983) <= layer2_outputs(2826);
    outputs(3984) <= not(layer2_outputs(4074));
    outputs(3985) <= not((layer2_outputs(490)) xor (layer2_outputs(2605)));
    outputs(3986) <= not(layer2_outputs(4400)) or (layer2_outputs(7969));
    outputs(3987) <= not((layer2_outputs(2546)) and (layer2_outputs(12)));
    outputs(3988) <= layer2_outputs(7509);
    outputs(3989) <= not((layer2_outputs(2452)) and (layer2_outputs(5985)));
    outputs(3990) <= not(layer2_outputs(5392));
    outputs(3991) <= not(layer2_outputs(10067));
    outputs(3992) <= not((layer2_outputs(7984)) or (layer2_outputs(8961)));
    outputs(3993) <= (layer2_outputs(7358)) xor (layer2_outputs(8125));
    outputs(3994) <= not(layer2_outputs(1222));
    outputs(3995) <= layer2_outputs(7049);
    outputs(3996) <= not((layer2_outputs(2253)) or (layer2_outputs(7845)));
    outputs(3997) <= not((layer2_outputs(2759)) xor (layer2_outputs(7364)));
    outputs(3998) <= layer2_outputs(9679);
    outputs(3999) <= not(layer2_outputs(7651));
    outputs(4000) <= layer2_outputs(6822);
    outputs(4001) <= layer2_outputs(2810);
    outputs(4002) <= not(layer2_outputs(8605));
    outputs(4003) <= not(layer2_outputs(1328));
    outputs(4004) <= (layer2_outputs(10231)) and (layer2_outputs(9152));
    outputs(4005) <= not((layer2_outputs(4450)) xor (layer2_outputs(7711)));
    outputs(4006) <= (layer2_outputs(10203)) xor (layer2_outputs(554));
    outputs(4007) <= layer2_outputs(25);
    outputs(4008) <= not(layer2_outputs(2073));
    outputs(4009) <= not((layer2_outputs(2757)) or (layer2_outputs(6642)));
    outputs(4010) <= not((layer2_outputs(4565)) xor (layer2_outputs(712)));
    outputs(4011) <= layer2_outputs(3099);
    outputs(4012) <= not(layer2_outputs(7628));
    outputs(4013) <= layer2_outputs(4130);
    outputs(4014) <= not(layer2_outputs(6926));
    outputs(4015) <= layer2_outputs(1029);
    outputs(4016) <= not(layer2_outputs(3676));
    outputs(4017) <= layer2_outputs(5603);
    outputs(4018) <= not(layer2_outputs(385)) or (layer2_outputs(7429));
    outputs(4019) <= (layer2_outputs(6924)) and not (layer2_outputs(606));
    outputs(4020) <= (layer2_outputs(898)) or (layer2_outputs(7115));
    outputs(4021) <= not((layer2_outputs(4677)) or (layer2_outputs(2603)));
    outputs(4022) <= (layer2_outputs(5800)) xor (layer2_outputs(5903));
    outputs(4023) <= not(layer2_outputs(4009));
    outputs(4024) <= not(layer2_outputs(1154));
    outputs(4025) <= layer2_outputs(8234);
    outputs(4026) <= (layer2_outputs(7121)) xor (layer2_outputs(3575));
    outputs(4027) <= layer2_outputs(2276);
    outputs(4028) <= layer2_outputs(263);
    outputs(4029) <= (layer2_outputs(9552)) and (layer2_outputs(1050));
    outputs(4030) <= (layer2_outputs(6600)) xor (layer2_outputs(2256));
    outputs(4031) <= not(layer2_outputs(6566));
    outputs(4032) <= (layer2_outputs(7538)) and not (layer2_outputs(8099));
    outputs(4033) <= (layer2_outputs(8213)) xor (layer2_outputs(2838));
    outputs(4034) <= not(layer2_outputs(90));
    outputs(4035) <= not(layer2_outputs(95));
    outputs(4036) <= not(layer2_outputs(5863));
    outputs(4037) <= layer2_outputs(651);
    outputs(4038) <= layer2_outputs(1813);
    outputs(4039) <= not((layer2_outputs(4959)) xor (layer2_outputs(5970)));
    outputs(4040) <= not((layer2_outputs(7213)) xor (layer2_outputs(6536)));
    outputs(4041) <= not(layer2_outputs(1322));
    outputs(4042) <= layer2_outputs(248);
    outputs(4043) <= (layer2_outputs(4957)) xor (layer2_outputs(1221));
    outputs(4044) <= (layer2_outputs(4089)) or (layer2_outputs(2333));
    outputs(4045) <= not(layer2_outputs(6380));
    outputs(4046) <= not(layer2_outputs(8316));
    outputs(4047) <= layer2_outputs(4381);
    outputs(4048) <= layer2_outputs(8884);
    outputs(4049) <= not(layer2_outputs(9615));
    outputs(4050) <= not(layer2_outputs(2664)) or (layer2_outputs(5399));
    outputs(4051) <= not(layer2_outputs(1220));
    outputs(4052) <= layer2_outputs(1422);
    outputs(4053) <= not(layer2_outputs(166));
    outputs(4054) <= layer2_outputs(5087);
    outputs(4055) <= not((layer2_outputs(7170)) xor (layer2_outputs(4820)));
    outputs(4056) <= not(layer2_outputs(4386));
    outputs(4057) <= (layer2_outputs(2772)) and not (layer2_outputs(10237));
    outputs(4058) <= (layer2_outputs(7241)) xor (layer2_outputs(5958));
    outputs(4059) <= layer2_outputs(9137);
    outputs(4060) <= (layer2_outputs(5656)) and (layer2_outputs(6512));
    outputs(4061) <= not((layer2_outputs(2318)) xor (layer2_outputs(10137)));
    outputs(4062) <= not(layer2_outputs(6412));
    outputs(4063) <= (layer2_outputs(1057)) and not (layer2_outputs(1639));
    outputs(4064) <= layer2_outputs(9291);
    outputs(4065) <= layer2_outputs(6565);
    outputs(4066) <= layer2_outputs(2625);
    outputs(4067) <= not(layer2_outputs(3758));
    outputs(4068) <= (layer2_outputs(4248)) and (layer2_outputs(7009));
    outputs(4069) <= (layer2_outputs(9649)) xor (layer2_outputs(2520));
    outputs(4070) <= not(layer2_outputs(7886));
    outputs(4071) <= layer2_outputs(886);
    outputs(4072) <= layer2_outputs(2994);
    outputs(4073) <= (layer2_outputs(3378)) and not (layer2_outputs(8145));
    outputs(4074) <= (layer2_outputs(1673)) xor (layer2_outputs(2876));
    outputs(4075) <= (layer2_outputs(7155)) and not (layer2_outputs(8308));
    outputs(4076) <= not((layer2_outputs(3700)) xor (layer2_outputs(8567)));
    outputs(4077) <= (layer2_outputs(9147)) and (layer2_outputs(9406));
    outputs(4078) <= not((layer2_outputs(5393)) xor (layer2_outputs(10168)));
    outputs(4079) <= not(layer2_outputs(51));
    outputs(4080) <= not(layer2_outputs(1308));
    outputs(4081) <= not(layer2_outputs(6220));
    outputs(4082) <= (layer2_outputs(5170)) xor (layer2_outputs(1619));
    outputs(4083) <= layer2_outputs(4312);
    outputs(4084) <= (layer2_outputs(920)) xor (layer2_outputs(5722));
    outputs(4085) <= (layer2_outputs(132)) xor (layer2_outputs(5419));
    outputs(4086) <= layer2_outputs(3352);
    outputs(4087) <= (layer2_outputs(4418)) and not (layer2_outputs(9489));
    outputs(4088) <= layer2_outputs(6069);
    outputs(4089) <= layer2_outputs(6342);
    outputs(4090) <= (layer2_outputs(2712)) xor (layer2_outputs(7871));
    outputs(4091) <= '1';
    outputs(4092) <= not((layer2_outputs(3135)) and (layer2_outputs(2859)));
    outputs(4093) <= not((layer2_outputs(437)) xor (layer2_outputs(1805)));
    outputs(4094) <= not(layer2_outputs(9286));
    outputs(4095) <= layer2_outputs(1232);
    outputs(4096) <= layer2_outputs(7125);
    outputs(4097) <= not(layer2_outputs(6018));
    outputs(4098) <= not((layer2_outputs(5949)) xor (layer2_outputs(343)));
    outputs(4099) <= not(layer2_outputs(4703));
    outputs(4100) <= not(layer2_outputs(6228));
    outputs(4101) <= (layer2_outputs(5179)) or (layer2_outputs(4149));
    outputs(4102) <= layer2_outputs(9371);
    outputs(4103) <= not(layer2_outputs(9360));
    outputs(4104) <= (layer2_outputs(3782)) xor (layer2_outputs(80));
    outputs(4105) <= not(layer2_outputs(6545)) or (layer2_outputs(9895));
    outputs(4106) <= layer2_outputs(5652);
    outputs(4107) <= (layer2_outputs(1657)) xor (layer2_outputs(7860));
    outputs(4108) <= not(layer2_outputs(9637));
    outputs(4109) <= not(layer2_outputs(2447));
    outputs(4110) <= layer2_outputs(3042);
    outputs(4111) <= layer2_outputs(2679);
    outputs(4112) <= layer2_outputs(3219);
    outputs(4113) <= not(layer2_outputs(8960));
    outputs(4114) <= not(layer2_outputs(8902));
    outputs(4115) <= (layer2_outputs(2269)) xor (layer2_outputs(4079));
    outputs(4116) <= not(layer2_outputs(4115));
    outputs(4117) <= layer2_outputs(9242);
    outputs(4118) <= (layer2_outputs(7659)) xor (layer2_outputs(1913));
    outputs(4119) <= (layer2_outputs(7864)) and not (layer2_outputs(8615));
    outputs(4120) <= not((layer2_outputs(2344)) and (layer2_outputs(7027)));
    outputs(4121) <= not(layer2_outputs(8297));
    outputs(4122) <= not((layer2_outputs(6387)) xor (layer2_outputs(5756)));
    outputs(4123) <= not(layer2_outputs(7709));
    outputs(4124) <= not(layer2_outputs(7865)) or (layer2_outputs(2652));
    outputs(4125) <= not((layer2_outputs(7711)) or (layer2_outputs(6982)));
    outputs(4126) <= (layer2_outputs(4077)) and not (layer2_outputs(6884));
    outputs(4127) <= not(layer2_outputs(9340)) or (layer2_outputs(9351));
    outputs(4128) <= not(layer2_outputs(2707));
    outputs(4129) <= (layer2_outputs(566)) and not (layer2_outputs(1891));
    outputs(4130) <= (layer2_outputs(5525)) xor (layer2_outputs(2940));
    outputs(4131) <= not(layer2_outputs(2972));
    outputs(4132) <= layer2_outputs(5244);
    outputs(4133) <= layer2_outputs(9917);
    outputs(4134) <= (layer2_outputs(6479)) and not (layer2_outputs(6165));
    outputs(4135) <= layer2_outputs(5310);
    outputs(4136) <= layer2_outputs(10049);
    outputs(4137) <= layer2_outputs(5414);
    outputs(4138) <= not((layer2_outputs(2328)) xor (layer2_outputs(4986)));
    outputs(4139) <= layer2_outputs(3390);
    outputs(4140) <= (layer2_outputs(5882)) xor (layer2_outputs(3844));
    outputs(4141) <= not(layer2_outputs(317));
    outputs(4142) <= layer2_outputs(7347);
    outputs(4143) <= layer2_outputs(4075);
    outputs(4144) <= (layer2_outputs(8006)) and not (layer2_outputs(7341));
    outputs(4145) <= layer2_outputs(5814);
    outputs(4146) <= not(layer2_outputs(1621));
    outputs(4147) <= layer2_outputs(4065);
    outputs(4148) <= (layer2_outputs(4485)) xor (layer2_outputs(3438));
    outputs(4149) <= not(layer2_outputs(9770));
    outputs(4150) <= not(layer2_outputs(7594));
    outputs(4151) <= layer2_outputs(8024);
    outputs(4152) <= not((layer2_outputs(5289)) xor (layer2_outputs(9431)));
    outputs(4153) <= not(layer2_outputs(8846));
    outputs(4154) <= not(layer2_outputs(8114));
    outputs(4155) <= (layer2_outputs(3811)) xor (layer2_outputs(3244));
    outputs(4156) <= not(layer2_outputs(6715));
    outputs(4157) <= not((layer2_outputs(8679)) xor (layer2_outputs(8008)));
    outputs(4158) <= (layer2_outputs(10110)) and (layer2_outputs(9432));
    outputs(4159) <= (layer2_outputs(4428)) or (layer2_outputs(1854));
    outputs(4160) <= not(layer2_outputs(10234));
    outputs(4161) <= not((layer2_outputs(2463)) xor (layer2_outputs(8116)));
    outputs(4162) <= (layer2_outputs(1338)) and not (layer2_outputs(724));
    outputs(4163) <= layer2_outputs(8789);
    outputs(4164) <= layer2_outputs(5509);
    outputs(4165) <= not(layer2_outputs(5518));
    outputs(4166) <= not(layer2_outputs(3583));
    outputs(4167) <= not(layer2_outputs(1160));
    outputs(4168) <= layer2_outputs(678);
    outputs(4169) <= not((layer2_outputs(9536)) xor (layer2_outputs(8518)));
    outputs(4170) <= layer2_outputs(4774);
    outputs(4171) <= (layer2_outputs(4611)) xor (layer2_outputs(3563));
    outputs(4172) <= layer2_outputs(2767);
    outputs(4173) <= (layer2_outputs(940)) or (layer2_outputs(8292));
    outputs(4174) <= not(layer2_outputs(1659));
    outputs(4175) <= (layer2_outputs(8119)) and not (layer2_outputs(375));
    outputs(4176) <= not(layer2_outputs(3548));
    outputs(4177) <= not(layer2_outputs(1191));
    outputs(4178) <= layer2_outputs(1682);
    outputs(4179) <= not(layer2_outputs(7607));
    outputs(4180) <= not((layer2_outputs(6667)) xor (layer2_outputs(2552)));
    outputs(4181) <= (layer2_outputs(4437)) xor (layer2_outputs(469));
    outputs(4182) <= not(layer2_outputs(5579));
    outputs(4183) <= not(layer2_outputs(5925));
    outputs(4184) <= not(layer2_outputs(9026));
    outputs(4185) <= not((layer2_outputs(8659)) xor (layer2_outputs(3010)));
    outputs(4186) <= layer2_outputs(1042);
    outputs(4187) <= layer2_outputs(3210);
    outputs(4188) <= layer2_outputs(3636);
    outputs(4189) <= layer2_outputs(6130);
    outputs(4190) <= layer2_outputs(5773);
    outputs(4191) <= not((layer2_outputs(161)) or (layer2_outputs(3820)));
    outputs(4192) <= not((layer2_outputs(10034)) xor (layer2_outputs(3238)));
    outputs(4193) <= not(layer2_outputs(3561));
    outputs(4194) <= not((layer2_outputs(7561)) xor (layer2_outputs(8487)));
    outputs(4195) <= not(layer2_outputs(2855));
    outputs(4196) <= not(layer2_outputs(4225));
    outputs(4197) <= layer2_outputs(1278);
    outputs(4198) <= layer2_outputs(6196);
    outputs(4199) <= not(layer2_outputs(7880));
    outputs(4200) <= layer2_outputs(4510);
    outputs(4201) <= (layer2_outputs(4779)) xor (layer2_outputs(10212));
    outputs(4202) <= (layer2_outputs(7597)) xor (layer2_outputs(2040));
    outputs(4203) <= (layer2_outputs(3225)) xor (layer2_outputs(5136));
    outputs(4204) <= layer2_outputs(7206);
    outputs(4205) <= not(layer2_outputs(2461));
    outputs(4206) <= not(layer2_outputs(6595));
    outputs(4207) <= layer2_outputs(5409);
    outputs(4208) <= not((layer2_outputs(3527)) or (layer2_outputs(1988)));
    outputs(4209) <= not(layer2_outputs(8825));
    outputs(4210) <= not(layer2_outputs(2699));
    outputs(4211) <= not(layer2_outputs(6901));
    outputs(4212) <= not((layer2_outputs(2293)) and (layer2_outputs(8074)));
    outputs(4213) <= not(layer2_outputs(3166));
    outputs(4214) <= (layer2_outputs(829)) xor (layer2_outputs(508));
    outputs(4215) <= (layer2_outputs(6877)) xor (layer2_outputs(9112));
    outputs(4216) <= not(layer2_outputs(4819)) or (layer2_outputs(5585));
    outputs(4217) <= not(layer2_outputs(9627));
    outputs(4218) <= not((layer2_outputs(4908)) xor (layer2_outputs(762)));
    outputs(4219) <= layer2_outputs(5921);
    outputs(4220) <= not(layer2_outputs(3492));
    outputs(4221) <= (layer2_outputs(6407)) or (layer2_outputs(442));
    outputs(4222) <= not(layer2_outputs(1981));
    outputs(4223) <= not(layer2_outputs(4885));
    outputs(4224) <= not(layer2_outputs(5524));
    outputs(4225) <= not(layer2_outputs(7562));
    outputs(4226) <= layer2_outputs(6742);
    outputs(4227) <= not(layer2_outputs(1356));
    outputs(4228) <= not(layer2_outputs(8841));
    outputs(4229) <= not(layer2_outputs(6165));
    outputs(4230) <= not(layer2_outputs(8048));
    outputs(4231) <= layer2_outputs(4713);
    outputs(4232) <= not(layer2_outputs(6189));
    outputs(4233) <= layer2_outputs(120);
    outputs(4234) <= (layer2_outputs(16)) xor (layer2_outputs(2834));
    outputs(4235) <= layer2_outputs(8992);
    outputs(4236) <= (layer2_outputs(6168)) and not (layer2_outputs(9972));
    outputs(4237) <= not((layer2_outputs(3562)) xor (layer2_outputs(2171)));
    outputs(4238) <= layer2_outputs(3659);
    outputs(4239) <= (layer2_outputs(9802)) xor (layer2_outputs(3931));
    outputs(4240) <= not(layer2_outputs(5566));
    outputs(4241) <= (layer2_outputs(7964)) xor (layer2_outputs(4727));
    outputs(4242) <= (layer2_outputs(6891)) xor (layer2_outputs(4228));
    outputs(4243) <= layer2_outputs(7974);
    outputs(4244) <= layer2_outputs(6794);
    outputs(4245) <= (layer2_outputs(7722)) and not (layer2_outputs(4958));
    outputs(4246) <= not((layer2_outputs(1863)) or (layer2_outputs(9110)));
    outputs(4247) <= not(layer2_outputs(67));
    outputs(4248) <= layer2_outputs(4871);
    outputs(4249) <= layer2_outputs(4742);
    outputs(4250) <= not((layer2_outputs(2106)) xor (layer2_outputs(2829)));
    outputs(4251) <= layer2_outputs(7483);
    outputs(4252) <= layer2_outputs(1408);
    outputs(4253) <= layer2_outputs(3859);
    outputs(4254) <= layer2_outputs(4100);
    outputs(4255) <= not(layer2_outputs(7412));
    outputs(4256) <= layer2_outputs(6721);
    outputs(4257) <= not(layer2_outputs(2856));
    outputs(4258) <= layer2_outputs(6367);
    outputs(4259) <= layer2_outputs(5379);
    outputs(4260) <= not((layer2_outputs(7975)) xor (layer2_outputs(837)));
    outputs(4261) <= (layer2_outputs(4522)) and not (layer2_outputs(453));
    outputs(4262) <= layer2_outputs(10030);
    outputs(4263) <= layer2_outputs(8129);
    outputs(4264) <= layer2_outputs(1898);
    outputs(4265) <= not(layer2_outputs(6110));
    outputs(4266) <= not(layer2_outputs(7555));
    outputs(4267) <= (layer2_outputs(5114)) xor (layer2_outputs(3608));
    outputs(4268) <= (layer2_outputs(2973)) and not (layer2_outputs(3826));
    outputs(4269) <= not(layer2_outputs(8965));
    outputs(4270) <= not(layer2_outputs(1373));
    outputs(4271) <= layer2_outputs(6259);
    outputs(4272) <= not((layer2_outputs(594)) xor (layer2_outputs(10134)));
    outputs(4273) <= not((layer2_outputs(578)) xor (layer2_outputs(5943)));
    outputs(4274) <= layer2_outputs(4499);
    outputs(4275) <= not(layer2_outputs(8684));
    outputs(4276) <= layer2_outputs(10099);
    outputs(4277) <= not((layer2_outputs(1227)) xor (layer2_outputs(7867)));
    outputs(4278) <= (layer2_outputs(6240)) xor (layer2_outputs(7793));
    outputs(4279) <= (layer2_outputs(7392)) xor (layer2_outputs(3953));
    outputs(4280) <= not((layer2_outputs(2355)) xor (layer2_outputs(1495)));
    outputs(4281) <= not((layer2_outputs(4669)) xor (layer2_outputs(4814)));
    outputs(4282) <= not((layer2_outputs(6930)) xor (layer2_outputs(8623)));
    outputs(4283) <= not(layer2_outputs(6345));
    outputs(4284) <= not(layer2_outputs(2658)) or (layer2_outputs(6939));
    outputs(4285) <= not(layer2_outputs(2497));
    outputs(4286) <= layer2_outputs(1885);
    outputs(4287) <= layer2_outputs(8096);
    outputs(4288) <= layer2_outputs(6086);
    outputs(4289) <= (layer2_outputs(1075)) and (layer2_outputs(6967));
    outputs(4290) <= layer2_outputs(6999);
    outputs(4291) <= not(layer2_outputs(1528));
    outputs(4292) <= layer2_outputs(4327);
    outputs(4293) <= not(layer2_outputs(18));
    outputs(4294) <= (layer2_outputs(7863)) xor (layer2_outputs(2550));
    outputs(4295) <= not(layer2_outputs(2348));
    outputs(4296) <= (layer2_outputs(10142)) xor (layer2_outputs(3589));
    outputs(4297) <= not(layer2_outputs(8029));
    outputs(4298) <= layer2_outputs(2663);
    outputs(4299) <= (layer2_outputs(5080)) xor (layer2_outputs(8552));
    outputs(4300) <= not((layer2_outputs(2388)) or (layer2_outputs(572)));
    outputs(4301) <= not(layer2_outputs(1518));
    outputs(4302) <= not((layer2_outputs(6733)) xor (layer2_outputs(2252)));
    outputs(4303) <= layer2_outputs(2700);
    outputs(4304) <= layer2_outputs(10153);
    outputs(4305) <= not((layer2_outputs(8272)) and (layer2_outputs(6100)));
    outputs(4306) <= not(layer2_outputs(5974));
    outputs(4307) <= layer2_outputs(2924);
    outputs(4308) <= layer2_outputs(3318);
    outputs(4309) <= layer2_outputs(919);
    outputs(4310) <= (layer2_outputs(7520)) xor (layer2_outputs(6003));
    outputs(4311) <= not((layer2_outputs(223)) xor (layer2_outputs(5082)));
    outputs(4312) <= not((layer2_outputs(8509)) xor (layer2_outputs(6043)));
    outputs(4313) <= layer2_outputs(1526);
    outputs(4314) <= not(layer2_outputs(6956));
    outputs(4315) <= layer2_outputs(3242);
    outputs(4316) <= layer2_outputs(3143);
    outputs(4317) <= not(layer2_outputs(1732));
    outputs(4318) <= (layer2_outputs(2257)) and (layer2_outputs(4245));
    outputs(4319) <= not((layer2_outputs(5664)) and (layer2_outputs(4315)));
    outputs(4320) <= layer2_outputs(1733);
    outputs(4321) <= layer2_outputs(4487);
    outputs(4322) <= (layer2_outputs(5942)) or (layer2_outputs(3687));
    outputs(4323) <= layer2_outputs(2642);
    outputs(4324) <= layer2_outputs(8871);
    outputs(4325) <= not(layer2_outputs(1959));
    outputs(4326) <= (layer2_outputs(5654)) and (layer2_outputs(3170));
    outputs(4327) <= not(layer2_outputs(6803));
    outputs(4328) <= layer2_outputs(6023);
    outputs(4329) <= not(layer2_outputs(4466));
    outputs(4330) <= not(layer2_outputs(8364));
    outputs(4331) <= not(layer2_outputs(8695));
    outputs(4332) <= layer2_outputs(6491);
    outputs(4333) <= layer2_outputs(7837);
    outputs(4334) <= not((layer2_outputs(7732)) and (layer2_outputs(3561)));
    outputs(4335) <= not(layer2_outputs(9095));
    outputs(4336) <= not(layer2_outputs(9301));
    outputs(4337) <= layer2_outputs(8998);
    outputs(4338) <= layer2_outputs(1687);
    outputs(4339) <= (layer2_outputs(3869)) xor (layer2_outputs(9055));
    outputs(4340) <= layer2_outputs(2744);
    outputs(4341) <= not(layer2_outputs(500));
    outputs(4342) <= layer2_outputs(3157);
    outputs(4343) <= not(layer2_outputs(1049));
    outputs(4344) <= layer2_outputs(6945);
    outputs(4345) <= not(layer2_outputs(1040));
    outputs(4346) <= not(layer2_outputs(8661));
    outputs(4347) <= layer2_outputs(4623);
    outputs(4348) <= (layer2_outputs(1579)) xor (layer2_outputs(4214));
    outputs(4349) <= (layer2_outputs(2876)) and not (layer2_outputs(6343));
    outputs(4350) <= (layer2_outputs(4974)) or (layer2_outputs(1229));
    outputs(4351) <= not(layer2_outputs(2173));
    outputs(4352) <= (layer2_outputs(5445)) xor (layer2_outputs(9597));
    outputs(4353) <= (layer2_outputs(9892)) and not (layer2_outputs(5243));
    outputs(4354) <= not(layer2_outputs(8507));
    outputs(4355) <= not(layer2_outputs(6382));
    outputs(4356) <= not(layer2_outputs(2335));
    outputs(4357) <= layer2_outputs(1710);
    outputs(4358) <= (layer2_outputs(807)) xor (layer2_outputs(2902));
    outputs(4359) <= not(layer2_outputs(10131));
    outputs(4360) <= not(layer2_outputs(4850));
    outputs(4361) <= (layer2_outputs(3613)) and not (layer2_outputs(5596));
    outputs(4362) <= (layer2_outputs(1650)) xor (layer2_outputs(7771));
    outputs(4363) <= layer2_outputs(7124);
    outputs(4364) <= not((layer2_outputs(3071)) xor (layer2_outputs(4676)));
    outputs(4365) <= not(layer2_outputs(125));
    outputs(4366) <= layer2_outputs(10037);
    outputs(4367) <= not(layer2_outputs(1147));
    outputs(4368) <= layer2_outputs(7721);
    outputs(4369) <= not(layer2_outputs(5343)) or (layer2_outputs(757));
    outputs(4370) <= layer2_outputs(2164);
    outputs(4371) <= (layer2_outputs(4758)) and (layer2_outputs(1562));
    outputs(4372) <= not((layer2_outputs(5457)) xor (layer2_outputs(6061)));
    outputs(4373) <= layer2_outputs(202);
    outputs(4374) <= not(layer2_outputs(1519));
    outputs(4375) <= (layer2_outputs(2987)) and not (layer2_outputs(8474));
    outputs(4376) <= (layer2_outputs(522)) and not (layer2_outputs(5303));
    outputs(4377) <= layer2_outputs(8030);
    outputs(4378) <= (layer2_outputs(9387)) xor (layer2_outputs(4222));
    outputs(4379) <= layer2_outputs(1123);
    outputs(4380) <= (layer2_outputs(9385)) and (layer2_outputs(9661));
    outputs(4381) <= (layer2_outputs(4727)) xor (layer2_outputs(7552));
    outputs(4382) <= not((layer2_outputs(1638)) xor (layer2_outputs(1761)));
    outputs(4383) <= (layer2_outputs(1209)) xor (layer2_outputs(9434));
    outputs(4384) <= (layer2_outputs(4486)) xor (layer2_outputs(5910));
    outputs(4385) <= layer2_outputs(7573);
    outputs(4386) <= not((layer2_outputs(8830)) xor (layer2_outputs(2883)));
    outputs(4387) <= layer2_outputs(5353);
    outputs(4388) <= not((layer2_outputs(3219)) xor (layer2_outputs(8085)));
    outputs(4389) <= not(layer2_outputs(4672));
    outputs(4390) <= not(layer2_outputs(5400));
    outputs(4391) <= not((layer2_outputs(7888)) or (layer2_outputs(9814)));
    outputs(4392) <= (layer2_outputs(7718)) xor (layer2_outputs(10001));
    outputs(4393) <= layer2_outputs(7706);
    outputs(4394) <= layer2_outputs(8938);
    outputs(4395) <= not(layer2_outputs(6113));
    outputs(4396) <= not(layer2_outputs(1584));
    outputs(4397) <= not((layer2_outputs(6651)) xor (layer2_outputs(5595)));
    outputs(4398) <= layer2_outputs(1100);
    outputs(4399) <= layer2_outputs(9799);
    outputs(4400) <= not((layer2_outputs(4759)) and (layer2_outputs(9221)));
    outputs(4401) <= (layer2_outputs(4747)) and (layer2_outputs(8339));
    outputs(4402) <= not(layer2_outputs(6760));
    outputs(4403) <= layer2_outputs(8012);
    outputs(4404) <= layer2_outputs(1274);
    outputs(4405) <= (layer2_outputs(4125)) xor (layer2_outputs(9839));
    outputs(4406) <= not(layer2_outputs(6762));
    outputs(4407) <= not(layer2_outputs(752));
    outputs(4408) <= not(layer2_outputs(1979)) or (layer2_outputs(8268));
    outputs(4409) <= not(layer2_outputs(3459));
    outputs(4410) <= layer2_outputs(7392);
    outputs(4411) <= not(layer2_outputs(1947));
    outputs(4412) <= not(layer2_outputs(267));
    outputs(4413) <= not((layer2_outputs(1375)) xor (layer2_outputs(8337)));
    outputs(4414) <= layer2_outputs(5999);
    outputs(4415) <= layer2_outputs(8233);
    outputs(4416) <= not((layer2_outputs(4375)) xor (layer2_outputs(2428)));
    outputs(4417) <= layer2_outputs(9708);
    outputs(4418) <= not(layer2_outputs(2599));
    outputs(4419) <= not(layer2_outputs(5113));
    outputs(4420) <= not((layer2_outputs(6641)) xor (layer2_outputs(8731)));
    outputs(4421) <= not(layer2_outputs(5866));
    outputs(4422) <= layer2_outputs(8073);
    outputs(4423) <= not(layer2_outputs(10231));
    outputs(4424) <= not((layer2_outputs(2666)) xor (layer2_outputs(4876)));
    outputs(4425) <= (layer2_outputs(9807)) xor (layer2_outputs(8352));
    outputs(4426) <= not((layer2_outputs(2190)) xor (layer2_outputs(1998)));
    outputs(4427) <= not(layer2_outputs(7436));
    outputs(4428) <= not(layer2_outputs(1875));
    outputs(4429) <= not((layer2_outputs(9366)) xor (layer2_outputs(59)));
    outputs(4430) <= not(layer2_outputs(5018)) or (layer2_outputs(9775));
    outputs(4431) <= layer2_outputs(2761);
    outputs(4432) <= layer2_outputs(26);
    outputs(4433) <= layer2_outputs(7238);
    outputs(4434) <= layer2_outputs(361);
    outputs(4435) <= (layer2_outputs(3212)) xor (layer2_outputs(2540));
    outputs(4436) <= not((layer2_outputs(8104)) or (layer2_outputs(1483)));
    outputs(4437) <= (layer2_outputs(6316)) xor (layer2_outputs(4943));
    outputs(4438) <= layer2_outputs(6181);
    outputs(4439) <= not(layer2_outputs(7668)) or (layer2_outputs(2874));
    outputs(4440) <= not(layer2_outputs(5705));
    outputs(4441) <= layer2_outputs(8648);
    outputs(4442) <= not(layer2_outputs(3094));
    outputs(4443) <= (layer2_outputs(2442)) and (layer2_outputs(24));
    outputs(4444) <= layer2_outputs(1324);
    outputs(4445) <= not(layer2_outputs(9077));
    outputs(4446) <= layer2_outputs(7537);
    outputs(4447) <= layer2_outputs(2515);
    outputs(4448) <= (layer2_outputs(6782)) and not (layer2_outputs(4760));
    outputs(4449) <= layer2_outputs(2383);
    outputs(4450) <= (layer2_outputs(3256)) xor (layer2_outputs(7153));
    outputs(4451) <= layer2_outputs(10025);
    outputs(4452) <= layer2_outputs(8845);
    outputs(4453) <= not(layer2_outputs(2968));
    outputs(4454) <= (layer2_outputs(4085)) and not (layer2_outputs(6743));
    outputs(4455) <= not((layer2_outputs(6236)) xor (layer2_outputs(1442)));
    outputs(4456) <= not(layer2_outputs(5540));
    outputs(4457) <= not(layer2_outputs(495));
    outputs(4458) <= layer2_outputs(7195);
    outputs(4459) <= layer2_outputs(3987);
    outputs(4460) <= layer2_outputs(1382);
    outputs(4461) <= layer2_outputs(7685);
    outputs(4462) <= (layer2_outputs(956)) and not (layer2_outputs(1277));
    outputs(4463) <= not(layer2_outputs(9737));
    outputs(4464) <= (layer2_outputs(7521)) xor (layer2_outputs(5489));
    outputs(4465) <= (layer2_outputs(5655)) xor (layer2_outputs(3188));
    outputs(4466) <= not(layer2_outputs(2613));
    outputs(4467) <= (layer2_outputs(6508)) and not (layer2_outputs(5894));
    outputs(4468) <= not(layer2_outputs(302));
    outputs(4469) <= (layer2_outputs(4664)) and not (layer2_outputs(9742));
    outputs(4470) <= (layer2_outputs(1410)) and not (layer2_outputs(399));
    outputs(4471) <= layer2_outputs(8973);
    outputs(4472) <= (layer2_outputs(5527)) xor (layer2_outputs(4528));
    outputs(4473) <= layer2_outputs(4366);
    outputs(4474) <= layer2_outputs(6215);
    outputs(4475) <= not(layer2_outputs(220)) or (layer2_outputs(7148));
    outputs(4476) <= not(layer2_outputs(218));
    outputs(4477) <= layer2_outputs(2128);
    outputs(4478) <= not(layer2_outputs(9942));
    outputs(4479) <= layer2_outputs(1953);
    outputs(4480) <= not(layer2_outputs(261));
    outputs(4481) <= not(layer2_outputs(7063));
    outputs(4482) <= layer2_outputs(2912);
    outputs(4483) <= layer2_outputs(2466);
    outputs(4484) <= not(layer2_outputs(8978));
    outputs(4485) <= layer2_outputs(5159);
    outputs(4486) <= (layer2_outputs(9927)) xor (layer2_outputs(6058));
    outputs(4487) <= not(layer2_outputs(96));
    outputs(4488) <= layer2_outputs(2314);
    outputs(4489) <= layer2_outputs(6677);
    outputs(4490) <= layer2_outputs(1302);
    outputs(4491) <= not(layer2_outputs(884));
    outputs(4492) <= (layer2_outputs(2880)) and not (layer2_outputs(6868));
    outputs(4493) <= (layer2_outputs(4826)) and not (layer2_outputs(4912));
    outputs(4494) <= not(layer2_outputs(306));
    outputs(4495) <= layer2_outputs(7652);
    outputs(4496) <= layer2_outputs(6086);
    outputs(4497) <= not(layer2_outputs(10010));
    outputs(4498) <= layer2_outputs(3201);
    outputs(4499) <= layer2_outputs(5075);
    outputs(4500) <= layer2_outputs(4182);
    outputs(4501) <= layer2_outputs(5895);
    outputs(4502) <= not(layer2_outputs(74));
    outputs(4503) <= not(layer2_outputs(5594));
    outputs(4504) <= not(layer2_outputs(9492)) or (layer2_outputs(680));
    outputs(4505) <= not(layer2_outputs(6175));
    outputs(4506) <= layer2_outputs(3501);
    outputs(4507) <= not((layer2_outputs(4083)) xor (layer2_outputs(3191)));
    outputs(4508) <= layer2_outputs(1642);
    outputs(4509) <= not(layer2_outputs(4401));
    outputs(4510) <= not(layer2_outputs(8829));
    outputs(4511) <= not(layer2_outputs(4279));
    outputs(4512) <= layer2_outputs(4645);
    outputs(4513) <= layer2_outputs(9205);
    outputs(4514) <= (layer2_outputs(7641)) and not (layer2_outputs(2272));
    outputs(4515) <= not((layer2_outputs(2816)) xor (layer2_outputs(4625)));
    outputs(4516) <= not(layer2_outputs(1289));
    outputs(4517) <= layer2_outputs(6312);
    outputs(4518) <= layer2_outputs(2772);
    outputs(4519) <= layer2_outputs(7610);
    outputs(4520) <= layer2_outputs(9749);
    outputs(4521) <= not(layer2_outputs(5073)) or (layer2_outputs(5529));
    outputs(4522) <= not(layer2_outputs(8827));
    outputs(4523) <= not((layer2_outputs(3884)) or (layer2_outputs(6262)));
    outputs(4524) <= not(layer2_outputs(7775));
    outputs(4525) <= layer2_outputs(42);
    outputs(4526) <= not(layer2_outputs(5904));
    outputs(4527) <= (layer2_outputs(7245)) xor (layer2_outputs(9762));
    outputs(4528) <= not(layer2_outputs(5681)) or (layer2_outputs(6785));
    outputs(4529) <= (layer2_outputs(3379)) xor (layer2_outputs(10011));
    outputs(4530) <= not(layer2_outputs(9716));
    outputs(4531) <= not(layer2_outputs(6755));
    outputs(4532) <= not(layer2_outputs(7181));
    outputs(4533) <= layer2_outputs(127);
    outputs(4534) <= layer2_outputs(3101);
    outputs(4535) <= layer2_outputs(1404);
    outputs(4536) <= (layer2_outputs(6177)) and (layer2_outputs(5630));
    outputs(4537) <= not(layer2_outputs(6703));
    outputs(4538) <= not(layer2_outputs(3914));
    outputs(4539) <= layer2_outputs(2606);
    outputs(4540) <= (layer2_outputs(3096)) and not (layer2_outputs(1859));
    outputs(4541) <= not((layer2_outputs(1964)) xor (layer2_outputs(1896)));
    outputs(4542) <= not((layer2_outputs(3040)) xor (layer2_outputs(2502)));
    outputs(4543) <= not(layer2_outputs(8382));
    outputs(4544) <= not(layer2_outputs(654));
    outputs(4545) <= not(layer2_outputs(7502));
    outputs(4546) <= not((layer2_outputs(2902)) or (layer2_outputs(4715)));
    outputs(4547) <= not(layer2_outputs(8217));
    outputs(4548) <= not((layer2_outputs(4532)) xor (layer2_outputs(5487)));
    outputs(4549) <= not(layer2_outputs(9230));
    outputs(4550) <= not(layer2_outputs(124));
    outputs(4551) <= layer2_outputs(10109);
    outputs(4552) <= not((layer2_outputs(2644)) and (layer2_outputs(1372)));
    outputs(4553) <= not(layer2_outputs(5793));
    outputs(4554) <= layer2_outputs(8924);
    outputs(4555) <= not(layer2_outputs(4379));
    outputs(4556) <= not(layer2_outputs(10162));
    outputs(4557) <= not(layer2_outputs(552));
    outputs(4558) <= layer2_outputs(6368);
    outputs(4559) <= not(layer2_outputs(5167));
    outputs(4560) <= not(layer2_outputs(5238));
    outputs(4561) <= layer2_outputs(1274);
    outputs(4562) <= layer2_outputs(1341);
    outputs(4563) <= layer2_outputs(9205);
    outputs(4564) <= not(layer2_outputs(9633));
    outputs(4565) <= not(layer2_outputs(8086)) or (layer2_outputs(6496));
    outputs(4566) <= not((layer2_outputs(1825)) xor (layer2_outputs(4405)));
    outputs(4567) <= layer2_outputs(7921);
    outputs(4568) <= not((layer2_outputs(3877)) xor (layer2_outputs(6957)));
    outputs(4569) <= layer2_outputs(5191);
    outputs(4570) <= not(layer2_outputs(6478));
    outputs(4571) <= layer2_outputs(5288);
    outputs(4572) <= not(layer2_outputs(4129));
    outputs(4573) <= not(layer2_outputs(8792));
    outputs(4574) <= not(layer2_outputs(1314));
    outputs(4575) <= not((layer2_outputs(9321)) or (layer2_outputs(9036)));
    outputs(4576) <= (layer2_outputs(2897)) xor (layer2_outputs(6534));
    outputs(4577) <= not((layer2_outputs(9437)) and (layer2_outputs(6718)));
    outputs(4578) <= not(layer2_outputs(5453));
    outputs(4579) <= not(layer2_outputs(7872));
    outputs(4580) <= (layer2_outputs(3598)) and not (layer2_outputs(1602));
    outputs(4581) <= not(layer2_outputs(1013));
    outputs(4582) <= layer2_outputs(3995);
    outputs(4583) <= (layer2_outputs(7996)) xor (layer2_outputs(6577));
    outputs(4584) <= (layer2_outputs(7419)) xor (layer2_outputs(8211));
    outputs(4585) <= layer2_outputs(6087);
    outputs(4586) <= layer2_outputs(2258);
    outputs(4587) <= not(layer2_outputs(8147));
    outputs(4588) <= not((layer2_outputs(4351)) xor (layer2_outputs(1382)));
    outputs(4589) <= not(layer2_outputs(8130));
    outputs(4590) <= layer2_outputs(5454);
    outputs(4591) <= layer2_outputs(4655);
    outputs(4592) <= not((layer2_outputs(10078)) xor (layer2_outputs(3569)));
    outputs(4593) <= layer2_outputs(6607);
    outputs(4594) <= layer2_outputs(7468);
    outputs(4595) <= not((layer2_outputs(8821)) xor (layer2_outputs(5257)));
    outputs(4596) <= not(layer2_outputs(5606));
    outputs(4597) <= (layer2_outputs(5007)) and not (layer2_outputs(9691));
    outputs(4598) <= layer2_outputs(4140);
    outputs(4599) <= not(layer2_outputs(5605));
    outputs(4600) <= layer2_outputs(133);
    outputs(4601) <= not(layer2_outputs(10056));
    outputs(4602) <= layer2_outputs(723);
    outputs(4603) <= not((layer2_outputs(4990)) xor (layer2_outputs(8288)));
    outputs(4604) <= (layer2_outputs(2883)) xor (layer2_outputs(1729));
    outputs(4605) <= not(layer2_outputs(10100));
    outputs(4606) <= (layer2_outputs(7414)) xor (layer2_outputs(8157));
    outputs(4607) <= not(layer2_outputs(2499));
    outputs(4608) <= (layer2_outputs(1663)) xor (layer2_outputs(5941));
    outputs(4609) <= not(layer2_outputs(2480));
    outputs(4610) <= not(layer2_outputs(9585));
    outputs(4611) <= (layer2_outputs(9035)) xor (layer2_outputs(7204));
    outputs(4612) <= (layer2_outputs(5466)) xor (layer2_outputs(7820));
    outputs(4613) <= not((layer2_outputs(5351)) xor (layer2_outputs(400)));
    outputs(4614) <= not(layer2_outputs(2803));
    outputs(4615) <= layer2_outputs(2995);
    outputs(4616) <= layer2_outputs(6057);
    outputs(4617) <= (layer2_outputs(7010)) xor (layer2_outputs(551));
    outputs(4618) <= (layer2_outputs(4353)) and not (layer2_outputs(931));
    outputs(4619) <= layer2_outputs(4167);
    outputs(4620) <= not(layer2_outputs(5246));
    outputs(4621) <= not((layer2_outputs(9933)) xor (layer2_outputs(1865)));
    outputs(4622) <= layer2_outputs(9087);
    outputs(4623) <= layer2_outputs(4903);
    outputs(4624) <= layer2_outputs(3164);
    outputs(4625) <= layer2_outputs(1172);
    outputs(4626) <= not(layer2_outputs(10220));
    outputs(4627) <= layer2_outputs(10044);
    outputs(4628) <= not((layer2_outputs(159)) xor (layer2_outputs(8851)));
    outputs(4629) <= layer2_outputs(1359);
    outputs(4630) <= not(layer2_outputs(3847));
    outputs(4631) <= layer2_outputs(6220);
    outputs(4632) <= layer2_outputs(8317);
    outputs(4633) <= (layer2_outputs(3250)) xor (layer2_outputs(7470));
    outputs(4634) <= '1';
    outputs(4635) <= layer2_outputs(2735);
    outputs(4636) <= layer2_outputs(6158);
    outputs(4637) <= layer2_outputs(4513);
    outputs(4638) <= not(layer2_outputs(491));
    outputs(4639) <= not(layer2_outputs(2480));
    outputs(4640) <= not(layer2_outputs(9425));
    outputs(4641) <= layer2_outputs(10099);
    outputs(4642) <= (layer2_outputs(4969)) and (layer2_outputs(310));
    outputs(4643) <= not((layer2_outputs(123)) xor (layer2_outputs(8241)));
    outputs(4644) <= layer2_outputs(1806);
    outputs(4645) <= (layer2_outputs(970)) xor (layer2_outputs(6010));
    outputs(4646) <= layer2_outputs(4899);
    outputs(4647) <= layer2_outputs(7094);
    outputs(4648) <= not(layer2_outputs(3302));
    outputs(4649) <= (layer2_outputs(10076)) and not (layer2_outputs(5444));
    outputs(4650) <= not(layer2_outputs(2699));
    outputs(4651) <= not((layer2_outputs(8183)) and (layer2_outputs(8745)));
    outputs(4652) <= not(layer2_outputs(9058)) or (layer2_outputs(9651));
    outputs(4653) <= not(layer2_outputs(7581));
    outputs(4654) <= not(layer2_outputs(7313));
    outputs(4655) <= not(layer2_outputs(292));
    outputs(4656) <= layer2_outputs(4884);
    outputs(4657) <= layer2_outputs(9676);
    outputs(4658) <= not(layer2_outputs(4609));
    outputs(4659) <= (layer2_outputs(6967)) xor (layer2_outputs(1927));
    outputs(4660) <= not(layer2_outputs(8132));
    outputs(4661) <= layer2_outputs(8814);
    outputs(4662) <= not(layer2_outputs(4281));
    outputs(4663) <= not(layer2_outputs(9479));
    outputs(4664) <= layer2_outputs(7046);
    outputs(4665) <= not(layer2_outputs(7562));
    outputs(4666) <= not(layer2_outputs(9081));
    outputs(4667) <= layer2_outputs(5648);
    outputs(4668) <= not((layer2_outputs(8960)) xor (layer2_outputs(8299)));
    outputs(4669) <= not(layer2_outputs(5855));
    outputs(4670) <= not(layer2_outputs(5079));
    outputs(4671) <= (layer2_outputs(8719)) xor (layer2_outputs(2048));
    outputs(4672) <= layer2_outputs(9450);
    outputs(4673) <= (layer2_outputs(8431)) and (layer2_outputs(2339));
    outputs(4674) <= (layer2_outputs(8467)) xor (layer2_outputs(8522));
    outputs(4675) <= not(layer2_outputs(8635));
    outputs(4676) <= (layer2_outputs(114)) xor (layer2_outputs(3052));
    outputs(4677) <= not(layer2_outputs(8359));
    outputs(4678) <= not(layer2_outputs(80));
    outputs(4679) <= layer2_outputs(2901);
    outputs(4680) <= (layer2_outputs(7746)) xor (layer2_outputs(1754));
    outputs(4681) <= not(layer2_outputs(10102));
    outputs(4682) <= not(layer2_outputs(9716));
    outputs(4683) <= not(layer2_outputs(3166));
    outputs(4684) <= not(layer2_outputs(6869));
    outputs(4685) <= not((layer2_outputs(5917)) xor (layer2_outputs(6995)));
    outputs(4686) <= layer2_outputs(4052);
    outputs(4687) <= layer2_outputs(9128);
    outputs(4688) <= layer2_outputs(8087);
    outputs(4689) <= not(layer2_outputs(7303));
    outputs(4690) <= not(layer2_outputs(5395));
    outputs(4691) <= layer2_outputs(6702);
    outputs(4692) <= not((layer2_outputs(2213)) xor (layer2_outputs(9661)));
    outputs(4693) <= not(layer2_outputs(4375));
    outputs(4694) <= (layer2_outputs(8125)) and (layer2_outputs(7432));
    outputs(4695) <= layer2_outputs(7041);
    outputs(4696) <= not((layer2_outputs(7554)) xor (layer2_outputs(9072)));
    outputs(4697) <= layer2_outputs(1043);
    outputs(4698) <= not(layer2_outputs(8173));
    outputs(4699) <= not(layer2_outputs(349)) or (layer2_outputs(2957));
    outputs(4700) <= not((layer2_outputs(1029)) and (layer2_outputs(7593)));
    outputs(4701) <= not((layer2_outputs(9154)) and (layer2_outputs(2104)));
    outputs(4702) <= not((layer2_outputs(5314)) xor (layer2_outputs(2918)));
    outputs(4703) <= (layer2_outputs(10115)) and not (layer2_outputs(9771));
    outputs(4704) <= (layer2_outputs(623)) xor (layer2_outputs(3464));
    outputs(4705) <= (layer2_outputs(8491)) or (layer2_outputs(840));
    outputs(4706) <= (layer2_outputs(1842)) xor (layer2_outputs(2483));
    outputs(4707) <= not(layer2_outputs(7314));
    outputs(4708) <= not(layer2_outputs(801)) or (layer2_outputs(9146));
    outputs(4709) <= layer2_outputs(3159);
    outputs(4710) <= layer2_outputs(8862);
    outputs(4711) <= not(layer2_outputs(419)) or (layer2_outputs(8515));
    outputs(4712) <= layer2_outputs(295);
    outputs(4713) <= layer2_outputs(7141);
    outputs(4714) <= not((layer2_outputs(1305)) or (layer2_outputs(558)));
    outputs(4715) <= not(layer2_outputs(8684));
    outputs(4716) <= layer2_outputs(1585);
    outputs(4717) <= (layer2_outputs(9445)) and (layer2_outputs(1035));
    outputs(4718) <= not(layer2_outputs(1293));
    outputs(4719) <= not(layer2_outputs(2426));
    outputs(4720) <= not((layer2_outputs(1589)) xor (layer2_outputs(1895)));
    outputs(4721) <= not(layer2_outputs(9070));
    outputs(4722) <= (layer2_outputs(1627)) and not (layer2_outputs(2309));
    outputs(4723) <= layer2_outputs(7525);
    outputs(4724) <= not(layer2_outputs(9851));
    outputs(4725) <= layer2_outputs(4038);
    outputs(4726) <= layer2_outputs(9993);
    outputs(4727) <= not(layer2_outputs(3756));
    outputs(4728) <= (layer2_outputs(2877)) and not (layer2_outputs(7690));
    outputs(4729) <= not(layer2_outputs(8332));
    outputs(4730) <= not(layer2_outputs(2192));
    outputs(4731) <= layer2_outputs(1418);
    outputs(4732) <= layer2_outputs(8041);
    outputs(4733) <= layer2_outputs(2148);
    outputs(4734) <= not(layer2_outputs(2482));
    outputs(4735) <= (layer2_outputs(430)) and (layer2_outputs(3083));
    outputs(4736) <= not(layer2_outputs(3491));
    outputs(4737) <= layer2_outputs(2324);
    outputs(4738) <= layer2_outputs(6152);
    outputs(4739) <= (layer2_outputs(3400)) xor (layer2_outputs(4572));
    outputs(4740) <= not(layer2_outputs(8109));
    outputs(4741) <= layer2_outputs(9303);
    outputs(4742) <= layer2_outputs(756);
    outputs(4743) <= layer2_outputs(3024);
    outputs(4744) <= not((layer2_outputs(3371)) xor (layer2_outputs(4007)));
    outputs(4745) <= layer2_outputs(476);
    outputs(4746) <= not(layer2_outputs(5671));
    outputs(4747) <= not(layer2_outputs(358));
    outputs(4748) <= not(layer2_outputs(5171));
    outputs(4749) <= not(layer2_outputs(4061));
    outputs(4750) <= not(layer2_outputs(4998));
    outputs(4751) <= not((layer2_outputs(2081)) xor (layer2_outputs(2582)));
    outputs(4752) <= not((layer2_outputs(8339)) or (layer2_outputs(2147)));
    outputs(4753) <= layer2_outputs(8593);
    outputs(4754) <= layer2_outputs(4412);
    outputs(4755) <= not((layer2_outputs(10059)) xor (layer2_outputs(2680)));
    outputs(4756) <= layer2_outputs(8008);
    outputs(4757) <= not((layer2_outputs(7773)) xor (layer2_outputs(570)));
    outputs(4758) <= not((layer2_outputs(2704)) xor (layer2_outputs(9243)));
    outputs(4759) <= (layer2_outputs(3450)) xor (layer2_outputs(6959));
    outputs(4760) <= layer2_outputs(1879);
    outputs(4761) <= layer2_outputs(5659);
    outputs(4762) <= not(layer2_outputs(3079));
    outputs(4763) <= (layer2_outputs(2289)) xor (layer2_outputs(4263));
    outputs(4764) <= not(layer2_outputs(124));
    outputs(4765) <= not((layer2_outputs(7869)) xor (layer2_outputs(1569)));
    outputs(4766) <= not((layer2_outputs(8141)) and (layer2_outputs(2169)));
    outputs(4767) <= (layer2_outputs(1328)) and (layer2_outputs(4111));
    outputs(4768) <= layer2_outputs(1432);
    outputs(4769) <= not((layer2_outputs(6458)) xor (layer2_outputs(3746)));
    outputs(4770) <= not((layer2_outputs(5718)) or (layer2_outputs(2974)));
    outputs(4771) <= (layer2_outputs(1271)) and (layer2_outputs(7432));
    outputs(4772) <= layer2_outputs(7584);
    outputs(4773) <= layer2_outputs(9096);
    outputs(4774) <= not(layer2_outputs(4559));
    outputs(4775) <= (layer2_outputs(5601)) xor (layer2_outputs(8013));
    outputs(4776) <= layer2_outputs(579);
    outputs(4777) <= layer2_outputs(7827);
    outputs(4778) <= not(layer2_outputs(6388));
    outputs(4779) <= not(layer2_outputs(10004));
    outputs(4780) <= not(layer2_outputs(7320));
    outputs(4781) <= not(layer2_outputs(3887));
    outputs(4782) <= layer2_outputs(9526);
    outputs(4783) <= not(layer2_outputs(2969));
    outputs(4784) <= (layer2_outputs(2493)) xor (layer2_outputs(9833));
    outputs(4785) <= layer2_outputs(1946);
    outputs(4786) <= layer2_outputs(9727);
    outputs(4787) <= layer2_outputs(2807);
    outputs(4788) <= (layer2_outputs(1913)) xor (layer2_outputs(5037));
    outputs(4789) <= layer2_outputs(8082);
    outputs(4790) <= not((layer2_outputs(3391)) xor (layer2_outputs(5537)));
    outputs(4791) <= (layer2_outputs(1641)) xor (layer2_outputs(2247));
    outputs(4792) <= not(layer2_outputs(1378));
    outputs(4793) <= layer2_outputs(6398);
    outputs(4794) <= layer2_outputs(4717);
    outputs(4795) <= not(layer2_outputs(5927));
    outputs(4796) <= (layer2_outputs(2033)) and not (layer2_outputs(2246));
    outputs(4797) <= not((layer2_outputs(6612)) xor (layer2_outputs(9007)));
    outputs(4798) <= not(layer2_outputs(1604));
    outputs(4799) <= (layer2_outputs(8274)) and not (layer2_outputs(3858));
    outputs(4800) <= not(layer2_outputs(3959));
    outputs(4801) <= (layer2_outputs(8887)) xor (layer2_outputs(3926));
    outputs(4802) <= not(layer2_outputs(9246)) or (layer2_outputs(3413));
    outputs(4803) <= (layer2_outputs(3975)) xor (layer2_outputs(4066));
    outputs(4804) <= layer2_outputs(2262);
    outputs(4805) <= not((layer2_outputs(4346)) xor (layer2_outputs(6863)));
    outputs(4806) <= (layer2_outputs(7023)) xor (layer2_outputs(1666));
    outputs(4807) <= not(layer2_outputs(9493));
    outputs(4808) <= layer2_outputs(7312);
    outputs(4809) <= (layer2_outputs(2860)) xor (layer2_outputs(3181));
    outputs(4810) <= layer2_outputs(1646);
    outputs(4811) <= (layer2_outputs(9174)) or (layer2_outputs(8571));
    outputs(4812) <= layer2_outputs(3822);
    outputs(4813) <= (layer2_outputs(2556)) xor (layer2_outputs(770));
    outputs(4814) <= not(layer2_outputs(242));
    outputs(4815) <= layer2_outputs(550);
    outputs(4816) <= (layer2_outputs(5812)) and not (layer2_outputs(6117));
    outputs(4817) <= layer2_outputs(1341);
    outputs(4818) <= (layer2_outputs(3030)) xor (layer2_outputs(743));
    outputs(4819) <= layer2_outputs(4633);
    outputs(4820) <= not(layer2_outputs(6134));
    outputs(4821) <= not(layer2_outputs(1559));
    outputs(4822) <= not(layer2_outputs(4453));
    outputs(4823) <= not(layer2_outputs(5842));
    outputs(4824) <= not(layer2_outputs(651));
    outputs(4825) <= not((layer2_outputs(6730)) xor (layer2_outputs(129)));
    outputs(4826) <= not(layer2_outputs(4924));
    outputs(4827) <= not(layer2_outputs(1916));
    outputs(4828) <= layer2_outputs(7334);
    outputs(4829) <= not(layer2_outputs(2313));
    outputs(4830) <= not(layer2_outputs(332));
    outputs(4831) <= not(layer2_outputs(8834)) or (layer2_outputs(3342));
    outputs(4832) <= (layer2_outputs(9243)) and not (layer2_outputs(3865));
    outputs(4833) <= not((layer2_outputs(7366)) xor (layer2_outputs(6353)));
    outputs(4834) <= not(layer2_outputs(6203));
    outputs(4835) <= not(layer2_outputs(1356));
    outputs(4836) <= not(layer2_outputs(955));
    outputs(4837) <= not(layer2_outputs(1589));
    outputs(4838) <= not(layer2_outputs(7750));
    outputs(4839) <= not(layer2_outputs(2405));
    outputs(4840) <= not(layer2_outputs(3399));
    outputs(4841) <= not(layer2_outputs(1133));
    outputs(4842) <= not(layer2_outputs(523));
    outputs(4843) <= not(layer2_outputs(6931));
    outputs(4844) <= (layer2_outputs(6094)) xor (layer2_outputs(493));
    outputs(4845) <= layer2_outputs(8238);
    outputs(4846) <= layer2_outputs(6215);
    outputs(4847) <= not(layer2_outputs(4792));
    outputs(4848) <= layer2_outputs(4264);
    outputs(4849) <= layer2_outputs(3897);
    outputs(4850) <= not(layer2_outputs(1581));
    outputs(4851) <= layer2_outputs(3537);
    outputs(4852) <= layer2_outputs(3014);
    outputs(4853) <= not(layer2_outputs(9313));
    outputs(4854) <= not((layer2_outputs(2796)) xor (layer2_outputs(7532)));
    outputs(4855) <= layer2_outputs(8404);
    outputs(4856) <= not(layer2_outputs(6548));
    outputs(4857) <= not((layer2_outputs(3182)) or (layer2_outputs(2710)));
    outputs(4858) <= layer2_outputs(2861);
    outputs(4859) <= not((layer2_outputs(3637)) or (layer2_outputs(7372)));
    outputs(4860) <= (layer2_outputs(783)) and not (layer2_outputs(4153));
    outputs(4861) <= not(layer2_outputs(1729));
    outputs(4862) <= not((layer2_outputs(2984)) xor (layer2_outputs(7864)));
    outputs(4863) <= (layer2_outputs(3222)) and not (layer2_outputs(8270));
    outputs(4864) <= not(layer2_outputs(9549));
    outputs(4865) <= layer2_outputs(3757);
    outputs(4866) <= layer2_outputs(4319);
    outputs(4867) <= not(layer2_outputs(1369));
    outputs(4868) <= (layer2_outputs(1742)) xor (layer2_outputs(8406));
    outputs(4869) <= layer2_outputs(5270);
    outputs(4870) <= (layer2_outputs(3017)) xor (layer2_outputs(932));
    outputs(4871) <= not((layer2_outputs(1563)) xor (layer2_outputs(2539)));
    outputs(4872) <= not(layer2_outputs(6725));
    outputs(4873) <= (layer2_outputs(353)) and not (layer2_outputs(9940));
    outputs(4874) <= layer2_outputs(1184);
    outputs(4875) <= (layer2_outputs(7917)) xor (layer2_outputs(9929));
    outputs(4876) <= layer2_outputs(3284);
    outputs(4877) <= not(layer2_outputs(3524));
    outputs(4878) <= not(layer2_outputs(2837));
    outputs(4879) <= layer2_outputs(1912);
    outputs(4880) <= layer2_outputs(4339);
    outputs(4881) <= not(layer2_outputs(2726));
    outputs(4882) <= not(layer2_outputs(1890));
    outputs(4883) <= not(layer2_outputs(6842));
    outputs(4884) <= layer2_outputs(5963);
    outputs(4885) <= (layer2_outputs(3747)) xor (layer2_outputs(8849));
    outputs(4886) <= layer2_outputs(2035);
    outputs(4887) <= not(layer2_outputs(5341));
    outputs(4888) <= layer2_outputs(2090);
    outputs(4889) <= not((layer2_outputs(3206)) or (layer2_outputs(4955)));
    outputs(4890) <= (layer2_outputs(9586)) xor (layer2_outputs(3170));
    outputs(4891) <= not(layer2_outputs(4894));
    outputs(4892) <= not(layer2_outputs(2952));
    outputs(4893) <= not((layer2_outputs(10101)) xor (layer2_outputs(1615)));
    outputs(4894) <= not(layer2_outputs(7768));
    outputs(4895) <= layer2_outputs(9174);
    outputs(4896) <= not(layer2_outputs(9722));
    outputs(4897) <= (layer2_outputs(5564)) xor (layer2_outputs(2053));
    outputs(4898) <= (layer2_outputs(4307)) and not (layer2_outputs(7844));
    outputs(4899) <= not(layer2_outputs(3199));
    outputs(4900) <= not(layer2_outputs(9587));
    outputs(4901) <= (layer2_outputs(3484)) and (layer2_outputs(9875));
    outputs(4902) <= (layer2_outputs(9247)) and (layer2_outputs(8778));
    outputs(4903) <= not(layer2_outputs(7973));
    outputs(4904) <= (layer2_outputs(929)) xor (layer2_outputs(2463));
    outputs(4905) <= not((layer2_outputs(900)) xor (layer2_outputs(9667)));
    outputs(4906) <= (layer2_outputs(5496)) and not (layer2_outputs(8032));
    outputs(4907) <= layer2_outputs(7308);
    outputs(4908) <= not(layer2_outputs(8866));
    outputs(4909) <= not(layer2_outputs(5752));
    outputs(4910) <= layer2_outputs(3273);
    outputs(4911) <= (layer2_outputs(9424)) and (layer2_outputs(8402));
    outputs(4912) <= (layer2_outputs(7941)) xor (layer2_outputs(8702));
    outputs(4913) <= not(layer2_outputs(9066));
    outputs(4914) <= layer2_outputs(4255);
    outputs(4915) <= layer2_outputs(8881);
    outputs(4916) <= not(layer2_outputs(7070));
    outputs(4917) <= not(layer2_outputs(8257));
    outputs(4918) <= layer2_outputs(3660);
    outputs(4919) <= (layer2_outputs(7079)) and not (layer2_outputs(7190));
    outputs(4920) <= layer2_outputs(7894);
    outputs(4921) <= not(layer2_outputs(9570));
    outputs(4922) <= not(layer2_outputs(9912));
    outputs(4923) <= layer2_outputs(9509);
    outputs(4924) <= not(layer2_outputs(4634));
    outputs(4925) <= not(layer2_outputs(3652));
    outputs(4926) <= not(layer2_outputs(9062));
    outputs(4927) <= layer2_outputs(2314);
    outputs(4928) <= not(layer2_outputs(2926));
    outputs(4929) <= layer2_outputs(1797);
    outputs(4930) <= not(layer2_outputs(3955));
    outputs(4931) <= (layer2_outputs(928)) xor (layer2_outputs(5295));
    outputs(4932) <= not((layer2_outputs(455)) xor (layer2_outputs(356)));
    outputs(4933) <= not(layer2_outputs(4126));
    outputs(4934) <= layer2_outputs(1667);
    outputs(4935) <= not(layer2_outputs(1715));
    outputs(4936) <= not(layer2_outputs(102)) or (layer2_outputs(3901));
    outputs(4937) <= not(layer2_outputs(3147));
    outputs(4938) <= layer2_outputs(6059);
    outputs(4939) <= layer2_outputs(7727);
    outputs(4940) <= not((layer2_outputs(9694)) and (layer2_outputs(1301)));
    outputs(4941) <= not(layer2_outputs(4145));
    outputs(4942) <= layer2_outputs(5585);
    outputs(4943) <= layer2_outputs(2638);
    outputs(4944) <= layer2_outputs(5233);
    outputs(4945) <= not(layer2_outputs(1607));
    outputs(4946) <= layer2_outputs(8059);
    outputs(4947) <= not(layer2_outputs(8930));
    outputs(4948) <= not(layer2_outputs(1055)) or (layer2_outputs(7901));
    outputs(4949) <= layer2_outputs(1218);
    outputs(4950) <= (layer2_outputs(8590)) xor (layer2_outputs(8367));
    outputs(4951) <= not((layer2_outputs(8995)) xor (layer2_outputs(8476)));
    outputs(4952) <= not(layer2_outputs(6983));
    outputs(4953) <= layer2_outputs(9971);
    outputs(4954) <= not((layer2_outputs(8244)) xor (layer2_outputs(5804)));
    outputs(4955) <= layer2_outputs(6491);
    outputs(4956) <= not(layer2_outputs(4324));
    outputs(4957) <= (layer2_outputs(2628)) and (layer2_outputs(4206));
    outputs(4958) <= (layer2_outputs(6877)) or (layer2_outputs(3790));
    outputs(4959) <= (layer2_outputs(6314)) xor (layer2_outputs(3941));
    outputs(4960) <= layer2_outputs(9721);
    outputs(4961) <= not(layer2_outputs(6925));
    outputs(4962) <= not(layer2_outputs(9420));
    outputs(4963) <= not(layer2_outputs(6336));
    outputs(4964) <= layer2_outputs(165);
    outputs(4965) <= not(layer2_outputs(3259));
    outputs(4966) <= not(layer2_outputs(782));
    outputs(4967) <= not(layer2_outputs(3027));
    outputs(4968) <= not(layer2_outputs(720));
    outputs(4969) <= layer2_outputs(8810);
    outputs(4970) <= layer2_outputs(7079);
    outputs(4971) <= layer2_outputs(2521);
    outputs(4972) <= layer2_outputs(746);
    outputs(4973) <= layer2_outputs(5301);
    outputs(4974) <= layer2_outputs(8229);
    outputs(4975) <= (layer2_outputs(6959)) xor (layer2_outputs(2));
    outputs(4976) <= not(layer2_outputs(1931)) or (layer2_outputs(23));
    outputs(4977) <= layer2_outputs(6000);
    outputs(4978) <= layer2_outputs(3242);
    outputs(4979) <= not(layer2_outputs(7716)) or (layer2_outputs(7945));
    outputs(4980) <= not(layer2_outputs(6338));
    outputs(4981) <= layer2_outputs(5951);
    outputs(4982) <= layer2_outputs(9853);
    outputs(4983) <= not(layer2_outputs(6659));
    outputs(4984) <= layer2_outputs(10214);
    outputs(4985) <= not(layer2_outputs(3011));
    outputs(4986) <= layer2_outputs(5967);
    outputs(4987) <= layer2_outputs(1720);
    outputs(4988) <= layer2_outputs(3783);
    outputs(4989) <= not(layer2_outputs(3678));
    outputs(4990) <= layer2_outputs(4331);
    outputs(4991) <= not(layer2_outputs(6362));
    outputs(4992) <= not(layer2_outputs(1787)) or (layer2_outputs(4058));
    outputs(4993) <= not(layer2_outputs(3623));
    outputs(4994) <= not(layer2_outputs(8594));
    outputs(4995) <= not((layer2_outputs(9325)) xor (layer2_outputs(3854)));
    outputs(4996) <= not(layer2_outputs(8494));
    outputs(4997) <= not(layer2_outputs(715));
    outputs(4998) <= not((layer2_outputs(5649)) or (layer2_outputs(7485)));
    outputs(4999) <= (layer2_outputs(6609)) and not (layer2_outputs(5926));
    outputs(5000) <= not(layer2_outputs(4734));
    outputs(5001) <= not((layer2_outputs(208)) xor (layer2_outputs(8498)));
    outputs(5002) <= not(layer2_outputs(9277));
    outputs(5003) <= (layer2_outputs(4728)) xor (layer2_outputs(8759));
    outputs(5004) <= layer2_outputs(2330);
    outputs(5005) <= not((layer2_outputs(2334)) xor (layer2_outputs(9951)));
    outputs(5006) <= layer2_outputs(9347);
    outputs(5007) <= not((layer2_outputs(8199)) xor (layer2_outputs(4243)));
    outputs(5008) <= not(layer2_outputs(5926));
    outputs(5009) <= not(layer2_outputs(5947)) or (layer2_outputs(9234));
    outputs(5010) <= layer2_outputs(3790);
    outputs(5011) <= not(layer2_outputs(3587));
    outputs(5012) <= not(layer2_outputs(810));
    outputs(5013) <= layer2_outputs(7894);
    outputs(5014) <= (layer2_outputs(6662)) or (layer2_outputs(364));
    outputs(5015) <= layer2_outputs(8972);
    outputs(5016) <= not(layer2_outputs(2537));
    outputs(5017) <= layer2_outputs(3766);
    outputs(5018) <= (layer2_outputs(9436)) xor (layer2_outputs(198));
    outputs(5019) <= layer2_outputs(10033);
    outputs(5020) <= layer2_outputs(9612);
    outputs(5021) <= not((layer2_outputs(8658)) or (layer2_outputs(4308)));
    outputs(5022) <= (layer2_outputs(5615)) xor (layer2_outputs(100));
    outputs(5023) <= not(layer2_outputs(3325));
    outputs(5024) <= layer2_outputs(6648);
    outputs(5025) <= layer2_outputs(8223);
    outputs(5026) <= layer2_outputs(4474);
    outputs(5027) <= not((layer2_outputs(2949)) xor (layer2_outputs(8767)));
    outputs(5028) <= not(layer2_outputs(7434));
    outputs(5029) <= not(layer2_outputs(660));
    outputs(5030) <= not(layer2_outputs(1922));
    outputs(5031) <= (layer2_outputs(8744)) or (layer2_outputs(8354));
    outputs(5032) <= layer2_outputs(918);
    outputs(5033) <= not(layer2_outputs(4144));
    outputs(5034) <= not(layer2_outputs(5050));
    outputs(5035) <= (layer2_outputs(6239)) and (layer2_outputs(7871));
    outputs(5036) <= (layer2_outputs(6879)) or (layer2_outputs(3461));
    outputs(5037) <= layer2_outputs(6375);
    outputs(5038) <= not((layer2_outputs(5876)) xor (layer2_outputs(4254)));
    outputs(5039) <= not(layer2_outputs(1401));
    outputs(5040) <= not(layer2_outputs(4839));
    outputs(5041) <= (layer2_outputs(8306)) and not (layer2_outputs(9337));
    outputs(5042) <= layer2_outputs(879);
    outputs(5043) <= not((layer2_outputs(3990)) xor (layer2_outputs(2727)));
    outputs(5044) <= layer2_outputs(6290);
    outputs(5045) <= layer2_outputs(9718);
    outputs(5046) <= not((layer2_outputs(8227)) xor (layer2_outputs(7665)));
    outputs(5047) <= not((layer2_outputs(3259)) or (layer2_outputs(5607)));
    outputs(5048) <= layer2_outputs(1168);
    outputs(5049) <= (layer2_outputs(8766)) and (layer2_outputs(8068));
    outputs(5050) <= layer2_outputs(367);
    outputs(5051) <= not(layer2_outputs(5620));
    outputs(5052) <= layer2_outputs(662);
    outputs(5053) <= layer2_outputs(7147);
    outputs(5054) <= not(layer2_outputs(4911));
    outputs(5055) <= not(layer2_outputs(9478));
    outputs(5056) <= not(layer2_outputs(8610));
    outputs(5057) <= not(layer2_outputs(8842));
    outputs(5058) <= layer2_outputs(5036);
    outputs(5059) <= not(layer2_outputs(2894));
    outputs(5060) <= not(layer2_outputs(4041));
    outputs(5061) <= not(layer2_outputs(1960)) or (layer2_outputs(6542));
    outputs(5062) <= layer2_outputs(7298);
    outputs(5063) <= not((layer2_outputs(7832)) xor (layer2_outputs(3620)));
    outputs(5064) <= not((layer2_outputs(4306)) and (layer2_outputs(1237)));
    outputs(5065) <= not(layer2_outputs(4598));
    outputs(5066) <= layer2_outputs(8563);
    outputs(5067) <= layer2_outputs(2162);
    outputs(5068) <= (layer2_outputs(9279)) and not (layer2_outputs(5126));
    outputs(5069) <= (layer2_outputs(893)) xor (layer2_outputs(4931));
    outputs(5070) <= layer2_outputs(5184);
    outputs(5071) <= not(layer2_outputs(8250));
    outputs(5072) <= not(layer2_outputs(5449));
    outputs(5073) <= not(layer2_outputs(7601));
    outputs(5074) <= layer2_outputs(2773);
    outputs(5075) <= layer2_outputs(1158);
    outputs(5076) <= layer2_outputs(3902);
    outputs(5077) <= not(layer2_outputs(6154));
    outputs(5078) <= layer2_outputs(2319);
    outputs(5079) <= (layer2_outputs(6985)) or (layer2_outputs(1565));
    outputs(5080) <= (layer2_outputs(3093)) and not (layer2_outputs(7905));
    outputs(5081) <= not(layer2_outputs(5141));
    outputs(5082) <= layer2_outputs(5066);
    outputs(5083) <= not((layer2_outputs(5453)) xor (layer2_outputs(453)));
    outputs(5084) <= (layer2_outputs(9412)) and (layer2_outputs(10163));
    outputs(5085) <= (layer2_outputs(7315)) and not (layer2_outputs(4197));
    outputs(5086) <= not((layer2_outputs(10182)) or (layer2_outputs(388)));
    outputs(5087) <= not(layer2_outputs(2312));
    outputs(5088) <= not(layer2_outputs(2013));
    outputs(5089) <= not(layer2_outputs(7149));
    outputs(5090) <= not((layer2_outputs(6666)) xor (layer2_outputs(7994)));
    outputs(5091) <= (layer2_outputs(2519)) xor (layer2_outputs(7804));
    outputs(5092) <= (layer2_outputs(5043)) xor (layer2_outputs(8886));
    outputs(5093) <= layer2_outputs(4764);
    outputs(5094) <= layer2_outputs(5720);
    outputs(5095) <= layer2_outputs(7885);
    outputs(5096) <= not(layer2_outputs(8367));
    outputs(5097) <= layer2_outputs(10029);
    outputs(5098) <= not(layer2_outputs(721));
    outputs(5099) <= not(layer2_outputs(2659));
    outputs(5100) <= (layer2_outputs(7453)) xor (layer2_outputs(2534));
    outputs(5101) <= not(layer2_outputs(3019));
    outputs(5102) <= (layer2_outputs(1217)) xor (layer2_outputs(7848));
    outputs(5103) <= (layer2_outputs(928)) and not (layer2_outputs(8764));
    outputs(5104) <= not(layer2_outputs(4642));
    outputs(5105) <= (layer2_outputs(4756)) and not (layer2_outputs(2905));
    outputs(5106) <= not((layer2_outputs(1588)) xor (layer2_outputs(8899)));
    outputs(5107) <= not(layer2_outputs(7191));
    outputs(5108) <= not((layer2_outputs(192)) xor (layer2_outputs(7637)));
    outputs(5109) <= (layer2_outputs(6679)) or (layer2_outputs(6748));
    outputs(5110) <= layer2_outputs(1296);
    outputs(5111) <= not(layer2_outputs(482));
    outputs(5112) <= (layer2_outputs(1252)) xor (layer2_outputs(182));
    outputs(5113) <= not(layer2_outputs(34));
    outputs(5114) <= not(layer2_outputs(4352));
    outputs(5115) <= layer2_outputs(5759);
    outputs(5116) <= not(layer2_outputs(4112));
    outputs(5117) <= not((layer2_outputs(9517)) or (layer2_outputs(6419)));
    outputs(5118) <= (layer2_outputs(9607)) xor (layer2_outputs(3763));
    outputs(5119) <= not(layer2_outputs(2557));
    outputs(5120) <= not(layer2_outputs(2337));
    outputs(5121) <= layer2_outputs(3737);
    outputs(5122) <= not(layer2_outputs(2971));
    outputs(5123) <= (layer2_outputs(9934)) and (layer2_outputs(811));
    outputs(5124) <= not(layer2_outputs(5317));
    outputs(5125) <= not(layer2_outputs(5610));
    outputs(5126) <= not(layer2_outputs(1492));
    outputs(5127) <= not(layer2_outputs(4348));
    outputs(5128) <= not((layer2_outputs(824)) xor (layer2_outputs(4040)));
    outputs(5129) <= layer2_outputs(7662);
    outputs(5130) <= not(layer2_outputs(4861));
    outputs(5131) <= not(layer2_outputs(7192));
    outputs(5132) <= not(layer2_outputs(1227));
    outputs(5133) <= not((layer2_outputs(2633)) xor (layer2_outputs(8548)));
    outputs(5134) <= layer2_outputs(7232);
    outputs(5135) <= (layer2_outputs(6023)) xor (layer2_outputs(4469));
    outputs(5136) <= layer2_outputs(8368);
    outputs(5137) <= (layer2_outputs(1543)) xor (layer2_outputs(6068));
    outputs(5138) <= (layer2_outputs(4144)) xor (layer2_outputs(188));
    outputs(5139) <= not(layer2_outputs(5287));
    outputs(5140) <= layer2_outputs(6066);
    outputs(5141) <= (layer2_outputs(238)) or (layer2_outputs(8218));
    outputs(5142) <= (layer2_outputs(2290)) or (layer2_outputs(8241));
    outputs(5143) <= layer2_outputs(9248);
    outputs(5144) <= (layer2_outputs(3468)) and not (layer2_outputs(2939));
    outputs(5145) <= (layer2_outputs(5650)) xor (layer2_outputs(8509));
    outputs(5146) <= layer2_outputs(9403);
    outputs(5147) <= not(layer2_outputs(9806));
    outputs(5148) <= (layer2_outputs(8417)) and (layer2_outputs(8572));
    outputs(5149) <= layer2_outputs(4728);
    outputs(5150) <= layer2_outputs(7061);
    outputs(5151) <= not(layer2_outputs(1491));
    outputs(5152) <= not((layer2_outputs(2036)) xor (layer2_outputs(2935)));
    outputs(5153) <= not((layer2_outputs(10122)) xor (layer2_outputs(416)));
    outputs(5154) <= not(layer2_outputs(2282));
    outputs(5155) <= layer2_outputs(9740);
    outputs(5156) <= (layer2_outputs(10154)) or (layer2_outputs(3118));
    outputs(5157) <= not((layer2_outputs(9869)) and (layer2_outputs(9159)));
    outputs(5158) <= not((layer2_outputs(373)) and (layer2_outputs(7390)));
    outputs(5159) <= layer2_outputs(8997);
    outputs(5160) <= layer2_outputs(9696);
    outputs(5161) <= not((layer2_outputs(2283)) xor (layer2_outputs(2339)));
    outputs(5162) <= not(layer2_outputs(7132));
    outputs(5163) <= layer2_outputs(7368);
    outputs(5164) <= not(layer2_outputs(2575));
    outputs(5165) <= not(layer2_outputs(2576));
    outputs(5166) <= (layer2_outputs(953)) and not (layer2_outputs(3829));
    outputs(5167) <= layer2_outputs(9629);
    outputs(5168) <= not((layer2_outputs(9865)) xor (layer2_outputs(5678)));
    outputs(5169) <= layer2_outputs(7678);
    outputs(5170) <= not((layer2_outputs(2365)) or (layer2_outputs(1828)));
    outputs(5171) <= not(layer2_outputs(2979));
    outputs(5172) <= layer2_outputs(8670);
    outputs(5173) <= not((layer2_outputs(1284)) or (layer2_outputs(4844)));
    outputs(5174) <= not(layer2_outputs(8668));
    outputs(5175) <= (layer2_outputs(6434)) and (layer2_outputs(9646));
    outputs(5176) <= (layer2_outputs(8376)) xor (layer2_outputs(2787));
    outputs(5177) <= not(layer2_outputs(71));
    outputs(5178) <= not(layer2_outputs(2462));
    outputs(5179) <= not(layer2_outputs(2285));
    outputs(5180) <= layer2_outputs(9843);
    outputs(5181) <= layer2_outputs(8944);
    outputs(5182) <= not((layer2_outputs(4859)) xor (layer2_outputs(3239)));
    outputs(5183) <= not((layer2_outputs(5627)) xor (layer2_outputs(8602)));
    outputs(5184) <= layer2_outputs(3937);
    outputs(5185) <= not((layer2_outputs(2761)) xor (layer2_outputs(3243)));
    outputs(5186) <= (layer2_outputs(4190)) and (layer2_outputs(9819));
    outputs(5187) <= not(layer2_outputs(9588)) or (layer2_outputs(1313));
    outputs(5188) <= layer2_outputs(9383);
    outputs(5189) <= (layer2_outputs(10145)) xor (layer2_outputs(9755));
    outputs(5190) <= (layer2_outputs(8739)) xor (layer2_outputs(2256));
    outputs(5191) <= (layer2_outputs(8064)) xor (layer2_outputs(4361));
    outputs(5192) <= not((layer2_outputs(4292)) and (layer2_outputs(821)));
    outputs(5193) <= layer2_outputs(8);
    outputs(5194) <= (layer2_outputs(3868)) or (layer2_outputs(6545));
    outputs(5195) <= not(layer2_outputs(4277));
    outputs(5196) <= not(layer2_outputs(4628));
    outputs(5197) <= not(layer2_outputs(8843));
    outputs(5198) <= layer2_outputs(3633);
    outputs(5199) <= (layer2_outputs(475)) or (layer2_outputs(7393));
    outputs(5200) <= not(layer2_outputs(7987));
    outputs(5201) <= (layer2_outputs(7625)) and (layer2_outputs(7224));
    outputs(5202) <= layer2_outputs(10202);
    outputs(5203) <= not(layer2_outputs(1482));
    outputs(5204) <= (layer2_outputs(7759)) and not (layer2_outputs(9290));
    outputs(5205) <= not((layer2_outputs(6941)) xor (layer2_outputs(3434)));
    outputs(5206) <= not((layer2_outputs(4093)) or (layer2_outputs(229)));
    outputs(5207) <= not(layer2_outputs(3264));
    outputs(5208) <= layer2_outputs(822);
    outputs(5209) <= layer2_outputs(2980);
    outputs(5210) <= (layer2_outputs(992)) xor (layer2_outputs(6778));
    outputs(5211) <= (layer2_outputs(5562)) and not (layer2_outputs(8836));
    outputs(5212) <= not(layer2_outputs(4258));
    outputs(5213) <= not(layer2_outputs(6171));
    outputs(5214) <= (layer2_outputs(10097)) and not (layer2_outputs(6719));
    outputs(5215) <= not(layer2_outputs(3026));
    outputs(5216) <= layer2_outputs(1083);
    outputs(5217) <= (layer2_outputs(5220)) xor (layer2_outputs(9171));
    outputs(5218) <= not((layer2_outputs(8371)) xor (layer2_outputs(1846)));
    outputs(5219) <= not(layer2_outputs(5726));
    outputs(5220) <= not(layer2_outputs(7577));
    outputs(5221) <= layer2_outputs(177);
    outputs(5222) <= layer2_outputs(2364);
    outputs(5223) <= (layer2_outputs(4116)) and (layer2_outputs(1817));
    outputs(5224) <= not(layer2_outputs(8976));
    outputs(5225) <= layer2_outputs(7680);
    outputs(5226) <= layer2_outputs(4725);
    outputs(5227) <= not(layer2_outputs(331));
    outputs(5228) <= layer2_outputs(1173);
    outputs(5229) <= layer2_outputs(8523);
    outputs(5230) <= layer2_outputs(10093);
    outputs(5231) <= layer2_outputs(9687);
    outputs(5232) <= not(layer2_outputs(8026));
    outputs(5233) <= layer2_outputs(608);
    outputs(5234) <= not(layer2_outputs(8507));
    outputs(5235) <= not((layer2_outputs(5383)) or (layer2_outputs(3460)));
    outputs(5236) <= not(layer2_outputs(1129));
    outputs(5237) <= layer2_outputs(6533);
    outputs(5238) <= not((layer2_outputs(8373)) xor (layer2_outputs(4286)));
    outputs(5239) <= not(layer2_outputs(3655));
    outputs(5240) <= not((layer2_outputs(3043)) xor (layer2_outputs(6206)));
    outputs(5241) <= (layer2_outputs(3804)) xor (layer2_outputs(3173));
    outputs(5242) <= not(layer2_outputs(4068));
    outputs(5243) <= layer2_outputs(7189);
    outputs(5244) <= (layer2_outputs(6318)) or (layer2_outputs(1838));
    outputs(5245) <= (layer2_outputs(3663)) xor (layer2_outputs(1762));
    outputs(5246) <= (layer2_outputs(6756)) xor (layer2_outputs(8501));
    outputs(5247) <= not((layer2_outputs(3966)) xor (layer2_outputs(7457)));
    outputs(5248) <= not(layer2_outputs(7555));
    outputs(5249) <= (layer2_outputs(5705)) xor (layer2_outputs(2626));
    outputs(5250) <= not(layer2_outputs(2932));
    outputs(5251) <= (layer2_outputs(1708)) xor (layer2_outputs(688));
    outputs(5252) <= not(layer2_outputs(1260));
    outputs(5253) <= layer2_outputs(4076);
    outputs(5254) <= not(layer2_outputs(6836));
    outputs(5255) <= not((layer2_outputs(5647)) xor (layer2_outputs(3165)));
    outputs(5256) <= not(layer2_outputs(2985));
    outputs(5257) <= not(layer2_outputs(1295));
    outputs(5258) <= not(layer2_outputs(118));
    outputs(5259) <= layer2_outputs(7175);
    outputs(5260) <= (layer2_outputs(4287)) xor (layer2_outputs(7168));
    outputs(5261) <= not(layer2_outputs(2591)) or (layer2_outputs(673));
    outputs(5262) <= (layer2_outputs(9543)) or (layer2_outputs(3002));
    outputs(5263) <= not((layer2_outputs(2692)) xor (layer2_outputs(2741)));
    outputs(5264) <= layer2_outputs(6708);
    outputs(5265) <= layer2_outputs(8538);
    outputs(5266) <= layer2_outputs(6861);
    outputs(5267) <= (layer2_outputs(1564)) xor (layer2_outputs(1127));
    outputs(5268) <= (layer2_outputs(3294)) or (layer2_outputs(8267));
    outputs(5269) <= not(layer2_outputs(2506));
    outputs(5270) <= layer2_outputs(1639);
    outputs(5271) <= layer2_outputs(1523);
    outputs(5272) <= not((layer2_outputs(4940)) xor (layer2_outputs(1358)));
    outputs(5273) <= not(layer2_outputs(7515));
    outputs(5274) <= (layer2_outputs(2458)) and not (layer2_outputs(4563));
    outputs(5275) <= layer2_outputs(4801);
    outputs(5276) <= layer2_outputs(5853);
    outputs(5277) <= layer2_outputs(3541);
    outputs(5278) <= layer2_outputs(838);
    outputs(5279) <= (layer2_outputs(3414)) and not (layer2_outputs(320));
    outputs(5280) <= not((layer2_outputs(8988)) xor (layer2_outputs(7714)));
    outputs(5281) <= (layer2_outputs(3025)) or (layer2_outputs(3156));
    outputs(5282) <= not((layer2_outputs(3394)) xor (layer2_outputs(3100)));
    outputs(5283) <= not((layer2_outputs(4740)) xor (layer2_outputs(2595)));
    outputs(5284) <= not(layer2_outputs(4852));
    outputs(5285) <= layer2_outputs(2113);
    outputs(5286) <= (layer2_outputs(6759)) or (layer2_outputs(6453));
    outputs(5287) <= not(layer2_outputs(2840));
    outputs(5288) <= not((layer2_outputs(6401)) xor (layer2_outputs(8512)));
    outputs(5289) <= layer2_outputs(6348);
    outputs(5290) <= not(layer2_outputs(5179));
    outputs(5291) <= not(layer2_outputs(5346));
    outputs(5292) <= layer2_outputs(6770);
    outputs(5293) <= (layer2_outputs(3777)) xor (layer2_outputs(7807));
    outputs(5294) <= not((layer2_outputs(1396)) xor (layer2_outputs(6570)));
    outputs(5295) <= not(layer2_outputs(8383)) or (layer2_outputs(9461));
    outputs(5296) <= (layer2_outputs(2870)) xor (layer2_outputs(9802));
    outputs(5297) <= not(layer2_outputs(3093));
    outputs(5298) <= layer2_outputs(10176);
    outputs(5299) <= not((layer2_outputs(1304)) and (layer2_outputs(1812)));
    outputs(5300) <= not(layer2_outputs(3221));
    outputs(5301) <= layer2_outputs(3316);
    outputs(5302) <= (layer2_outputs(10184)) and not (layer2_outputs(3035));
    outputs(5303) <= not((layer2_outputs(5685)) xor (layer2_outputs(9906)));
    outputs(5304) <= (layer2_outputs(3013)) or (layer2_outputs(790));
    outputs(5305) <= not((layer2_outputs(3504)) xor (layer2_outputs(4530)));
    outputs(5306) <= (layer2_outputs(8326)) and not (layer2_outputs(3751));
    outputs(5307) <= (layer2_outputs(5939)) xor (layer2_outputs(2622));
    outputs(5308) <= not((layer2_outputs(8171)) xor (layer2_outputs(6106)));
    outputs(5309) <= (layer2_outputs(2362)) and (layer2_outputs(3168));
    outputs(5310) <= not(layer2_outputs(4371));
    outputs(5311) <= layer2_outputs(7524);
    outputs(5312) <= layer2_outputs(10113);
    outputs(5313) <= not(layer2_outputs(4222));
    outputs(5314) <= (layer2_outputs(2417)) xor (layer2_outputs(5591));
    outputs(5315) <= not((layer2_outputs(5524)) and (layer2_outputs(5975)));
    outputs(5316) <= not(layer2_outputs(2609));
    outputs(5317) <= (layer2_outputs(5224)) xor (layer2_outputs(4749));
    outputs(5318) <= not((layer2_outputs(1628)) xor (layer2_outputs(5610)));
    outputs(5319) <= (layer2_outputs(7690)) xor (layer2_outputs(2071));
    outputs(5320) <= not(layer2_outputs(5765));
    outputs(5321) <= not(layer2_outputs(3221));
    outputs(5322) <= layer2_outputs(9388);
    outputs(5323) <= layer2_outputs(7936);
    outputs(5324) <= not((layer2_outputs(1897)) xor (layer2_outputs(1139)));
    outputs(5325) <= not((layer2_outputs(9820)) xor (layer2_outputs(3114)));
    outputs(5326) <= layer2_outputs(9391);
    outputs(5327) <= not(layer2_outputs(1466));
    outputs(5328) <= layer2_outputs(2494);
    outputs(5329) <= (layer2_outputs(9926)) xor (layer2_outputs(6359));
    outputs(5330) <= layer2_outputs(2264);
    outputs(5331) <= not(layer2_outputs(10144)) or (layer2_outputs(8282));
    outputs(5332) <= not(layer2_outputs(180));
    outputs(5333) <= not(layer2_outputs(2533));
    outputs(5334) <= layer2_outputs(8160);
    outputs(5335) <= not(layer2_outputs(10214));
    outputs(5336) <= (layer2_outputs(7102)) and not (layer2_outputs(8537));
    outputs(5337) <= layer2_outputs(3262);
    outputs(5338) <= not(layer2_outputs(4948)) or (layer2_outputs(5354));
    outputs(5339) <= not(layer2_outputs(6006));
    outputs(5340) <= not(layer2_outputs(46));
    outputs(5341) <= (layer2_outputs(7316)) xor (layer2_outputs(8737));
    outputs(5342) <= not(layer2_outputs(2559));
    outputs(5343) <= not((layer2_outputs(7726)) xor (layer2_outputs(4605)));
    outputs(5344) <= layer2_outputs(5516);
    outputs(5345) <= (layer2_outputs(999)) xor (layer2_outputs(7858));
    outputs(5346) <= layer2_outputs(7898);
    outputs(5347) <= not(layer2_outputs(9267)) or (layer2_outputs(2794));
    outputs(5348) <= layer2_outputs(1362);
    outputs(5349) <= not(layer2_outputs(9147));
    outputs(5350) <= not(layer2_outputs(1085));
    outputs(5351) <= not(layer2_outputs(593));
    outputs(5352) <= not(layer2_outputs(8185));
    outputs(5353) <= (layer2_outputs(281)) xor (layer2_outputs(8001));
    outputs(5354) <= not(layer2_outputs(6442));
    outputs(5355) <= layer2_outputs(4056);
    outputs(5356) <= not((layer2_outputs(6463)) xor (layer2_outputs(346)));
    outputs(5357) <= not(layer2_outputs(5030));
    outputs(5358) <= not(layer2_outputs(9005));
    outputs(5359) <= not((layer2_outputs(3252)) xor (layer2_outputs(3109)));
    outputs(5360) <= not(layer2_outputs(4783));
    outputs(5361) <= not(layer2_outputs(4607));
    outputs(5362) <= (layer2_outputs(3181)) xor (layer2_outputs(3969));
    outputs(5363) <= not((layer2_outputs(6979)) xor (layer2_outputs(6264)));
    outputs(5364) <= not(layer2_outputs(4472));
    outputs(5365) <= layer2_outputs(7904);
    outputs(5366) <= not((layer2_outputs(2371)) xor (layer2_outputs(3685)));
    outputs(5367) <= layer2_outputs(9534);
    outputs(5368) <= (layer2_outputs(7614)) xor (layer2_outputs(7670));
    outputs(5369) <= layer2_outputs(1696);
    outputs(5370) <= not((layer2_outputs(5677)) xor (layer2_outputs(3506)));
    outputs(5371) <= not((layer2_outputs(9038)) xor (layer2_outputs(2703)));
    outputs(5372) <= layer2_outputs(1059);
    outputs(5373) <= not(layer2_outputs(4904));
    outputs(5374) <= layer2_outputs(6245);
    outputs(5375) <= not((layer2_outputs(554)) xor (layer2_outputs(2200)));
    outputs(5376) <= not(layer2_outputs(2820));
    outputs(5377) <= not(layer2_outputs(1749)) or (layer2_outputs(4780));
    outputs(5378) <= (layer2_outputs(909)) xor (layer2_outputs(4989));
    outputs(5379) <= layer2_outputs(985);
    outputs(5380) <= layer2_outputs(9097);
    outputs(5381) <= not((layer2_outputs(8586)) xor (layer2_outputs(595)));
    outputs(5382) <= (layer2_outputs(745)) and (layer2_outputs(2165));
    outputs(5383) <= not(layer2_outputs(2722));
    outputs(5384) <= not(layer2_outputs(8088));
    outputs(5385) <= not(layer2_outputs(1667));
    outputs(5386) <= layer2_outputs(3291);
    outputs(5387) <= not(layer2_outputs(1126));
    outputs(5388) <= layer2_outputs(3278);
    outputs(5389) <= not(layer2_outputs(6882));
    outputs(5390) <= layer2_outputs(9825);
    outputs(5391) <= (layer2_outputs(8800)) and not (layer2_outputs(7493));
    outputs(5392) <= not((layer2_outputs(1444)) xor (layer2_outputs(62)));
    outputs(5393) <= not(layer2_outputs(3340));
    outputs(5394) <= not(layer2_outputs(9412));
    outputs(5395) <= layer2_outputs(4500);
    outputs(5396) <= not((layer2_outputs(6351)) xor (layer2_outputs(130)));
    outputs(5397) <= not(layer2_outputs(5644));
    outputs(5398) <= not(layer2_outputs(4032));
    outputs(5399) <= layer2_outputs(5670);
    outputs(5400) <= not(layer2_outputs(3711));
    outputs(5401) <= not((layer2_outputs(3354)) xor (layer2_outputs(5842)));
    outputs(5402) <= not((layer2_outputs(8196)) xor (layer2_outputs(3496)));
    outputs(5403) <= not((layer2_outputs(734)) xor (layer2_outputs(7613)));
    outputs(5404) <= layer2_outputs(2192);
    outputs(5405) <= not(layer2_outputs(7909));
    outputs(5406) <= not(layer2_outputs(4201));
    outputs(5407) <= not(layer2_outputs(9398));
    outputs(5408) <= layer2_outputs(960);
    outputs(5409) <= not(layer2_outputs(2946));
    outputs(5410) <= not(layer2_outputs(6970)) or (layer2_outputs(9068));
    outputs(5411) <= (layer2_outputs(271)) and not (layer2_outputs(3311));
    outputs(5412) <= not((layer2_outputs(261)) xor (layer2_outputs(1098)));
    outputs(5413) <= not((layer2_outputs(5822)) xor (layer2_outputs(4761)));
    outputs(5414) <= not(layer2_outputs(4212));
    outputs(5415) <= not(layer2_outputs(789));
    outputs(5416) <= not((layer2_outputs(9275)) xor (layer2_outputs(4452)));
    outputs(5417) <= not((layer2_outputs(2817)) and (layer2_outputs(5254)));
    outputs(5418) <= not((layer2_outputs(3719)) xor (layer2_outputs(10013)));
    outputs(5419) <= not(layer2_outputs(1616));
    outputs(5420) <= not((layer2_outputs(4447)) xor (layer2_outputs(3158)));
    outputs(5421) <= layer2_outputs(2715);
    outputs(5422) <= not(layer2_outputs(159)) or (layer2_outputs(1567));
    outputs(5423) <= not(layer2_outputs(2732));
    outputs(5424) <= (layer2_outputs(1718)) or (layer2_outputs(4832));
    outputs(5425) <= (layer2_outputs(9787)) xor (layer2_outputs(1244));
    outputs(5426) <= not((layer2_outputs(383)) xor (layer2_outputs(7047)));
    outputs(5427) <= layer2_outputs(271);
    outputs(5428) <= not(layer2_outputs(9518)) or (layer2_outputs(1125));
    outputs(5429) <= (layer2_outputs(7791)) and (layer2_outputs(2792));
    outputs(5430) <= layer2_outputs(3423);
    outputs(5431) <= not(layer2_outputs(5808));
    outputs(5432) <= (layer2_outputs(5065)) xor (layer2_outputs(4961));
    outputs(5433) <= not(layer2_outputs(9067));
    outputs(5434) <= not((layer2_outputs(7007)) and (layer2_outputs(2034)));
    outputs(5435) <= (layer2_outputs(663)) and (layer2_outputs(8770));
    outputs(5436) <= (layer2_outputs(5245)) and not (layer2_outputs(4036));
    outputs(5437) <= not((layer2_outputs(423)) and (layer2_outputs(5119)));
    outputs(5438) <= not((layer2_outputs(3037)) xor (layer2_outputs(8807)));
    outputs(5439) <= not(layer2_outputs(866));
    outputs(5440) <= layer2_outputs(6377);
    outputs(5441) <= layer2_outputs(5624);
    outputs(5442) <= (layer2_outputs(8108)) and (layer2_outputs(502));
    outputs(5443) <= not(layer2_outputs(1835));
    outputs(5444) <= not(layer2_outputs(5028)) or (layer2_outputs(5745));
    outputs(5445) <= layer2_outputs(426);
    outputs(5446) <= (layer2_outputs(8982)) xor (layer2_outputs(2273));
    outputs(5447) <= layer2_outputs(2288);
    outputs(5448) <= (layer2_outputs(6826)) or (layer2_outputs(7259));
    outputs(5449) <= not(layer2_outputs(4631));
    outputs(5450) <= layer2_outputs(6265);
    outputs(5451) <= (layer2_outputs(3717)) or (layer2_outputs(1930));
    outputs(5452) <= not(layer2_outputs(8455));
    outputs(5453) <= layer2_outputs(3497);
    outputs(5454) <= not(layer2_outputs(4659));
    outputs(5455) <= not((layer2_outputs(9282)) xor (layer2_outputs(2352)));
    outputs(5456) <= layer2_outputs(7356);
    outputs(5457) <= not((layer2_outputs(1094)) xor (layer2_outputs(646)));
    outputs(5458) <= layer2_outputs(7016);
    outputs(5459) <= (layer2_outputs(1212)) xor (layer2_outputs(5123));
    outputs(5460) <= layer2_outputs(4796);
    outputs(5461) <= layer2_outputs(4041);
    outputs(5462) <= not(layer2_outputs(1086));
    outputs(5463) <= not(layer2_outputs(7544));
    outputs(5464) <= not((layer2_outputs(3130)) and (layer2_outputs(9732)));
    outputs(5465) <= layer2_outputs(5522);
    outputs(5466) <= not(layer2_outputs(6752));
    outputs(5467) <= (layer2_outputs(5066)) xor (layer2_outputs(1673));
    outputs(5468) <= not((layer2_outputs(5576)) xor (layer2_outputs(1288)));
    outputs(5469) <= not(layer2_outputs(5029));
    outputs(5470) <= layer2_outputs(2418);
    outputs(5471) <= (layer2_outputs(3313)) xor (layer2_outputs(1855));
    outputs(5472) <= (layer2_outputs(4017)) xor (layer2_outputs(9782));
    outputs(5473) <= not(layer2_outputs(10209));
    outputs(5474) <= (layer2_outputs(4362)) xor (layer2_outputs(3434));
    outputs(5475) <= not(layer2_outputs(2768));
    outputs(5476) <= layer2_outputs(8216);
    outputs(5477) <= not(layer2_outputs(4926));
    outputs(5478) <= not((layer2_outputs(3177)) xor (layer2_outputs(7406)));
    outputs(5479) <= not(layer2_outputs(5302));
    outputs(5480) <= (layer2_outputs(5387)) xor (layer2_outputs(742));
    outputs(5481) <= layer2_outputs(2416);
    outputs(5482) <= (layer2_outputs(4535)) and not (layer2_outputs(6565));
    outputs(5483) <= not(layer2_outputs(5143));
    outputs(5484) <= layer2_outputs(3377);
    outputs(5485) <= (layer2_outputs(2392)) and not (layer2_outputs(7011));
    outputs(5486) <= layer2_outputs(6394);
    outputs(5487) <= layer2_outputs(9334);
    outputs(5488) <= not((layer2_outputs(8338)) xor (layer2_outputs(4826)));
    outputs(5489) <= layer2_outputs(6085);
    outputs(5490) <= layer2_outputs(3212);
    outputs(5491) <= layer2_outputs(344);
    outputs(5492) <= not((layer2_outputs(1386)) and (layer2_outputs(8664)));
    outputs(5493) <= not(layer2_outputs(6383));
    outputs(5494) <= not((layer2_outputs(3106)) or (layer2_outputs(6566)));
    outputs(5495) <= (layer2_outputs(1205)) or (layer2_outputs(2491));
    outputs(5496) <= not((layer2_outputs(7216)) or (layer2_outputs(894)));
    outputs(5497) <= layer2_outputs(10229);
    outputs(5498) <= layer2_outputs(7547);
    outputs(5499) <= (layer2_outputs(3643)) xor (layer2_outputs(3506));
    outputs(5500) <= (layer2_outputs(4257)) xor (layer2_outputs(3895));
    outputs(5501) <= not(layer2_outputs(3185)) or (layer2_outputs(2644));
    outputs(5502) <= layer2_outputs(6773);
    outputs(5503) <= not((layer2_outputs(7681)) xor (layer2_outputs(681)));
    outputs(5504) <= not((layer2_outputs(10)) or (layer2_outputs(145)));
    outputs(5505) <= not(layer2_outputs(126)) or (layer2_outputs(5948));
    outputs(5506) <= not(layer2_outputs(9807));
    outputs(5507) <= layer2_outputs(7176);
    outputs(5508) <= (layer2_outputs(6433)) xor (layer2_outputs(1300));
    outputs(5509) <= not(layer2_outputs(7053));
    outputs(5510) <= not(layer2_outputs(4562));
    outputs(5511) <= (layer2_outputs(10191)) xor (layer2_outputs(7096));
    outputs(5512) <= not(layer2_outputs(7350));
    outputs(5513) <= layer2_outputs(8034);
    outputs(5514) <= (layer2_outputs(2338)) xor (layer2_outputs(7036));
    outputs(5515) <= not((layer2_outputs(296)) xor (layer2_outputs(5434)));
    outputs(5516) <= not(layer2_outputs(1715));
    outputs(5517) <= layer2_outputs(3418);
    outputs(5518) <= not((layer2_outputs(4001)) xor (layer2_outputs(9700)));
    outputs(5519) <= not((layer2_outputs(7702)) xor (layer2_outputs(2753)));
    outputs(5520) <= layer2_outputs(7986);
    outputs(5521) <= not((layer2_outputs(7646)) xor (layer2_outputs(8520)));
    outputs(5522) <= not(layer2_outputs(7443));
    outputs(5523) <= layer2_outputs(1062);
    outputs(5524) <= layer2_outputs(7847);
    outputs(5525) <= not(layer2_outputs(8637));
    outputs(5526) <= not((layer2_outputs(634)) xor (layer2_outputs(9965)));
    outputs(5527) <= layer2_outputs(1180);
    outputs(5528) <= not(layer2_outputs(3892)) or (layer2_outputs(5413));
    outputs(5529) <= layer2_outputs(5039);
    outputs(5530) <= not(layer2_outputs(9102));
    outputs(5531) <= layer2_outputs(8957);
    outputs(5532) <= layer2_outputs(2343);
    outputs(5533) <= layer2_outputs(9362);
    outputs(5534) <= layer2_outputs(4025);
    outputs(5535) <= layer2_outputs(7302);
    outputs(5536) <= layer2_outputs(4923);
    outputs(5537) <= (layer2_outputs(4460)) and (layer2_outputs(6485));
    outputs(5538) <= not((layer2_outputs(5090)) xor (layer2_outputs(7535)));
    outputs(5539) <= (layer2_outputs(691)) or (layer2_outputs(9381));
    outputs(5540) <= not(layer2_outputs(7149));
    outputs(5541) <= layer2_outputs(1120);
    outputs(5542) <= (layer2_outputs(9615)) and not (layer2_outputs(8167));
    outputs(5543) <= (layer2_outputs(4719)) xor (layer2_outputs(92));
    outputs(5544) <= layer2_outputs(3580);
    outputs(5545) <= (layer2_outputs(3486)) xor (layer2_outputs(6055));
    outputs(5546) <= not((layer2_outputs(8728)) xor (layer2_outputs(9283)));
    outputs(5547) <= layer2_outputs(1583);
    outputs(5548) <= layer2_outputs(9458);
    outputs(5549) <= not(layer2_outputs(2654)) or (layer2_outputs(1315));
    outputs(5550) <= layer2_outputs(1613);
    outputs(5551) <= (layer2_outputs(386)) and not (layer2_outputs(1369));
    outputs(5552) <= (layer2_outputs(5145)) xor (layer2_outputs(2955));
    outputs(5553) <= layer2_outputs(5748);
    outputs(5554) <= layer2_outputs(886);
    outputs(5555) <= (layer2_outputs(6305)) xor (layer2_outputs(9947));
    outputs(5556) <= layer2_outputs(1206);
    outputs(5557) <= layer2_outputs(9723);
    outputs(5558) <= not((layer2_outputs(162)) and (layer2_outputs(1108)));
    outputs(5559) <= not(layer2_outputs(2055));
    outputs(5560) <= (layer2_outputs(6852)) or (layer2_outputs(1743));
    outputs(5561) <= (layer2_outputs(9600)) xor (layer2_outputs(5965));
    outputs(5562) <= not(layer2_outputs(4477));
    outputs(5563) <= not((layer2_outputs(2833)) and (layer2_outputs(2636)));
    outputs(5564) <= (layer2_outputs(791)) and (layer2_outputs(9803));
    outputs(5565) <= (layer2_outputs(7935)) xor (layer2_outputs(263));
    outputs(5566) <= layer2_outputs(1807);
    outputs(5567) <= layer2_outputs(230);
    outputs(5568) <= not((layer2_outputs(9914)) xor (layer2_outputs(8034)));
    outputs(5569) <= (layer2_outputs(1567)) xor (layer2_outputs(9294));
    outputs(5570) <= not(layer2_outputs(3618));
    outputs(5571) <= not(layer2_outputs(967));
    outputs(5572) <= layer2_outputs(4765);
    outputs(5573) <= layer2_outputs(9630);
    outputs(5574) <= (layer2_outputs(2849)) xor (layer2_outputs(2848));
    outputs(5575) <= (layer2_outputs(5612)) xor (layer2_outputs(620));
    outputs(5576) <= layer2_outputs(7045);
    outputs(5577) <= not(layer2_outputs(8204));
    outputs(5578) <= not(layer2_outputs(1549));
    outputs(5579) <= (layer2_outputs(9363)) and (layer2_outputs(5796));
    outputs(5580) <= not((layer2_outputs(7396)) xor (layer2_outputs(210)));
    outputs(5581) <= (layer2_outputs(7387)) xor (layer2_outputs(8529));
    outputs(5582) <= layer2_outputs(6052);
    outputs(5583) <= not(layer2_outputs(4900));
    outputs(5584) <= not(layer2_outputs(3978));
    outputs(5585) <= not((layer2_outputs(1376)) xor (layer2_outputs(8624)));
    outputs(5586) <= not(layer2_outputs(6002)) or (layer2_outputs(6864));
    outputs(5587) <= layer2_outputs(6739);
    outputs(5588) <= not(layer2_outputs(1506));
    outputs(5589) <= layer2_outputs(1286);
    outputs(5590) <= layer2_outputs(5903);
    outputs(5591) <= layer2_outputs(2921);
    outputs(5592) <= (layer2_outputs(9221)) and not (layer2_outputs(8826));
    outputs(5593) <= (layer2_outputs(10041)) xor (layer2_outputs(8288));
    outputs(5594) <= not(layer2_outputs(6098));
    outputs(5595) <= not(layer2_outputs(1770));
    outputs(5596) <= layer2_outputs(8754);
    outputs(5597) <= not(layer2_outputs(1427));
    outputs(5598) <= layer2_outputs(2241);
    outputs(5599) <= not(layer2_outputs(3397)) or (layer2_outputs(7494));
    outputs(5600) <= not(layer2_outputs(9155));
    outputs(5601) <= (layer2_outputs(9599)) or (layer2_outputs(3634));
    outputs(5602) <= layer2_outputs(9602);
    outputs(5603) <= not((layer2_outputs(2260)) xor (layer2_outputs(9998)));
    outputs(5604) <= layer2_outputs(615);
    outputs(5605) <= not(layer2_outputs(2089)) or (layer2_outputs(8269));
    outputs(5606) <= not(layer2_outputs(4662));
    outputs(5607) <= not(layer2_outputs(297));
    outputs(5608) <= layer2_outputs(8653);
    outputs(5609) <= not((layer2_outputs(6830)) or (layer2_outputs(3353)));
    outputs(5610) <= not(layer2_outputs(3493));
    outputs(5611) <= not(layer2_outputs(477)) or (layer2_outputs(1254));
    outputs(5612) <= (layer2_outputs(3458)) xor (layer2_outputs(1533));
    outputs(5613) <= layer2_outputs(7143);
    outputs(5614) <= (layer2_outputs(542)) xor (layer2_outputs(2278));
    outputs(5615) <= layer2_outputs(2066);
    outputs(5616) <= not(layer2_outputs(8688));
    outputs(5617) <= layer2_outputs(1582);
    outputs(5618) <= (layer2_outputs(212)) xor (layer2_outputs(2163));
    outputs(5619) <= (layer2_outputs(6776)) xor (layer2_outputs(2749));
    outputs(5620) <= layer2_outputs(3492);
    outputs(5621) <= layer2_outputs(8698);
    outputs(5622) <= not((layer2_outputs(6547)) or (layer2_outputs(5560)));
    outputs(5623) <= not(layer2_outputs(3812));
    outputs(5624) <= not((layer2_outputs(1810)) xor (layer2_outputs(6784)));
    outputs(5625) <= layer2_outputs(8757);
    outputs(5626) <= not(layer2_outputs(3544));
    outputs(5627) <= layer2_outputs(2327);
    outputs(5628) <= layer2_outputs(1850);
    outputs(5629) <= not(layer2_outputs(9386));
    outputs(5630) <= not(layer2_outputs(2657));
    outputs(5631) <= not(layer2_outputs(6879));
    outputs(5632) <= not(layer2_outputs(6624));
    outputs(5633) <= layer2_outputs(141);
    outputs(5634) <= not(layer2_outputs(4243));
    outputs(5635) <= not(layer2_outputs(1504)) or (layer2_outputs(3417));
    outputs(5636) <= not(layer2_outputs(309)) or (layer2_outputs(5677));
    outputs(5637) <= not((layer2_outputs(2103)) xor (layer2_outputs(395)));
    outputs(5638) <= not(layer2_outputs(3296));
    outputs(5639) <= not((layer2_outputs(4697)) xor (layer2_outputs(7477)));
    outputs(5640) <= not(layer2_outputs(6871));
    outputs(5641) <= (layer2_outputs(8682)) xor (layer2_outputs(1562));
    outputs(5642) <= not((layer2_outputs(1503)) xor (layer2_outputs(7664)));
    outputs(5643) <= not(layer2_outputs(4439));
    outputs(5644) <= (layer2_outputs(2077)) or (layer2_outputs(8915));
    outputs(5645) <= layer2_outputs(4818);
    outputs(5646) <= layer2_outputs(6663);
    outputs(5647) <= not(layer2_outputs(9268));
    outputs(5648) <= layer2_outputs(4532);
    outputs(5649) <= not((layer2_outputs(5741)) xor (layer2_outputs(128)));
    outputs(5650) <= not(layer2_outputs(6278));
    outputs(5651) <= layer2_outputs(10107);
    outputs(5652) <= layer2_outputs(638);
    outputs(5653) <= not(layer2_outputs(7519));
    outputs(5654) <= layer2_outputs(48);
    outputs(5655) <= (layer2_outputs(4916)) xor (layer2_outputs(7203));
    outputs(5656) <= not(layer2_outputs(8208));
    outputs(5657) <= not((layer2_outputs(7551)) or (layer2_outputs(285)));
    outputs(5658) <= (layer2_outputs(512)) xor (layer2_outputs(6890));
    outputs(5659) <= layer2_outputs(9602);
    outputs(5660) <= (layer2_outputs(758)) and not (layer2_outputs(6527));
    outputs(5661) <= layer2_outputs(1006);
    outputs(5662) <= not(layer2_outputs(8665));
    outputs(5663) <= not(layer2_outputs(3437));
    outputs(5664) <= not(layer2_outputs(8805));
    outputs(5665) <= not((layer2_outputs(7388)) xor (layer2_outputs(3552)));
    outputs(5666) <= not(layer2_outputs(5004));
    outputs(5667) <= layer2_outputs(2301);
    outputs(5668) <= not(layer2_outputs(7085));
    outputs(5669) <= layer2_outputs(9250);
    outputs(5670) <= not((layer2_outputs(10135)) xor (layer2_outputs(1563)));
    outputs(5671) <= not(layer2_outputs(7988)) or (layer2_outputs(733));
    outputs(5672) <= layer2_outputs(3979);
    outputs(5673) <= (layer2_outputs(1657)) xor (layer2_outputs(8118));
    outputs(5674) <= not(layer2_outputs(6356));
    outputs(5675) <= not(layer2_outputs(5580));
    outputs(5676) <= not((layer2_outputs(1769)) xor (layer2_outputs(1452)));
    outputs(5677) <= (layer2_outputs(7556)) xor (layer2_outputs(10005));
    outputs(5678) <= not((layer2_outputs(1298)) or (layer2_outputs(2571)));
    outputs(5679) <= (layer2_outputs(9040)) xor (layer2_outputs(5685));
    outputs(5680) <= not(layer2_outputs(1389));
    outputs(5681) <= (layer2_outputs(7222)) or (layer2_outputs(4496));
    outputs(5682) <= not((layer2_outputs(9711)) and (layer2_outputs(10109)));
    outputs(5683) <= not(layer2_outputs(5983));
    outputs(5684) <= (layer2_outputs(3929)) and not (layer2_outputs(8205));
    outputs(5685) <= (layer2_outputs(2166)) or (layer2_outputs(2027));
    outputs(5686) <= layer2_outputs(7878);
    outputs(5687) <= layer2_outputs(6918);
    outputs(5688) <= (layer2_outputs(7672)) and not (layer2_outputs(7007));
    outputs(5689) <= not(layer2_outputs(764)) or (layer2_outputs(9769));
    outputs(5690) <= not((layer2_outputs(2951)) xor (layer2_outputs(4605)));
    outputs(5691) <= (layer2_outputs(632)) xor (layer2_outputs(8821));
    outputs(5692) <= layer2_outputs(7439);
    outputs(5693) <= not((layer2_outputs(7205)) or (layer2_outputs(6306)));
    outputs(5694) <= not(layer2_outputs(2849));
    outputs(5695) <= not(layer2_outputs(6414));
    outputs(5696) <= not(layer2_outputs(3190));
    outputs(5697) <= layer2_outputs(2222);
    outputs(5698) <= (layer2_outputs(8908)) and not (layer2_outputs(6764));
    outputs(5699) <= layer2_outputs(8179);
    outputs(5700) <= (layer2_outputs(4107)) xor (layer2_outputs(2252));
    outputs(5701) <= layer2_outputs(1602);
    outputs(5702) <= (layer2_outputs(10227)) xor (layer2_outputs(8830));
    outputs(5703) <= (layer2_outputs(5511)) or (layer2_outputs(350));
    outputs(5704) <= layer2_outputs(3707);
    outputs(5705) <= not(layer2_outputs(2965));
    outputs(5706) <= not(layer2_outputs(8079));
    outputs(5707) <= layer2_outputs(4331);
    outputs(5708) <= not(layer2_outputs(2185));
    outputs(5709) <= layer2_outputs(3468);
    outputs(5710) <= not(layer2_outputs(3280));
    outputs(5711) <= not(layer2_outputs(3426));
    outputs(5712) <= not(layer2_outputs(6291));
    outputs(5713) <= not(layer2_outputs(6887)) or (layer2_outputs(774));
    outputs(5714) <= not(layer2_outputs(5340));
    outputs(5715) <= (layer2_outputs(3124)) xor (layer2_outputs(2565));
    outputs(5716) <= not(layer2_outputs(1553));
    outputs(5717) <= not(layer2_outputs(1153));
    outputs(5718) <= layer2_outputs(5505);
    outputs(5719) <= layer2_outputs(8474);
    outputs(5720) <= not(layer2_outputs(2879));
    outputs(5721) <= (layer2_outputs(8038)) xor (layer2_outputs(9778));
    outputs(5722) <= layer2_outputs(4213);
    outputs(5723) <= layer2_outputs(9538);
    outputs(5724) <= not((layer2_outputs(8562)) xor (layer2_outputs(3553)));
    outputs(5725) <= layer2_outputs(6488);
    outputs(5726) <= not(layer2_outputs(3005));
    outputs(5727) <= not(layer2_outputs(3353));
    outputs(5728) <= (layer2_outputs(4537)) and not (layer2_outputs(3072));
    outputs(5729) <= not((layer2_outputs(4644)) xor (layer2_outputs(8388)));
    outputs(5730) <= not(layer2_outputs(7856));
    outputs(5731) <= (layer2_outputs(7486)) and not (layer2_outputs(10080));
    outputs(5732) <= not((layer2_outputs(6247)) and (layer2_outputs(7035)));
    outputs(5733) <= not(layer2_outputs(5017));
    outputs(5734) <= not(layer2_outputs(114));
    outputs(5735) <= not(layer2_outputs(3131));
    outputs(5736) <= (layer2_outputs(8703)) and (layer2_outputs(4399));
    outputs(5737) <= layer2_outputs(278);
    outputs(5738) <= (layer2_outputs(7152)) xor (layer2_outputs(9811));
    outputs(5739) <= (layer2_outputs(1532)) xor (layer2_outputs(6486));
    outputs(5740) <= layer2_outputs(1299);
    outputs(5741) <= layer2_outputs(4420);
    outputs(5742) <= (layer2_outputs(2023)) and (layer2_outputs(9863));
    outputs(5743) <= not((layer2_outputs(3951)) xor (layer2_outputs(9215)));
    outputs(5744) <= not(layer2_outputs(2001));
    outputs(5745) <= not((layer2_outputs(2575)) xor (layer2_outputs(4027)));
    outputs(5746) <= layer2_outputs(4086);
    outputs(5747) <= not(layer2_outputs(832));
    outputs(5748) <= not((layer2_outputs(3474)) xor (layer2_outputs(663)));
    outputs(5749) <= not(layer2_outputs(77));
    outputs(5750) <= (layer2_outputs(5487)) xor (layer2_outputs(3306));
    outputs(5751) <= not(layer2_outputs(4619));
    outputs(5752) <= not(layer2_outputs(7491));
    outputs(5753) <= layer2_outputs(756);
    outputs(5754) <= layer2_outputs(3192);
    outputs(5755) <= layer2_outputs(6213);
    outputs(5756) <= not(layer2_outputs(17));
    outputs(5757) <= not(layer2_outputs(1171));
    outputs(5758) <= layer2_outputs(9765);
    outputs(5759) <= layer2_outputs(6416);
    outputs(5760) <= not(layer2_outputs(9708));
    outputs(5761) <= layer2_outputs(5182);
    outputs(5762) <= layer2_outputs(2095);
    outputs(5763) <= layer2_outputs(9845);
    outputs(5764) <= not((layer2_outputs(1736)) xor (layer2_outputs(635)));
    outputs(5765) <= not(layer2_outputs(2160));
    outputs(5766) <= not((layer2_outputs(8266)) or (layer2_outputs(52)));
    outputs(5767) <= layer2_outputs(7363);
    outputs(5768) <= not(layer2_outputs(3600));
    outputs(5769) <= not((layer2_outputs(7280)) xor (layer2_outputs(3529)));
    outputs(5770) <= not(layer2_outputs(10106));
    outputs(5771) <= layer2_outputs(73);
    outputs(5772) <= not(layer2_outputs(7365));
    outputs(5773) <= not(layer2_outputs(4852));
    outputs(5774) <= not(layer2_outputs(1198));
    outputs(5775) <= layer2_outputs(4875);
    outputs(5776) <= not(layer2_outputs(5058));
    outputs(5777) <= not(layer2_outputs(2160));
    outputs(5778) <= not(layer2_outputs(7786));
    outputs(5779) <= not((layer2_outputs(6089)) xor (layer2_outputs(5840)));
    outputs(5780) <= not((layer2_outputs(115)) and (layer2_outputs(5469)));
    outputs(5781) <= (layer2_outputs(5264)) and not (layer2_outputs(2137));
    outputs(5782) <= not((layer2_outputs(8881)) or (layer2_outputs(4602)));
    outputs(5783) <= layer2_outputs(7137);
    outputs(5784) <= not((layer2_outputs(6429)) and (layer2_outputs(5558)));
    outputs(5785) <= not(layer2_outputs(6423));
    outputs(5786) <= not(layer2_outputs(8462));
    outputs(5787) <= (layer2_outputs(861)) and (layer2_outputs(2237));
    outputs(5788) <= layer2_outputs(4232);
    outputs(5789) <= not(layer2_outputs(7163));
    outputs(5790) <= layer2_outputs(752);
    outputs(5791) <= not(layer2_outputs(6774));
    outputs(5792) <= not(layer2_outputs(6421)) or (layer2_outputs(2720));
    outputs(5793) <= not(layer2_outputs(1034));
    outputs(5794) <= not(layer2_outputs(778));
    outputs(5795) <= layer2_outputs(1035);
    outputs(5796) <= not((layer2_outputs(5443)) xor (layer2_outputs(7362)));
    outputs(5797) <= not(layer2_outputs(283));
    outputs(5798) <= not(layer2_outputs(6406));
    outputs(5799) <= not(layer2_outputs(7164));
    outputs(5800) <= layer2_outputs(7692);
    outputs(5801) <= not((layer2_outputs(5069)) or (layer2_outputs(3728)));
    outputs(5802) <= not((layer2_outputs(5280)) xor (layer2_outputs(5391)));
    outputs(5803) <= layer2_outputs(500);
    outputs(5804) <= not(layer2_outputs(6695));
    outputs(5805) <= not(layer2_outputs(6827));
    outputs(5806) <= not((layer2_outputs(10050)) or (layer2_outputs(5653)));
    outputs(5807) <= layer2_outputs(7700);
    outputs(5808) <= layer2_outputs(8197);
    outputs(5809) <= (layer2_outputs(2228)) xor (layer2_outputs(10095));
    outputs(5810) <= layer2_outputs(6118);
    outputs(5811) <= not((layer2_outputs(8219)) or (layer2_outputs(8487)));
    outputs(5812) <= not(layer2_outputs(8356));
    outputs(5813) <= layer2_outputs(2621);
    outputs(5814) <= layer2_outputs(1552);
    outputs(5815) <= not(layer2_outputs(2279)) or (layer2_outputs(7444));
    outputs(5816) <= not(layer2_outputs(3834));
    outputs(5817) <= not((layer2_outputs(3103)) xor (layer2_outputs(223)));
    outputs(5818) <= not(layer2_outputs(4776));
    outputs(5819) <= not((layer2_outputs(3533)) xor (layer2_outputs(3075)));
    outputs(5820) <= not(layer2_outputs(5497));
    outputs(5821) <= not((layer2_outputs(5498)) xor (layer2_outputs(4187)));
    outputs(5822) <= not((layer2_outputs(4675)) and (layer2_outputs(3835)));
    outputs(5823) <= (layer2_outputs(518)) xor (layer2_outputs(9030));
    outputs(5824) <= not(layer2_outputs(9969));
    outputs(5825) <= layer2_outputs(2684);
    outputs(5826) <= not(layer2_outputs(1661));
    outputs(5827) <= (layer2_outputs(2863)) and not (layer2_outputs(7200));
    outputs(5828) <= (layer2_outputs(1307)) xor (layer2_outputs(10151));
    outputs(5829) <= not(layer2_outputs(9495));
    outputs(5830) <= not(layer2_outputs(4114)) or (layer2_outputs(7076));
    outputs(5831) <= layer2_outputs(303);
    outputs(5832) <= not(layer2_outputs(5117));
    outputs(5833) <= layer2_outputs(7001);
    outputs(5834) <= layer2_outputs(1821);
    outputs(5835) <= not((layer2_outputs(2802)) xor (layer2_outputs(3211)));
    outputs(5836) <= not((layer2_outputs(1869)) xor (layer2_outputs(9988)));
    outputs(5837) <= layer2_outputs(3511);
    outputs(5838) <= layer2_outputs(7114);
    outputs(5839) <= not(layer2_outputs(10141));
    outputs(5840) <= not(layer2_outputs(1471));
    outputs(5841) <= layer2_outputs(7783);
    outputs(5842) <= not(layer2_outputs(6511));
    outputs(5843) <= layer2_outputs(6751);
    outputs(5844) <= not(layer2_outputs(949));
    outputs(5845) <= (layer2_outputs(8429)) or (layer2_outputs(8392));
    outputs(5846) <= not(layer2_outputs(1827));
    outputs(5847) <= not((layer2_outputs(3148)) and (layer2_outputs(8581)));
    outputs(5848) <= layer2_outputs(9578);
    outputs(5849) <= not(layer2_outputs(430)) or (layer2_outputs(5467));
    outputs(5850) <= not(layer2_outputs(4550)) or (layer2_outputs(1872));
    outputs(5851) <= not(layer2_outputs(7699));
    outputs(5852) <= not((layer2_outputs(9729)) xor (layer2_outputs(7227)));
    outputs(5853) <= not(layer2_outputs(1957));
    outputs(5854) <= not(layer2_outputs(6625));
    outputs(5855) <= not((layer2_outputs(4483)) xor (layer2_outputs(4503)));
    outputs(5856) <= layer2_outputs(2422);
    outputs(5857) <= not(layer2_outputs(3642));
    outputs(5858) <= layer2_outputs(6273);
    outputs(5859) <= not(layer2_outputs(4320)) or (layer2_outputs(10072));
    outputs(5860) <= (layer2_outputs(2007)) and not (layer2_outputs(2687));
    outputs(5861) <= layer2_outputs(498);
    outputs(5862) <= not(layer2_outputs(1975));
    outputs(5863) <= layer2_outputs(8263);
    outputs(5864) <= layer2_outputs(9758);
    outputs(5865) <= not(layer2_outputs(3361)) or (layer2_outputs(14));
    outputs(5866) <= not((layer2_outputs(7254)) xor (layer2_outputs(938)));
    outputs(5867) <= layer2_outputs(4686);
    outputs(5868) <= layer2_outputs(1234);
    outputs(5869) <= not(layer2_outputs(9871));
    outputs(5870) <= layer2_outputs(5979);
    outputs(5871) <= not((layer2_outputs(5769)) xor (layer2_outputs(6646)));
    outputs(5872) <= layer2_outputs(7028);
    outputs(5873) <= not((layer2_outputs(7021)) xor (layer2_outputs(8578)));
    outputs(5874) <= layer2_outputs(7552);
    outputs(5875) <= (layer2_outputs(9087)) xor (layer2_outputs(1992));
    outputs(5876) <= not(layer2_outputs(10071));
    outputs(5877) <= layer2_outputs(7222);
    outputs(5878) <= layer2_outputs(481);
    outputs(5879) <= (layer2_outputs(2582)) xor (layer2_outputs(2239));
    outputs(5880) <= (layer2_outputs(2631)) and not (layer2_outputs(4251));
    outputs(5881) <= not(layer2_outputs(1429));
    outputs(5882) <= layer2_outputs(1645);
    outputs(5883) <= not(layer2_outputs(9743));
    outputs(5884) <= (layer2_outputs(4121)) xor (layer2_outputs(4332));
    outputs(5885) <= (layer2_outputs(8772)) and not (layer2_outputs(4137));
    outputs(5886) <= layer2_outputs(603);
    outputs(5887) <= (layer2_outputs(7320)) and not (layer2_outputs(590));
    outputs(5888) <= not((layer2_outputs(9251)) xor (layer2_outputs(1076)));
    outputs(5889) <= not(layer2_outputs(2460));
    outputs(5890) <= (layer2_outputs(1636)) xor (layer2_outputs(6073));
    outputs(5891) <= (layer2_outputs(5416)) xor (layer2_outputs(4002));
    outputs(5892) <= (layer2_outputs(972)) xor (layer2_outputs(9449));
    outputs(5893) <= not(layer2_outputs(3263)) or (layer2_outputs(5663));
    outputs(5894) <= layer2_outputs(6289);
    outputs(5895) <= not((layer2_outputs(9428)) xor (layer2_outputs(1349)));
    outputs(5896) <= not((layer2_outputs(2338)) xor (layer2_outputs(7492)));
    outputs(5897) <= not((layer2_outputs(4542)) xor (layer2_outputs(3978)));
    outputs(5898) <= not((layer2_outputs(3056)) xor (layer2_outputs(8997)));
    outputs(5899) <= (layer2_outputs(8251)) xor (layer2_outputs(9767));
    outputs(5900) <= (layer2_outputs(7605)) or (layer2_outputs(6452));
    outputs(5901) <= layer2_outputs(4824);
    outputs(5902) <= layer2_outputs(4229);
    outputs(5903) <= (layer2_outputs(1808)) or (layer2_outputs(6843));
    outputs(5904) <= (layer2_outputs(6265)) and not (layer2_outputs(10166));
    outputs(5905) <= layer2_outputs(6333);
    outputs(5906) <= layer2_outputs(9850);
    outputs(5907) <= not(layer2_outputs(4926));
    outputs(5908) <= not(layer2_outputs(4681));
    outputs(5909) <= layer2_outputs(8350);
    outputs(5910) <= not((layer2_outputs(6216)) and (layer2_outputs(8789)));
    outputs(5911) <= not(layer2_outputs(4996)) or (layer2_outputs(445));
    outputs(5912) <= layer2_outputs(363);
    outputs(5913) <= layer2_outputs(10091);
    outputs(5914) <= not(layer2_outputs(7518));
    outputs(5915) <= layer2_outputs(7136);
    outputs(5916) <= layer2_outputs(8273);
    outputs(5917) <= layer2_outputs(4128);
    outputs(5918) <= layer2_outputs(667);
    outputs(5919) <= layer2_outputs(9653);
    outputs(5920) <= not(layer2_outputs(1389));
    outputs(5921) <= layer2_outputs(457);
    outputs(5922) <= (layer2_outputs(8801)) and (layer2_outputs(351));
    outputs(5923) <= not((layer2_outputs(5676)) or (layer2_outputs(5455)));
    outputs(5924) <= not(layer2_outputs(10122));
    outputs(5925) <= not(layer2_outputs(1919));
    outputs(5926) <= (layer2_outputs(3092)) xor (layer2_outputs(9136));
    outputs(5927) <= not((layer2_outputs(3279)) xor (layer2_outputs(8102)));
    outputs(5928) <= not((layer2_outputs(4396)) xor (layer2_outputs(7428)));
    outputs(5929) <= not(layer2_outputs(7812));
    outputs(5930) <= not(layer2_outputs(8385));
    outputs(5931) <= not(layer2_outputs(6672));
    outputs(5932) <= (layer2_outputs(4389)) xor (layer2_outputs(4377));
    outputs(5933) <= layer2_outputs(1537);
    outputs(5934) <= not(layer2_outputs(7879));
    outputs(5935) <= layer2_outputs(8048);
    outputs(5936) <= not(layer2_outputs(10123));
    outputs(5937) <= not(layer2_outputs(7237));
    outputs(5938) <= not((layer2_outputs(4344)) or (layer2_outputs(6709)));
    outputs(5939) <= layer2_outputs(8017);
    outputs(5940) <= not(layer2_outputs(1889));
    outputs(5941) <= (layer2_outputs(717)) xor (layer2_outputs(4370));
    outputs(5942) <= (layer2_outputs(1665)) xor (layer2_outputs(8069));
    outputs(5943) <= not(layer2_outputs(9069));
    outputs(5944) <= not((layer2_outputs(7406)) xor (layer2_outputs(7360)));
    outputs(5945) <= layer2_outputs(2173);
    outputs(5946) <= (layer2_outputs(5247)) and (layer2_outputs(2134));
    outputs(5947) <= not((layer2_outputs(8925)) and (layer2_outputs(2529)));
    outputs(5948) <= layer2_outputs(3404);
    outputs(5949) <= not(layer2_outputs(7454));
    outputs(5950) <= not(layer2_outputs(5094));
    outputs(5951) <= not((layer2_outputs(4118)) xor (layer2_outputs(2948)));
    outputs(5952) <= not((layer2_outputs(5421)) xor (layer2_outputs(8449)));
    outputs(5953) <= not(layer2_outputs(7029));
    outputs(5954) <= not(layer2_outputs(174));
    outputs(5955) <= not(layer2_outputs(5472));
    outputs(5956) <= not(layer2_outputs(8101));
    outputs(5957) <= not(layer2_outputs(9488));
    outputs(5958) <= (layer2_outputs(6144)) xor (layer2_outputs(7103));
    outputs(5959) <= (layer2_outputs(11)) xor (layer2_outputs(3310));
    outputs(5960) <= layer2_outputs(8530);
    outputs(5961) <= not((layer2_outputs(7960)) and (layer2_outputs(7676)));
    outputs(5962) <= layer2_outputs(10085);
    outputs(5963) <= (layer2_outputs(3284)) xor (layer2_outputs(6198));
    outputs(5964) <= layer2_outputs(4097);
    outputs(5965) <= (layer2_outputs(226)) xor (layer2_outputs(7037));
    outputs(5966) <= (layer2_outputs(5588)) xor (layer2_outputs(8638));
    outputs(5967) <= not(layer2_outputs(3603));
    outputs(5968) <= not((layer2_outputs(5638)) xor (layer2_outputs(2210)));
    outputs(5969) <= not(layer2_outputs(4507));
    outputs(5970) <= not(layer2_outputs(1680));
    outputs(5971) <= not((layer2_outputs(1578)) and (layer2_outputs(4616)));
    outputs(5972) <= not((layer2_outputs(242)) xor (layer2_outputs(8832)));
    outputs(5973) <= not(layer2_outputs(5483));
    outputs(5974) <= (layer2_outputs(1453)) and not (layer2_outputs(3320));
    outputs(5975) <= layer2_outputs(4726);
    outputs(5976) <= layer2_outputs(4225);
    outputs(5977) <= not(layer2_outputs(1839));
    outputs(5978) <= layer2_outputs(3993);
    outputs(5979) <= layer2_outputs(8907);
    outputs(5980) <= not((layer2_outputs(5802)) xor (layer2_outputs(8191)));
    outputs(5981) <= (layer2_outputs(3773)) and not (layer2_outputs(6892));
    outputs(5982) <= not((layer2_outputs(8174)) xor (layer2_outputs(2310)));
    outputs(5983) <= layer2_outputs(7915);
    outputs(5984) <= layer2_outputs(1170);
    outputs(5985) <= layer2_outputs(5366);
    outputs(5986) <= not(layer2_outputs(1364));
    outputs(5987) <= not((layer2_outputs(4956)) or (layer2_outputs(4186)));
    outputs(5988) <= layer2_outputs(7378);
    outputs(5989) <= not(layer2_outputs(7794));
    outputs(5990) <= not((layer2_outputs(6400)) or (layer2_outputs(2118)));
    outputs(5991) <= (layer2_outputs(8232)) xor (layer2_outputs(5068));
    outputs(5992) <= layer2_outputs(7713);
    outputs(5993) <= (layer2_outputs(9521)) and (layer2_outputs(2431));
    outputs(5994) <= not(layer2_outputs(9090));
    outputs(5995) <= layer2_outputs(9455);
    outputs(5996) <= layer2_outputs(8638);
    outputs(5997) <= layer2_outputs(5435);
    outputs(5998) <= layer2_outputs(6833);
    outputs(5999) <= not(layer2_outputs(4721));
    outputs(6000) <= not((layer2_outputs(10053)) xor (layer2_outputs(6299)));
    outputs(6001) <= not(layer2_outputs(739));
    outputs(6002) <= not((layer2_outputs(7810)) xor (layer2_outputs(5622)));
    outputs(6003) <= (layer2_outputs(7968)) xor (layer2_outputs(7535));
    outputs(6004) <= not(layer2_outputs(3938));
    outputs(6005) <= not(layer2_outputs(145)) or (layer2_outputs(6054));
    outputs(6006) <= not(layer2_outputs(8665));
    outputs(6007) <= not((layer2_outputs(5289)) and (layer2_outputs(5348)));
    outputs(6008) <= (layer2_outputs(813)) and (layer2_outputs(1686));
    outputs(6009) <= not(layer2_outputs(5543)) or (layer2_outputs(9886));
    outputs(6010) <= layer2_outputs(3956);
    outputs(6011) <= (layer2_outputs(10075)) xor (layer2_outputs(1755));
    outputs(6012) <= not((layer2_outputs(3354)) and (layer2_outputs(7658)));
    outputs(6013) <= not(layer2_outputs(3713)) or (layer2_outputs(2857));
    outputs(6014) <= (layer2_outputs(5700)) xor (layer2_outputs(6036));
    outputs(6015) <= layer2_outputs(7843);
    outputs(6016) <= layer2_outputs(2782);
    outputs(6017) <= (layer2_outputs(2865)) or (layer2_outputs(7356));
    outputs(6018) <= layer2_outputs(4072);
    outputs(6019) <= (layer2_outputs(1650)) xor (layer2_outputs(8548));
    outputs(6020) <= not(layer2_outputs(4864));
    outputs(6021) <= not(layer2_outputs(5016)) or (layer2_outputs(8342));
    outputs(6022) <= not(layer2_outputs(824));
    outputs(6023) <= layer2_outputs(341);
    outputs(6024) <= not(layer2_outputs(6518));
    outputs(6025) <= layer2_outputs(6354);
    outputs(6026) <= layer2_outputs(8304);
    outputs(6027) <= layer2_outputs(7269);
    outputs(6028) <= not(layer2_outputs(9882));
    outputs(6029) <= layer2_outputs(2952);
    outputs(6030) <= layer2_outputs(1535);
    outputs(6031) <= (layer2_outputs(5583)) xor (layer2_outputs(7266));
    outputs(6032) <= (layer2_outputs(204)) xor (layer2_outputs(4614));
    outputs(6033) <= not(layer2_outputs(7354));
    outputs(6034) <= layer2_outputs(7889);
    outputs(6035) <= layer2_outputs(6544);
    outputs(6036) <= layer2_outputs(9175);
    outputs(6037) <= layer2_outputs(6078);
    outputs(6038) <= not(layer2_outputs(10190));
    outputs(6039) <= not((layer2_outputs(6822)) xor (layer2_outputs(7828)));
    outputs(6040) <= not(layer2_outputs(5060));
    outputs(6041) <= layer2_outputs(9803);
    outputs(6042) <= layer2_outputs(9256);
    outputs(6043) <= (layer2_outputs(2893)) xor (layer2_outputs(1986));
    outputs(6044) <= layer2_outputs(7604);
    outputs(6045) <= not((layer2_outputs(115)) xor (layer2_outputs(2428)));
    outputs(6046) <= layer2_outputs(5431);
    outputs(6047) <= not((layer2_outputs(992)) xor (layer2_outputs(5308)));
    outputs(6048) <= (layer2_outputs(7781)) xor (layer2_outputs(1402));
    outputs(6049) <= not(layer2_outputs(6744));
    outputs(6050) <= layer2_outputs(3818);
    outputs(6051) <= (layer2_outputs(8296)) xor (layer2_outputs(1179));
    outputs(6052) <= layer2_outputs(2249);
    outputs(6053) <= not(layer2_outputs(5361));
    outputs(6054) <= not(layer2_outputs(8660));
    outputs(6055) <= not(layer2_outputs(3298));
    outputs(6056) <= layer2_outputs(5093);
    outputs(6057) <= not(layer2_outputs(7196));
    outputs(6058) <= not((layer2_outputs(7972)) and (layer2_outputs(1896)));
    outputs(6059) <= (layer2_outputs(463)) xor (layer2_outputs(3463));
    outputs(6060) <= not((layer2_outputs(486)) xor (layer2_outputs(876)));
    outputs(6061) <= not((layer2_outputs(1765)) xor (layer2_outputs(2730)));
    outputs(6062) <= layer2_outputs(7449);
    outputs(6063) <= not((layer2_outputs(1796)) xor (layer2_outputs(3038)));
    outputs(6064) <= not(layer2_outputs(7443));
    outputs(6065) <= not((layer2_outputs(5757)) xor (layer2_outputs(63)));
    outputs(6066) <= (layer2_outputs(3545)) xor (layer2_outputs(2172));
    outputs(6067) <= not(layer2_outputs(8817)) or (layer2_outputs(467));
    outputs(6068) <= not((layer2_outputs(2819)) xor (layer2_outputs(3670)));
    outputs(6069) <= layer2_outputs(5298);
    outputs(6070) <= not(layer2_outputs(1721));
    outputs(6071) <= not(layer2_outputs(6051));
    outputs(6072) <= layer2_outputs(3351);
    outputs(6073) <= (layer2_outputs(9707)) and (layer2_outputs(1406));
    outputs(6074) <= not((layer2_outputs(1833)) or (layer2_outputs(1677)));
    outputs(6075) <= layer2_outputs(8347);
    outputs(6076) <= layer2_outputs(4711);
    outputs(6077) <= not((layer2_outputs(2317)) xor (layer2_outputs(4900)));
    outputs(6078) <= layer2_outputs(4537);
    outputs(6079) <= not((layer2_outputs(7074)) and (layer2_outputs(9715)));
    outputs(6080) <= (layer2_outputs(601)) or (layer2_outputs(6519));
    outputs(6081) <= not(layer2_outputs(3062));
    outputs(6082) <= layer2_outputs(6544);
    outputs(6083) <= not(layer2_outputs(4556));
    outputs(6084) <= (layer2_outputs(6461)) and not (layer2_outputs(840));
    outputs(6085) <= (layer2_outputs(2459)) and not (layer2_outputs(2261));
    outputs(6086) <= not((layer2_outputs(6386)) xor (layer2_outputs(930)));
    outputs(6087) <= layer2_outputs(5790);
    outputs(6088) <= not(layer2_outputs(6128));
    outputs(6089) <= layer2_outputs(6345);
    outputs(6090) <= not((layer2_outputs(6163)) xor (layer2_outputs(9254)));
    outputs(6091) <= not(layer2_outputs(1437));
    outputs(6092) <= (layer2_outputs(3602)) xor (layer2_outputs(9650));
    outputs(6093) <= (layer2_outputs(3508)) and not (layer2_outputs(2716));
    outputs(6094) <= not((layer2_outputs(8591)) or (layer2_outputs(6766)));
    outputs(6095) <= layer2_outputs(6031);
    outputs(6096) <= layer2_outputs(9733);
    outputs(6097) <= layer2_outputs(5684);
    outputs(6098) <= layer2_outputs(8370);
    outputs(6099) <= layer2_outputs(3878);
    outputs(6100) <= not((layer2_outputs(1015)) xor (layer2_outputs(7937)));
    outputs(6101) <= (layer2_outputs(1725)) xor (layer2_outputs(2592));
    outputs(6102) <= not(layer2_outputs(6252)) or (layer2_outputs(7119));
    outputs(6103) <= not(layer2_outputs(4344));
    outputs(6104) <= (layer2_outputs(3875)) and not (layer2_outputs(9045));
    outputs(6105) <= (layer2_outputs(6463)) xor (layer2_outputs(8053));
    outputs(6106) <= not(layer2_outputs(7262));
    outputs(6107) <= not((layer2_outputs(4882)) xor (layer2_outputs(3765)));
    outputs(6108) <= not(layer2_outputs(8303));
    outputs(6109) <= (layer2_outputs(79)) or (layer2_outputs(1698));
    outputs(6110) <= not(layer2_outputs(2526));
    outputs(6111) <= layer2_outputs(4262);
    outputs(6112) <= (layer2_outputs(9345)) and not (layer2_outputs(3453));
    outputs(6113) <= not((layer2_outputs(1297)) and (layer2_outputs(3161)));
    outputs(6114) <= not(layer2_outputs(9595));
    outputs(6115) <= layer2_outputs(138);
    outputs(6116) <= not(layer2_outputs(6927));
    outputs(6117) <= not(layer2_outputs(5855)) or (layer2_outputs(1242));
    outputs(6118) <= not(layer2_outputs(1978));
    outputs(6119) <= not(layer2_outputs(7760));
    outputs(6120) <= layer2_outputs(7800);
    outputs(6121) <= layer2_outputs(8927);
    outputs(6122) <= (layer2_outputs(350)) and not (layer2_outputs(2266));
    outputs(6123) <= not((layer2_outputs(4799)) xor (layer2_outputs(1739)));
    outputs(6124) <= layer2_outputs(5204);
    outputs(6125) <= (layer2_outputs(7911)) xor (layer2_outputs(86));
    outputs(6126) <= not(layer2_outputs(5933));
    outputs(6127) <= not(layer2_outputs(3558));
    outputs(6128) <= not(layer2_outputs(769));
    outputs(6129) <= (layer2_outputs(3228)) or (layer2_outputs(8539));
    outputs(6130) <= not((layer2_outputs(6254)) xor (layer2_outputs(556)));
    outputs(6131) <= not(layer2_outputs(7979));
    outputs(6132) <= not(layer2_outputs(6179));
    outputs(6133) <= layer2_outputs(3415);
    outputs(6134) <= not((layer2_outputs(4713)) xor (layer2_outputs(10026)));
    outputs(6135) <= not(layer2_outputs(6083));
    outputs(6136) <= layer2_outputs(10192);
    outputs(6137) <= (layer2_outputs(8076)) xor (layer2_outputs(6971));
    outputs(6138) <= not(layer2_outputs(235));
    outputs(6139) <= layer2_outputs(4696);
    outputs(6140) <= not(layer2_outputs(823));
    outputs(6141) <= layer2_outputs(10148);
    outputs(6142) <= layer2_outputs(3865);
    outputs(6143) <= (layer2_outputs(7435)) xor (layer2_outputs(5871));
    outputs(6144) <= (layer2_outputs(3155)) and not (layer2_outputs(8205));
    outputs(6145) <= not(layer2_outputs(4582));
    outputs(6146) <= layer2_outputs(3531);
    outputs(6147) <= not(layer2_outputs(6750));
    outputs(6148) <= not(layer2_outputs(7649));
    outputs(6149) <= not(layer2_outputs(4460)) or (layer2_outputs(4694));
    outputs(6150) <= layer2_outputs(3709);
    outputs(6151) <= not(layer2_outputs(8755));
    outputs(6152) <= not(layer2_outputs(10169));
    outputs(6153) <= (layer2_outputs(7713)) and (layer2_outputs(5641));
    outputs(6154) <= not((layer2_outputs(10062)) xor (layer2_outputs(3685)));
    outputs(6155) <= layer2_outputs(2652);
    outputs(6156) <= not(layer2_outputs(5300));
    outputs(6157) <= not(layer2_outputs(8224));
    outputs(6158) <= layer2_outputs(8807);
    outputs(6159) <= not(layer2_outputs(8093));
    outputs(6160) <= not((layer2_outputs(8731)) xor (layer2_outputs(9191)));
    outputs(6161) <= not(layer2_outputs(4458));
    outputs(6162) <= not(layer2_outputs(7151));
    outputs(6163) <= not(layer2_outputs(1421));
    outputs(6164) <= (layer2_outputs(5342)) and (layer2_outputs(3509));
    outputs(6165) <= not(layer2_outputs(3202));
    outputs(6166) <= not(layer2_outputs(441));
    outputs(6167) <= not((layer2_outputs(4768)) xor (layer2_outputs(1778)));
    outputs(6168) <= not(layer2_outputs(9130));
    outputs(6169) <= not((layer2_outputs(3813)) xor (layer2_outputs(1858)));
    outputs(6170) <= (layer2_outputs(784)) or (layer2_outputs(6618));
    outputs(6171) <= not(layer2_outputs(7330));
    outputs(6172) <= (layer2_outputs(414)) and not (layer2_outputs(916));
    outputs(6173) <= layer2_outputs(9149);
    outputs(6174) <= not(layer2_outputs(7266));
    outputs(6175) <= layer2_outputs(58);
    outputs(6176) <= layer2_outputs(9319);
    outputs(6177) <= not(layer2_outputs(7451));
    outputs(6178) <= layer2_outputs(7508);
    outputs(6179) <= not(layer2_outputs(2618));
    outputs(6180) <= layer2_outputs(7615);
    outputs(6181) <= layer2_outputs(7461);
    outputs(6182) <= not(layer2_outputs(1166));
    outputs(6183) <= layer2_outputs(9772);
    outputs(6184) <= not(layer2_outputs(1966));
    outputs(6185) <= not((layer2_outputs(655)) xor (layer2_outputs(3309)));
    outputs(6186) <= layer2_outputs(6526);
    outputs(6187) <= (layer2_outputs(2432)) xor (layer2_outputs(2240));
    outputs(6188) <= not(layer2_outputs(6267));
    outputs(6189) <= layer2_outputs(4393);
    outputs(6190) <= not((layer2_outputs(6)) or (layer2_outputs(3076)));
    outputs(6191) <= not(layer2_outputs(6661));
    outputs(6192) <= not(layer2_outputs(5300));
    outputs(6193) <= layer2_outputs(743);
    outputs(6194) <= layer2_outputs(5234);
    outputs(6195) <= not(layer2_outputs(1595));
    outputs(6196) <= not(layer2_outputs(5869));
    outputs(6197) <= (layer2_outputs(4733)) and not (layer2_outputs(6934));
    outputs(6198) <= layer2_outputs(8965);
    outputs(6199) <= (layer2_outputs(7271)) xor (layer2_outputs(2561));
    outputs(6200) <= not(layer2_outputs(6824));
    outputs(6201) <= layer2_outputs(4447);
    outputs(6202) <= layer2_outputs(1606);
    outputs(6203) <= not(layer2_outputs(343));
    outputs(6204) <= not((layer2_outputs(1399)) xor (layer2_outputs(10067)));
    outputs(6205) <= layer2_outputs(1093);
    outputs(6206) <= not(layer2_outputs(2090));
    outputs(6207) <= not(layer2_outputs(3248));
    outputs(6208) <= layer2_outputs(521);
    outputs(6209) <= not(layer2_outputs(8319));
    outputs(6210) <= layer2_outputs(61);
    outputs(6211) <= (layer2_outputs(3293)) and not (layer2_outputs(4356));
    outputs(6212) <= (layer2_outputs(1781)) xor (layer2_outputs(6900));
    outputs(6213) <= layer2_outputs(5262);
    outputs(6214) <= not(layer2_outputs(8163));
    outputs(6215) <= not(layer2_outputs(5332)) or (layer2_outputs(1904));
    outputs(6216) <= not(layer2_outputs(1078));
    outputs(6217) <= not(layer2_outputs(6839));
    outputs(6218) <= layer2_outputs(6498);
    outputs(6219) <= not(layer2_outputs(8986));
    outputs(6220) <= layer2_outputs(1101);
    outputs(6221) <= not(layer2_outputs(6789));
    outputs(6222) <= layer2_outputs(33);
    outputs(6223) <= not(layer2_outputs(217));
    outputs(6224) <= not(layer2_outputs(362));
    outputs(6225) <= layer2_outputs(4283);
    outputs(6226) <= not(layer2_outputs(2914));
    outputs(6227) <= layer2_outputs(3840);
    outputs(6228) <= (layer2_outputs(8460)) and not (layer2_outputs(85));
    outputs(6229) <= layer2_outputs(5850);
    outputs(6230) <= not(layer2_outputs(9673));
    outputs(6231) <= layer2_outputs(2967);
    outputs(6232) <= not(layer2_outputs(6506));
    outputs(6233) <= layer2_outputs(6182);
    outputs(6234) <= not(layer2_outputs(2342));
    outputs(6235) <= layer2_outputs(872);
    outputs(6236) <= (layer2_outputs(2232)) and not (layer2_outputs(4818));
    outputs(6237) <= (layer2_outputs(6730)) and not (layer2_outputs(6574));
    outputs(6238) <= not((layer2_outputs(5158)) or (layer2_outputs(3798)));
    outputs(6239) <= not((layer2_outputs(3050)) or (layer2_outputs(9866)));
    outputs(6240) <= not(layer2_outputs(243));
    outputs(6241) <= not(layer2_outputs(7503));
    outputs(6242) <= layer2_outputs(8344);
    outputs(6243) <= not(layer2_outputs(8526));
    outputs(6244) <= not((layer2_outputs(349)) xor (layer2_outputs(6936)));
    outputs(6245) <= layer2_outputs(7300);
    outputs(6246) <= (layer2_outputs(10055)) xor (layer2_outputs(313));
    outputs(6247) <= (layer2_outputs(8568)) and (layer2_outputs(9744));
    outputs(6248) <= layer2_outputs(6103);
    outputs(6249) <= not(layer2_outputs(7445)) or (layer2_outputs(1359));
    outputs(6250) <= not(layer2_outputs(4972));
    outputs(6251) <= not(layer2_outputs(4284));
    outputs(6252) <= (layer2_outputs(1865)) xor (layer2_outputs(5133));
    outputs(6253) <= not(layer2_outputs(5844)) or (layer2_outputs(4343));
    outputs(6254) <= not(layer2_outputs(5809));
    outputs(6255) <= layer2_outputs(3592);
    outputs(6256) <= layer2_outputs(1878);
    outputs(6257) <= layer2_outputs(5415);
    outputs(6258) <= layer2_outputs(8639);
    outputs(6259) <= (layer2_outputs(2426)) and not (layer2_outputs(5231));
    outputs(6260) <= layer2_outputs(7378);
    outputs(6261) <= not(layer2_outputs(944));
    outputs(6262) <= (layer2_outputs(286)) xor (layer2_outputs(1063));
    outputs(6263) <= not(layer2_outputs(3358));
    outputs(6264) <= not(layer2_outputs(5130));
    outputs(6265) <= not(layer2_outputs(317));
    outputs(6266) <= not(layer2_outputs(6589)) or (layer2_outputs(3724));
    outputs(6267) <= layer2_outputs(4154);
    outputs(6268) <= not((layer2_outputs(4013)) or (layer2_outputs(2598)));
    outputs(6269) <= (layer2_outputs(5048)) xor (layer2_outputs(2311));
    outputs(6270) <= not(layer2_outputs(4993));
    outputs(6271) <= layer2_outputs(5327);
    outputs(6272) <= layer2_outputs(136);
    outputs(6273) <= not(layer2_outputs(4618));
    outputs(6274) <= layer2_outputs(6395);
    outputs(6275) <= not(layer2_outputs(5730));
    outputs(6276) <= not(layer2_outputs(3338));
    outputs(6277) <= layer2_outputs(78);
    outputs(6278) <= not(layer2_outputs(8877));
    outputs(6279) <= layer2_outputs(1642);
    outputs(6280) <= layer2_outputs(3325);
    outputs(6281) <= not(layer2_outputs(669));
    outputs(6282) <= not(layer2_outputs(8582));
    outputs(6283) <= not((layer2_outputs(4252)) or (layer2_outputs(7630)));
    outputs(6284) <= not(layer2_outputs(8187));
    outputs(6285) <= layer2_outputs(6409);
    outputs(6286) <= (layer2_outputs(4021)) xor (layer2_outputs(1056));
    outputs(6287) <= layer2_outputs(8901);
    outputs(6288) <= layer2_outputs(7884);
    outputs(6289) <= layer2_outputs(9790);
    outputs(6290) <= not(layer2_outputs(4449));
    outputs(6291) <= layer2_outputs(1186);
    outputs(6292) <= layer2_outputs(228);
    outputs(6293) <= layer2_outputs(4205);
    outputs(6294) <= (layer2_outputs(8766)) and not (layer2_outputs(1000));
    outputs(6295) <= layer2_outputs(10072);
    outputs(6296) <= layer2_outputs(2656);
    outputs(6297) <= not(layer2_outputs(5689));
    outputs(6298) <= not(layer2_outputs(6363));
    outputs(6299) <= not(layer2_outputs(595));
    outputs(6300) <= not(layer2_outputs(6235));
    outputs(6301) <= not(layer2_outputs(7697));
    outputs(6302) <= (layer2_outputs(8985)) xor (layer2_outputs(5549));
    outputs(6303) <= not(layer2_outputs(10006));
    outputs(6304) <= (layer2_outputs(6184)) or (layer2_outputs(9212));
    outputs(6305) <= layer2_outputs(6246);
    outputs(6306) <= not(layer2_outputs(1942));
    outputs(6307) <= not(layer2_outputs(9924));
    outputs(6308) <= (layer2_outputs(2315)) xor (layer2_outputs(4561));
    outputs(6309) <= not(layer2_outputs(8912));
    outputs(6310) <= not(layer2_outputs(6099));
    outputs(6311) <= layer2_outputs(4329);
    outputs(6312) <= not(layer2_outputs(8146));
    outputs(6313) <= (layer2_outputs(7033)) xor (layer2_outputs(2737));
    outputs(6314) <= not((layer2_outputs(3098)) and (layer2_outputs(5833)));
    outputs(6315) <= not((layer2_outputs(481)) xor (layer2_outputs(6341)));
    outputs(6316) <= layer2_outputs(4024);
    outputs(6317) <= not(layer2_outputs(2811));
    outputs(6318) <= layer2_outputs(8524);
    outputs(6319) <= (layer2_outputs(3571)) xor (layer2_outputs(3060));
    outputs(6320) <= layer2_outputs(4320);
    outputs(6321) <= not(layer2_outputs(3301));
    outputs(6322) <= layer2_outputs(2673);
    outputs(6323) <= not(layer2_outputs(8148));
    outputs(6324) <= not(layer2_outputs(9105));
    outputs(6325) <= layer2_outputs(6065);
    outputs(6326) <= not(layer2_outputs(8103));
    outputs(6327) <= not((layer2_outputs(903)) or (layer2_outputs(7782)));
    outputs(6328) <= not(layer2_outputs(7990)) or (layer2_outputs(2650));
    outputs(6329) <= not((layer2_outputs(7462)) or (layer2_outputs(1711)));
    outputs(6330) <= not(layer2_outputs(9571));
    outputs(6331) <= not(layer2_outputs(5833));
    outputs(6332) <= layer2_outputs(4231);
    outputs(6333) <= layer2_outputs(9640);
    outputs(6334) <= layer2_outputs(2255);
    outputs(6335) <= layer2_outputs(9902);
    outputs(6336) <= not(layer2_outputs(1649));
    outputs(6337) <= layer2_outputs(9197);
    outputs(6338) <= (layer2_outputs(10061)) xor (layer2_outputs(9899));
    outputs(6339) <= layer2_outputs(9068);
    outputs(6340) <= not(layer2_outputs(1443));
    outputs(6341) <= (layer2_outputs(4487)) and (layer2_outputs(984));
    outputs(6342) <= layer2_outputs(8441);
    outputs(6343) <= layer2_outputs(7249);
    outputs(6344) <= layer2_outputs(7034);
    outputs(6345) <= layer2_outputs(2908);
    outputs(6346) <= not((layer2_outputs(434)) and (layer2_outputs(1287)));
    outputs(6347) <= (layer2_outputs(3484)) xor (layer2_outputs(7296));
    outputs(6348) <= layer2_outputs(5351);
    outputs(6349) <= not((layer2_outputs(10086)) and (layer2_outputs(1942)));
    outputs(6350) <= not(layer2_outputs(6851));
    outputs(6351) <= not(layer2_outputs(8658));
    outputs(6352) <= layer2_outputs(5439);
    outputs(6353) <= layer2_outputs(8302);
    outputs(6354) <= (layer2_outputs(3954)) and (layer2_outputs(9201));
    outputs(6355) <= layer2_outputs(8712);
    outputs(6356) <= not(layer2_outputs(1075));
    outputs(6357) <= not(layer2_outputs(585)) or (layer2_outputs(591));
    outputs(6358) <= layer2_outputs(4147);
    outputs(6359) <= layer2_outputs(6400);
    outputs(6360) <= not((layer2_outputs(5000)) xor (layer2_outputs(454)));
    outputs(6361) <= layer2_outputs(2402);
    outputs(6362) <= (layer2_outputs(3408)) or (layer2_outputs(178));
    outputs(6363) <= layer2_outputs(9564);
    outputs(6364) <= not(layer2_outputs(182));
    outputs(6365) <= (layer2_outputs(2229)) xor (layer2_outputs(9061));
    outputs(6366) <= (layer2_outputs(9042)) and (layer2_outputs(5156));
    outputs(6367) <= not(layer2_outputs(2251));
    outputs(6368) <= not(layer2_outputs(4803));
    outputs(6369) <= not(layer2_outputs(6636));
    outputs(6370) <= (layer2_outputs(6960)) xor (layer2_outputs(9403));
    outputs(6371) <= (layer2_outputs(6314)) and not (layer2_outputs(8904));
    outputs(6372) <= layer2_outputs(555);
    outputs(6373) <= not((layer2_outputs(7370)) and (layer2_outputs(4700)));
    outputs(6374) <= (layer2_outputs(4910)) xor (layer2_outputs(3113));
    outputs(6375) <= layer2_outputs(3161);
    outputs(6376) <= not(layer2_outputs(4263));
    outputs(6377) <= layer2_outputs(2536);
    outputs(6378) <= not((layer2_outputs(10071)) xor (layer2_outputs(7715)));
    outputs(6379) <= not((layer2_outputs(3008)) xor (layer2_outputs(9781)));
    outputs(6380) <= layer2_outputs(3982);
    outputs(6381) <= layer2_outputs(6547);
    outputs(6382) <= (layer2_outputs(3467)) and not (layer2_outputs(9346));
    outputs(6383) <= not(layer2_outputs(3906));
    outputs(6384) <= not(layer2_outputs(2077)) or (layer2_outputs(8201));
    outputs(6385) <= layer2_outputs(2068);
    outputs(6386) <= not(layer2_outputs(2468));
    outputs(6387) <= not((layer2_outputs(2693)) xor (layer2_outputs(9293)));
    outputs(6388) <= layer2_outputs(808);
    outputs(6389) <= not((layer2_outputs(8545)) or (layer2_outputs(5384)));
    outputs(6390) <= layer2_outputs(9132);
    outputs(6391) <= not(layer2_outputs(9316));
    outputs(6392) <= layer2_outputs(2936);
    outputs(6393) <= layer2_outputs(3627);
    outputs(6394) <= not(layer2_outputs(268));
    outputs(6395) <= not(layer2_outputs(3119));
    outputs(6396) <= not(layer2_outputs(7374));
    outputs(6397) <= (layer2_outputs(6257)) xor (layer2_outputs(8272));
    outputs(6398) <= (layer2_outputs(8039)) xor (layer2_outputs(8176));
    outputs(6399) <= not(layer2_outputs(9017));
    outputs(6400) <= (layer2_outputs(896)) xor (layer2_outputs(10082));
    outputs(6401) <= not(layer2_outputs(8011));
    outputs(6402) <= not(layer2_outputs(10098));
    outputs(6403) <= not(layer2_outputs(7949));
    outputs(6404) <= not((layer2_outputs(7566)) xor (layer2_outputs(1019)));
    outputs(6405) <= layer2_outputs(3687);
    outputs(6406) <= layer2_outputs(3440);
    outputs(6407) <= layer2_outputs(8222);
    outputs(6408) <= (layer2_outputs(5026)) xor (layer2_outputs(2332));
    outputs(6409) <= not(layer2_outputs(1003));
    outputs(6410) <= layer2_outputs(3656);
    outputs(6411) <= (layer2_outputs(4412)) xor (layer2_outputs(10053));
    outputs(6412) <= not(layer2_outputs(8209));
    outputs(6413) <= (layer2_outputs(6915)) xor (layer2_outputs(8350));
    outputs(6414) <= layer2_outputs(7093);
    outputs(6415) <= layer2_outputs(994);
    outputs(6416) <= not(layer2_outputs(4584));
    outputs(6417) <= layer2_outputs(9915);
    outputs(6418) <= not(layer2_outputs(2350)) or (layer2_outputs(8788));
    outputs(6419) <= (layer2_outputs(7118)) and not (layer2_outputs(728));
    outputs(6420) <= layer2_outputs(2227);
    outputs(6421) <= layer2_outputs(7038);
    outputs(6422) <= not(layer2_outputs(1527));
    outputs(6423) <= not(layer2_outputs(2535));
    outputs(6424) <= not(layer2_outputs(8151));
    outputs(6425) <= not(layer2_outputs(2614));
    outputs(6426) <= layer2_outputs(6128);
    outputs(6427) <= layer2_outputs(5870);
    outputs(6428) <= (layer2_outputs(6246)) and (layer2_outputs(6653));
    outputs(6429) <= not((layer2_outputs(330)) or (layer2_outputs(4008)));
    outputs(6430) <= (layer2_outputs(5623)) xor (layer2_outputs(575));
    outputs(6431) <= not(layer2_outputs(3589));
    outputs(6432) <= (layer2_outputs(9678)) or (layer2_outputs(7240));
    outputs(6433) <= layer2_outputs(3276);
    outputs(6434) <= layer2_outputs(6850);
    outputs(6435) <= not(layer2_outputs(4414));
    outputs(6436) <= not(layer2_outputs(2721));
    outputs(6437) <= not(layer2_outputs(272)) or (layer2_outputs(2617));
    outputs(6438) <= not(layer2_outputs(9188));
    outputs(6439) <= not((layer2_outputs(4124)) xor (layer2_outputs(5235)));
    outputs(6440) <= not((layer2_outputs(1335)) xor (layer2_outputs(5713)));
    outputs(6441) <= layer2_outputs(789);
    outputs(6442) <= not(layer2_outputs(6383)) or (layer2_outputs(7815));
    outputs(6443) <= (layer2_outputs(4162)) and not (layer2_outputs(3688));
    outputs(6444) <= not(layer2_outputs(8448));
    outputs(6445) <= not(layer2_outputs(5658));
    outputs(6446) <= (layer2_outputs(913)) or (layer2_outputs(2574));
    outputs(6447) <= (layer2_outputs(1507)) xor (layer2_outputs(1599));
    outputs(6448) <= not(layer2_outputs(6633));
    outputs(6449) <= not(layer2_outputs(498));
    outputs(6450) <= not(layer2_outputs(1204));
    outputs(6451) <= not(layer2_outputs(2632));
    outputs(6452) <= layer2_outputs(8883);
    outputs(6453) <= not(layer2_outputs(1325));
    outputs(6454) <= not(layer2_outputs(4564));
    outputs(6455) <= not((layer2_outputs(8873)) xor (layer2_outputs(3387)));
    outputs(6456) <= not(layer2_outputs(9098));
    outputs(6457) <= not(layer2_outputs(6559));
    outputs(6458) <= not(layer2_outputs(9645));
    outputs(6459) <= not((layer2_outputs(4104)) xor (layer2_outputs(395)));
    outputs(6460) <= layer2_outputs(2011);
    outputs(6461) <= not(layer2_outputs(1943));
    outputs(6462) <= (layer2_outputs(9805)) and (layer2_outputs(9298));
    outputs(6463) <= not(layer2_outputs(6460));
    outputs(6464) <= not(layer2_outputs(10012));
    outputs(6465) <= (layer2_outputs(2791)) and (layer2_outputs(1070));
    outputs(6466) <= not(layer2_outputs(1681));
    outputs(6467) <= not(layer2_outputs(6084));
    outputs(6468) <= not(layer2_outputs(1746));
    outputs(6469) <= not((layer2_outputs(5148)) xor (layer2_outputs(8885)));
    outputs(6470) <= (layer2_outputs(6905)) xor (layer2_outputs(3888));
    outputs(6471) <= not(layer2_outputs(2464));
    outputs(6472) <= not((layer2_outputs(7909)) xor (layer2_outputs(9927)));
    outputs(6473) <= not(layer2_outputs(158));
    outputs(6474) <= not(layer2_outputs(6316));
    outputs(6475) <= not(layer2_outputs(4214));
    outputs(6476) <= not(layer2_outputs(577));
    outputs(6477) <= layer2_outputs(9573);
    outputs(6478) <= not(layer2_outputs(5737));
    outputs(6479) <= not(layer2_outputs(7559));
    outputs(6480) <= not(layer2_outputs(4789));
    outputs(6481) <= not(layer2_outputs(75));
    outputs(6482) <= layer2_outputs(7953);
    outputs(6483) <= (layer2_outputs(509)) xor (layer2_outputs(1273));
    outputs(6484) <= (layer2_outputs(6969)) xor (layer2_outputs(2316));
    outputs(6485) <= layer2_outputs(3292);
    outputs(6486) <= layer2_outputs(222);
    outputs(6487) <= layer2_outputs(1842);
    outputs(6488) <= layer2_outputs(5556);
    outputs(6489) <= layer2_outputs(941);
    outputs(6490) <= not(layer2_outputs(6062)) or (layer2_outputs(1142));
    outputs(6491) <= not(layer2_outputs(1950));
    outputs(6492) <= layer2_outputs(4006);
    outputs(6493) <= layer2_outputs(2323);
    outputs(6494) <= not(layer2_outputs(5680));
    outputs(6495) <= not(layer2_outputs(7315));
    outputs(6496) <= not(layer2_outputs(516)) or (layer2_outputs(691));
    outputs(6497) <= (layer2_outputs(6444)) and (layer2_outputs(7304));
    outputs(6498) <= not(layer2_outputs(5033));
    outputs(6499) <= layer2_outputs(3015);
    outputs(6500) <= not((layer2_outputs(915)) xor (layer2_outputs(4003)));
    outputs(6501) <= (layer2_outputs(9024)) and not (layer2_outputs(9907));
    outputs(6502) <= layer2_outputs(8849);
    outputs(6503) <= not(layer2_outputs(5336));
    outputs(6504) <= not((layer2_outputs(6269)) xor (layer2_outputs(5214)));
    outputs(6505) <= layer2_outputs(6708);
    outputs(6506) <= layer2_outputs(8458);
    outputs(6507) <= (layer2_outputs(4433)) xor (layer2_outputs(1554));
    outputs(6508) <= layer2_outputs(310);
    outputs(6509) <= (layer2_outputs(5010)) and not (layer2_outputs(7260));
    outputs(6510) <= layer2_outputs(2906);
    outputs(6511) <= layer2_outputs(3162);
    outputs(6512) <= layer2_outputs(6192);
    outputs(6513) <= not(layer2_outputs(6295));
    outputs(6514) <= not(layer2_outputs(8578));
    outputs(6515) <= layer2_outputs(7878);
    outputs(6516) <= not(layer2_outputs(9373));
    outputs(6517) <= not(layer2_outputs(7054));
    outputs(6518) <= not(layer2_outputs(6876));
    outputs(6519) <= not(layer2_outputs(3466));
    outputs(6520) <= layer2_outputs(560);
    outputs(6521) <= layer2_outputs(329);
    outputs(6522) <= not(layer2_outputs(8465));
    outputs(6523) <= not(layer2_outputs(8706));
    outputs(6524) <= not(layer2_outputs(1674));
    outputs(6525) <= (layer2_outputs(3297)) xor (layer2_outputs(6075));
    outputs(6526) <= layer2_outputs(7905);
    outputs(6527) <= not(layer2_outputs(5830));
    outputs(6528) <= not((layer2_outputs(8572)) or (layer2_outputs(5229)));
    outputs(6529) <= not(layer2_outputs(211));
    outputs(6530) <= not(layer2_outputs(2679));
    outputs(6531) <= layer2_outputs(9522);
    outputs(6532) <= not(layer2_outputs(2516));
    outputs(6533) <= layer2_outputs(8284);
    outputs(6534) <= not(layer2_outputs(2324));
    outputs(6535) <= not(layer2_outputs(3732));
    outputs(6536) <= not(layer2_outputs(3374));
    outputs(6537) <= layer2_outputs(2016);
    outputs(6538) <= not(layer2_outputs(9587));
    outputs(6539) <= layer2_outputs(7305);
    outputs(6540) <= (layer2_outputs(3594)) and not (layer2_outputs(5368));
    outputs(6541) <= not(layer2_outputs(1952));
    outputs(6542) <= layer2_outputs(4941);
    outputs(6543) <= not(layer2_outputs(2025));
    outputs(6544) <= layer2_outputs(2220);
    outputs(6545) <= (layer2_outputs(5470)) and not (layer2_outputs(2332));
    outputs(6546) <= not((layer2_outputs(3039)) and (layer2_outputs(7128)));
    outputs(6547) <= not((layer2_outputs(851)) xor (layer2_outputs(9521)));
    outputs(6548) <= not((layer2_outputs(8557)) and (layer2_outputs(9004)));
    outputs(6549) <= layer2_outputs(7825);
    outputs(6550) <= not(layer2_outputs(4416));
    outputs(6551) <= not(layer2_outputs(7156));
    outputs(6552) <= (layer2_outputs(1011)) xor (layer2_outputs(679));
    outputs(6553) <= layer2_outputs(5154);
    outputs(6554) <= layer2_outputs(627);
    outputs(6555) <= not(layer2_outputs(3842));
    outputs(6556) <= not(layer2_outputs(9034));
    outputs(6557) <= not(layer2_outputs(9897));
    outputs(6558) <= not(layer2_outputs(1915));
    outputs(6559) <= not(layer2_outputs(3077));
    outputs(6560) <= not(layer2_outputs(5889));
    outputs(6561) <= not(layer2_outputs(9808));
    outputs(6562) <= not(layer2_outputs(4132));
    outputs(6563) <= not(layer2_outputs(1047));
    outputs(6564) <= layer2_outputs(298);
    outputs(6565) <= layer2_outputs(10201);
    outputs(6566) <= layer2_outputs(757);
    outputs(6567) <= not((layer2_outputs(9747)) xor (layer2_outputs(7032)));
    outputs(6568) <= not(layer2_outputs(2729));
    outputs(6569) <= not(layer2_outputs(10046));
    outputs(6570) <= not(layer2_outputs(4098));
    outputs(6571) <= layer2_outputs(10091);
    outputs(6572) <= (layer2_outputs(6810)) xor (layer2_outputs(2307));
    outputs(6573) <= layer2_outputs(7065);
    outputs(6574) <= layer2_outputs(8229);
    outputs(6575) <= not(layer2_outputs(5864));
    outputs(6576) <= layer2_outputs(1790);
    outputs(6577) <= not((layer2_outputs(3615)) xor (layer2_outputs(1487)));
    outputs(6578) <= not(layer2_outputs(3983));
    outputs(6579) <= not(layer2_outputs(4736));
    outputs(6580) <= not(layer2_outputs(2062));
    outputs(6581) <= (layer2_outputs(4474)) xor (layer2_outputs(926));
    outputs(6582) <= layer2_outputs(4385);
    outputs(6583) <= not(layer2_outputs(4124));
    outputs(6584) <= (layer2_outputs(1409)) and (layer2_outputs(3518));
    outputs(6585) <= not(layer2_outputs(9452));
    outputs(6586) <= layer2_outputs(27);
    outputs(6587) <= layer2_outputs(7017);
    outputs(6588) <= not(layer2_outputs(3769));
    outputs(6589) <= not(layer2_outputs(2598));
    outputs(6590) <= layer2_outputs(8120);
    outputs(6591) <= not(layer2_outputs(6285));
    outputs(6592) <= layer2_outputs(1820);
    outputs(6593) <= not(layer2_outputs(811));
    outputs(6594) <= layer2_outputs(934);
    outputs(6595) <= not((layer2_outputs(4407)) xor (layer2_outputs(8096)));
    outputs(6596) <= not(layer2_outputs(5332));
    outputs(6597) <= not(layer2_outputs(286));
    outputs(6598) <= layer2_outputs(10150);
    outputs(6599) <= layer2_outputs(278);
    outputs(6600) <= not(layer2_outputs(722));
    outputs(6601) <= layer2_outputs(8357);
    outputs(6602) <= (layer2_outputs(4021)) or (layer2_outputs(1773));
    outputs(6603) <= not(layer2_outputs(381));
    outputs(6604) <= not((layer2_outputs(2272)) xor (layer2_outputs(2714)));
    outputs(6605) <= layer2_outputs(3403);
    outputs(6606) <= not(layer2_outputs(9164));
    outputs(6607) <= not(layer2_outputs(3669));
    outputs(6608) <= layer2_outputs(2551);
    outputs(6609) <= not(layer2_outputs(10217));
    outputs(6610) <= (layer2_outputs(5684)) xor (layer2_outputs(7333));
    outputs(6611) <= layer2_outputs(2920);
    outputs(6612) <= layer2_outputs(622);
    outputs(6613) <= not(layer2_outputs(9001));
    outputs(6614) <= not(layer2_outputs(1257));
    outputs(6615) <= layer2_outputs(7835);
    outputs(6616) <= not(layer2_outputs(4039));
    outputs(6617) <= layer2_outputs(2441);
    outputs(6618) <= (layer2_outputs(8620)) xor (layer2_outputs(3436));
    outputs(6619) <= not((layer2_outputs(6143)) xor (layer2_outputs(3307)));
    outputs(6620) <= layer2_outputs(6910);
    outputs(6621) <= (layer2_outputs(873)) and (layer2_outputs(7747));
    outputs(6622) <= (layer2_outputs(8066)) xor (layer2_outputs(7653));
    outputs(6623) <= layer2_outputs(2448);
    outputs(6624) <= not(layer2_outputs(2543));
    outputs(6625) <= layer2_outputs(9859);
    outputs(6626) <= layer2_outputs(5281);
    outputs(6627) <= (layer2_outputs(5305)) and (layer2_outputs(7682));
    outputs(6628) <= (layer2_outputs(6732)) and not (layer2_outputs(2858));
    outputs(6629) <= layer2_outputs(6575);
    outputs(6630) <= (layer2_outputs(525)) xor (layer2_outputs(8443));
    outputs(6631) <= layer2_outputs(8921);
    outputs(6632) <= not(layer2_outputs(3072));
    outputs(6633) <= (layer2_outputs(5185)) xor (layer2_outputs(5795));
    outputs(6634) <= not(layer2_outputs(6014));
    outputs(6635) <= (layer2_outputs(4355)) and not (layer2_outputs(7));
    outputs(6636) <= layer2_outputs(3366);
    outputs(6637) <= not(layer2_outputs(6235));
    outputs(6638) <= not(layer2_outputs(1047));
    outputs(6639) <= layer2_outputs(6373);
    outputs(6640) <= layer2_outputs(6167);
    outputs(6641) <= (layer2_outputs(8417)) and not (layer2_outputs(4711));
    outputs(6642) <= layer2_outputs(7989);
    outputs(6643) <= layer2_outputs(354);
    outputs(6644) <= layer2_outputs(2372);
    outputs(6645) <= layer2_outputs(4112);
    outputs(6646) <= layer2_outputs(1323);
    outputs(6647) <= layer2_outputs(2351);
    outputs(6648) <= layer2_outputs(5642);
    outputs(6649) <= not(layer2_outputs(10068));
    outputs(6650) <= not((layer2_outputs(9510)) xor (layer2_outputs(1206)));
    outputs(6651) <= not(layer2_outputs(2132));
    outputs(6652) <= not(layer2_outputs(6168));
    outputs(6653) <= not(layer2_outputs(8510));
    outputs(6654) <= (layer2_outputs(7600)) and (layer2_outputs(3823));
    outputs(6655) <= layer2_outputs(3684);
    outputs(6656) <= not(layer2_outputs(6710));
    outputs(6657) <= not(layer2_outputs(5102));
    outputs(6658) <= (layer2_outputs(8165)) and (layer2_outputs(10194));
    outputs(6659) <= layer2_outputs(4262);
    outputs(6660) <= not(layer2_outputs(8369));
    outputs(6661) <= layer2_outputs(4722);
    outputs(6662) <= not(layer2_outputs(5322));
    outputs(6663) <= not(layer2_outputs(9425));
    outputs(6664) <= layer2_outputs(9606);
    outputs(6665) <= layer2_outputs(3894);
    outputs(6666) <= layer2_outputs(8695);
    outputs(6667) <= layer2_outputs(3049);
    outputs(6668) <= '0';
    outputs(6669) <= layer2_outputs(1424);
    outputs(6670) <= layer2_outputs(10110);
    outputs(6671) <= not(layer2_outputs(4951));
    outputs(6672) <= not(layer2_outputs(5768));
    outputs(6673) <= layer2_outputs(2110);
    outputs(6674) <= not(layer2_outputs(10088)) or (layer2_outputs(8262));
    outputs(6675) <= (layer2_outputs(2172)) and (layer2_outputs(9895));
    outputs(6676) <= layer2_outputs(3956);
    outputs(6677) <= not(layer2_outputs(4087));
    outputs(6678) <= not((layer2_outputs(5142)) and (layer2_outputs(3718)));
    outputs(6679) <= not(layer2_outputs(3623));
    outputs(6680) <= layer2_outputs(6425);
    outputs(6681) <= not(layer2_outputs(3699));
    outputs(6682) <= not(layer2_outputs(7265));
    outputs(6683) <= not(layer2_outputs(9623));
    outputs(6684) <= not(layer2_outputs(6586));
    outputs(6685) <= not(layer2_outputs(4651));
    outputs(6686) <= not(layer2_outputs(5883));
    outputs(6687) <= not(layer2_outputs(6887));
    outputs(6688) <= not((layer2_outputs(8452)) xor (layer2_outputs(10216)));
    outputs(6689) <= not(layer2_outputs(8492));
    outputs(6690) <= not(layer2_outputs(2988));
    outputs(6691) <= not(layer2_outputs(5582));
    outputs(6692) <= not((layer2_outputs(6510)) or (layer2_outputs(6915)));
    outputs(6693) <= layer2_outputs(2710);
    outputs(6694) <= not(layer2_outputs(8783));
    outputs(6695) <= not((layer2_outputs(2336)) or (layer2_outputs(129)));
    outputs(6696) <= not(layer2_outputs(6422));
    outputs(6697) <= (layer2_outputs(1217)) and not (layer2_outputs(9143));
    outputs(6698) <= not((layer2_outputs(4431)) or (layer2_outputs(9332)));
    outputs(6699) <= (layer2_outputs(3037)) and (layer2_outputs(2950));
    outputs(6700) <= layer2_outputs(4163);
    outputs(6701) <= not((layer2_outputs(1711)) or (layer2_outputs(933)));
    outputs(6702) <= not(layer2_outputs(9788));
    outputs(6703) <= layer2_outputs(3271);
    outputs(6704) <= layer2_outputs(88);
    outputs(6705) <= not(layer2_outputs(6343));
    outputs(6706) <= layer2_outputs(4804);
    outputs(6707) <= not(layer2_outputs(441));
    outputs(6708) <= layer2_outputs(3630);
    outputs(6709) <= not(layer2_outputs(1272));
    outputs(6710) <= not(layer2_outputs(10012));
    outputs(6711) <= layer2_outputs(8616);
    outputs(6712) <= not((layer2_outputs(4213)) or (layer2_outputs(9999)));
    outputs(6713) <= layer2_outputs(8897);
    outputs(6714) <= layer2_outputs(9192);
    outputs(6715) <= layer2_outputs(10226);
    outputs(6716) <= layer2_outputs(1654);
    outputs(6717) <= layer2_outputs(9048);
    outputs(6718) <= not(layer2_outputs(907));
    outputs(6719) <= layer2_outputs(4881);
    outputs(6720) <= not(layer2_outputs(10015));
    outputs(6721) <= layer2_outputs(2091);
    outputs(6722) <= not(layer2_outputs(1956));
    outputs(6723) <= layer2_outputs(9390);
    outputs(6724) <= not(layer2_outputs(7317));
    outputs(6725) <= (layer2_outputs(5357)) xor (layer2_outputs(8981));
    outputs(6726) <= (layer2_outputs(6232)) and not (layer2_outputs(7936));
    outputs(6727) <= layer2_outputs(3451);
    outputs(6728) <= (layer2_outputs(3254)) xor (layer2_outputs(10027));
    outputs(6729) <= layer2_outputs(9405);
    outputs(6730) <= not(layer2_outputs(6004));
    outputs(6731) <= not(layer2_outputs(2619));
    outputs(6732) <= layer2_outputs(5076);
    outputs(6733) <= (layer2_outputs(6989)) and not (layer2_outputs(2151));
    outputs(6734) <= not((layer2_outputs(8026)) xor (layer2_outputs(7861)));
    outputs(6735) <= not(layer2_outputs(5740));
    outputs(6736) <= layer2_outputs(1486);
    outputs(6737) <= not(layer2_outputs(4767));
    outputs(6738) <= (layer2_outputs(566)) and not (layer2_outputs(6626));
    outputs(6739) <= layer2_outputs(2783);
    outputs(6740) <= not(layer2_outputs(1985));
    outputs(6741) <= layer2_outputs(1827);
    outputs(6742) <= not(layer2_outputs(1671));
    outputs(6743) <= layer2_outputs(106);
    outputs(6744) <= layer2_outputs(3738);
    outputs(6745) <= layer2_outputs(7461);
    outputs(6746) <= not(layer2_outputs(4538));
    outputs(6747) <= layer2_outputs(2444);
    outputs(6748) <= layer2_outputs(1685);
    outputs(6749) <= not(layer2_outputs(7247));
    outputs(6750) <= layer2_outputs(2223);
    outputs(6751) <= layer2_outputs(583);
    outputs(6752) <= not(layer2_outputs(7180));
    outputs(6753) <= not(layer2_outputs(2576));
    outputs(6754) <= not(layer2_outputs(1014));
    outputs(6755) <= (layer2_outputs(4864)) and not (layer2_outputs(2832));
    outputs(6756) <= layer2_outputs(4242);
    outputs(6757) <= not(layer2_outputs(5339));
    outputs(6758) <= not(layer2_outputs(4914));
    outputs(6759) <= layer2_outputs(8323);
    outputs(6760) <= layer2_outputs(6008);
    outputs(6761) <= not(layer2_outputs(4858));
    outputs(6762) <= layer2_outputs(6582);
    outputs(6763) <= layer2_outputs(7853);
    outputs(6764) <= not(layer2_outputs(6824));
    outputs(6765) <= not(layer2_outputs(4888));
    outputs(6766) <= not(layer2_outputs(6994));
    outputs(6767) <= not(layer2_outputs(1653));
    outputs(6768) <= layer2_outputs(53);
    outputs(6769) <= not(layer2_outputs(8364));
    outputs(6770) <= layer2_outputs(8872);
    outputs(6771) <= layer2_outputs(10020);
    outputs(6772) <= layer2_outputs(9319);
    outputs(6773) <= not(layer2_outputs(9203));
    outputs(6774) <= not(layer2_outputs(5587));
    outputs(6775) <= not(layer2_outputs(6689));
    outputs(6776) <= not(layer2_outputs(865));
    outputs(6777) <= not(layer2_outputs(5491)) or (layer2_outputs(2959));
    outputs(6778) <= not(layer2_outputs(9271));
    outputs(6779) <= layer2_outputs(4463);
    outputs(6780) <= layer2_outputs(1874);
    outputs(6781) <= not(layer2_outputs(7993));
    outputs(6782) <= not(layer2_outputs(4788));
    outputs(6783) <= layer2_outputs(4527);
    outputs(6784) <= layer2_outputs(2513);
    outputs(6785) <= (layer2_outputs(4971)) and not (layer2_outputs(319));
    outputs(6786) <= not(layer2_outputs(7066));
    outputs(6787) <= layer2_outputs(3488);
    outputs(6788) <= layer2_outputs(6539);
    outputs(6789) <= not((layer2_outputs(1304)) and (layer2_outputs(1368)));
    outputs(6790) <= not((layer2_outputs(698)) xor (layer2_outputs(6097)));
    outputs(6791) <= not((layer2_outputs(10027)) xor (layer2_outputs(10155)));
    outputs(6792) <= layer2_outputs(6130);
    outputs(6793) <= (layer2_outputs(596)) xor (layer2_outputs(7685));
    outputs(6794) <= (layer2_outputs(8245)) and (layer2_outputs(7176));
    outputs(6795) <= not(layer2_outputs(10139));
    outputs(6796) <= not(layer2_outputs(6599));
    outputs(6797) <= not(layer2_outputs(4571));
    outputs(6798) <= not(layer2_outputs(3268));
    outputs(6799) <= (layer2_outputs(8389)) and not (layer2_outputs(9930));
    outputs(6800) <= not(layer2_outputs(2898)) or (layer2_outputs(5871));
    outputs(6801) <= not(layer2_outputs(6697));
    outputs(6802) <= layer2_outputs(1904);
    outputs(6803) <= not(layer2_outputs(6457));
    outputs(6804) <= (layer2_outputs(6034)) xor (layer2_outputs(7108));
    outputs(6805) <= (layer2_outputs(9347)) and not (layer2_outputs(7958));
    outputs(6806) <= not((layer2_outputs(1938)) xor (layer2_outputs(7533)));
    outputs(6807) <= layer2_outputs(333);
    outputs(6808) <= not(layer2_outputs(6445));
    outputs(6809) <= not((layer2_outputs(1223)) xor (layer2_outputs(6347)));
    outputs(6810) <= not(layer2_outputs(2187));
    outputs(6811) <= not(layer2_outputs(4732));
    outputs(6812) <= not(layer2_outputs(1118));
    outputs(6813) <= not(layer2_outputs(3900));
    outputs(6814) <= not(layer2_outputs(9692));
    outputs(6815) <= not(layer2_outputs(2811));
    outputs(6816) <= layer2_outputs(5397);
    outputs(6817) <= not(layer2_outputs(5303)) or (layer2_outputs(1576));
    outputs(6818) <= layer2_outputs(3599);
    outputs(6819) <= not(layer2_outputs(4939));
    outputs(6820) <= layer2_outputs(5528);
    outputs(6821) <= layer2_outputs(1971);
    outputs(6822) <= not(layer2_outputs(4831)) or (layer2_outputs(2958));
    outputs(6823) <= not(layer2_outputs(213));
    outputs(6824) <= layer2_outputs(1101);
    outputs(6825) <= not(layer2_outputs(3770));
    outputs(6826) <= layer2_outputs(7072);
    outputs(6827) <= layer2_outputs(3804);
    outputs(6828) <= not(layer2_outputs(2112));
    outputs(6829) <= (layer2_outputs(9985)) and (layer2_outputs(5253));
    outputs(6830) <= layer2_outputs(6726);
    outputs(6831) <= (layer2_outputs(3736)) and not (layer2_outputs(1279));
    outputs(6832) <= layer2_outputs(4269);
    outputs(6833) <= not(layer2_outputs(2062));
    outputs(6834) <= layer2_outputs(3481);
    outputs(6835) <= layer2_outputs(8372);
    outputs(6836) <= layer2_outputs(1879);
    outputs(6837) <= not((layer2_outputs(36)) xor (layer2_outputs(6031)));
    outputs(6838) <= not(layer2_outputs(2502));
    outputs(6839) <= not(layer2_outputs(7275));
    outputs(6840) <= layer2_outputs(93);
    outputs(6841) <= (layer2_outputs(1935)) xor (layer2_outputs(4613));
    outputs(6842) <= layer2_outputs(5584);
    outputs(6843) <= not(layer2_outputs(9021));
    outputs(6844) <= layer2_outputs(8372);
    outputs(6845) <= layer2_outputs(2905);
    outputs(6846) <= not(layer2_outputs(8280));
    outputs(6847) <= layer2_outputs(4035);
    outputs(6848) <= not(layer2_outputs(9812));
    outputs(6849) <= not(layer2_outputs(4165));
    outputs(6850) <= not(layer2_outputs(1214));
    outputs(6851) <= not((layer2_outputs(9946)) or (layer2_outputs(6506)));
    outputs(6852) <= layer2_outputs(2209);
    outputs(6853) <= layer2_outputs(8883);
    outputs(6854) <= not(layer2_outputs(5240));
    outputs(6855) <= not(layer2_outputs(1851));
    outputs(6856) <= not(layer2_outputs(5777));
    outputs(6857) <= not(layer2_outputs(4250));
    outputs(6858) <= not((layer2_outputs(6522)) xor (layer2_outputs(5499)));
    outputs(6859) <= layer2_outputs(10181);
    outputs(6860) <= layer2_outputs(2136);
    outputs(6861) <= layer2_outputs(464);
    outputs(6862) <= not(layer2_outputs(1803));
    outputs(6863) <= not((layer2_outputs(3585)) xor (layer2_outputs(5018)));
    outputs(6864) <= not(layer2_outputs(8385));
    outputs(6865) <= not(layer2_outputs(9946));
    outputs(6866) <= not(layer2_outputs(1656));
    outputs(6867) <= layer2_outputs(5333);
    outputs(6868) <= layer2_outputs(3599);
    outputs(6869) <= layer2_outputs(7900);
    outputs(6870) <= not(layer2_outputs(5228));
    outputs(6871) <= layer2_outputs(9977);
    outputs(6872) <= layer2_outputs(6392);
    outputs(6873) <= not(layer2_outputs(2419));
    outputs(6874) <= not(layer2_outputs(6063));
    outputs(6875) <= layer2_outputs(5311);
    outputs(6876) <= layer2_outputs(4369);
    outputs(6877) <= not(layer2_outputs(7811));
    outputs(6878) <= not(layer2_outputs(3819));
    outputs(6879) <= layer2_outputs(8143);
    outputs(6880) <= layer2_outputs(1385);
    outputs(6881) <= layer2_outputs(8430);
    outputs(6882) <= not(layer2_outputs(5320));
    outputs(6883) <= not((layer2_outputs(8934)) xor (layer2_outputs(8514)));
    outputs(6884) <= (layer2_outputs(4867)) or (layer2_outputs(9738));
    outputs(6885) <= not(layer2_outputs(2096));
    outputs(6886) <= not((layer2_outputs(2440)) xor (layer2_outputs(3825)));
    outputs(6887) <= (layer2_outputs(5665)) xor (layer2_outputs(9262));
    outputs(6888) <= not((layer2_outputs(7400)) or (layer2_outputs(1144)));
    outputs(6889) <= layer2_outputs(2237);
    outputs(6890) <= layer2_outputs(8911);
    outputs(6891) <= not(layer2_outputs(9996));
    outputs(6892) <= (layer2_outputs(7185)) xor (layer2_outputs(9313));
    outputs(6893) <= layer2_outputs(2500);
    outputs(6894) <= layer2_outputs(982);
    outputs(6895) <= not(layer2_outputs(8318));
    outputs(6896) <= layer2_outputs(1246);
    outputs(6897) <= layer2_outputs(1474);
    outputs(6898) <= not(layer2_outputs(7502));
    outputs(6899) <= layer2_outputs(8383);
    outputs(6900) <= not(layer2_outputs(2842)) or (layer2_outputs(2821));
    outputs(6901) <= not(layer2_outputs(6793));
    outputs(6902) <= layer2_outputs(8616);
    outputs(6903) <= not(layer2_outputs(3692));
    outputs(6904) <= not(layer2_outputs(6740));
    outputs(6905) <= layer2_outputs(7295);
    outputs(6906) <= (layer2_outputs(452)) or (layer2_outputs(5505));
    outputs(6907) <= not((layer2_outputs(2317)) and (layer2_outputs(4408)));
    outputs(6908) <= not(layer2_outputs(3759));
    outputs(6909) <= not(layer2_outputs(1509));
    outputs(6910) <= not((layer2_outputs(1730)) xor (layer2_outputs(10146)));
    outputs(6911) <= (layer2_outputs(8746)) and (layer2_outputs(1475));
    outputs(6912) <= not(layer2_outputs(2935)) or (layer2_outputs(5290));
    outputs(6913) <= not((layer2_outputs(7950)) xor (layer2_outputs(1079)));
    outputs(6914) <= not(layer2_outputs(7117));
    outputs(6915) <= layer2_outputs(8633);
    outputs(6916) <= (layer2_outputs(8746)) and not (layer2_outputs(1069));
    outputs(6917) <= layer2_outputs(260);
    outputs(6918) <= layer2_outputs(5845);
    outputs(6919) <= not(layer2_outputs(3770));
    outputs(6920) <= not(layer2_outputs(6423));
    outputs(6921) <= not(layer2_outputs(883));
    outputs(6922) <= layer2_outputs(2541);
    outputs(6923) <= not(layer2_outputs(5542)) or (layer2_outputs(6738));
    outputs(6924) <= (layer2_outputs(2054)) xor (layer2_outputs(1090));
    outputs(6925) <= layer2_outputs(3540);
    outputs(6926) <= layer2_outputs(2962);
    outputs(6927) <= not(layer2_outputs(4473));
    outputs(6928) <= (layer2_outputs(2102)) and not (layer2_outputs(172));
    outputs(6929) <= (layer2_outputs(1076)) xor (layer2_outputs(9051));
    outputs(6930) <= not(layer2_outputs(5123));
    outputs(6931) <= (layer2_outputs(10161)) xor (layer2_outputs(8938));
    outputs(6932) <= layer2_outputs(2111);
    outputs(6933) <= (layer2_outputs(4690)) and not (layer2_outputs(4497));
    outputs(6934) <= not(layer2_outputs(64));
    outputs(6935) <= layer2_outputs(1149);
    outputs(6936) <= layer2_outputs(3432);
    outputs(6937) <= layer2_outputs(3728);
    outputs(6938) <= not(layer2_outputs(8325));
    outputs(6939) <= layer2_outputs(5462);
    outputs(6940) <= layer2_outputs(8963);
    outputs(6941) <= layer2_outputs(3045);
    outputs(6942) <= not(layer2_outputs(5837));
    outputs(6943) <= not(layer2_outputs(1219));
    outputs(6944) <= layer2_outputs(2762);
    outputs(6945) <= not(layer2_outputs(2250));
    outputs(6946) <= (layer2_outputs(4847)) xor (layer2_outputs(612));
    outputs(6947) <= not(layer2_outputs(6849));
    outputs(6948) <= (layer2_outputs(2881)) and not (layer2_outputs(7754));
    outputs(6949) <= not(layer2_outputs(1527));
    outputs(6950) <= not(layer2_outputs(3119));
    outputs(6951) <= not(layer2_outputs(5175));
    outputs(6952) <= layer2_outputs(8717);
    outputs(6953) <= not(layer2_outputs(1327));
    outputs(6954) <= not(layer2_outputs(6282)) or (layer2_outputs(3564));
    outputs(6955) <= (layer2_outputs(9903)) and not (layer2_outputs(3175));
    outputs(6956) <= layer2_outputs(6488);
    outputs(6957) <= (layer2_outputs(754)) xor (layer2_outputs(1398));
    outputs(6958) <= layer2_outputs(6990);
    outputs(6959) <= layer2_outputs(8356);
    outputs(6960) <= layer2_outputs(8463);
    outputs(6961) <= layer2_outputs(5982);
    outputs(6962) <= layer2_outputs(10);
    outputs(6963) <= layer2_outputs(9015);
    outputs(6964) <= layer2_outputs(3042);
    outputs(6965) <= (layer2_outputs(1282)) or (layer2_outputs(1235));
    outputs(6966) <= not(layer2_outputs(6221));
    outputs(6967) <= layer2_outputs(8213);
    outputs(6968) <= (layer2_outputs(7548)) and not (layer2_outputs(6244));
    outputs(6969) <= layer2_outputs(822);
    outputs(6970) <= not(layer2_outputs(9518));
    outputs(6971) <= (layer2_outputs(6872)) and (layer2_outputs(8044));
    outputs(6972) <= not(layer2_outputs(5176));
    outputs(6973) <= layer2_outputs(3733);
    outputs(6974) <= (layer2_outputs(872)) and (layer2_outputs(3851));
    outputs(6975) <= layer2_outputs(1253);
    outputs(6976) <= not(layer2_outputs(9413));
    outputs(6977) <= layer2_outputs(2816);
    outputs(6978) <= layer2_outputs(3970);
    outputs(6979) <= layer2_outputs(4802);
    outputs(6980) <= layer2_outputs(1615);
    outputs(6981) <= not(layer2_outputs(4481));
    outputs(6982) <= not(layer2_outputs(798));
    outputs(6983) <= not((layer2_outputs(5135)) or (layer2_outputs(8036)));
    outputs(6984) <= not(layer2_outputs(9684));
    outputs(6985) <= not((layer2_outputs(1815)) xor (layer2_outputs(3984)));
    outputs(6986) <= not((layer2_outputs(9904)) or (layer2_outputs(6616)));
    outputs(6987) <= not(layer2_outputs(10054));
    outputs(6988) <= not(layer2_outputs(6851));
    outputs(6989) <= layer2_outputs(6701);
    outputs(6990) <= not((layer2_outputs(5702)) and (layer2_outputs(6924)));
    outputs(6991) <= layer2_outputs(1478);
    outputs(6992) <= (layer2_outputs(9186)) and (layer2_outputs(9915));
    outputs(6993) <= not(layer2_outputs(9804));
    outputs(6994) <= layer2_outputs(9548);
    outputs(6995) <= layer2_outputs(7489);
    outputs(6996) <= (layer2_outputs(6178)) xor (layer2_outputs(3478));
    outputs(6997) <= not(layer2_outputs(2490));
    outputs(6998) <= not(layer2_outputs(5408)) or (layer2_outputs(7897));
    outputs(6999) <= not(layer2_outputs(8974));
    outputs(7000) <= not(layer2_outputs(2612));
    outputs(7001) <= layer2_outputs(5867);
    outputs(7002) <= layer2_outputs(2340);
    outputs(7003) <= layer2_outputs(7576);
    outputs(7004) <= not(layer2_outputs(8745));
    outputs(7005) <= not(layer2_outputs(6883));
    outputs(7006) <= layer2_outputs(5530);
    outputs(7007) <= layer2_outputs(8570);
    outputs(7008) <= layer2_outputs(4183);
    outputs(7009) <= not(layer2_outputs(7584));
    outputs(7010) <= not(layer2_outputs(6540));
    outputs(7011) <= layer2_outputs(989);
    outputs(7012) <= (layer2_outputs(7524)) and not (layer2_outputs(5056));
    outputs(7013) <= not(layer2_outputs(5085));
    outputs(7014) <= not(layer2_outputs(7255));
    outputs(7015) <= not(layer2_outputs(6668));
    outputs(7016) <= not(layer2_outputs(10048));
    outputs(7017) <= not((layer2_outputs(6026)) xor (layer2_outputs(2918)));
    outputs(7018) <= layer2_outputs(1330);
    outputs(7019) <= not(layer2_outputs(351));
    outputs(7020) <= not(layer2_outputs(4198)) or (layer2_outputs(4689));
    outputs(7021) <= layer2_outputs(1016);
    outputs(7022) <= layer2_outputs(3186);
    outputs(7023) <= layer2_outputs(4402);
    outputs(7024) <= not(layer2_outputs(9561));
    outputs(7025) <= (layer2_outputs(2694)) and (layer2_outputs(7912));
    outputs(7026) <= not((layer2_outputs(1525)) xor (layer2_outputs(3753)));
    outputs(7027) <= layer2_outputs(6076);
    outputs(7028) <= (layer2_outputs(2182)) and not (layer2_outputs(8900));
    outputs(7029) <= layer2_outputs(9709);
    outputs(7030) <= not(layer2_outputs(6497)) or (layer2_outputs(8838));
    outputs(7031) <= not(layer2_outputs(1746)) or (layer2_outputs(8313));
    outputs(7032) <= not(layer2_outputs(9182));
    outputs(7033) <= not(layer2_outputs(1185)) or (layer2_outputs(4042));
    outputs(7034) <= layer2_outputs(4587);
    outputs(7035) <= not(layer2_outputs(9814));
    outputs(7036) <= not(layer2_outputs(508));
    outputs(7037) <= not(layer2_outputs(217));
    outputs(7038) <= layer2_outputs(4488);
    outputs(7039) <= (layer2_outputs(5538)) xor (layer2_outputs(3414));
    outputs(7040) <= not((layer2_outputs(3536)) or (layer2_outputs(6490)));
    outputs(7041) <= layer2_outputs(6464);
    outputs(7042) <= not(layer2_outputs(7593));
    outputs(7043) <= layer2_outputs(8525);
    outputs(7044) <= layer2_outputs(853);
    outputs(7045) <= (layer2_outputs(9902)) xor (layer2_outputs(8619));
    outputs(7046) <= not(layer2_outputs(4609)) or (layer2_outputs(7971));
    outputs(7047) <= not((layer2_outputs(2585)) xor (layer2_outputs(701)));
    outputs(7048) <= (layer2_outputs(6984)) xor (layer2_outputs(1735));
    outputs(7049) <= not(layer2_outputs(4817));
    outputs(7050) <= not((layer2_outputs(9202)) xor (layer2_outputs(5432)));
    outputs(7051) <= not(layer2_outputs(9350));
    outputs(7052) <= layer2_outputs(685);
    outputs(7053) <= not(layer2_outputs(2887));
    outputs(7054) <= not((layer2_outputs(4469)) or (layer2_outputs(1791)));
    outputs(7055) <= layer2_outputs(4887);
    outputs(7056) <= not((layer2_outputs(9258)) and (layer2_outputs(57)));
    outputs(7057) <= layer2_outputs(4049);
    outputs(7058) <= not(layer2_outputs(2378));
    outputs(7059) <= not(layer2_outputs(9470)) or (layer2_outputs(2845));
    outputs(7060) <= not(layer2_outputs(8644)) or (layer2_outputs(9576));
    outputs(7061) <= (layer2_outputs(5611)) and not (layer2_outputs(7039));
    outputs(7062) <= layer2_outputs(2398);
    outputs(7063) <= not(layer2_outputs(9218));
    outputs(7064) <= not(layer2_outputs(2637));
    outputs(7065) <= layer2_outputs(3574);
    outputs(7066) <= (layer2_outputs(4265)) and not (layer2_outputs(3085));
    outputs(7067) <= layer2_outputs(7437);
    outputs(7068) <= not(layer2_outputs(3140));
    outputs(7069) <= not(layer2_outputs(9375));
    outputs(7070) <= layer2_outputs(2978);
    outputs(7071) <= not(layer2_outputs(1608));
    outputs(7072) <= layer2_outputs(2060);
    outputs(7073) <= (layer2_outputs(6212)) xor (layer2_outputs(1254));
    outputs(7074) <= layer2_outputs(5905);
    outputs(7075) <= not((layer2_outputs(385)) and (layer2_outputs(8154)));
    outputs(7076) <= layer2_outputs(4738);
    outputs(7077) <= not((layer2_outputs(3550)) or (layer2_outputs(2343)));
    outputs(7078) <= not(layer2_outputs(6994));
    outputs(7079) <= not(layer2_outputs(7088));
    outputs(7080) <= layer2_outputs(1505);
    outputs(7081) <= layer2_outputs(3069);
    outputs(7082) <= layer2_outputs(1723);
    outputs(7083) <= layer2_outputs(8435);
    outputs(7084) <= not((layer2_outputs(7441)) and (layer2_outputs(10158)));
    outputs(7085) <= layer2_outputs(4444);
    outputs(7086) <= not(layer2_outputs(7569));
    outputs(7087) <= layer2_outputs(6761);
    outputs(7088) <= (layer2_outputs(8574)) xor (layer2_outputs(3029));
    outputs(7089) <= not(layer2_outputs(1133));
    outputs(7090) <= layer2_outputs(3873);
    outputs(7091) <= layer2_outputs(7233);
    outputs(7092) <= layer2_outputs(8159);
    outputs(7093) <= not(layer2_outputs(426));
    outputs(7094) <= layer2_outputs(5551);
    outputs(7095) <= not((layer2_outputs(677)) xor (layer2_outputs(4671)));
    outputs(7096) <= layer2_outputs(5691);
    outputs(7097) <= not(layer2_outputs(2599));
    outputs(7098) <= layer2_outputs(8303);
    outputs(7099) <= not(layer2_outputs(8297));
    outputs(7100) <= layer2_outputs(5564);
    outputs(7101) <= not(layer2_outputs(9438));
    outputs(7102) <= not(layer2_outputs(7169));
    outputs(7103) <= layer2_outputs(2052);
    outputs(7104) <= not((layer2_outputs(7547)) and (layer2_outputs(6435)));
    outputs(7105) <= layer2_outputs(9119);
    outputs(7106) <= layer2_outputs(2762);
    outputs(7107) <= not((layer2_outputs(9128)) or (layer2_outputs(4316)));
    outputs(7108) <= layer2_outputs(2269);
    outputs(7109) <= not(layer2_outputs(1248));
    outputs(7110) <= layer2_outputs(685);
    outputs(7111) <= not(layer2_outputs(4809));
    outputs(7112) <= (layer2_outputs(59)) xor (layer2_outputs(4942));
    outputs(7113) <= layer2_outputs(7124);
    outputs(7114) <= layer2_outputs(8460);
    outputs(7115) <= not(layer2_outputs(3742));
    outputs(7116) <= not(layer2_outputs(1948));
    outputs(7117) <= not(layer2_outputs(5189));
    outputs(7118) <= (layer2_outputs(3710)) and not (layer2_outputs(6964));
    outputs(7119) <= layer2_outputs(9315);
    outputs(7120) <= not((layer2_outputs(7269)) or (layer2_outputs(4766)));
    outputs(7121) <= (layer2_outputs(5868)) xor (layer2_outputs(7671));
    outputs(7122) <= (layer2_outputs(9659)) and not (layer2_outputs(815));
    outputs(7123) <= not(layer2_outputs(1353));
    outputs(7124) <= layer2_outputs(5397);
    outputs(7125) <= layer2_outputs(2233);
    outputs(7126) <= not(layer2_outputs(176));
    outputs(7127) <= (layer2_outputs(3398)) xor (layer2_outputs(8739));
    outputs(7128) <= not(layer2_outputs(1270)) or (layer2_outputs(2501));
    outputs(7129) <= not(layer2_outputs(3016));
    outputs(7130) <= layer2_outputs(842);
    outputs(7131) <= not(layer2_outputs(4917)) or (layer2_outputs(10196));
    outputs(7132) <= layer2_outputs(5256);
    outputs(7133) <= not(layer2_outputs(626));
    outputs(7134) <= layer2_outputs(3785);
    outputs(7135) <= layer2_outputs(2045);
    outputs(7136) <= layer2_outputs(3386);
    outputs(7137) <= layer2_outputs(4168);
    outputs(7138) <= not(layer2_outputs(5715));
    outputs(7139) <= layer2_outputs(5914);
    outputs(7140) <= not(layer2_outputs(5668));
    outputs(7141) <= not(layer2_outputs(5779));
    outputs(7142) <= layer2_outputs(799);
    outputs(7143) <= layer2_outputs(9791);
    outputs(7144) <= (layer2_outputs(6835)) xor (layer2_outputs(1268));
    outputs(7145) <= layer2_outputs(466);
    outputs(7146) <= (layer2_outputs(4612)) and not (layer2_outputs(1283));
    outputs(7147) <= layer2_outputs(6076);
    outputs(7148) <= layer2_outputs(9581);
    outputs(7149) <= not(layer2_outputs(9730));
    outputs(7150) <= layer2_outputs(5568);
    outputs(7151) <= (layer2_outputs(1618)) xor (layer2_outputs(9709));
    outputs(7152) <= not((layer2_outputs(209)) xor (layer2_outputs(2201)));
    outputs(7153) <= layer2_outputs(421);
    outputs(7154) <= not(layer2_outputs(6113));
    outputs(7155) <= layer2_outputs(9335);
    outputs(7156) <= layer2_outputs(2921);
    outputs(7157) <= not(layer2_outputs(2619));
    outputs(7158) <= layer2_outputs(6075);
    outputs(7159) <= layer2_outputs(2653);
    outputs(7160) <= not((layer2_outputs(3169)) or (layer2_outputs(9436)));
    outputs(7161) <= layer2_outputs(5001);
    outputs(7162) <= (layer2_outputs(4714)) xor (layer2_outputs(3659));
    outputs(7163) <= not(layer2_outputs(1945));
    outputs(7164) <= not(layer2_outputs(5896));
    outputs(7165) <= layer2_outputs(3123);
    outputs(7166) <= not(layer2_outputs(6315));
    outputs(7167) <= layer2_outputs(9540);
    outputs(7168) <= layer2_outputs(5098);
    outputs(7169) <= not((layer2_outputs(7059)) xor (layer2_outputs(3105)));
    outputs(7170) <= layer2_outputs(5430);
    outputs(7171) <= (layer2_outputs(3146)) and not (layer2_outputs(3132));
    outputs(7172) <= not(layer2_outputs(1502));
    outputs(7173) <= not(layer2_outputs(466)) or (layer2_outputs(4879));
    outputs(7174) <= (layer2_outputs(9409)) and not (layer2_outputs(2444));
    outputs(7175) <= layer2_outputs(5370);
    outputs(7176) <= (layer2_outputs(5404)) and (layer2_outputs(2843));
    outputs(7177) <= (layer2_outputs(4135)) and not (layer2_outputs(1049));
    outputs(7178) <= layer2_outputs(3048);
    outputs(7179) <= layer2_outputs(2606);
    outputs(7180) <= not(layer2_outputs(7946));
    outputs(7181) <= layer2_outputs(5224);
    outputs(7182) <= layer2_outputs(3462);
    outputs(7183) <= layer2_outputs(8035);
    outputs(7184) <= not(layer2_outputs(6743));
    outputs(7185) <= layer2_outputs(9919);
    outputs(7186) <= not(layer2_outputs(5881));
    outputs(7187) <= not(layer2_outputs(6686));
    outputs(7188) <= not(layer2_outputs(8805));
    outputs(7189) <= not(layer2_outputs(7914));
    outputs(7190) <= (layer2_outputs(2094)) xor (layer2_outputs(6564));
    outputs(7191) <= not(layer2_outputs(4369));
    outputs(7192) <= not(layer2_outputs(7389));
    outputs(7193) <= layer2_outputs(3838);
    outputs(7194) <= layer2_outputs(7949);
    outputs(7195) <= layer2_outputs(5293);
    outputs(7196) <= not(layer2_outputs(6263));
    outputs(7197) <= not((layer2_outputs(126)) xor (layer2_outputs(1238)));
    outputs(7198) <= (layer2_outputs(6214)) xor (layer2_outputs(3882));
    outputs(7199) <= not(layer2_outputs(326));
    outputs(7200) <= layer2_outputs(378);
    outputs(7201) <= (layer2_outputs(1154)) and not (layer2_outputs(7999));
    outputs(7202) <= (layer2_outputs(7893)) and (layer2_outputs(5237));
    outputs(7203) <= layer2_outputs(5786);
    outputs(7204) <= not(layer2_outputs(3944));
    outputs(7205) <= not(layer2_outputs(1601));
    outputs(7206) <= not(layer2_outputs(3575));
    outputs(7207) <= (layer2_outputs(2859)) xor (layer2_outputs(3107));
    outputs(7208) <= layer2_outputs(1693);
    outputs(7209) <= not(layer2_outputs(6872));
    outputs(7210) <= not(layer2_outputs(9262));
    outputs(7211) <= layer2_outputs(8558);
    outputs(7212) <= layer2_outputs(409);
    outputs(7213) <= not(layer2_outputs(5139));
    outputs(7214) <= not((layer2_outputs(1124)) xor (layer2_outputs(4987)));
    outputs(7215) <= layer2_outputs(1490);
    outputs(7216) <= layer2_outputs(6005);
    outputs(7217) <= layer2_outputs(9539);
    outputs(7218) <= not(layer2_outputs(6411));
    outputs(7219) <= layer2_outputs(4768);
    outputs(7220) <= layer2_outputs(9220);
    outputs(7221) <= layer2_outputs(536);
    outputs(7222) <= layer2_outputs(4972);
    outputs(7223) <= layer2_outputs(5353);
    outputs(7224) <= not(layer2_outputs(4173));
    outputs(7225) <= not((layer2_outputs(4406)) and (layer2_outputs(1244)));
    outputs(7226) <= layer2_outputs(3789);
    outputs(7227) <= layer2_outputs(9333);
    outputs(7228) <= (layer2_outputs(6412)) and (layer2_outputs(5900));
    outputs(7229) <= not((layer2_outputs(6403)) or (layer2_outputs(5280)));
    outputs(7230) <= layer2_outputs(3638);
    outputs(7231) <= not(layer2_outputs(8723));
    outputs(7232) <= layer2_outputs(6678);
    outputs(7233) <= not(layer2_outputs(8220));
    outputs(7234) <= not(layer2_outputs(6587));
    outputs(7235) <= not(layer2_outputs(2853));
    outputs(7236) <= (layer2_outputs(342)) and (layer2_outputs(9188));
    outputs(7237) <= not((layer2_outputs(878)) xor (layer2_outputs(3078)));
    outputs(7238) <= not((layer2_outputs(9138)) xor (layer2_outputs(954)));
    outputs(7239) <= not((layer2_outputs(5767)) xor (layer2_outputs(4012)));
    outputs(7240) <= not(layer2_outputs(9833));
    outputs(7241) <= not(layer2_outputs(9125)) or (layer2_outputs(8542));
    outputs(7242) <= not((layer2_outputs(8928)) or (layer2_outputs(7069)));
    outputs(7243) <= not(layer2_outputs(5334));
    outputs(7244) <= not(layer2_outputs(9532));
    outputs(7245) <= layer2_outputs(8736);
    outputs(7246) <= not(layer2_outputs(8237));
    outputs(7247) <= (layer2_outputs(3732)) and (layer2_outputs(2848));
    outputs(7248) <= layer2_outputs(9152);
    outputs(7249) <= (layer2_outputs(7010)) xor (layer2_outputs(9826));
    outputs(7250) <= not(layer2_outputs(9745));
    outputs(7251) <= (layer2_outputs(903)) xor (layer2_outputs(6592));
    outputs(7252) <= layer2_outputs(5983);
    outputs(7253) <= not(layer2_outputs(45));
    outputs(7254) <= layer2_outputs(7681);
    outputs(7255) <= not(layer2_outputs(9584));
    outputs(7256) <= (layer2_outputs(7925)) and not (layer2_outputs(6323));
    outputs(7257) <= layer2_outputs(7569);
    outputs(7258) <= (layer2_outputs(9217)) xor (layer2_outputs(742));
    outputs(7259) <= layer2_outputs(7282);
    outputs(7260) <= not((layer2_outputs(7998)) xor (layer2_outputs(3577)));
    outputs(7261) <= layer2_outputs(9892);
    outputs(7262) <= layer2_outputs(5578);
    outputs(7263) <= layer2_outputs(6860);
    outputs(7264) <= not(layer2_outputs(3269));
    outputs(7265) <= not(layer2_outputs(5014));
    outputs(7266) <= not(layer2_outputs(6029));
    outputs(7267) <= not(layer2_outputs(8401));
    outputs(7268) <= not(layer2_outputs(4753));
    outputs(7269) <= (layer2_outputs(1889)) or (layer2_outputs(3553));
    outputs(7270) <= not(layer2_outputs(10111));
    outputs(7271) <= layer2_outputs(5239);
    outputs(7272) <= not(layer2_outputs(5022));
    outputs(7273) <= layer2_outputs(8892);
    outputs(7274) <= not(layer2_outputs(4751));
    outputs(7275) <= layer2_outputs(4739);
    outputs(7276) <= (layer2_outputs(6713)) xor (layer2_outputs(1008));
    outputs(7277) <= layer2_outputs(7405);
    outputs(7278) <= (layer2_outputs(1950)) xor (layer2_outputs(2903));
    outputs(7279) <= layer2_outputs(1591);
    outputs(7280) <= not(layer2_outputs(3898));
    outputs(7281) <= not(layer2_outputs(95));
    outputs(7282) <= not((layer2_outputs(7316)) xor (layer2_outputs(4863)));
    outputs(7283) <= layer2_outputs(975);
    outputs(7284) <= layer2_outputs(4547);
    outputs(7285) <= not(layer2_outputs(2717));
    outputs(7286) <= layer2_outputs(4543);
    outputs(7287) <= layer2_outputs(9593);
    outputs(7288) <= layer2_outputs(273);
    outputs(7289) <= not(layer2_outputs(9051));
    outputs(7290) <= layer2_outputs(3104);
    outputs(7291) <= (layer2_outputs(5202)) and not (layer2_outputs(4325));
    outputs(7292) <= not((layer2_outputs(5635)) xor (layer2_outputs(5049)));
    outputs(7293) <= layer2_outputs(9957);
    outputs(7294) <= not(layer2_outputs(4278));
    outputs(7295) <= not(layer2_outputs(7885));
    outputs(7296) <= not(layer2_outputs(150));
    outputs(7297) <= not(layer2_outputs(6832));
    outputs(7298) <= layer2_outputs(4321);
    outputs(7299) <= not((layer2_outputs(7105)) or (layer2_outputs(9192)));
    outputs(7300) <= not(layer2_outputs(7998));
    outputs(7301) <= not((layer2_outputs(7528)) xor (layer2_outputs(479)));
    outputs(7302) <= not((layer2_outputs(3695)) or (layer2_outputs(7271)));
    outputs(7303) <= not(layer2_outputs(5338));
    outputs(7304) <= layer2_outputs(7887);
    outputs(7305) <= not(layer2_outputs(4047));
    outputs(7306) <= (layer2_outputs(3250)) and (layer2_outputs(5647));
    outputs(7307) <= layer2_outputs(5629);
    outputs(7308) <= layer2_outputs(5592);
    outputs(7309) <= not(layer2_outputs(451));
    outputs(7310) <= layer2_outputs(5422);
    outputs(7311) <= layer2_outputs(8547);
    outputs(7312) <= not((layer2_outputs(8064)) xor (layer2_outputs(8530)));
    outputs(7313) <= (layer2_outputs(7753)) and not (layer2_outputs(5835));
    outputs(7314) <= layer2_outputs(8730);
    outputs(7315) <= not(layer2_outputs(6022)) or (layer2_outputs(9331));
    outputs(7316) <= layer2_outputs(9739);
    outputs(7317) <= layer2_outputs(6760);
    outputs(7318) <= not(layer2_outputs(4189));
    outputs(7319) <= layer2_outputs(6668);
    outputs(7320) <= not(layer2_outputs(3961));
    outputs(7321) <= '1';
    outputs(7322) <= layer2_outputs(8184);
    outputs(7323) <= not(layer2_outputs(1784));
    outputs(7324) <= layer2_outputs(3844);
    outputs(7325) <= (layer2_outputs(2320)) xor (layer2_outputs(2976));
    outputs(7326) <= (layer2_outputs(8343)) and not (layer2_outputs(9419));
    outputs(7327) <= (layer2_outputs(6859)) xor (layer2_outputs(2371));
    outputs(7328) <= not(layer2_outputs(7904));
    outputs(7329) <= not(layer2_outputs(4385));
    outputs(7330) <= layer2_outputs(9263);
    outputs(7331) <= layer2_outputs(10183);
    outputs(7332) <= not(layer2_outputs(4411));
    outputs(7333) <= not(layer2_outputs(2080));
    outputs(7334) <= not(layer2_outputs(1161));
    outputs(7335) <= not(layer2_outputs(6201));
    outputs(7336) <= layer2_outputs(1458);
    outputs(7337) <= layer2_outputs(6905);
    outputs(7338) <= layer2_outputs(7383);
    outputs(7339) <= not((layer2_outputs(7731)) and (layer2_outputs(562)));
    outputs(7340) <= layer2_outputs(7742);
    outputs(7341) <= layer2_outputs(4601);
    outputs(7342) <= not(layer2_outputs(8236));
    outputs(7343) <= layer2_outputs(7169);
    outputs(7344) <= not(layer2_outputs(6507));
    outputs(7345) <= (layer2_outputs(2286)) xor (layer2_outputs(371));
    outputs(7346) <= not(layer2_outputs(9699));
    outputs(7347) <= not(layer2_outputs(1379));
    outputs(7348) <= not((layer2_outputs(5219)) xor (layer2_outputs(7976)));
    outputs(7349) <= (layer2_outputs(1680)) xor (layer2_outputs(429));
    outputs(7350) <= layer2_outputs(5134);
    outputs(7351) <= (layer2_outputs(6914)) xor (layer2_outputs(5553));
    outputs(7352) <= layer2_outputs(1570);
    outputs(7353) <= not((layer2_outputs(1103)) xor (layer2_outputs(3185)));
    outputs(7354) <= layer2_outputs(4037);
    outputs(7355) <= layer2_outputs(2201);
    outputs(7356) <= not(layer2_outputs(3184));
    outputs(7357) <= not(layer2_outputs(5557));
    outputs(7358) <= (layer2_outputs(4771)) or (layer2_outputs(3473));
    outputs(7359) <= (layer2_outputs(4023)) and not (layer2_outputs(4904));
    outputs(7360) <= (layer2_outputs(189)) xor (layer2_outputs(6627));
    outputs(7361) <= (layer2_outputs(9632)) and not (layer2_outputs(7152));
    outputs(7362) <= not(layer2_outputs(501)) or (layer2_outputs(8539));
    outputs(7363) <= layer2_outputs(2825);
    outputs(7364) <= not(layer2_outputs(1970));
    outputs(7365) <= (layer2_outputs(8674)) and (layer2_outputs(5251));
    outputs(7366) <= layer2_outputs(865);
    outputs(7367) <= (layer2_outputs(4408)) xor (layer2_outputs(3294));
    outputs(7368) <= layer2_outputs(8882);
    outputs(7369) <= layer2_outputs(7966);
    outputs(7370) <= layer2_outputs(3701);
    outputs(7371) <= layer2_outputs(4443);
    outputs(7372) <= not((layer2_outputs(246)) and (layer2_outputs(9701)));
    outputs(7373) <= layer2_outputs(3976);
    outputs(7374) <= layer2_outputs(4176);
    outputs(7375) <= layer2_outputs(5776);
    outputs(7376) <= not((layer2_outputs(3327)) xor (layer2_outputs(27)));
    outputs(7377) <= layer2_outputs(9824);
    outputs(7378) <= not(layer2_outputs(8668));
    outputs(7379) <= not(layer2_outputs(1747));
    outputs(7380) <= (layer2_outputs(2140)) xor (layer2_outputs(8154));
    outputs(7381) <= (layer2_outputs(1329)) xor (layer2_outputs(1325));
    outputs(7382) <= layer2_outputs(5451);
    outputs(7383) <= not(layer2_outputs(7197));
    outputs(7384) <= (layer2_outputs(9520)) xor (layer2_outputs(6276));
    outputs(7385) <= (layer2_outputs(5606)) and not (layer2_outputs(5930));
    outputs(7386) <= not(layer2_outputs(10224));
    outputs(7387) <= (layer2_outputs(2810)) and not (layer2_outputs(6056));
    outputs(7388) <= layer2_outputs(7587);
    outputs(7389) <= not((layer2_outputs(960)) xor (layer2_outputs(4413)));
    outputs(7390) <= not(layer2_outputs(1267));
    outputs(7391) <= layer2_outputs(7670);
    outputs(7392) <= not(layer2_outputs(4845));
    outputs(7393) <= not(layer2_outputs(5569));
    outputs(7394) <= layer2_outputs(2889);
    outputs(7395) <= layer2_outputs(1110);
    outputs(7396) <= not((layer2_outputs(5989)) xor (layer2_outputs(4324)));
    outputs(7397) <= layer2_outputs(2553);
    outputs(7398) <= not(layer2_outputs(5881));
    outputs(7399) <= layer2_outputs(1551);
    outputs(7400) <= layer2_outputs(8584);
    outputs(7401) <= layer2_outputs(9783);
    outputs(7402) <= layer2_outputs(4507);
    outputs(7403) <= layer2_outputs(3388);
    outputs(7404) <= not(layer2_outputs(1530)) or (layer2_outputs(2607));
    outputs(7405) <= layer2_outputs(5593);
    outputs(7406) <= not(layer2_outputs(9468));
    outputs(7407) <= (layer2_outputs(10207)) and not (layer2_outputs(9443));
    outputs(7408) <= layer2_outputs(8276);
    outputs(7409) <= not(layer2_outputs(3143));
    outputs(7410) <= not(layer2_outputs(7353));
    outputs(7411) <= layer2_outputs(4077);
    outputs(7412) <= not(layer2_outputs(1672));
    outputs(7413) <= not(layer2_outputs(4169));
    outputs(7414) <= not((layer2_outputs(7030)) or (layer2_outputs(6690)));
    outputs(7415) <= not(layer2_outputs(1759));
    outputs(7416) <= not((layer2_outputs(2739)) xor (layer2_outputs(4805)));
    outputs(7417) <= (layer2_outputs(7488)) xor (layer2_outputs(31));
    outputs(7418) <= layer2_outputs(9385);
    outputs(7419) <= (layer2_outputs(869)) and not (layer2_outputs(4461));
    outputs(7420) <= not((layer2_outputs(8039)) or (layer2_outputs(1648)));
    outputs(7421) <= layer2_outputs(1858);
    outputs(7422) <= not(layer2_outputs(2831));
    outputs(7423) <= (layer2_outputs(1331)) and not (layer2_outputs(7016));
    outputs(7424) <= not((layer2_outputs(4637)) and (layer2_outputs(5423)));
    outputs(7425) <= layer2_outputs(5621);
    outputs(7426) <= (layer2_outputs(7684)) xor (layer2_outputs(7924));
    outputs(7427) <= not(layer2_outputs(2031));
    outputs(7428) <= (layer2_outputs(5706)) xor (layer2_outputs(8399));
    outputs(7429) <= not((layer2_outputs(8420)) xor (layer2_outputs(3731)));
    outputs(7430) <= not(layer2_outputs(9228));
    outputs(7431) <= layer2_outputs(2098);
    outputs(7432) <= not(layer2_outputs(2705)) or (layer2_outputs(1345));
    outputs(7433) <= layer2_outputs(3469);
    outputs(7434) <= not((layer2_outputs(845)) xor (layer2_outputs(6844)));
    outputs(7435) <= layer2_outputs(1263);
    outputs(7436) <= (layer2_outputs(428)) xor (layer2_outputs(1061));
    outputs(7437) <= layer2_outputs(726);
    outputs(7438) <= layer2_outputs(4157);
    outputs(7439) <= layer2_outputs(10041);
    outputs(7440) <= layer2_outputs(5385);
    outputs(7441) <= layer2_outputs(9388);
    outputs(7442) <= (layer2_outputs(3406)) xor (layer2_outputs(1727));
    outputs(7443) <= layer2_outputs(644);
    outputs(7444) <= layer2_outputs(539);
    outputs(7445) <= not(layer2_outputs(4009));
    outputs(7446) <= not((layer2_outputs(10154)) or (layer2_outputs(8863)));
    outputs(7447) <= not(layer2_outputs(6792));
    outputs(7448) <= layer2_outputs(7290);
    outputs(7449) <= layer2_outputs(1512);
    outputs(7450) <= not((layer2_outputs(8139)) xor (layer2_outputs(469)));
    outputs(7451) <= (layer2_outputs(3022)) or (layer2_outputs(200));
    outputs(7452) <= not((layer2_outputs(4588)) xor (layer2_outputs(2487)));
    outputs(7453) <= (layer2_outputs(10159)) xor (layer2_outputs(8444));
    outputs(7454) <= (layer2_outputs(1946)) xor (layer2_outputs(6112));
    outputs(7455) <= not((layer2_outputs(2488)) xor (layer2_outputs(1595)));
    outputs(7456) <= not((layer2_outputs(3068)) xor (layer2_outputs(1821)));
    outputs(7457) <= not(layer2_outputs(4592));
    outputs(7458) <= layer2_outputs(2366);
    outputs(7459) <= not(layer2_outputs(568));
    outputs(7460) <= layer2_outputs(3767);
    outputs(7461) <= not(layer2_outputs(6153));
    outputs(7462) <= not(layer2_outputs(5568));
    outputs(7463) <= layer2_outputs(3472);
    outputs(7464) <= not(layer2_outputs(4251));
    outputs(7465) <= (layer2_outputs(3700)) and not (layer2_outputs(7040));
    outputs(7466) <= layer2_outputs(3276);
    outputs(7467) <= (layer2_outputs(2871)) and not (layer2_outputs(9658));
    outputs(7468) <= layer2_outputs(5816);
    outputs(7469) <= (layer2_outputs(487)) and not (layer2_outputs(8420));
    outputs(7470) <= layer2_outputs(6381);
    outputs(7471) <= layer2_outputs(10232);
    outputs(7472) <= not(layer2_outputs(2423));
    outputs(7473) <= not((layer2_outputs(3895)) or (layer2_outputs(8588)));
    outputs(7474) <= not((layer2_outputs(2019)) xor (layer2_outputs(5854)));
    outputs(7475) <= layer2_outputs(8558);
    outputs(7476) <= not(layer2_outputs(7639));
    outputs(7477) <= not(layer2_outputs(8291));
    outputs(7478) <= not(layer2_outputs(1365));
    outputs(7479) <= not(layer2_outputs(5203)) or (layer2_outputs(3808));
    outputs(7480) <= not(layer2_outputs(4472)) or (layer2_outputs(6101));
    outputs(7481) <= (layer2_outputs(10117)) and (layer2_outputs(9510));
    outputs(7482) <= layer2_outputs(9010);
    outputs(7483) <= not(layer2_outputs(369));
    outputs(7484) <= not(layer2_outputs(10186));
    outputs(7485) <= layer2_outputs(3087);
    outputs(7486) <= (layer2_outputs(8323)) xor (layer2_outputs(7214));
    outputs(7487) <= not(layer2_outputs(8396)) or (layer2_outputs(9694));
    outputs(7488) <= (layer2_outputs(8063)) xor (layer2_outputs(3144));
    outputs(7489) <= not(layer2_outputs(1048));
    outputs(7490) <= (layer2_outputs(8519)) xor (layer2_outputs(6205));
    outputs(7491) <= layer2_outputs(10145);
    outputs(7492) <= (layer2_outputs(378)) and not (layer2_outputs(6754));
    outputs(7493) <= (layer2_outputs(6260)) xor (layer2_outputs(5165));
    outputs(7494) <= not(layer2_outputs(7881));
    outputs(7495) <= (layer2_outputs(9839)) xor (layer2_outputs(4109));
    outputs(7496) <= (layer2_outputs(3283)) and (layer2_outputs(5243));
    outputs(7497) <= not((layer2_outputs(2213)) xor (layer2_outputs(8781)));
    outputs(7498) <= not(layer2_outputs(9982));
    outputs(7499) <= (layer2_outputs(6916)) and not (layer2_outputs(5373));
    outputs(7500) <= not(layer2_outputs(6907));
    outputs(7501) <= not(layer2_outputs(4535));
    outputs(7502) <= not(layer2_outputs(9497));
    outputs(7503) <= not(layer2_outputs(5725));
    outputs(7504) <= layer2_outputs(4471);
    outputs(7505) <= layer2_outputs(4431);
    outputs(7506) <= not((layer2_outputs(5071)) or (layer2_outputs(3359)));
    outputs(7507) <= not(layer2_outputs(5687));
    outputs(7508) <= layer2_outputs(3550);
    outputs(7509) <= not(layer2_outputs(2622));
    outputs(7510) <= layer2_outputs(5400);
    outputs(7511) <= not(layer2_outputs(1107));
    outputs(7512) <= not(layer2_outputs(3755));
    outputs(7513) <= layer2_outputs(4679);
    outputs(7514) <= layer2_outputs(2157);
    outputs(7515) <= layer2_outputs(4893);
    outputs(7516) <= layer2_outputs(8804);
    outputs(7517) <= layer2_outputs(3447);
    outputs(7518) <= not(layer2_outputs(7779));
    outputs(7519) <= not((layer2_outputs(10045)) xor (layer2_outputs(10205)));
    outputs(7520) <= not(layer2_outputs(2203));
    outputs(7521) <= layer2_outputs(1999);
    outputs(7522) <= not(layer2_outputs(2091));
    outputs(7523) <= not((layer2_outputs(1383)) and (layer2_outputs(9228)));
    outputs(7524) <= not(layer2_outputs(1557));
    outputs(7525) <= layer2_outputs(8920);
    outputs(7526) <= not(layer2_outputs(8607));
    outputs(7527) <= (layer2_outputs(8865)) and not (layer2_outputs(1738));
    outputs(7528) <= (layer2_outputs(5309)) and not (layer2_outputs(9528));
    outputs(7529) <= layer2_outputs(4290);
    outputs(7530) <= layer2_outputs(7138);
    outputs(7531) <= not(layer2_outputs(5405));
    outputs(7532) <= not((layer2_outputs(1247)) and (layer2_outputs(4554)));
    outputs(7533) <= layer2_outputs(1547);
    outputs(7534) <= not(layer2_outputs(335));
    outputs(7535) <= layer2_outputs(9407);
    outputs(7536) <= not(layer2_outputs(6156));
    outputs(7537) <= (layer2_outputs(9928)) and (layer2_outputs(5197));
    outputs(7538) <= not(layer2_outputs(5107));
    outputs(7539) <= (layer2_outputs(1869)) and not (layer2_outputs(4581));
    outputs(7540) <= (layer2_outputs(7961)) and (layer2_outputs(4989));
    outputs(7541) <= not(layer2_outputs(1141));
    outputs(7542) <= layer2_outputs(4209);
    outputs(7543) <= (layer2_outputs(7488)) xor (layer2_outputs(4142));
    outputs(7544) <= (layer2_outputs(4781)) and (layer2_outputs(4637));
    outputs(7545) <= layer2_outputs(5258);
    outputs(7546) <= layer2_outputs(8397);
    outputs(7547) <= layer2_outputs(3662);
    outputs(7548) <= not(layer2_outputs(5696));
    outputs(7549) <= layer2_outputs(4482);
    outputs(7550) <= layer2_outputs(6911);
    outputs(7551) <= not(layer2_outputs(7517));
    outputs(7552) <= not((layer2_outputs(611)) xor (layer2_outputs(291)));
    outputs(7553) <= (layer2_outputs(1753)) xor (layer2_outputs(10065));
    outputs(7554) <= not(layer2_outputs(4475));
    outputs(7555) <= (layer2_outputs(2150)) and not (layer2_outputs(8116));
    outputs(7556) <= (layer2_outputs(5539)) and (layer2_outputs(3747));
    outputs(7557) <= layer2_outputs(2629);
    outputs(7558) <= not(layer2_outputs(1099));
    outputs(7559) <= (layer2_outputs(9657)) and (layer2_outputs(5389));
    outputs(7560) <= layer2_outputs(213);
    outputs(7561) <= layer2_outputs(1430);
    outputs(7562) <= not(layer2_outputs(3944));
    outputs(7563) <= not(layer2_outputs(8717));
    outputs(7564) <= not(layer2_outputs(6208));
    outputs(7565) <= not((layer2_outputs(2156)) or (layer2_outputs(3843)));
    outputs(7566) <= not(layer2_outputs(1759));
    outputs(7567) <= layer2_outputs(7177);
    outputs(7568) <= not(layer2_outputs(2560));
    outputs(7569) <= layer2_outputs(887);
    outputs(7570) <= not(layer2_outputs(7780));
    outputs(7571) <= layer2_outputs(716);
    outputs(7572) <= layer2_outputs(4534);
    outputs(7573) <= '0';
    outputs(7574) <= layer2_outputs(5055);
    outputs(7575) <= (layer2_outputs(2244)) and not (layer2_outputs(5982));
    outputs(7576) <= not(layer2_outputs(3556));
    outputs(7577) <= not(layer2_outputs(1630)) or (layer2_outputs(339));
    outputs(7578) <= not(layer2_outputs(4322));
    outputs(7579) <= (layer2_outputs(5787)) xor (layer2_outputs(7677));
    outputs(7580) <= not(layer2_outputs(7577));
    outputs(7581) <= layer2_outputs(361);
    outputs(7582) <= not(layer2_outputs(1763));
    outputs(7583) <= not(layer2_outputs(1266));
    outputs(7584) <= layer2_outputs(8431);
    outputs(7585) <= not(layer2_outputs(9304));
    outputs(7586) <= not(layer2_outputs(4678));
    outputs(7587) <= (layer2_outputs(7159)) xor (layer2_outputs(8726));
    outputs(7588) <= layer2_outputs(6605);
    outputs(7589) <= not(layer2_outputs(10036));
    outputs(7590) <= layer2_outputs(684);
    outputs(7591) <= (layer2_outputs(365)) and not (layer2_outputs(6392));
    outputs(7592) <= not(layer2_outputs(599)) or (layer2_outputs(6019));
    outputs(7593) <= layer2_outputs(6873);
    outputs(7594) <= not(layer2_outputs(2235));
    outputs(7595) <= (layer2_outputs(4566)) xor (layer2_outputs(9818));
    outputs(7596) <= not(layer2_outputs(2668));
    outputs(7597) <= '0';
    outputs(7598) <= layer2_outputs(8411);
    outputs(7599) <= not(layer2_outputs(1162));
    outputs(7600) <= not(layer2_outputs(9160));
    outputs(7601) <= not(layer2_outputs(1180)) or (layer2_outputs(7649));
    outputs(7602) <= not(layer2_outputs(1020));
    outputs(7603) <= not(layer2_outputs(226));
    outputs(7604) <= layer2_outputs(9879);
    outputs(7605) <= not(layer2_outputs(282));
    outputs(7606) <= layer2_outputs(850);
    outputs(7607) <= not((layer2_outputs(600)) xor (layer2_outputs(6524)));
    outputs(7608) <= (layer2_outputs(5221)) and (layer2_outputs(5780));
    outputs(7609) <= (layer2_outputs(8815)) and (layer2_outputs(2377));
    outputs(7610) <= not(layer2_outputs(7675));
    outputs(7611) <= not(layer2_outputs(4663));
    outputs(7612) <= not((layer2_outputs(8461)) xor (layer2_outputs(8854)));
    outputs(7613) <= layer2_outputs(9537);
    outputs(7614) <= not(layer2_outputs(5632));
    outputs(7615) <= not(layer2_outputs(5701));
    outputs(7616) <= layer2_outputs(7312);
    outputs(7617) <= not((layer2_outputs(1967)) or (layer2_outputs(9270)));
    outputs(7618) <= not((layer2_outputs(1679)) or (layer2_outputs(5950)));
    outputs(7619) <= not(layer2_outputs(9410));
    outputs(7620) <= not((layer2_outputs(9393)) xor (layer2_outputs(6120)));
    outputs(7621) <= not(layer2_outputs(7968));
    outputs(7622) <= not(layer2_outputs(3741));
    outputs(7623) <= not((layer2_outputs(8940)) xor (layer2_outputs(6694)));
    outputs(7624) <= not(layer2_outputs(4078));
    outputs(7625) <= (layer2_outputs(10002)) xor (layer2_outputs(5777));
    outputs(7626) <= not(layer2_outputs(7305));
    outputs(7627) <= not(layer2_outputs(3947));
    outputs(7628) <= not(layer2_outputs(7869));
    outputs(7629) <= (layer2_outputs(1144)) and not (layer2_outputs(4090));
    outputs(7630) <= layer2_outputs(5922);
    outputs(7631) <= layer2_outputs(6363);
    outputs(7632) <= not((layer2_outputs(8932)) or (layer2_outputs(9598)));
    outputs(7633) <= layer2_outputs(3469);
    outputs(7634) <= layer2_outputs(9569);
    outputs(7635) <= layer2_outputs(7184);
    outputs(7636) <= not((layer2_outputs(384)) xor (layer2_outputs(4983)));
    outputs(7637) <= layer2_outputs(7189);
    outputs(7638) <= not(layer2_outputs(693));
    outputs(7639) <= not(layer2_outputs(1162)) or (layer2_outputs(9173));
    outputs(7640) <= not(layer2_outputs(6938));
    outputs(7641) <= not(layer2_outputs(755));
    outputs(7642) <= not(layer2_outputs(6769));
    outputs(7643) <= (layer2_outputs(4119)) and not (layer2_outputs(8642));
    outputs(7644) <= not(layer2_outputs(9609));
    outputs(7645) <= layer2_outputs(5859);
    outputs(7646) <= (layer2_outputs(76)) and (layer2_outputs(8579));
    outputs(7647) <= not(layer2_outputs(3666));
    outputs(7648) <= not(layer2_outputs(6301)) or (layer2_outputs(7148));
    outputs(7649) <= layer2_outputs(3485);
    outputs(7650) <= (layer2_outputs(7553)) xor (layer2_outputs(8243));
    outputs(7651) <= not(layer2_outputs(8869));
    outputs(7652) <= not(layer2_outputs(9430));
    outputs(7653) <= layer2_outputs(4383);
    outputs(7654) <= not((layer2_outputs(7942)) xor (layer2_outputs(7134)));
    outputs(7655) <= not(layer2_outputs(6535)) or (layer2_outputs(7630));
    outputs(7656) <= layer2_outputs(4914);
    outputs(7657) <= not(layer2_outputs(8602));
    outputs(7658) <= not(layer2_outputs(3824));
    outputs(7659) <= layer2_outputs(5577);
    outputs(7660) <= (layer2_outputs(6801)) and not (layer2_outputs(7770));
    outputs(7661) <= not(layer2_outputs(84));
    outputs(7662) <= not(layer2_outputs(5081));
    outputs(7663) <= layer2_outputs(7492);
    outputs(7664) <= (layer2_outputs(7797)) xor (layer2_outputs(2686));
    outputs(7665) <= not(layer2_outputs(9314));
    outputs(7666) <= (layer2_outputs(1058)) xor (layer2_outputs(8168));
    outputs(7667) <= layer2_outputs(6687);
    outputs(7668) <= not((layer2_outputs(6090)) xor (layer2_outputs(2139)));
    outputs(7669) <= layer2_outputs(1114);
    outputs(7670) <= layer2_outputs(3668);
    outputs(7671) <= not(layer2_outputs(8400));
    outputs(7672) <= not((layer2_outputs(4912)) or (layer2_outputs(234)));
    outputs(7673) <= not(layer2_outputs(6498));
    outputs(7674) <= (layer2_outputs(9906)) and not (layer2_outputs(1526));
    outputs(7675) <= layer2_outputs(1651);
    outputs(7676) <= (layer2_outputs(4057)) and (layer2_outputs(1561));
    outputs(7677) <= layer2_outputs(7490);
    outputs(7678) <= layer2_outputs(4440);
    outputs(7679) <= not((layer2_outputs(6738)) xor (layer2_outputs(2944)));
    outputs(7680) <= not(layer2_outputs(7854));
    outputs(7681) <= (layer2_outputs(7634)) xor (layer2_outputs(6490));
    outputs(7682) <= not(layer2_outputs(3684));
    outputs(7683) <= (layer2_outputs(3370)) and not (layer2_outputs(9482));
    outputs(7684) <= not(layer2_outputs(4014));
    outputs(7685) <= layer2_outputs(8225);
    outputs(7686) <= not(layer2_outputs(2231));
    outputs(7687) <= not(layer2_outputs(5781));
    outputs(7688) <= layer2_outputs(1017);
    outputs(7689) <= layer2_outputs(7427);
    outputs(7690) <= (layer2_outputs(2188)) and not (layer2_outputs(9638));
    outputs(7691) <= layer2_outputs(2492);
    outputs(7692) <= not(layer2_outputs(228));
    outputs(7693) <= layer2_outputs(1479);
    outputs(7694) <= (layer2_outputs(9355)) xor (layer2_outputs(389));
    outputs(7695) <= layer2_outputs(2133);
    outputs(7696) <= (layer2_outputs(6258)) xor (layer2_outputs(3888));
    outputs(7697) <= not((layer2_outputs(7510)) xor (layer2_outputs(653)));
    outputs(7698) <= not(layer2_outputs(5388));
    outputs(7699) <= not(layer2_outputs(8943));
    outputs(7700) <= (layer2_outputs(244)) and (layer2_outputs(5117));
    outputs(7701) <= layer2_outputs(4829);
    outputs(7702) <= not((layer2_outputs(3691)) xor (layer2_outputs(1772)));
    outputs(7703) <= not(layer2_outputs(2609));
    outputs(7704) <= (layer2_outputs(3788)) xor (layer2_outputs(9943));
    outputs(7705) <= not(layer2_outputs(6209));
    outputs(7706) <= (layer2_outputs(7414)) xor (layer2_outputs(8427));
    outputs(7707) <= (layer2_outputs(4779)) and (layer2_outputs(10003));
    outputs(7708) <= layer2_outputs(1326);
    outputs(7709) <= not((layer2_outputs(3653)) xor (layer2_outputs(6661)));
    outputs(7710) <= (layer2_outputs(2071)) xor (layer2_outputs(9956));
    outputs(7711) <= not(layer2_outputs(197));
    outputs(7712) <= (layer2_outputs(5382)) and not (layer2_outputs(3395));
    outputs(7713) <= not(layer2_outputs(9402));
    outputs(7714) <= not(layer2_outputs(8358));
    outputs(7715) <= (layer2_outputs(5128)) or (layer2_outputs(6462));
    outputs(7716) <= layer2_outputs(5002);
    outputs(7717) <= not(layer2_outputs(8632)) or (layer2_outputs(3207));
    outputs(7718) <= not((layer2_outputs(7194)) xor (layer2_outputs(503)));
    outputs(7719) <= not(layer2_outputs(6191));
    outputs(7720) <= layer2_outputs(8689);
    outputs(7721) <= (layer2_outputs(6962)) and not (layer2_outputs(1041));
    outputs(7722) <= not((layer2_outputs(9217)) xor (layer2_outputs(9498)));
    outputs(7723) <= layer2_outputs(7219);
    outputs(7724) <= (layer2_outputs(2320)) and not (layer2_outputs(3279));
    outputs(7725) <= not((layer2_outputs(1565)) xor (layer2_outputs(7281)));
    outputs(7726) <= (layer2_outputs(700)) xor (layer2_outputs(6964));
    outputs(7727) <= not(layer2_outputs(1873));
    outputs(7728) <= not((layer2_outputs(8080)) and (layer2_outputs(3740)));
    outputs(7729) <= (layer2_outputs(8803)) xor (layer2_outputs(10087));
    outputs(7730) <= not((layer2_outputs(7106)) or (layer2_outputs(9986)));
    outputs(7731) <= not(layer2_outputs(8090));
    outputs(7732) <= layer2_outputs(8587);
    outputs(7733) <= layer2_outputs(2133);
    outputs(7734) <= layer2_outputs(9103);
    outputs(7735) <= not(layer2_outputs(3006)) or (layer2_outputs(3858));
    outputs(7736) <= layer2_outputs(6324);
    outputs(7737) <= layer2_outputs(5190);
    outputs(7738) <= layer2_outputs(9657);
    outputs(7739) <= (layer2_outputs(10000)) and (layer2_outputs(6374));
    outputs(7740) <= (layer2_outputs(842)) and not (layer2_outputs(187));
    outputs(7741) <= not(layer2_outputs(1700));
    outputs(7742) <= not(layer2_outputs(2411)) or (layer2_outputs(3523));
    outputs(7743) <= (layer2_outputs(10179)) xor (layer2_outputs(1156));
    outputs(7744) <= layer2_outputs(7769);
    outputs(7745) <= not(layer2_outputs(2588));
    outputs(7746) <= not(layer2_outputs(6917));
    outputs(7747) <= layer2_outputs(6300);
    outputs(7748) <= not((layer2_outputs(10182)) or (layer2_outputs(5417)));
    outputs(7749) <= layer2_outputs(661);
    outputs(7750) <= not(layer2_outputs(6608));
    outputs(7751) <= layer2_outputs(7755);
    outputs(7752) <= not((layer2_outputs(2302)) or (layer2_outputs(10004)));
    outputs(7753) <= not(layer2_outputs(805)) or (layer2_outputs(7272));
    outputs(7754) <= not(layer2_outputs(5794));
    outputs(7755) <= not(layer2_outputs(3287)) or (layer2_outputs(6090));
    outputs(7756) <= not((layer2_outputs(62)) and (layer2_outputs(5594)));
    outputs(7757) <= not(layer2_outputs(604));
    outputs(7758) <= (layer2_outputs(6072)) and (layer2_outputs(3943));
    outputs(7759) <= (layer2_outputs(5722)) xor (layer2_outputs(1634));
    outputs(7760) <= layer2_outputs(3205);
    outputs(7761) <= not(layer2_outputs(9599));
    outputs(7762) <= (layer2_outputs(6922)) and (layer2_outputs(7107));
    outputs(7763) <= not(layer2_outputs(9244));
    outputs(7764) <= not(layer2_outputs(3410));
    outputs(7765) <= not(layer2_outputs(7303));
    outputs(7766) <= not((layer2_outputs(3120)) or (layer2_outputs(4790)));
    outputs(7767) <= not(layer2_outputs(2827));
    outputs(7768) <= not((layer2_outputs(136)) xor (layer2_outputs(9921)));
    outputs(7769) <= not(layer2_outputs(2501));
    outputs(7770) <= not(layer2_outputs(8031));
    outputs(7771) <= not((layer2_outputs(8204)) or (layer2_outputs(6518)));
    outputs(7772) <= not(layer2_outputs(3003));
    outputs(7773) <= (layer2_outputs(1709)) xor (layer2_outputs(2373));
    outputs(7774) <= layer2_outputs(9597);
    outputs(7775) <= layer2_outputs(8803);
    outputs(7776) <= layer2_outputs(8790);
    outputs(7777) <= layer2_outputs(1832);
    outputs(7778) <= not(layer2_outputs(1725));
    outputs(7779) <= (layer2_outputs(153)) and not (layer2_outputs(1724));
    outputs(7780) <= layer2_outputs(4793);
    outputs(7781) <= (layer2_outputs(3456)) xor (layer2_outputs(3810));
    outputs(7782) <= (layer2_outputs(5322)) and (layer2_outputs(9291));
    outputs(7783) <= (layer2_outputs(1003)) and not (layer2_outputs(2915));
    outputs(7784) <= not(layer2_outputs(8534));
    outputs(7785) <= (layer2_outputs(8696)) xor (layer2_outputs(3864));
    outputs(7786) <= layer2_outputs(2732);
    outputs(7787) <= not((layer2_outputs(6424)) xor (layer2_outputs(5236)));
    outputs(7788) <= not(layer2_outputs(6515));
    outputs(7789) <= not(layer2_outputs(6778));
    outputs(7790) <= layer2_outputs(6472);
    outputs(7791) <= (layer2_outputs(8386)) and not (layer2_outputs(8596));
    outputs(7792) <= not((layer2_outputs(4231)) xor (layer2_outputs(474)));
    outputs(7793) <= layer2_outputs(6758);
    outputs(7794) <= layer2_outputs(1203);
    outputs(7795) <= not(layer2_outputs(4921));
    outputs(7796) <= not(layer2_outputs(5550));
    outputs(7797) <= layer2_outputs(6751);
    outputs(7798) <= layer2_outputs(1845);
    outputs(7799) <= layer2_outputs(1581);
    outputs(7800) <= not(layer2_outputs(5956));
    outputs(7801) <= (layer2_outputs(5459)) xor (layer2_outputs(2615));
    outputs(7802) <= (layer2_outputs(2204)) and (layer2_outputs(3165));
    outputs(7803) <= layer2_outputs(5920);
    outputs(7804) <= (layer2_outputs(2565)) xor (layer2_outputs(7629));
    outputs(7805) <= not(layer2_outputs(7682));
    outputs(7806) <= (layer2_outputs(683)) and not (layer2_outputs(6495));
    outputs(7807) <= not(layer2_outputs(4569));
    outputs(7808) <= layer2_outputs(7361);
    outputs(7809) <= not(layer2_outputs(1044));
    outputs(7810) <= not(layer2_outputs(9481)) or (layer2_outputs(8502));
    outputs(7811) <= not((layer2_outputs(4860)) xor (layer2_outputs(761)));
    outputs(7812) <= not(layer2_outputs(6919));
    outputs(7813) <= not((layer2_outputs(4751)) or (layer2_outputs(9614)));
    outputs(7814) <= layer2_outputs(1271);
    outputs(7815) <= layer2_outputs(9589);
    outputs(7816) <= layer2_outputs(8495);
    outputs(7817) <= layer2_outputs(8673);
    outputs(7818) <= layer2_outputs(9208);
    outputs(7819) <= (layer2_outputs(65)) xor (layer2_outputs(709));
    outputs(7820) <= layer2_outputs(3664);
    outputs(7821) <= (layer2_outputs(9085)) xor (layer2_outputs(6906));
    outputs(7822) <= layer2_outputs(10213);
    outputs(7823) <= (layer2_outputs(7860)) xor (layer2_outputs(6329));
    outputs(7824) <= (layer2_outputs(2286)) xor (layer2_outputs(1659));
    outputs(7825) <= layer2_outputs(6285);
    outputs(7826) <= not(layer2_outputs(1039));
    outputs(7827) <= not(layer2_outputs(1492));
    outputs(7828) <= not((layer2_outputs(8335)) or (layer2_outputs(5762)));
    outputs(7829) <= not(layer2_outputs(630));
    outputs(7830) <= not((layer2_outputs(3424)) xor (layer2_outputs(8966)));
    outputs(7831) <= (layer2_outputs(5711)) and not (layer2_outputs(5824));
    outputs(7832) <= layer2_outputs(8086);
    outputs(7833) <= not((layer2_outputs(1643)) xor (layer2_outputs(1476)));
    outputs(7834) <= not((layer2_outputs(9356)) xor (layer2_outputs(7761)));
    outputs(7835) <= not(layer2_outputs(9851));
    outputs(7836) <= layer2_outputs(9577);
    outputs(7837) <= layer2_outputs(5180);
    outputs(7838) <= not(layer2_outputs(8488));
    outputs(7839) <= not(layer2_outputs(8029));
    outputs(7840) <= not(layer2_outputs(1213));
    outputs(7841) <= layer2_outputs(2328);
    outputs(7842) <= layer2_outputs(1506);
    outputs(7843) <= not(layer2_outputs(3825));
    outputs(7844) <= layer2_outputs(4895);
    outputs(7845) <= not((layer2_outputs(1238)) xor (layer2_outputs(5122)));
    outputs(7846) <= not(layer2_outputs(3400)) or (layer2_outputs(6720));
    outputs(7847) <= layer2_outputs(4261);
    outputs(7848) <= (layer2_outputs(2367)) and not (layer2_outputs(9322));
    outputs(7849) <= (layer2_outputs(116)) xor (layer2_outputs(6045));
    outputs(7850) <= not(layer2_outputs(3735));
    outputs(7851) <= not(layer2_outputs(316));
    outputs(7852) <= layer2_outputs(4799);
    outputs(7853) <= not(layer2_outputs(9241));
    outputs(7854) <= (layer2_outputs(4982)) xor (layer2_outputs(123));
    outputs(7855) <= (layer2_outputs(3495)) xor (layer2_outputs(5140));
    outputs(7856) <= not((layer2_outputs(2466)) xor (layer2_outputs(2635)));
    outputs(7857) <= not(layer2_outputs(8471));
    outputs(7858) <= layer2_outputs(7268);
    outputs(7859) <= (layer2_outputs(10177)) and (layer2_outputs(4358));
    outputs(7860) <= not(layer2_outputs(6685));
    outputs(7861) <= layer2_outputs(7993);
    outputs(7862) <= (layer2_outputs(7043)) and not (layer2_outputs(1963));
    outputs(7863) <= not(layer2_outputs(4944));
    outputs(7864) <= not((layer2_outputs(1704)) and (layer2_outputs(8606)));
    outputs(7865) <= not(layer2_outputs(9463));
    outputs(7866) <= layer2_outputs(5783);
    outputs(7867) <= not(layer2_outputs(2499));
    outputs(7868) <= (layer2_outputs(4390)) and not (layer2_outputs(4656));
    outputs(7869) <= not(layer2_outputs(1407));
    outputs(7870) <= layer2_outputs(8419);
    outputs(7871) <= layer2_outputs(2465);
    outputs(7872) <= not((layer2_outputs(2839)) and (layer2_outputs(3738)));
    outputs(7873) <= layer2_outputs(10207);
    outputs(7874) <= not(layer2_outputs(9940));
    outputs(7875) <= layer2_outputs(4433);
    outputs(7876) <= (layer2_outputs(9356)) and not (layer2_outputs(3303));
    outputs(7877) <= layer2_outputs(7952);
    outputs(7878) <= layer2_outputs(3591);
    outputs(7879) <= not(layer2_outputs(9515));
    outputs(7880) <= (layer2_outputs(4195)) or (layer2_outputs(1336));
    outputs(7881) <= not((layer2_outputs(9828)) or (layer2_outputs(1635)));
    outputs(7882) <= not(layer2_outputs(106)) or (layer2_outputs(8643));
    outputs(7883) <= layer2_outputs(8657);
    outputs(7884) <= layer2_outputs(597);
    outputs(7885) <= not((layer2_outputs(9210)) or (layer2_outputs(9326)));
    outputs(7886) <= (layer2_outputs(2553)) and not (layer2_outputs(1703));
    outputs(7887) <= not((layer2_outputs(128)) xor (layer2_outputs(6376)));
    outputs(7888) <= (layer2_outputs(4817)) and not (layer2_outputs(2479));
    outputs(7889) <= not((layer2_outputs(4361)) or (layer2_outputs(1722)));
    outputs(7890) <= not(layer2_outputs(2591));
    outputs(7891) <= not(layer2_outputs(6116));
    outputs(7892) <= layer2_outputs(683);
    outputs(7893) <= not(layer2_outputs(231));
    outputs(7894) <= (layer2_outputs(4968)) xor (layer2_outputs(6337));
    outputs(7895) <= not((layer2_outputs(2738)) or (layer2_outputs(4129)));
    outputs(7896) <= not((layer2_outputs(8737)) and (layer2_outputs(5283)));
    outputs(7897) <= not((layer2_outputs(4257)) xor (layer2_outputs(2196)));
    outputs(7898) <= not(layer2_outputs(9831));
    outputs(7899) <= layer2_outputs(7221);
    outputs(7900) <= (layer2_outputs(7200)) and (layer2_outputs(6935));
    outputs(7901) <= not(layer2_outputs(1727));
    outputs(7902) <= layer2_outputs(8287);
    outputs(7903) <= layer2_outputs(2387);
    outputs(7904) <= (layer2_outputs(2892)) xor (layer2_outputs(4557));
    outputs(7905) <= layer2_outputs(8798);
    outputs(7906) <= not(layer2_outputs(8853));
    outputs(7907) <= (layer2_outputs(8403)) and not (layer2_outputs(5548));
    outputs(7908) <= not(layer2_outputs(6817));
    outputs(7909) <= not((layer2_outputs(3856)) or (layer2_outputs(7230)));
    outputs(7910) <= (layer2_outputs(6196)) and (layer2_outputs(7326));
    outputs(7911) <= layer2_outputs(7418);
    outputs(7912) <= (layer2_outputs(7466)) and not (layer2_outputs(5210));
    outputs(7913) <= not(layer2_outputs(1182)) or (layer2_outputs(122));
    outputs(7914) <= layer2_outputs(3053);
    outputs(7915) <= not((layer2_outputs(8289)) or (layer2_outputs(9358)));
    outputs(7916) <= layer2_outputs(2119);
    outputs(7917) <= layer2_outputs(7277);
    outputs(7918) <= not(layer2_outputs(2938));
    outputs(7919) <= not((layer2_outputs(6605)) xor (layer2_outputs(9746)));
    outputs(7920) <= (layer2_outputs(5349)) and not (layer2_outputs(5773));
    outputs(7921) <= layer2_outputs(4131);
    outputs(7922) <= not(layer2_outputs(5064)) or (layer2_outputs(5995));
    outputs(7923) <= not(layer2_outputs(2991));
    outputs(7924) <= layer2_outputs(3100);
    outputs(7925) <= not((layer2_outputs(3974)) xor (layer2_outputs(5807)));
    outputs(7926) <= (layer2_outputs(4685)) and not (layer2_outputs(6972));
    outputs(7927) <= not(layer2_outputs(4076));
    outputs(7928) <= layer2_outputs(3792);
    outputs(7929) <= not(layer2_outputs(8267));
    outputs(7930) <= layer2_outputs(1027);
    outputs(7931) <= layer2_outputs(9922);
    outputs(7932) <= layer2_outputs(9269);
    outputs(7933) <= layer2_outputs(7174);
    outputs(7934) <= layer2_outputs(9983);
    outputs(7935) <= not(layer2_outputs(1541));
    outputs(7936) <= layer2_outputs(9621);
    outputs(7937) <= not((layer2_outputs(6716)) xor (layer2_outputs(5451)));
    outputs(7938) <= not((layer2_outputs(2451)) and (layer2_outputs(8158)));
    outputs(7939) <= layer2_outputs(6555);
    outputs(7940) <= layer2_outputs(731);
    outputs(7941) <= not(layer2_outputs(3));
    outputs(7942) <= not((layer2_outputs(6448)) xor (layer2_outputs(1072)));
    outputs(7943) <= not((layer2_outputs(3235)) xor (layer2_outputs(6834)));
    outputs(7944) <= not((layer2_outputs(8691)) or (layer2_outputs(8890)));
    outputs(7945) <= not(layer2_outputs(8874));
    outputs(7946) <= layer2_outputs(9056);
    outputs(7947) <= (layer2_outputs(3102)) and not (layer2_outputs(3415));
    outputs(7948) <= not(layer2_outputs(5498));
    outputs(7949) <= not(layer2_outputs(2290));
    outputs(7950) <= not((layer2_outputs(5989)) xor (layer2_outputs(2218)));
    outputs(7951) <= not(layer2_outputs(1995));
    outputs(7952) <= layer2_outputs(9199);
    outputs(7953) <= layer2_outputs(3626);
    outputs(7954) <= layer2_outputs(1368);
    outputs(7955) <= layer2_outputs(4832);
    outputs(7956) <= not(layer2_outputs(6622));
    outputs(7957) <= layer2_outputs(292);
    outputs(7958) <= not(layer2_outputs(2604));
    outputs(7959) <= layer2_outputs(370);
    outputs(7960) <= (layer2_outputs(614)) xor (layer2_outputs(5937));
    outputs(7961) <= layer2_outputs(8097);
    outputs(7962) <= not(layer2_outputs(3644));
    outputs(7963) <= (layer2_outputs(3528)) xor (layer2_outputs(118));
    outputs(7964) <= not(layer2_outputs(7554));
    outputs(7965) <= layer2_outputs(3117);
    outputs(7966) <= not(layer2_outputs(6790));
    outputs(7967) <= not((layer2_outputs(905)) and (layer2_outputs(1554)));
    outputs(7968) <= not((layer2_outputs(6952)) xor (layer2_outputs(6713)));
    outputs(7969) <= layer2_outputs(5392);
    outputs(7970) <= layer2_outputs(1921);
    outputs(7971) <= (layer2_outputs(4113)) xor (layer2_outputs(5437));
    outputs(7972) <= not((layer2_outputs(8354)) xor (layer2_outputs(4132)));
    outputs(7973) <= not(layer2_outputs(1475));
    outputs(7974) <= (layer2_outputs(6195)) and not (layer2_outputs(3455));
    outputs(7975) <= not((layer2_outputs(8278)) and (layer2_outputs(4182)));
    outputs(7976) <= not(layer2_outputs(8263));
    outputs(7977) <= not((layer2_outputs(4234)) xor (layer2_outputs(1266)));
    outputs(7978) <= layer2_outputs(4039);
    outputs(7979) <= layer2_outputs(5733);
    outputs(7980) <= not((layer2_outputs(1929)) or (layer2_outputs(6465)));
    outputs(7981) <= not((layer2_outputs(2521)) xor (layer2_outputs(4279)));
    outputs(7982) <= not((layer2_outputs(3901)) xor (layer2_outputs(507)));
    outputs(7983) <= layer2_outputs(661);
    outputs(7984) <= layer2_outputs(1288);
    outputs(7985) <= layer2_outputs(4961);
    outputs(7986) <= layer2_outputs(5225);
    outputs(7987) <= layer2_outputs(8493);
    outputs(7988) <= not((layer2_outputs(8690)) xor (layer2_outputs(9213)));
    outputs(7989) <= layer2_outputs(5134);
    outputs(7990) <= not(layer2_outputs(6733));
    outputs(7991) <= not(layer2_outputs(2791));
    outputs(7992) <= layer2_outputs(5160);
    outputs(7993) <= (layer2_outputs(9567)) xor (layer2_outputs(6030));
    outputs(7994) <= not(layer2_outputs(8738)) or (layer2_outputs(6281));
    outputs(7995) <= layer2_outputs(9459);
    outputs(7996) <= (layer2_outputs(7890)) xor (layer2_outputs(7801));
    outputs(7997) <= layer2_outputs(2638);
    outputs(7998) <= layer2_outputs(3878);
    outputs(7999) <= not(layer2_outputs(4557));
    outputs(8000) <= layer2_outputs(8092);
    outputs(8001) <= not(layer2_outputs(5396));
    outputs(8002) <= layer2_outputs(5165);
    outputs(8003) <= not(layer2_outputs(9197));
    outputs(8004) <= layer2_outputs(446);
    outputs(8005) <= not((layer2_outputs(7212)) xor (layer2_outputs(7731)));
    outputs(8006) <= not(layer2_outputs(63));
    outputs(8007) <= layer2_outputs(9810);
    outputs(8008) <= (layer2_outputs(7679)) xor (layer2_outputs(1692));
    outputs(8009) <= not(layer2_outputs(171));
    outputs(8010) <= (layer2_outputs(5588)) xor (layer2_outputs(7931));
    outputs(8011) <= not(layer2_outputs(8111));
    outputs(8012) <= (layer2_outputs(7926)) and (layer2_outputs(6589));
    outputs(8013) <= not(layer2_outputs(6384));
    outputs(8014) <= layer2_outputs(3789);
    outputs(8015) <= not((layer2_outputs(5575)) xor (layer2_outputs(800)));
    outputs(8016) <= not(layer2_outputs(251));
    outputs(8017) <= not((layer2_outputs(3300)) xor (layer2_outputs(9392)));
    outputs(8018) <= not(layer2_outputs(9868));
    outputs(8019) <= not(layer2_outputs(7005));
    outputs(8020) <= layer2_outputs(5924);
    outputs(8021) <= not(layer2_outputs(1676));
    outputs(8022) <= (layer2_outputs(6470)) and not (layer2_outputs(6469));
    outputs(8023) <= layer2_outputs(3281);
    outputs(8024) <= not(layer2_outputs(4630));
    outputs(8025) <= not(layer2_outputs(4219));
    outputs(8026) <= not(layer2_outputs(4757));
    outputs(8027) <= (layer2_outputs(8098)) and not (layer2_outputs(1678));
    outputs(8028) <= not(layer2_outputs(6189));
    outputs(8029) <= not(layer2_outputs(1338));
    outputs(8030) <= layer2_outputs(2944);
    outputs(8031) <= not(layer2_outputs(1145));
    outputs(8032) <= not((layer2_outputs(9212)) and (layer2_outputs(10151)));
    outputs(8033) <= layer2_outputs(7384);
    outputs(8034) <= (layer2_outputs(5377)) and (layer2_outputs(3343));
    outputs(8035) <= not(layer2_outputs(2931));
    outputs(8036) <= not(layer2_outputs(9565));
    outputs(8037) <= not((layer2_outputs(82)) xor (layer2_outputs(7430)));
    outputs(8038) <= not(layer2_outputs(2448));
    outputs(8039) <= (layer2_outputs(9161)) and (layer2_outputs(3633));
    outputs(8040) <= not(layer2_outputs(9533));
    outputs(8041) <= layer2_outputs(3248);
    outputs(8042) <= layer2_outputs(5221);
    outputs(8043) <= (layer2_outputs(9337)) xor (layer2_outputs(5847));
    outputs(8044) <= (layer2_outputs(7081)) xor (layer2_outputs(3624));
    outputs(8045) <= not(layer2_outputs(10078));
    outputs(8046) <= (layer2_outputs(1965)) and not (layer2_outputs(7644));
    outputs(8047) <= layer2_outputs(10161);
    outputs(8048) <= not(layer2_outputs(4581));
    outputs(8049) <= layer2_outputs(3299);
    outputs(8050) <= layer2_outputs(4610);
    outputs(8051) <= not((layer2_outputs(3503)) xor (layer2_outputs(9142)));
    outputs(8052) <= layer2_outputs(1549);
    outputs(8053) <= not((layer2_outputs(7100)) xor (layer2_outputs(4623)));
    outputs(8054) <= not(layer2_outputs(2402));
    outputs(8055) <= not(layer2_outputs(7249)) or (layer2_outputs(1573));
    outputs(8056) <= not((layer2_outputs(567)) xor (layer2_outputs(4150)));
    outputs(8057) <= not(layer2_outputs(3196));
    outputs(8058) <= not(layer2_outputs(7127));
    outputs(8059) <= (layer2_outputs(1608)) and (layer2_outputs(2815));
    outputs(8060) <= not(layer2_outputs(970));
    outputs(8061) <= not(layer2_outputs(1734));
    outputs(8062) <= layer2_outputs(2215);
    outputs(8063) <= (layer2_outputs(8309)) xor (layer2_outputs(8294));
    outputs(8064) <= (layer2_outputs(1092)) and (layer2_outputs(7659));
    outputs(8065) <= (layer2_outputs(5219)) and (layer2_outputs(956));
    outputs(8066) <= not(layer2_outputs(5337)) or (layer2_outputs(6890));
    outputs(8067) <= layer2_outputs(1546);
    outputs(8068) <= not(layer2_outputs(4486));
    outputs(8069) <= layer2_outputs(5459);
    outputs(8070) <= (layer2_outputs(6349)) and not (layer2_outputs(8051));
    outputs(8071) <= layer2_outputs(7976);
    outputs(8072) <= not(layer2_outputs(5691));
    outputs(8073) <= layer2_outputs(714);
    outputs(8074) <= (layer2_outputs(4874)) xor (layer2_outputs(851));
    outputs(8075) <= (layer2_outputs(8649)) xor (layer2_outputs(3683));
    outputs(8076) <= not(layer2_outputs(7167));
    outputs(8077) <= layer2_outputs(4854);
    outputs(8078) <= layer2_outputs(2632);
    outputs(8079) <= not(layer2_outputs(4299));
    outputs(8080) <= (layer2_outputs(7293)) xor (layer2_outputs(4278));
    outputs(8081) <= not(layer2_outputs(9650));
    outputs(8082) <= (layer2_outputs(7868)) and not (layer2_outputs(5509));
    outputs(8083) <= layer2_outputs(9970);
    outputs(8084) <= layer2_outputs(6482);
    outputs(8085) <= not(layer2_outputs(8872)) or (layer2_outputs(8982));
    outputs(8086) <= layer2_outputs(5006);
    outputs(8087) <= not(layer2_outputs(390));
    outputs(8088) <= (layer2_outputs(631)) and (layer2_outputs(1714));
    outputs(8089) <= (layer2_outputs(8433)) and (layer2_outputs(3421));
    outputs(8090) <= not((layer2_outputs(5182)) xor (layer2_outputs(4138)));
    outputs(8091) <= not((layer2_outputs(1756)) xor (layer2_outputs(6245)));
    outputs(8092) <= layer2_outputs(6909);
    outputs(8093) <= (layer2_outputs(1150)) and not (layer2_outputs(7877));
    outputs(8094) <= not(layer2_outputs(2756));
    outputs(8095) <= not(layer2_outputs(1314));
    outputs(8096) <= not((layer2_outputs(9258)) xor (layer2_outputs(1406)));
    outputs(8097) <= layer2_outputs(5102);
    outputs(8098) <= (layer2_outputs(2961)) and (layer2_outputs(5143));
    outputs(8099) <= layer2_outputs(4089);
    outputs(8100) <= layer2_outputs(2627);
    outputs(8101) <= layer2_outputs(2236);
    outputs(8102) <= not(layer2_outputs(1157));
    outputs(8103) <= (layer2_outputs(8414)) and (layer2_outputs(6157));
    outputs(8104) <= (layer2_outputs(5598)) xor (layer2_outputs(828));
    outputs(8105) <= not(layer2_outputs(6273));
    outputs(8106) <= layer2_outputs(6939);
    outputs(8107) <= not((layer2_outputs(9429)) and (layer2_outputs(9963)));
    outputs(8108) <= not(layer2_outputs(1428));
    outputs(8109) <= layer2_outputs(3662);
    outputs(8110) <= (layer2_outputs(10229)) and not (layer2_outputs(5535));
    outputs(8111) <= layer2_outputs(2451);
    outputs(8112) <= layer2_outputs(1603);
    outputs(8113) <= not(layer2_outputs(3667));
    outputs(8114) <= not(layer2_outputs(1413));
    outputs(8115) <= layer2_outputs(10149);
    outputs(8116) <= layer2_outputs(8081);
    outputs(8117) <= (layer2_outputs(3392)) or (layer2_outputs(5209));
    outputs(8118) <= (layer2_outputs(4336)) xor (layer2_outputs(9089));
    outputs(8119) <= layer2_outputs(9121);
    outputs(8120) <= layer2_outputs(8526);
    outputs(8121) <= (layer2_outputs(3134)) and not (layer2_outputs(3651));
    outputs(8122) <= layer2_outputs(1597);
    outputs(8123) <= not(layer2_outputs(6170));
    outputs(8124) <= not(layer2_outputs(6944)) or (layer2_outputs(1339));
    outputs(8125) <= layer2_outputs(8392);
    outputs(8126) <= layer2_outputs(158);
    outputs(8127) <= not((layer2_outputs(9002)) xor (layer2_outputs(3151)));
    outputs(8128) <= not(layer2_outputs(7657));
    outputs(8129) <= not((layer2_outputs(9666)) xor (layer2_outputs(2095)));
    outputs(8130) <= not(layer2_outputs(8678));
    outputs(8131) <= not(layer2_outputs(5146));
    outputs(8132) <= not((layer2_outputs(7246)) xor (layer2_outputs(4271)));
    outputs(8133) <= not(layer2_outputs(551));
    outputs(8134) <= layer2_outputs(6169);
    outputs(8135) <= (layer2_outputs(5648)) and (layer2_outputs(4196));
    outputs(8136) <= layer2_outputs(5798);
    outputs(8137) <= (layer2_outputs(4834)) xor (layer2_outputs(6261));
    outputs(8138) <= layer2_outputs(1400);
    outputs(8139) <= layer2_outputs(7061);
    outputs(8140) <= layer2_outputs(1309);
    outputs(8141) <= not(layer2_outputs(488));
    outputs(8142) <= (layer2_outputs(894)) and not (layer2_outputs(5015));
    outputs(8143) <= layer2_outputs(8425);
    outputs(8144) <= not((layer2_outputs(8582)) xor (layer2_outputs(1887)));
    outputs(8145) <= layer2_outputs(5267);
    outputs(8146) <= (layer2_outputs(1001)) and (layer2_outputs(3246));
    outputs(8147) <= layer2_outputs(5753);
    outputs(8148) <= not((layer2_outputs(9930)) xor (layer2_outputs(1342)));
    outputs(8149) <= layer2_outputs(995);
    outputs(8150) <= not(layer2_outputs(8836));
    outputs(8151) <= not(layer2_outputs(4378));
    outputs(8152) <= not(layer2_outputs(674)) or (layer2_outputs(7208));
    outputs(8153) <= layer2_outputs(1156);
    outputs(8154) <= not((layer2_outputs(5642)) xor (layer2_outputs(10223)));
    outputs(8155) <= not((layer2_outputs(8451)) and (layer2_outputs(8361)));
    outputs(8156) <= layer2_outputs(6187);
    outputs(8157) <= layer2_outputs(7219);
    outputs(8158) <= not((layer2_outputs(9363)) xor (layer2_outputs(484)));
    outputs(8159) <= not(layer2_outputs(2012));
    outputs(8160) <= not(layer2_outputs(8568));
    outputs(8161) <= not(layer2_outputs(2510));
    outputs(8162) <= not((layer2_outputs(2806)) xor (layer2_outputs(1115)));
    outputs(8163) <= not(layer2_outputs(2714));
    outputs(8164) <= (layer2_outputs(4179)) and not (layer2_outputs(3494));
    outputs(8165) <= not((layer2_outputs(9230)) and (layer2_outputs(6533)));
    outputs(8166) <= not(layer2_outputs(3530));
    outputs(8167) <= not(layer2_outputs(8314));
    outputs(8168) <= (layer2_outputs(107)) xor (layer2_outputs(4656));
    outputs(8169) <= layer2_outputs(1256);
    outputs(8170) <= layer2_outputs(4949);
    outputs(8171) <= (layer2_outputs(9143)) xor (layer2_outputs(3586));
    outputs(8172) <= (layer2_outputs(3780)) xor (layer2_outputs(200));
    outputs(8173) <= not(layer2_outputs(9236));
    outputs(8174) <= not(layer2_outputs(5928));
    outputs(8175) <= not(layer2_outputs(9293));
    outputs(8176) <= (layer2_outputs(1611)) and (layer2_outputs(233));
    outputs(8177) <= not((layer2_outputs(460)) xor (layer2_outputs(1622)));
    outputs(8178) <= layer2_outputs(4837);
    outputs(8179) <= not(layer2_outputs(7944));
    outputs(8180) <= not(layer2_outputs(3985));
    outputs(8181) <= not(layer2_outputs(7862));
    outputs(8182) <= not(layer2_outputs(7763)) or (layer2_outputs(3341));
    outputs(8183) <= layer2_outputs(8366);
    outputs(8184) <= layer2_outputs(5206);
    outputs(8185) <= not(layer2_outputs(1187));
    outputs(8186) <= layer2_outputs(9438);
    outputs(8187) <= not(layer2_outputs(10031));
    outputs(8188) <= (layer2_outputs(8927)) xor (layer2_outputs(3736));
    outputs(8189) <= not(layer2_outputs(2103));
    outputs(8190) <= not(layer2_outputs(8941));
    outputs(8191) <= layer2_outputs(2573);
    outputs(8192) <= not((layer2_outputs(10030)) xor (layer2_outputs(6936)));
    outputs(8193) <= not((layer2_outputs(3464)) xor (layer2_outputs(5418)));
    outputs(8194) <= not((layer2_outputs(6740)) xor (layer2_outputs(3365)));
    outputs(8195) <= not((layer2_outputs(2110)) xor (layer2_outputs(7398)));
    outputs(8196) <= layer2_outputs(8714);
    outputs(8197) <= layer2_outputs(8055);
    outputs(8198) <= (layer2_outputs(4228)) xor (layer2_outputs(4702));
    outputs(8199) <= (layer2_outputs(8300)) and not (layer2_outputs(8071));
    outputs(8200) <= not(layer2_outputs(3138));
    outputs(8201) <= layer2_outputs(1116);
    outputs(8202) <= not((layer2_outputs(5105)) xor (layer2_outputs(381)));
    outputs(8203) <= (layer2_outputs(7472)) xor (layer2_outputs(1151));
    outputs(8204) <= not(layer2_outputs(5526));
    outputs(8205) <= not(layer2_outputs(9956));
    outputs(8206) <= not((layer2_outputs(1264)) xor (layer2_outputs(98)));
    outputs(8207) <= layer2_outputs(1914);
    outputs(8208) <= layer2_outputs(174);
    outputs(8209) <= not(layer2_outputs(8652));
    outputs(8210) <= not(layer2_outputs(5633)) or (layer2_outputs(5746));
    outputs(8211) <= not((layer2_outputs(4909)) xor (layer2_outputs(8795)));
    outputs(8212) <= not((layer2_outputs(5042)) xor (layer2_outputs(8219)));
    outputs(8213) <= not(layer2_outputs(10193));
    outputs(8214) <= not(layer2_outputs(9526)) or (layer2_outputs(3803));
    outputs(8215) <= layer2_outputs(3920);
    outputs(8216) <= layer2_outputs(8550);
    outputs(8217) <= layer2_outputs(9532);
    outputs(8218) <= not((layer2_outputs(4730)) xor (layer2_outputs(5566)));
    outputs(8219) <= layer2_outputs(9464);
    outputs(8220) <= (layer2_outputs(264)) xor (layer2_outputs(7962));
    outputs(8221) <= not(layer2_outputs(1228));
    outputs(8222) <= not(layer2_outputs(2025));
    outputs(8223) <= layer2_outputs(729);
    outputs(8224) <= layer2_outputs(6556);
    outputs(8225) <= layer2_outputs(5378);
    outputs(8226) <= not(layer2_outputs(849));
    outputs(8227) <= (layer2_outputs(6176)) xor (layer2_outputs(6462));
    outputs(8228) <= layer2_outputs(3807);
    outputs(8229) <= not((layer2_outputs(3307)) and (layer2_outputs(6237)));
    outputs(8230) <= not(layer2_outputs(4931));
    outputs(8231) <= not(layer2_outputs(6532));
    outputs(8232) <= not((layer2_outputs(3379)) and (layer2_outputs(9216)));
    outputs(8233) <= '1';
    outputs(8234) <= layer2_outputs(4296);
    outputs(8235) <= not((layer2_outputs(9756)) xor (layer2_outputs(1018)));
    outputs(8236) <= layer2_outputs(2414);
    outputs(8237) <= layer2_outputs(9126);
    outputs(8238) <= not(layer2_outputs(7185));
    outputs(8239) <= not(layer2_outputs(8345)) or (layer2_outputs(8384));
    outputs(8240) <= not((layer2_outputs(5742)) and (layer2_outputs(9277)));
    outputs(8241) <= not((layer2_outputs(4143)) xor (layer2_outputs(5012)));
    outputs(8242) <= not((layer2_outputs(2148)) xor (layer2_outputs(3627)));
    outputs(8243) <= layer2_outputs(10228);
    outputs(8244) <= not(layer2_outputs(9576));
    outputs(8245) <= not(layer2_outputs(7381));
    outputs(8246) <= not(layer2_outputs(2563)) or (layer2_outputs(4886));
    outputs(8247) <= layer2_outputs(5428);
    outputs(8248) <= not(layer2_outputs(8741));
    outputs(8249) <= not((layer2_outputs(3531)) xor (layer2_outputs(4803)));
    outputs(8250) <= not(layer2_outputs(3639));
    outputs(8251) <= layer2_outputs(84);
    outputs(8252) <= not((layer2_outputs(2698)) xor (layer2_outputs(4253)));
    outputs(8253) <= layer2_outputs(2562);
    outputs(8254) <= not(layer2_outputs(1793));
    outputs(8255) <= not(layer2_outputs(8802)) or (layer2_outputs(6510));
    outputs(8256) <= layer2_outputs(5496);
    outputs(8257) <= layer2_outputs(1964);
    outputs(8258) <= layer2_outputs(8505);
    outputs(8259) <= not(layer2_outputs(379));
    outputs(8260) <= layer2_outputs(8506);
    outputs(8261) <= not(layer2_outputs(5651));
    outputs(8262) <= not(layer2_outputs(1860)) or (layer2_outputs(2960));
    outputs(8263) <= layer2_outputs(998);
    outputs(8264) <= not(layer2_outputs(4750)) or (layer2_outputs(3598));
    outputs(8265) <= not(layer2_outputs(7202));
    outputs(8266) <= layer2_outputs(4055);
    outputs(8267) <= layer2_outputs(9836);
    outputs(8268) <= (layer2_outputs(9047)) and (layer2_outputs(5020));
    outputs(8269) <= not((layer2_outputs(2963)) and (layer2_outputs(9033)));
    outputs(8270) <= layer2_outputs(2455);
    outputs(8271) <= layer2_outputs(8301);
    outputs(8272) <= layer2_outputs(2020);
    outputs(8273) <= not(layer2_outputs(8258)) or (layer2_outputs(4872));
    outputs(8274) <= layer2_outputs(816);
    outputs(8275) <= not((layer2_outputs(397)) xor (layer2_outputs(5180)));
    outputs(8276) <= not((layer2_outputs(32)) xor (layer2_outputs(2751)));
    outputs(8277) <= (layer2_outputs(9993)) xor (layer2_outputs(1445));
    outputs(8278) <= (layer2_outputs(151)) xor (layer2_outputs(7482));
    outputs(8279) <= not(layer2_outputs(751));
    outputs(8280) <= not(layer2_outputs(5393));
    outputs(8281) <= not((layer2_outputs(4639)) xor (layer2_outputs(4513)));
    outputs(8282) <= layer2_outputs(7699);
    outputs(8283) <= layer2_outputs(8666);
    outputs(8284) <= not(layer2_outputs(6451));
    outputs(8285) <= (layer2_outputs(10195)) and not (layer2_outputs(8157));
    outputs(8286) <= not((layer2_outputs(2082)) and (layer2_outputs(9045)));
    outputs(8287) <= layer2_outputs(966);
    outputs(8288) <= layer2_outputs(4299);
    outputs(8289) <= not(layer2_outputs(37));
    outputs(8290) <= not(layer2_outputs(3927));
    outputs(8291) <= layer2_outputs(6116);
    outputs(8292) <= (layer2_outputs(4632)) and (layer2_outputs(2731));
    outputs(8293) <= layer2_outputs(8724);
    outputs(8294) <= not((layer2_outputs(9280)) xor (layer2_outputs(6752)));
    outputs(8295) <= layer2_outputs(2359);
    outputs(8296) <= layer2_outputs(6505);
    outputs(8297) <= not(layer2_outputs(5931));
    outputs(8298) <= not(layer2_outputs(3501));
    outputs(8299) <= not((layer2_outputs(1901)) xor (layer2_outputs(7929)));
    outputs(8300) <= not((layer2_outputs(1519)) xor (layer2_outputs(2356)));
    outputs(8301) <= layer2_outputs(8400);
    outputs(8302) <= (layer2_outputs(2701)) xor (layer2_outputs(7616));
    outputs(8303) <= not((layer2_outputs(3591)) xor (layer2_outputs(8132)));
    outputs(8304) <= not(layer2_outputs(1149));
    outputs(8305) <= not((layer2_outputs(1566)) xor (layer2_outputs(8696)));
    outputs(8306) <= (layer2_outputs(8458)) xor (layer2_outputs(4172));
    outputs(8307) <= not((layer2_outputs(4394)) xor (layer2_outputs(6071)));
    outputs(8308) <= not((layer2_outputs(14)) xor (layer2_outputs(7060)));
    outputs(8309) <= layer2_outputs(239);
    outputs(8310) <= not((layer2_outputs(1007)) xor (layer2_outputs(2421)));
    outputs(8311) <= not(layer2_outputs(9200)) or (layer2_outputs(225));
    outputs(8312) <= not(layer2_outputs(1067)) or (layer2_outputs(1774));
    outputs(8313) <= not(layer2_outputs(2075));
    outputs(8314) <= not((layer2_outputs(9611)) xor (layer2_outputs(9476)));
    outputs(8315) <= layer2_outputs(5928);
    outputs(8316) <= (layer2_outputs(6714)) and not (layer2_outputs(9677));
    outputs(8317) <= (layer2_outputs(2208)) xor (layer2_outputs(4968));
    outputs(8318) <= (layer2_outputs(7331)) xor (layer2_outputs(10008));
    outputs(8319) <= '1';
    outputs(8320) <= not((layer2_outputs(4591)) xor (layer2_outputs(6576)));
    outputs(8321) <= layer2_outputs(8775);
    outputs(8322) <= (layer2_outputs(1788)) xor (layer2_outputs(3300));
    outputs(8323) <= not(layer2_outputs(2305));
    outputs(8324) <= layer2_outputs(971);
    outputs(8325) <= layer2_outputs(8319);
    outputs(8326) <= not(layer2_outputs(9020)) or (layer2_outputs(6421));
    outputs(8327) <= (layer2_outputs(6126)) and not (layer2_outputs(6827));
    outputs(8328) <= not((layer2_outputs(6443)) xor (layer2_outputs(4667)));
    outputs(8329) <= (layer2_outputs(3352)) or (layer2_outputs(4578));
    outputs(8330) <= not(layer2_outputs(4619)) or (layer2_outputs(4350));
    outputs(8331) <= (layer2_outputs(3362)) xor (layer2_outputs(1351));
    outputs(8332) <= layer2_outputs(2385);
    outputs(8333) <= layer2_outputs(7763);
    outputs(8334) <= (layer2_outputs(8832)) xor (layer2_outputs(9739));
    outputs(8335) <= not(layer2_outputs(7707)) or (layer2_outputs(724));
    outputs(8336) <= not(layer2_outputs(9211)) or (layer2_outputs(5407));
    outputs(8337) <= (layer2_outputs(5936)) and not (layer2_outputs(8758));
    outputs(8338) <= (layer2_outputs(8224)) or (layer2_outputs(3486));
    outputs(8339) <= not(layer2_outputs(7919));
    outputs(8340) <= not((layer2_outputs(6369)) xor (layer2_outputs(1935)));
    outputs(8341) <= layer2_outputs(4673);
    outputs(8342) <= not(layer2_outputs(9386)) or (layer2_outputs(7503));
    outputs(8343) <= layer2_outputs(8072);
    outputs(8344) <= (layer2_outputs(5130)) xor (layer2_outputs(346));
    outputs(8345) <= not((layer2_outputs(8987)) and (layer2_outputs(185)));
    outputs(8346) <= not((layer2_outputs(9973)) xor (layer2_outputs(6969)));
    outputs(8347) <= not(layer2_outputs(8195)) or (layer2_outputs(5131));
    outputs(8348) <= not(layer2_outputs(328));
    outputs(8349) <= not(layer2_outputs(4108));
    outputs(8350) <= not((layer2_outputs(6706)) or (layer2_outputs(2168)));
    outputs(8351) <= not(layer2_outputs(9166));
    outputs(8352) <= not(layer2_outputs(9073)) or (layer2_outputs(8680));
    outputs(8353) <= (layer2_outputs(7321)) xor (layer2_outputs(7270));
    outputs(8354) <= (layer2_outputs(7252)) or (layer2_outputs(3585));
    outputs(8355) <= (layer2_outputs(37)) xor (layer2_outputs(7127));
    outputs(8356) <= (layer2_outputs(1969)) xor (layer2_outputs(9481));
    outputs(8357) <= (layer2_outputs(1929)) xor (layer2_outputs(3768));
    outputs(8358) <= not(layer2_outputs(862)) or (layer2_outputs(4868));
    outputs(8359) <= not((layer2_outputs(9675)) and (layer2_outputs(2989)));
    outputs(8360) <= not((layer2_outputs(10135)) xor (layer2_outputs(585)));
    outputs(8361) <= (layer2_outputs(5307)) xor (layer2_outputs(1358));
    outputs(8362) <= layer2_outputs(6419);
    outputs(8363) <= not(layer2_outputs(7094));
    outputs(8364) <= (layer2_outputs(6012)) and not (layer2_outputs(3227));
    outputs(8365) <= layer2_outputs(3848);
    outputs(8366) <= not((layer2_outputs(3245)) and (layer2_outputs(3650)));
    outputs(8367) <= layer2_outputs(9628);
    outputs(8368) <= (layer2_outputs(5946)) xor (layer2_outputs(1684));
    outputs(8369) <= not(layer2_outputs(9371));
    outputs(8370) <= (layer2_outputs(7238)) xor (layer2_outputs(7423));
    outputs(8371) <= (layer2_outputs(844)) xor (layer2_outputs(8467));
    outputs(8372) <= (layer2_outputs(120)) and (layer2_outputs(6066));
    outputs(8373) <= layer2_outputs(6378);
    outputs(8374) <= (layer2_outputs(10175)) xor (layer2_outputs(6321));
    outputs(8375) <= not(layer2_outputs(7762)) or (layer2_outputs(2206));
    outputs(8376) <= not((layer2_outputs(7870)) or (layer2_outputs(6870)));
    outputs(8377) <= not(layer2_outputs(529));
    outputs(8378) <= layer2_outputs(5441);
    outputs(8379) <= (layer2_outputs(4435)) xor (layer2_outputs(622));
    outputs(8380) <= not(layer2_outputs(8043));
    outputs(8381) <= (layer2_outputs(2596)) xor (layer2_outputs(1323));
    outputs(8382) <= layer2_outputs(843);
    outputs(8383) <= layer2_outputs(8396);
    outputs(8384) <= layer2_outputs(4869);
    outputs(8385) <= (layer2_outputs(7146)) xor (layer2_outputs(10212));
    outputs(8386) <= layer2_outputs(9487);
    outputs(8387) <= (layer2_outputs(9352)) and (layer2_outputs(8663));
    outputs(8388) <= (layer2_outputs(2099)) and not (layer2_outputs(209));
    outputs(8389) <= not(layer2_outputs(4902));
    outputs(8390) <= not(layer2_outputs(4218));
    outputs(8391) <= not((layer2_outputs(1812)) xor (layer2_outputs(7876)));
    outputs(8392) <= not(layer2_outputs(367));
    outputs(8393) <= layer2_outputs(800);
    outputs(8394) <= not((layer2_outputs(3990)) xor (layer2_outputs(138)));
    outputs(8395) <= (layer2_outputs(3055)) xor (layer2_outputs(7395));
    outputs(8396) <= not((layer2_outputs(10233)) xor (layer2_outputs(9180)));
    outputs(8397) <= not(layer2_outputs(9503));
    outputs(8398) <= (layer2_outputs(2631)) or (layer2_outputs(2574));
    outputs(8399) <= not((layer2_outputs(1688)) xor (layer2_outputs(5245)));
    outputs(8400) <= (layer2_outputs(9546)) and (layer2_outputs(8246));
    outputs(8401) <= layer2_outputs(7588);
    outputs(8402) <= layer2_outputs(4659);
    outputs(8403) <= (layer2_outputs(8725)) and not (layer2_outputs(2180));
    outputs(8404) <= layer2_outputs(6529);
    outputs(8405) <= layer2_outputs(2242);
    outputs(8406) <= layer2_outputs(3951);
    outputs(8407) <= not(layer2_outputs(7452)) or (layer2_outputs(5875));
    outputs(8408) <= (layer2_outputs(520)) and not (layer2_outputs(6003));
    outputs(8409) <= not(layer2_outputs(942)) or (layer2_outputs(9764));
    outputs(8410) <= layer2_outputs(6672);
    outputs(8411) <= (layer2_outputs(7618)) xor (layer2_outputs(1002));
    outputs(8412) <= not((layer2_outputs(9981)) xor (layer2_outputs(8733)));
    outputs(8413) <= layer2_outputs(1690);
    outputs(8414) <= not(layer2_outputs(131)) or (layer2_outputs(1452));
    outputs(8415) <= layer2_outputs(4110);
    outputs(8416) <= (layer2_outputs(9719)) xor (layer2_outputs(862));
    outputs(8417) <= not(layer2_outputs(6980));
    outputs(8418) <= (layer2_outputs(9422)) xor (layer2_outputs(3373));
    outputs(8419) <= not(layer2_outputs(7756)) or (layer2_outputs(3254));
    outputs(8420) <= (layer2_outputs(7131)) xor (layer2_outputs(7212));
    outputs(8421) <= layer2_outputs(7654);
    outputs(8422) <= not(layer2_outputs(917)) or (layer2_outputs(3605));
    outputs(8423) <= not((layer2_outputs(6561)) xor (layer2_outputs(7258)));
    outputs(8424) <= not(layer2_outputs(4545));
    outputs(8425) <= layer2_outputs(7540);
    outputs(8426) <= layer2_outputs(7517);
    outputs(8427) <= layer2_outputs(9843);
    outputs(8428) <= (layer2_outputs(7261)) xor (layer2_outputs(1463));
    outputs(8429) <= not(layer2_outputs(9970));
    outputs(8430) <= not(layer2_outputs(8023));
    outputs(8431) <= layer2_outputs(2207);
    outputs(8432) <= (layer2_outputs(3081)) xor (layer2_outputs(4966));
    outputs(8433) <= not(layer2_outputs(9949));
    outputs(8434) <= not(layer2_outputs(8405)) or (layer2_outputs(2156));
    outputs(8435) <= not((layer2_outputs(184)) and (layer2_outputs(1584)));
    outputs(8436) <= not(layer2_outputs(1829));
    outputs(8437) <= not(layer2_outputs(9804));
    outputs(8438) <= not(layer2_outputs(6160)) or (layer2_outputs(8254));
    outputs(8439) <= layer2_outputs(2747);
    outputs(8440) <= layer2_outputs(296);
    outputs(8441) <= (layer2_outputs(678)) xor (layer2_outputs(4446));
    outputs(8442) <= not((layer2_outputs(9269)) or (layer2_outputs(4396)));
    outputs(8443) <= layer2_outputs(9777);
    outputs(8444) <= not(layer2_outputs(4700)) or (layer2_outputs(932));
    outputs(8445) <= not((layer2_outputs(7567)) xor (layer2_outputs(7230)));
    outputs(8446) <= not(layer2_outputs(4981));
    outputs(8447) <= not(layer2_outputs(7762));
    outputs(8448) <= not((layer2_outputs(7820)) xor (layer2_outputs(7231)));
    outputs(8449) <= not(layer2_outputs(4573));
    outputs(8450) <= not((layer2_outputs(3581)) xor (layer2_outputs(5730)));
    outputs(8451) <= '1';
    outputs(8452) <= layer2_outputs(4544);
    outputs(8453) <= not((layer2_outputs(6953)) xor (layer2_outputs(4070)));
    outputs(8454) <= layer2_outputs(9541);
    outputs(8455) <= layer2_outputs(506);
    outputs(8456) <= layer2_outputs(669);
    outputs(8457) <= not(layer2_outputs(6362));
    outputs(8458) <= not((layer2_outputs(5111)) and (layer2_outputs(7231)));
    outputs(8459) <= layer2_outputs(5600);
    outputs(8460) <= (layer2_outputs(1207)) xor (layer2_outputs(4495));
    outputs(8461) <= layer2_outputs(5464);
    outputs(8462) <= layer2_outputs(8206);
    outputs(8463) <= not(layer2_outputs(5824));
    outputs(8464) <= not(layer2_outputs(7748));
    outputs(8465) <= not(layer2_outputs(4691));
    outputs(8466) <= not(layer2_outputs(642)) or (layer2_outputs(83));
    outputs(8467) <= layer2_outputs(5508);
    outputs(8468) <= not(layer2_outputs(841));
    outputs(8469) <= (layer2_outputs(3327)) and not (layer2_outputs(9972));
    outputs(8470) <= layer2_outputs(4567);
    outputs(8471) <= layer2_outputs(1177);
    outputs(8472) <= layer2_outputs(4354);
    outputs(8473) <= not(layer2_outputs(6377)) or (layer2_outputs(4313));
    outputs(8474) <= layer2_outputs(6030);
    outputs(8475) <= not((layer2_outputs(7147)) xor (layer2_outputs(1594)));
    outputs(8476) <= (layer2_outputs(4322)) xor (layer2_outputs(625));
    outputs(8477) <= layer2_outputs(771);
    outputs(8478) <= layer2_outputs(6865);
    outputs(8479) <= not(layer2_outputs(207));
    outputs(8480) <= not(layer2_outputs(1999));
    outputs(8481) <= not(layer2_outputs(8920));
    outputs(8482) <= (layer2_outputs(5624)) or (layer2_outputs(2904));
    outputs(8483) <= not((layer2_outputs(4621)) or (layer2_outputs(9514)));
    outputs(8484) <= not(layer2_outputs(3385));
    outputs(8485) <= not(layer2_outputs(10060));
    outputs(8486) <= not(layer2_outputs(6437));
    outputs(8487) <= not((layer2_outputs(6604)) xor (layer2_outputs(7158)));
    outputs(8488) <= layer2_outputs(144);
    outputs(8489) <= (layer2_outputs(750)) and not (layer2_outputs(3257));
    outputs(8490) <= (layer2_outputs(5161)) and not (layer2_outputs(5491));
    outputs(8491) <= not(layer2_outputs(6855));
    outputs(8492) <= not(layer2_outputs(8128));
    outputs(8493) <= layer2_outputs(6366);
    outputs(8494) <= not((layer2_outputs(2123)) or (layer2_outputs(3711)));
    outputs(8495) <= not(layer2_outputs(3846));
    outputs(8496) <= not((layer2_outputs(3039)) xor (layer2_outputs(6082)));
    outputs(8497) <= layer2_outputs(9785);
    outputs(8498) <= layer2_outputs(8078);
    outputs(8499) <= not(layer2_outputs(4720));
    outputs(8500) <= not(layer2_outputs(5792));
    outputs(8501) <= not(layer2_outputs(9406));
    outputs(8502) <= (layer2_outputs(7766)) or (layer2_outputs(250));
    outputs(8503) <= not(layer2_outputs(9817)) or (layer2_outputs(1446));
    outputs(8504) <= not(layer2_outputs(2261));
    outputs(8505) <= (layer2_outputs(3876)) or (layer2_outputs(1412));
    outputs(8506) <= not(layer2_outputs(4499)) or (layer2_outputs(2803));
    outputs(8507) <= layer2_outputs(3123);
    outputs(8508) <= layer2_outputs(5503);
    outputs(8509) <= not((layer2_outputs(8449)) and (layer2_outputs(7021)));
    outputs(8510) <= not(layer2_outputs(1934));
    outputs(8511) <= not(layer2_outputs(6203));
    outputs(8512) <= (layer2_outputs(8410)) xor (layer2_outputs(9402));
    outputs(8513) <= layer2_outputs(2092);
    outputs(8514) <= not((layer2_outputs(7338)) xor (layer2_outputs(4679)));
    outputs(8515) <= not(layer2_outputs(6457));
    outputs(8516) <= (layer2_outputs(7525)) and not (layer2_outputs(3245));
    outputs(8517) <= not((layer2_outputs(2930)) xor (layer2_outputs(5538)));
    outputs(8518) <= not(layer2_outputs(3603));
    outputs(8519) <= (layer2_outputs(4640)) xor (layer2_outputs(3708));
    outputs(8520) <= not(layer2_outputs(9225));
    outputs(8521) <= not((layer2_outputs(5925)) xor (layer2_outputs(945)));
    outputs(8522) <= layer2_outputs(3267);
    outputs(8523) <= not(layer2_outputs(3786));
    outputs(8524) <= not((layer2_outputs(8387)) xor (layer2_outputs(8512)));
    outputs(8525) <= not(layer2_outputs(5970));
    outputs(8526) <= not((layer2_outputs(6554)) xor (layer2_outputs(976)));
    outputs(8527) <= not((layer2_outputs(1947)) xor (layer2_outputs(6649)));
    outputs(8528) <= not(layer2_outputs(2998));
    outputs(8529) <= layer2_outputs(6098);
    outputs(8530) <= layer2_outputs(3795);
    outputs(8531) <= (layer2_outputs(1230)) xor (layer2_outputs(5507));
    outputs(8532) <= (layer2_outputs(5797)) xor (layer2_outputs(2548));
    outputs(8533) <= layer2_outputs(4929);
    outputs(8534) <= not(layer2_outputs(4427));
    outputs(8535) <= not((layer2_outputs(2820)) xor (layer2_outputs(2755)));
    outputs(8536) <= not(layer2_outputs(7313));
    outputs(8537) <= not(layer2_outputs(4665)) or (layer2_outputs(6429));
    outputs(8538) <= not((layer2_outputs(7264)) xor (layer2_outputs(4312)));
    outputs(8539) <= not(layer2_outputs(4365));
    outputs(8540) <= not(layer2_outputs(8932));
    outputs(8541) <= not(layer2_outputs(8047)) or (layer2_outputs(7383));
    outputs(8542) <= (layer2_outputs(10104)) or (layer2_outputs(6351));
    outputs(8543) <= layer2_outputs(6410);
    outputs(8544) <= (layer2_outputs(7413)) xor (layer2_outputs(6483));
    outputs(8545) <= not((layer2_outputs(6370)) xor (layer2_outputs(7413)));
    outputs(8546) <= not(layer2_outputs(8790));
    outputs(8547) <= not(layer2_outputs(4275)) or (layer2_outputs(5565));
    outputs(8548) <= not((layer2_outputs(1148)) xor (layer2_outputs(665)));
    outputs(8549) <= (layer2_outputs(1892)) or (layer2_outputs(2636));
    outputs(8550) <= not((layer2_outputs(7550)) xor (layer2_outputs(7371)));
    outputs(8551) <= layer2_outputs(9515);
    outputs(8552) <= not((layer2_outputs(2701)) xor (layer2_outputs(4920)));
    outputs(8553) <= (layer2_outputs(6658)) xor (layer2_outputs(8380));
    outputs(8554) <= layer2_outputs(1861);
    outputs(8555) <= not((layer2_outputs(8661)) xor (layer2_outputs(4329)));
    outputs(8556) <= not(layer2_outputs(2028));
    outputs(8557) <= not(layer2_outputs(9298));
    outputs(8558) <= not(layer2_outputs(4970));
    outputs(8559) <= (layer2_outputs(5205)) xor (layer2_outputs(5017));
    outputs(8560) <= not((layer2_outputs(3214)) and (layer2_outputs(9081)));
    outputs(8561) <= not(layer2_outputs(3090));
    outputs(8562) <= layer2_outputs(714);
    outputs(8563) <= not(layer2_outputs(2460));
    outputs(8564) <= not(layer2_outputs(4603)) or (layer2_outputs(5225));
    outputs(8565) <= layer2_outputs(284);
    outputs(8566) <= not(layer2_outputs(9408));
    outputs(8567) <= not(layer2_outputs(2797));
    outputs(8568) <= not((layer2_outputs(3754)) and (layer2_outputs(6978)));
    outputs(8569) <= not(layer2_outputs(1691));
    outputs(8570) <= not(layer2_outputs(10010));
    outputs(8571) <= not((layer2_outputs(9506)) and (layer2_outputs(8685)));
    outputs(8572) <= not(layer2_outputs(2685));
    outputs(8573) <= layer2_outputs(4856);
    outputs(8574) <= layer2_outputs(8604);
    outputs(8575) <= not(layer2_outputs(9172)) or (layer2_outputs(5));
    outputs(8576) <= not(layer2_outputs(6183));
    outputs(8577) <= layer2_outputs(703);
    outputs(8578) <= not(layer2_outputs(6006));
    outputs(8579) <= layer2_outputs(2988);
    outputs(8580) <= not((layer2_outputs(6178)) and (layer2_outputs(5543)));
    outputs(8581) <= (layer2_outputs(4780)) xor (layer2_outputs(3795));
    outputs(8582) <= not((layer2_outputs(8478)) xor (layer2_outputs(5262)));
    outputs(8583) <= layer2_outputs(5007);
    outputs(8584) <= layer2_outputs(6408);
    outputs(8585) <= not(layer2_outputs(6742));
    outputs(8586) <= not((layer2_outputs(2564)) and (layer2_outputs(4927)));
    outputs(8587) <= (layer2_outputs(6080)) xor (layer2_outputs(4216));
    outputs(8588) <= not(layer2_outputs(4658)) or (layer2_outputs(9075));
    outputs(8589) <= (layer2_outputs(1548)) xor (layer2_outputs(5837));
    outputs(8590) <= not((layer2_outputs(3074)) xor (layer2_outputs(4878)));
    outputs(8591) <= not((layer2_outputs(1832)) and (layer2_outputs(7051)));
    outputs(8592) <= layer2_outputs(4618);
    outputs(8593) <= layer2_outputs(6091);
    outputs(8594) <= layer2_outputs(6815);
    outputs(8595) <= not(layer2_outputs(6074)) or (layer2_outputs(1037));
    outputs(8596) <= not(layer2_outputs(3820));
    outputs(8597) <= layer2_outputs(9495);
    outputs(8598) <= not((layer2_outputs(9224)) xor (layer2_outputs(2074)));
    outputs(8599) <= layer2_outputs(1308);
    outputs(8600) <= (layer2_outputs(7160)) xor (layer2_outputs(3920));
    outputs(8601) <= not(layer2_outputs(8551));
    outputs(8602) <= not(layer2_outputs(7248)) or (layer2_outputs(8961));
    outputs(8603) <= not(layer2_outputs(5211));
    outputs(8604) <= layer2_outputs(2417);
    outputs(8605) <= layer2_outputs(4546);
    outputs(8606) <= layer2_outputs(29);
    outputs(8607) <= layer2_outputs(9535);
    outputs(8608) <= layer2_outputs(404);
    outputs(8609) <= (layer2_outputs(299)) and not (layer2_outputs(6812));
    outputs(8610) <= not(layer2_outputs(3976));
    outputs(8611) <= (layer2_outputs(7609)) xor (layer2_outputs(4343));
    outputs(8612) <= not(layer2_outputs(5011)) or (layer2_outputs(4171));
    outputs(8613) <= not(layer2_outputs(4239));
    outputs(8614) <= not(layer2_outputs(6974));
    outputs(8615) <= (layer2_outputs(85)) xor (layer2_outputs(1864));
    outputs(8616) <= (layer2_outputs(9896)) xor (layer2_outputs(2805));
    outputs(8617) <= layer2_outputs(5670);
    outputs(8618) <= layer2_outputs(3937);
    outputs(8619) <= layer2_outputs(8614);
    outputs(8620) <= not(layer2_outputs(492));
    outputs(8621) <= (layer2_outputs(6010)) xor (layer2_outputs(2718));
    outputs(8622) <= (layer2_outputs(7595)) or (layer2_outputs(1327));
    outputs(8623) <= not(layer2_outputs(9745));
    outputs(8624) <= not(layer2_outputs(2114)) or (layer2_outputs(108));
    outputs(8625) <= not(layer2_outputs(786));
    outputs(8626) <= not((layer2_outputs(9328)) and (layer2_outputs(3106)));
    outputs(8627) <= not((layer2_outputs(6361)) xor (layer2_outputs(7318)));
    outputs(8628) <= not(layer2_outputs(8200));
    outputs(8629) <= not(layer2_outputs(9013));
    outputs(8630) <= not(layer2_outputs(818));
    outputs(8631) <= layer2_outputs(3162);
    outputs(8632) <= not((layer2_outputs(3673)) xor (layer2_outputs(7965)));
    outputs(8633) <= not((layer2_outputs(9512)) xor (layer2_outputs(3628)));
    outputs(8634) <= (layer2_outputs(1891)) xor (layer2_outputs(9714));
    outputs(8635) <= '1';
    outputs(8636) <= (layer2_outputs(2945)) xor (layer2_outputs(10111));
    outputs(8637) <= not((layer2_outputs(6329)) xor (layer2_outputs(3774)));
    outputs(8638) <= not(layer2_outputs(6226));
    outputs(8639) <= not((layer2_outputs(8147)) xor (layer2_outputs(6677)));
    outputs(8640) <= layer2_outputs(4878);
    outputs(8641) <= layer2_outputs(2452);
    outputs(8642) <= not(layer2_outputs(5729)) or (layer2_outputs(7190));
    outputs(8643) <= not((layer2_outputs(9737)) xor (layer2_outputs(4349)));
    outputs(8644) <= not(layer2_outputs(7447));
    outputs(8645) <= layer2_outputs(6474);
    outputs(8646) <= not(layer2_outputs(2142));
    outputs(8647) <= layer2_outputs(10218);
    outputs(8648) <= (layer2_outputs(3652)) xor (layer2_outputs(3393));
    outputs(8649) <= not(layer2_outputs(2138));
    outputs(8650) <= (layer2_outputs(9634)) or (layer2_outputs(4249));
    outputs(8651) <= layer2_outputs(9353);
    outputs(8652) <= layer2_outputs(5249);
    outputs(8653) <= not(layer2_outputs(5260));
    outputs(8654) <= not(layer2_outputs(1464));
    outputs(8655) <= not((layer2_outputs(4103)) and (layer2_outputs(3015)));
    outputs(8656) <= not((layer2_outputs(3032)) xor (layer2_outputs(3249)));
    outputs(8657) <= (layer2_outputs(4000)) xor (layer2_outputs(2547));
    outputs(8658) <= layer2_outputs(6268);
    outputs(8659) <= not(layer2_outputs(10026));
    outputs(8660) <= not(layer2_outputs(7455));
    outputs(8661) <= layer2_outputs(2954);
    outputs(8662) <= (layer2_outputs(4964)) or (layer2_outputs(3577));
    outputs(8663) <= not(layer2_outputs(4326));
    outputs(8664) <= not(layer2_outputs(3860));
    outputs(8665) <= layer2_outputs(1760);
    outputs(8666) <= layer2_outputs(318);
    outputs(8667) <= layer2_outputs(2162);
    outputs(8668) <= (layer2_outputs(7812)) xor (layer2_outputs(9728));
    outputs(8669) <= not((layer2_outputs(1121)) xor (layer2_outputs(5614)));
    outputs(8670) <= not(layer2_outputs(5349));
    outputs(8671) <= (layer2_outputs(121)) and not (layer2_outputs(3487));
    outputs(8672) <= '0';
    outputs(8673) <= not(layer2_outputs(5256));
    outputs(8674) <= not(layer2_outputs(1750));
    outputs(8675) <= not(layer2_outputs(9938));
    outputs(8676) <= layer2_outputs(1578);
    outputs(8677) <= not((layer2_outputs(2442)) or (layer2_outputs(472)));
    outputs(8678) <= not(layer2_outputs(6382));
    outputs(8679) <= layer2_outputs(8045);
    outputs(8680) <= not((layer2_outputs(1841)) xor (layer2_outputs(3213)));
    outputs(8681) <= (layer2_outputs(2306)) xor (layer2_outputs(9617));
    outputs(8682) <= (layer2_outputs(160)) xor (layer2_outputs(6818));
    outputs(8683) <= layer2_outputs(5259);
    outputs(8684) <= not((layer2_outputs(4853)) xor (layer2_outputs(561)));
    outputs(8685) <= not((layer2_outputs(7410)) xor (layer2_outputs(2707)));
    outputs(8686) <= not(layer2_outputs(4555));
    outputs(8687) <= layer2_outputs(6494);
    outputs(8688) <= not((layer2_outputs(2415)) or (layer2_outputs(6456)));
    outputs(8689) <= not(layer2_outputs(7953));
    outputs(8690) <= layer2_outputs(9157);
    outputs(8691) <= layer2_outputs(7833);
    outputs(8692) <= not((layer2_outputs(1876)) xor (layer2_outputs(4934)));
    outputs(8693) <= not(layer2_outputs(4304));
    outputs(8694) <= not((layer2_outputs(4052)) and (layer2_outputs(8625)));
    outputs(8695) <= not(layer2_outputs(2082));
    outputs(8696) <= not((layer2_outputs(1852)) xor (layer2_outputs(916)));
    outputs(8697) <= not(layer2_outputs(9635));
    outputs(8698) <= not(layer2_outputs(6928));
    outputs(8699) <= not(layer2_outputs(4333));
    outputs(8700) <= not((layer2_outputs(8675)) xor (layer2_outputs(8104)));
    outputs(8701) <= not(layer2_outputs(10160));
    outputs(8702) <= not(layer2_outputs(472));
    outputs(8703) <= not(layer2_outputs(10046));
    outputs(8704) <= (layer2_outputs(3256)) and not (layer2_outputs(5267));
    outputs(8705) <= not((layer2_outputs(2895)) xor (layer2_outputs(4655)));
    outputs(8706) <= not(layer2_outputs(5862));
    outputs(8707) <= not(layer2_outputs(9647)) or (layer2_outputs(6468));
    outputs(8708) <= not(layer2_outputs(2235));
    outputs(8709) <= layer2_outputs(912);
    outputs(8710) <= not(layer2_outputs(7719));
    outputs(8711) <= not(layer2_outputs(682)) or (layer2_outputs(923));
    outputs(8712) <= not((layer2_outputs(8787)) xor (layer2_outputs(1972)));
    outputs(8713) <= not((layer2_outputs(4034)) xor (layer2_outputs(964)));
    outputs(8714) <= not(layer2_outputs(5274));
    outputs(8715) <= not((layer2_outputs(1183)) xor (layer2_outputs(1233)));
    outputs(8716) <= not(layer2_outputs(709));
    outputs(8717) <= (layer2_outputs(9725)) xor (layer2_outputs(6578));
    outputs(8718) <= (layer2_outputs(1178)) xor (layer2_outputs(1071));
    outputs(8719) <= layer2_outputs(1007);
    outputs(8720) <= layer2_outputs(2203);
    outputs(8721) <= not((layer2_outputs(4238)) and (layer2_outputs(704)));
    outputs(8722) <= not(layer2_outputs(7504));
    outputs(8723) <= not(layer2_outputs(2003));
    outputs(8724) <= not((layer2_outputs(4488)) xor (layer2_outputs(5731)));
    outputs(8725) <= (layer2_outputs(2747)) and not (layer2_outputs(8239));
    outputs(8726) <= layer2_outputs(4663);
    outputs(8727) <= layer2_outputs(8215);
    outputs(8728) <= layer2_outputs(513);
    outputs(8729) <= layer2_outputs(5041);
    outputs(8730) <= not(layer2_outputs(6517));
    outputs(8731) <= layer2_outputs(7714);
    outputs(8732) <= not(layer2_outputs(4895));
    outputs(8733) <= not(layer2_outputs(1426));
    outputs(8734) <= (layer2_outputs(4413)) xor (layer2_outputs(1501));
    outputs(8735) <= layer2_outputs(47);
    outputs(8736) <= layer2_outputs(9114);
    outputs(8737) <= layer2_outputs(5192);
    outputs(8738) <= not(layer2_outputs(4984));
    outputs(8739) <= layer2_outputs(3359);
    outputs(8740) <= not(layer2_outputs(10070));
    outputs(8741) <= not(layer2_outputs(4536));
    outputs(8742) <= not(layer2_outputs(860));
    outputs(8743) <= not((layer2_outputs(5961)) and (layer2_outputs(8631)));
    outputs(8744) <= (layer2_outputs(7833)) or (layer2_outputs(4195));
    outputs(8745) <= layer2_outputs(5879);
    outputs(8746) <= not(layer2_outputs(8779)) or (layer2_outputs(7119));
    outputs(8747) <= (layer2_outputs(4)) xor (layer2_outputs(9891));
    outputs(8748) <= not(layer2_outputs(157));
    outputs(8749) <= not(layer2_outputs(2815));
    outputs(8750) <= (layer2_outputs(8977)) xor (layer2_outputs(725));
    outputs(8751) <= not(layer2_outputs(5912));
    outputs(8752) <= (layer2_outputs(7653)) xor (layer2_outputs(7586));
    outputs(8753) <= (layer2_outputs(7563)) or (layer2_outputs(8353));
    outputs(8754) <= (layer2_outputs(6299)) and not (layer2_outputs(9885));
    outputs(8755) <= not(layer2_outputs(366));
    outputs(8756) <= not(layer2_outputs(8761));
    outputs(8757) <= not(layer2_outputs(7642));
    outputs(8758) <= layer2_outputs(8513);
    outputs(8759) <= (layer2_outputs(10007)) xor (layer2_outputs(1448));
    outputs(8760) <= not(layer2_outputs(1384));
    outputs(8761) <= (layer2_outputs(747)) or (layer2_outputs(7274));
    outputs(8762) <= (layer2_outputs(10020)) xor (layer2_outputs(2572));
    outputs(8763) <= not((layer2_outputs(3097)) xor (layer2_outputs(4629)));
    outputs(8764) <= not(layer2_outputs(9075)) or (layer2_outputs(1607));
    outputs(8765) <= not(layer2_outputs(4026));
    outputs(8766) <= (layer2_outputs(885)) xor (layer2_outputs(909));
    outputs(8767) <= (layer2_outputs(6948)) and (layer2_outputs(4913));
    outputs(8768) <= not(layer2_outputs(4555));
    outputs(8769) <= not(layer2_outputs(3913));
    outputs(8770) <= layer2_outputs(1319);
    outputs(8771) <= not((layer2_outputs(8884)) xor (layer2_outputs(4680)));
    outputs(8772) <= not((layer2_outputs(8305)) and (layer2_outputs(657)));
    outputs(8773) <= (layer2_outputs(8355)) xor (layer2_outputs(6543));
    outputs(8774) <= layer2_outputs(256);
    outputs(8775) <= (layer2_outputs(8362)) xor (layer2_outputs(4199));
    outputs(8776) <= layer2_outputs(7776);
    outputs(8777) <= (layer2_outputs(9471)) xor (layer2_outputs(8457));
    outputs(8778) <= (layer2_outputs(3286)) xor (layer2_outputs(3208));
    outputs(8779) <= not((layer2_outputs(4919)) xor (layer2_outputs(7922)));
    outputs(8780) <= (layer2_outputs(99)) and not (layer2_outputs(5634));
    outputs(8781) <= (layer2_outputs(7674)) or (layer2_outputs(6997));
    outputs(8782) <= '0';
    outputs(8783) <= (layer2_outputs(4018)) xor (layer2_outputs(8156));
    outputs(8784) <= not(layer2_outputs(5100));
    outputs(8785) <= layer2_outputs(8072);
    outputs(8786) <= not(layer2_outputs(9604)) or (layer2_outputs(1363));
    outputs(8787) <= (layer2_outputs(7071)) or (layer2_outputs(5138));
    outputs(8788) <= not((layer2_outputs(6141)) xor (layer2_outputs(6662)));
    outputs(8789) <= layer2_outputs(6505);
    outputs(8790) <= not(layer2_outputs(4737));
    outputs(8791) <= not((layer2_outputs(9214)) xor (layer2_outputs(9274)));
    outputs(8792) <= layer2_outputs(3328);
    outputs(8793) <= not(layer2_outputs(4484));
    outputs(8794) <= not(layer2_outputs(3130));
    outputs(8795) <= not(layer2_outputs(9186));
    outputs(8796) <= layer2_outputs(325);
    outputs(8797) <= (layer2_outputs(8276)) and not (layer2_outputs(9111));
    outputs(8798) <= (layer2_outputs(6903)) xor (layer2_outputs(6210));
    outputs(8799) <= not(layer2_outputs(7724)) or (layer2_outputs(6138));
    outputs(8800) <= layer2_outputs(312);
    outputs(8801) <= not((layer2_outputs(8859)) xor (layer2_outputs(5306)));
    outputs(8802) <= not((layer2_outputs(8989)) xor (layer2_outputs(9813)));
    outputs(8803) <= not(layer2_outputs(3195));
    outputs(8804) <= layer2_outputs(9239);
    outputs(8805) <= not(layer2_outputs(3198)) or (layer2_outputs(6571));
    outputs(8806) <= layer2_outputs(5693);
    outputs(8807) <= (layer2_outputs(7218)) xor (layer2_outputs(3681));
    outputs(8808) <= not(layer2_outputs(4520));
    outputs(8809) <= not(layer2_outputs(6480));
    outputs(8810) <= not(layer2_outputs(9822));
    outputs(8811) <= not(layer2_outputs(5943));
    outputs(8812) <= not((layer2_outputs(4242)) or (layer2_outputs(252)));
    outputs(8813) <= layer2_outputs(877);
    outputs(8814) <= (layer2_outputs(5964)) xor (layer2_outputs(2321));
    outputs(8815) <= layer2_outputs(6021);
    outputs(8816) <= (layer2_outputs(7084)) and not (layer2_outputs(3347));
    outputs(8817) <= (layer2_outputs(3807)) or (layer2_outputs(4822));
    outputs(8818) <= not(layer2_outputs(4313)) or (layer2_outputs(1494));
    outputs(8819) <= not(layer2_outputs(9185));
    outputs(8820) <= not((layer2_outputs(7409)) xor (layer2_outputs(9417)));
    outputs(8821) <= layer2_outputs(4494);
    outputs(8822) <= '1';
    outputs(8823) <= not(layer2_outputs(1371));
    outputs(8824) <= layer2_outputs(5504);
    outputs(8825) <= not(layer2_outputs(4196));
    outputs(8826) <= not((layer2_outputs(194)) or (layer2_outputs(9731)));
    outputs(8827) <= not(layer2_outputs(1372));
    outputs(8828) <= not((layer2_outputs(6355)) xor (layer2_outputs(5166)));
    outputs(8829) <= not(layer2_outputs(2378));
    outputs(8830) <= not(layer2_outputs(9424));
    outputs(8831) <= layer2_outputs(9244);
    outputs(8832) <= layer2_outputs(3192);
    outputs(8833) <= layer2_outputs(981);
    outputs(8834) <= not((layer2_outputs(10018)) xor (layer2_outputs(2060)));
    outputs(8835) <= (layer2_outputs(38)) and (layer2_outputs(4194));
    outputs(8836) <= not(layer2_outputs(8784));
    outputs(8837) <= (layer2_outputs(4966)) or (layer2_outputs(2850));
    outputs(8838) <= not((layer2_outputs(2049)) or (layer2_outputs(536)));
    outputs(8839) <= (layer2_outputs(4582)) xor (layer2_outputs(6327));
    outputs(8840) <= not(layer2_outputs(1906));
    outputs(8841) <= layer2_outputs(9198);
    outputs(8842) <= layer2_outputs(7701);
    outputs(8843) <= not(layer2_outputs(4387));
    outputs(8844) <= layer2_outputs(4473);
    outputs(8845) <= not(layer2_outputs(7787));
    outputs(8846) <= not(layer2_outputs(4461)) or (layer2_outputs(6675));
    outputs(8847) <= layer2_outputs(3091);
    outputs(8848) <= layer2_outputs(1370);
    outputs(8849) <= layer2_outputs(2567);
    outputs(8850) <= not((layer2_outputs(1505)) xor (layer2_outputs(9127)));
    outputs(8851) <= not(layer2_outputs(4877));
    outputs(8852) <= (layer2_outputs(3889)) and not (layer2_outputs(6229));
    outputs(8853) <= (layer2_outputs(3160)) xor (layer2_outputs(5878));
    outputs(8854) <= not(layer2_outputs(6266));
    outputs(8855) <= layer2_outputs(10120);
    outputs(8856) <= not(layer2_outputs(5753));
    outputs(8857) <= not((layer2_outputs(2303)) xor (layer2_outputs(2275)));
    outputs(8858) <= not((layer2_outputs(9848)) and (layer2_outputs(3587)));
    outputs(8859) <= layer2_outputs(4175);
    outputs(8860) <= (layer2_outputs(4640)) xor (layer2_outputs(2209));
    outputs(8861) <= layer2_outputs(6769);
    outputs(8862) <= (layer2_outputs(8824)) xor (layer2_outputs(7880));
    outputs(8863) <= not((layer2_outputs(7065)) or (layer2_outputs(991)));
    outputs(8864) <= not(layer2_outputs(5350));
    outputs(8865) <= layer2_outputs(7839);
    outputs(8866) <= not(layer2_outputs(5045));
    outputs(8867) <= layer2_outputs(8809);
    outputs(8868) <= (layer2_outputs(3800)) and (layer2_outputs(71));
    outputs(8869) <= not((layer2_outputs(311)) xor (layer2_outputs(666)));
    outputs(8870) <= not(layer2_outputs(671));
    outputs(8871) <= layer2_outputs(9723);
    outputs(8872) <= not(layer2_outputs(1941));
    outputs(8873) <= not(layer2_outputs(1830)) or (layer2_outputs(6067));
    outputs(8874) <= layer2_outputs(806);
    outputs(8875) <= '1';
    outputs(8876) <= not(layer2_outputs(7560));
    outputs(8877) <= not(layer2_outputs(1775));
    outputs(8878) <= layer2_outputs(9878);
    outputs(8879) <= layer2_outputs(2891);
    outputs(8880) <= not((layer2_outputs(9446)) xor (layer2_outputs(5667)));
    outputs(8881) <= (layer2_outputs(2292)) xor (layer2_outputs(4988));
    outputs(8882) <= layer2_outputs(5667);
    outputs(8883) <= layer2_outputs(7794);
    outputs(8884) <= not(layer2_outputs(3218));
    outputs(8885) <= layer2_outputs(9236);
    outputs(8886) <= layer2_outputs(7201);
    outputs(8887) <= layer2_outputs(1972);
    outputs(8888) <= not(layer2_outputs(10024));
    outputs(8889) <= layer2_outputs(7607);
    outputs(8890) <= not(layer2_outputs(6293));
    outputs(8891) <= not((layer2_outputs(7346)) xor (layer2_outputs(1402)));
    outputs(8892) <= (layer2_outputs(2522)) xor (layer2_outputs(10032));
    outputs(8893) <= not((layer2_outputs(7585)) and (layer2_outputs(4538)));
    outputs(8894) <= not(layer2_outputs(9794));
    outputs(8895) <= layer2_outputs(4492);
    outputs(8896) <= not(layer2_outputs(7184));
    outputs(8897) <= layer2_outputs(1952);
    outputs(8898) <= layer2_outputs(3007);
    outputs(8899) <= not((layer2_outputs(4437)) and (layer2_outputs(1706)));
    outputs(8900) <= not(layer2_outputs(9116)) or (layer2_outputs(8140));
    outputs(8901) <= layer2_outputs(4939);
    outputs(8902) <= not(layer2_outputs(510));
    outputs(8903) <= not(layer2_outputs(3425));
    outputs(8904) <= layer2_outputs(8574);
    outputs(8905) <= (layer2_outputs(5313)) and (layer2_outputs(1352));
    outputs(8906) <= not((layer2_outputs(3252)) and (layer2_outputs(3426)));
    outputs(8907) <= layer2_outputs(3739);
    outputs(8908) <= not((layer2_outputs(3818)) xor (layer2_outputs(10008)));
    outputs(8909) <= (layer2_outputs(1376)) and (layer2_outputs(4403));
    outputs(8910) <= layer2_outputs(5545);
    outputs(8911) <= not((layer2_outputs(8662)) and (layer2_outputs(5268)));
    outputs(8912) <= layer2_outputs(2942);
    outputs(8913) <= (layer2_outputs(9565)) or (layer2_outputs(4441));
    outputs(8914) <= (layer2_outputs(4615)) and not (layer2_outputs(884));
    outputs(8915) <= not(layer2_outputs(8828));
    outputs(8916) <= not((layer2_outputs(996)) and (layer2_outputs(1063)));
    outputs(8917) <= not(layer2_outputs(10174));
    outputs(8918) <= not((layer2_outputs(7247)) and (layer2_outputs(4067)));
    outputs(8919) <= (layer2_outputs(5821)) and not (layer2_outputs(2013));
    outputs(8920) <= layer2_outputs(4617);
    outputs(8921) <= not(layer2_outputs(5514));
    outputs(8922) <= layer2_outputs(3948);
    outputs(8923) <= not(layer2_outputs(6954)) or (layer2_outputs(1652));
    outputs(8924) <= not(layer2_outputs(1209)) or (layer2_outputs(810));
    outputs(8925) <= not((layer2_outputs(5858)) xor (layer2_outputs(8567)));
    outputs(8926) <= layer2_outputs(9867);
    outputs(8927) <= layer2_outputs(9022);
    outputs(8928) <= not(layer2_outputs(6847)) or (layer2_outputs(5105));
    outputs(8929) <= (layer2_outputs(9962)) xor (layer2_outputs(4031));
    outputs(8930) <= layer2_outputs(6921);
    outputs(8931) <= layer2_outputs(6212);
    outputs(8932) <= layer2_outputs(5707);
    outputs(8933) <= layer2_outputs(3996);
    outputs(8934) <= (layer2_outputs(2489)) xor (layer2_outputs(1776));
    outputs(8935) <= not(layer2_outputs(6562));
    outputs(8936) <= not(layer2_outputs(21));
    outputs(8937) <= layer2_outputs(5693);
    outputs(8938) <= not((layer2_outputs(489)) xor (layer2_outputs(9057)));
    outputs(8939) <= not((layer2_outputs(1393)) xor (layer2_outputs(231)));
    outputs(8940) <= not(layer2_outputs(44));
    outputs(8941) <= layer2_outputs(3054);
    outputs(8942) <= layer2_outputs(369);
    outputs(8943) <= not((layer2_outputs(7643)) or (layer2_outputs(9426)));
    outputs(8944) <= not(layer2_outputs(2532));
    outputs(8945) <= not(layer2_outputs(6147));
    outputs(8946) <= not(layer2_outputs(10202));
    outputs(8947) <= not(layer2_outputs(1848));
    outputs(8948) <= not(layer2_outputs(8846)) or (layer2_outputs(6297));
    outputs(8949) <= not(layer2_outputs(2669)) or (layer2_outputs(10188));
    outputs(8950) <= layer2_outputs(9808);
    outputs(8951) <= not(layer2_outputs(1699));
    outputs(8952) <= (layer2_outputs(649)) xor (layer2_outputs(9748));
    outputs(8953) <= not(layer2_outputs(9551)) or (layer2_outputs(6798));
    outputs(8954) <= (layer2_outputs(10188)) xor (layer2_outputs(1991));
    outputs(8955) <= (layer2_outputs(8549)) xor (layer2_outputs(1468));
    outputs(8956) <= layer2_outputs(2301);
    outputs(8957) <= not(layer2_outputs(7680));
    outputs(8958) <= not(layer2_outputs(4130)) or (layer2_outputs(9053));
    outputs(8959) <= layer2_outputs(374);
    outputs(8960) <= not((layer2_outputs(2506)) xor (layer2_outputs(2503)));
    outputs(8961) <= (layer2_outputs(518)) xor (layer2_outputs(9980));
    outputs(8962) <= layer2_outputs(3305);
    outputs(8963) <= (layer2_outputs(3605)) or (layer2_outputs(9530));
    outputs(8964) <= layer2_outputs(7666);
    outputs(8965) <= not((layer2_outputs(8615)) xor (layer2_outputs(2176)));
    outputs(8966) <= (layer2_outputs(4719)) or (layer2_outputs(7641));
    outputs(8967) <= layer2_outputs(2108);
    outputs(8968) <= not(layer2_outputs(3217));
    outputs(8969) <= layer2_outputs(5402);
    outputs(8970) <= (layer2_outputs(10023)) and (layer2_outputs(5095));
    outputs(8971) <= (layer2_outputs(5732)) xor (layer2_outputs(5418));
    outputs(8972) <= (layer2_outputs(7380)) xor (layer2_outputs(1134));
    outputs(8973) <= not(layer2_outputs(2361));
    outputs(8974) <= layer2_outputs(2861);
    outputs(8975) <= layer2_outputs(4937);
    outputs(8976) <= layer2_outputs(7248);
    outputs(8977) <= (layer2_outputs(874)) xor (layer2_outputs(6702));
    outputs(8978) <= not((layer2_outputs(3247)) xor (layer2_outputs(5356)));
    outputs(8979) <= not(layer2_outputs(7977));
    outputs(8980) <= (layer2_outputs(1655)) xor (layer2_outputs(6059));
    outputs(8981) <= not(layer2_outputs(3515));
    outputs(8982) <= layer2_outputs(2705);
    outputs(8983) <= not((layer2_outputs(2692)) xor (layer2_outputs(2867)));
    outputs(8984) <= layer2_outputs(587);
    outputs(8985) <= (layer2_outputs(6644)) xor (layer2_outputs(5743));
    outputs(8986) <= (layer2_outputs(3333)) xor (layer2_outputs(1081));
    outputs(8987) <= not(layer2_outputs(9052));
    outputs(8988) <= not(layer2_outputs(7957));
    outputs(8989) <= layer2_outputs(6961);
    outputs(8990) <= not((layer2_outputs(2337)) and (layer2_outputs(3607)));
    outputs(8991) <= not((layer2_outputs(5581)) xor (layer2_outputs(7549)));
    outputs(8992) <= layer2_outputs(10236);
    outputs(8993) <= layer2_outputs(9462);
    outputs(8994) <= not((layer2_outputs(5195)) xor (layer2_outputs(6812)));
    outputs(8995) <= layer2_outputs(7933);
    outputs(8996) <= not(layer2_outputs(7626));
    outputs(8997) <= not(layer2_outputs(43)) or (layer2_outputs(2005));
    outputs(8998) <= not(layer2_outputs(3334)) or (layer2_outputs(8563));
    outputs(8999) <= layer2_outputs(1653);
    outputs(9000) <= layer2_outputs(10077);
    outputs(9001) <= (layer2_outputs(9679)) or (layer2_outputs(1210));
    outputs(9002) <= not(layer2_outputs(7631)) or (layer2_outputs(2202));
    outputs(9003) <= not(layer2_outputs(1609));
    outputs(9004) <= layer2_outputs(4568);
    outputs(9005) <= not(layer2_outputs(2179)) or (layer2_outputs(8708));
    outputs(9006) <= layer2_outputs(1631);
    outputs(9007) <= not(layer2_outputs(1944));
    outputs(9008) <= not((layer2_outputs(8119)) and (layer2_outputs(3077)));
    outputs(9009) <= layer2_outputs(7340);
    outputs(9010) <= layer2_outputs(9003);
    outputs(9011) <= layer2_outputs(1064);
    outputs(9012) <= not((layer2_outputs(4185)) xor (layer2_outputs(9966)));
    outputs(9013) <= layer2_outputs(8079);
    outputs(9014) <= not((layer2_outputs(6921)) xor (layer2_outputs(6406)));
    outputs(9015) <= not((layer2_outputs(6947)) and (layer2_outputs(10028)));
    outputs(9016) <= (layer2_outputs(7487)) and not (layer2_outputs(4092));
    outputs(9017) <= (layer2_outputs(5238)) xor (layer2_outputs(6937));
    outputs(9018) <= layer2_outputs(1072);
    outputs(9019) <= not(layer2_outputs(8408)) or (layer2_outputs(5764));
    outputs(9020) <= layer2_outputs(10227);
    outputs(9021) <= not(layer2_outputs(643));
    outputs(9022) <= (layer2_outputs(9264)) xor (layer2_outputs(7695));
    outputs(9023) <= not((layer2_outputs(7940)) xor (layer2_outputs(9264)));
    outputs(9024) <= layer2_outputs(9460);
    outputs(9025) <= not(layer2_outputs(6154)) or (layer2_outputs(5315));
    outputs(9026) <= not((layer2_outputs(1793)) or (layer2_outputs(6873)));
    outputs(9027) <= not(layer2_outputs(3722));
    outputs(9028) <= not(layer2_outputs(6557));
    outputs(9029) <= layer2_outputs(2299);
    outputs(9030) <= not(layer2_outputs(8994)) or (layer2_outputs(2578));
    outputs(9031) <= not((layer2_outputs(5994)) or (layer2_outputs(9887)));
    outputs(9032) <= layer2_outputs(1175);
    outputs(9033) <= not((layer2_outputs(6011)) and (layer2_outputs(3459)));
    outputs(9034) <= (layer2_outputs(3881)) xor (layer2_outputs(5069));
    outputs(9035) <= (layer2_outputs(5263)) or (layer2_outputs(1480));
    outputs(9036) <= not(layer2_outputs(8525)) or (layer2_outputs(8825));
    outputs(9037) <= layer2_outputs(2567);
    outputs(9038) <= layer2_outputs(8859);
    outputs(9039) <= not((layer2_outputs(1442)) or (layer2_outputs(9591)));
    outputs(9040) <= not(layer2_outputs(6241));
    outputs(9041) <= not(layer2_outputs(5168));
    outputs(9042) <= layer2_outputs(3690);
    outputs(9043) <= not(layer2_outputs(1951));
    outputs(9044) <= (layer2_outputs(7062)) xor (layer2_outputs(3578));
    outputs(9045) <= layer2_outputs(2854);
    outputs(9046) <= not(layer2_outputs(6259));
    outputs(9047) <= not(layer2_outputs(882));
    outputs(9048) <= (layer2_outputs(5021)) xor (layer2_outputs(6736));
    outputs(9049) <= (layer2_outputs(5299)) xor (layer2_outputs(5986));
    outputs(9050) <= (layer2_outputs(6556)) xor (layer2_outputs(2029));
    outputs(9051) <= layer2_outputs(9905);
    outputs(9052) <= (layer2_outputs(3430)) xor (layer2_outputs(8189));
    outputs(9053) <= not((layer2_outputs(5073)) xor (layer2_outputs(3781)));
    outputs(9054) <= not(layer2_outputs(5342)) or (layer2_outputs(249));
    outputs(9055) <= '0';
    outputs(9056) <= (layer2_outputs(3360)) xor (layer2_outputs(101));
    outputs(9057) <= not((layer2_outputs(5804)) xor (layer2_outputs(10200)));
    outputs(9058) <= (layer2_outputs(676)) and (layer2_outputs(6792));
    outputs(9059) <= not(layer2_outputs(260));
    outputs(9060) <= not(layer2_outputs(751));
    outputs(9061) <= layer2_outputs(9261);
    outputs(9062) <= not(layer2_outputs(8917));
    outputs(9063) <= layer2_outputs(8799);
    outputs(9064) <= not(layer2_outputs(5620));
    outputs(9065) <= layer2_outputs(7798);
    outputs(9066) <= not(layer2_outputs(995));
    outputs(9067) <= layer2_outputs(480);
    outputs(9068) <= not(layer2_outputs(6862));
    outputs(9069) <= not((layer2_outputs(6211)) xor (layer2_outputs(2808)));
    outputs(9070) <= not(layer2_outputs(7112)) or (layer2_outputs(4347));
    outputs(9071) <= not(layer2_outputs(6279));
    outputs(9072) <= not(layer2_outputs(7643));
    outputs(9073) <= not(layer2_outputs(4194)) or (layer2_outputs(7513));
    outputs(9074) <= not(layer2_outputs(1490));
    outputs(9075) <= layer2_outputs(2023);
    outputs(9076) <= not(layer2_outputs(7556));
    outputs(9077) <= layer2_outputs(7015);
    outputs(9078) <= layer2_outputs(2909);
    outputs(9079) <= (layer2_outputs(6803)) or (layer2_outputs(4178));
    outputs(9080) <= not(layer2_outputs(6444));
    outputs(9081) <= not((layer2_outputs(7956)) and (layer2_outputs(347)));
    outputs(9082) <= layer2_outputs(9334);
    outputs(9083) <= not(layer2_outputs(2486));
    outputs(9084) <= not(layer2_outputs(5714)) or (layer2_outputs(4273));
    outputs(9085) <= (layer2_outputs(5275)) and not (layer2_outputs(3425));
    outputs(9086) <= not((layer2_outputs(6893)) xor (layer2_outputs(895)));
    outputs(9087) <= not(layer2_outputs(1749));
    outputs(9088) <= not((layer2_outputs(5801)) xor (layer2_outputs(9799)));
    outputs(9089) <= not(layer2_outputs(9225)) or (layer2_outputs(163));
    outputs(9090) <= not(layer2_outputs(5092));
    outputs(9091) <= not((layer2_outputs(4593)) xor (layer2_outputs(1644)));
    outputs(9092) <= (layer2_outputs(5274)) xor (layer2_outputs(4615));
    outputs(9093) <= layer2_outputs(3224);
    outputs(9094) <= not(layer2_outputs(5251));
    outputs(9095) <= layer2_outputs(5658);
    outputs(9096) <= not(layer2_outputs(6888));
    outputs(9097) <= (layer2_outputs(989)) xor (layer2_outputs(2047));
    outputs(9098) <= (layer2_outputs(4216)) xor (layer2_outputs(9923));
    outputs(9099) <= not((layer2_outputs(911)) and (layer2_outputs(6292)));
    outputs(9100) <= layer2_outputs(5319);
    outputs(9101) <= (layer2_outputs(6551)) xor (layer2_outputs(8457));
    outputs(9102) <= not(layer2_outputs(7031));
    outputs(9103) <= not((layer2_outputs(5264)) xor (layer2_outputs(8393)));
    outputs(9104) <= not(layer2_outputs(3914)) or (layer2_outputs(5330));
    outputs(9105) <= layer2_outputs(6476);
    outputs(9106) <= not((layer2_outputs(9501)) xor (layer2_outputs(2429)));
    outputs(9107) <= not(layer2_outputs(8363));
    outputs(9108) <= layer2_outputs(4357);
    outputs(9109) <= not((layer2_outputs(5371)) xor (layer2_outputs(708)));
    outputs(9110) <= layer2_outputs(7226);
    outputs(9111) <= (layer2_outputs(8950)) xor (layer2_outputs(3903));
    outputs(9112) <= (layer2_outputs(4376)) xor (layer2_outputs(8106));
    outputs(9113) <= layer2_outputs(5364);
    outputs(9114) <= (layer2_outputs(9329)) xor (layer2_outputs(9032));
    outputs(9115) <= not(layer2_outputs(6866));
    outputs(9116) <= layer2_outputs(6185);
    outputs(9117) <= (layer2_outputs(5020)) xor (layer2_outputs(5515));
    outputs(9118) <= not(layer2_outputs(4858));
    outputs(9119) <= not(layer2_outputs(4236));
    outputs(9120) <= not(layer2_outputs(6971)) or (layer2_outputs(10196));
    outputs(9121) <= not((layer2_outputs(9389)) xor (layer2_outputs(4811)));
    outputs(9122) <= layer2_outputs(8778);
    outputs(9123) <= not(layer2_outputs(6313));
    outputs(9124) <= (layer2_outputs(9591)) xor (layer2_outputs(6587));
    outputs(9125) <= layer2_outputs(7399);
    outputs(9126) <= (layer2_outputs(2065)) and not (layer2_outputs(3733));
    outputs(9127) <= not((layer2_outputs(8634)) xor (layer2_outputs(2443)));
    outputs(9128) <= layer2_outputs(3466);
    outputs(9129) <= layer2_outputs(307);
    outputs(9130) <= not((layer2_outputs(6093)) xor (layer2_outputs(9365)));
    outputs(9131) <= layer2_outputs(1403);
    outputs(9132) <= not((layer2_outputs(1374)) xor (layer2_outputs(9995)));
    outputs(9133) <= (layer2_outputs(376)) xor (layer2_outputs(1911));
    outputs(9134) <= not(layer2_outputs(5463));
    outputs(9135) <= not(layer2_outputs(9630));
    outputs(9136) <= not((layer2_outputs(2625)) xor (layer2_outputs(1428)));
    outputs(9137) <= not(layer2_outputs(3620));
    outputs(9138) <= (layer2_outputs(4677)) or (layer2_outputs(5851));
    outputs(9139) <= not((layer2_outputs(8838)) xor (layer2_outputs(9112)));
    outputs(9140) <= not(layer2_outputs(4397));
    outputs(9141) <= not((layer2_outputs(1783)) xor (layer2_outputs(2550)));
    outputs(9142) <= layer2_outputs(2980);
    outputs(9143) <= layer2_outputs(548);
    outputs(9144) <= (layer2_outputs(8483)) or (layer2_outputs(7228));
    outputs(9145) <= not(layer2_outputs(7645));
    outputs(9146) <= layer2_outputs(6896);
    outputs(9147) <= (layer2_outputs(9701)) and (layer2_outputs(2896));
    outputs(9148) <= not(layer2_outputs(5829));
    outputs(9149) <= not(layer2_outputs(5125));
    outputs(9150) <= not(layer2_outputs(2982));
    outputs(9151) <= layer2_outputs(8328);
    outputs(9152) <= layer2_outputs(7650);
    outputs(9153) <= (layer2_outputs(7514)) xor (layer2_outputs(8757));
    outputs(9154) <= layer2_outputs(3396);
    outputs(9155) <= not(layer2_outputs(327));
    outputs(9156) <= layer2_outputs(4568);
    outputs(9157) <= not((layer2_outputs(626)) xor (layer2_outputs(206)));
    outputs(9158) <= not(layer2_outputs(9484));
    outputs(9159) <= not(layer2_outputs(10211)) or (layer2_outputs(10197));
    outputs(9160) <= layer2_outputs(9307);
    outputs(9161) <= not(layer2_outputs(8014)) or (layer2_outputs(6881));
    outputs(9162) <= layer2_outputs(5284);
    outputs(9163) <= (layer2_outputs(2078)) or (layer2_outputs(3376));
    outputs(9164) <= not(layer2_outputs(8899)) or (layer2_outputs(2197));
    outputs(9165) <= layer2_outputs(4246);
    outputs(9166) <= not(layer2_outputs(89)) or (layer2_outputs(374));
    outputs(9167) <= not(layer2_outputs(929));
    outputs(9168) <= layer2_outputs(1794);
    outputs(9169) <= (layer2_outputs(2493)) xor (layer2_outputs(1084));
    outputs(9170) <= (layer2_outputs(3337)) and not (layer2_outputs(8646));
    outputs(9171) <= (layer2_outputs(8756)) and not (layer2_outputs(8442));
    outputs(9172) <= layer2_outputs(6042);
    outputs(9173) <= (layer2_outputs(4099)) or (layer2_outputs(4884));
    outputs(9174) <= (layer2_outputs(9015)) xor (layer2_outputs(2620));
    outputs(9175) <= not(layer2_outputs(7787));
    outputs(9176) <= not(layer2_outputs(3773));
    outputs(9177) <= not(layer2_outputs(7217));
    outputs(9178) <= not(layer2_outputs(10000)) or (layer2_outputs(1516));
    outputs(9179) <= layer2_outputs(5669);
    outputs(9180) <= (layer2_outputs(7605)) or (layer2_outputs(9553));
    outputs(9181) <= not((layer2_outputs(8949)) and (layer2_outputs(8970)));
    outputs(9182) <= not(layer2_outputs(6496));
    outputs(9183) <= not((layer2_outputs(5401)) xor (layer2_outputs(9954)));
    outputs(9184) <= not(layer2_outputs(3669));
    outputs(9185) <= layer2_outputs(2394);
    outputs(9186) <= (layer2_outputs(990)) xor (layer2_outputs(5809));
    outputs(9187) <= not((layer2_outputs(2057)) xor (layer2_outputs(2245)));
    outputs(9188) <= layer2_outputs(3845);
    outputs(9189) <= (layer2_outputs(7604)) xor (layer2_outputs(5374));
    outputs(9190) <= not(layer2_outputs(7745));
    outputs(9191) <= not((layer2_outputs(4364)) xor (layer2_outputs(1500)));
    outputs(9192) <= layer2_outputs(7445);
    outputs(9193) <= not(layer2_outputs(1880));
    outputs(9194) <= (layer2_outputs(2964)) or (layer2_outputs(6631));
    outputs(9195) <= not(layer2_outputs(6635)) or (layer2_outputs(656));
    outputs(9196) <= (layer2_outputs(8291)) and not (layer2_outputs(10140));
    outputs(9197) <= layer2_outputs(6684);
    outputs(9198) <= layer2_outputs(2459);
    outputs(9199) <= layer2_outputs(2374);
    outputs(9200) <= not(layer2_outputs(6755));
    outputs(9201) <= (layer2_outputs(2042)) xor (layer2_outputs(7589));
    outputs(9202) <= layer2_outputs(427);
    outputs(9203) <= (layer2_outputs(2847)) xor (layer2_outputs(1604));
    outputs(9204) <= layer2_outputs(5435);
    outputs(9205) <= layer2_outputs(6590);
    outputs(9206) <= (layer2_outputs(2785)) xor (layer2_outputs(8222));
    outputs(9207) <= (layer2_outputs(5099)) or (layer2_outputs(8861));
    outputs(9208) <= (layer2_outputs(5034)) xor (layer2_outputs(8620));
    outputs(9209) <= layer2_outputs(948);
    outputs(9210) <= (layer2_outputs(10115)) xor (layer2_outputs(7741));
    outputs(9211) <= not(layer2_outputs(8353)) or (layer2_outputs(9589));
    outputs(9212) <= layer2_outputs(8324);
    outputs(9213) <= layer2_outputs(517);
    outputs(9214) <= layer2_outputs(10167);
    outputs(9215) <= (layer2_outputs(936)) xor (layer2_outputs(6394));
    outputs(9216) <= not(layer2_outputs(1484));
    outputs(9217) <= not((layer2_outputs(8471)) xor (layer2_outputs(6193)));
    outputs(9218) <= layer2_outputs(183);
    outputs(9219) <= not(layer2_outputs(1557));
    outputs(9220) <= layer2_outputs(1470);
    outputs(9221) <= layer2_outputs(7656);
    outputs(9222) <= not(layer2_outputs(616));
    outputs(9223) <= not(layer2_outputs(3925));
    outputs(9224) <= (layer2_outputs(5747)) xor (layer2_outputs(4923));
    outputs(9225) <= not((layer2_outputs(4502)) and (layer2_outputs(4855)));
    outputs(9226) <= not(layer2_outputs(3849));
    outputs(9227) <= not(layer2_outputs(4098));
    outputs(9228) <= layer2_outputs(1933);
    outputs(9229) <= not(layer2_outputs(4224));
    outputs(9230) <= not(layer2_outputs(3559));
    outputs(9231) <= not(layer2_outputs(8102));
    outputs(9232) <= not((layer2_outputs(5151)) xor (layer2_outputs(6358)));
    outputs(9233) <= not(layer2_outputs(2136));
    outputs(9234) <= not(layer2_outputs(4380));
    outputs(9235) <= (layer2_outputs(9908)) or (layer2_outputs(2618));
    outputs(9236) <= not(layer2_outputs(8089));
    outputs(9237) <= layer2_outputs(1087);
    outputs(9238) <= not((layer2_outputs(1318)) xor (layer2_outputs(8606)));
    outputs(9239) <= not(layer2_outputs(852));
    outputs(9240) <= (layer2_outputs(2353)) xor (layer2_outputs(1826));
    outputs(9241) <= not(layer2_outputs(3292));
    outputs(9242) <= layer2_outputs(5657);
    outputs(9243) <= not(layer2_outputs(6011));
    outputs(9244) <= not(layer2_outputs(3601));
    outputs(9245) <= not(layer2_outputs(140));
    outputs(9246) <= not(layer2_outputs(8351));
    outputs(9247) <= layer2_outputs(4345);
    outputs(9248) <= not((layer2_outputs(2006)) or (layer2_outputs(7235)));
    outputs(9249) <= not(layer2_outputs(9241));
    outputs(9250) <= not(layer2_outputs(6932));
    outputs(9251) <= layer2_outputs(8705);
    outputs(9252) <= layer2_outputs(8290);
    outputs(9253) <= (layer2_outputs(547)) or (layer2_outputs(771));
    outputs(9254) <= not((layer2_outputs(3948)) xor (layer2_outputs(9016)));
    outputs(9255) <= layer2_outputs(153);
    outputs(9256) <= layer2_outputs(2603);
    outputs(9257) <= not(layer2_outputs(5839));
    outputs(9258) <= layer2_outputs(5094);
    outputs(9259) <= not(layer2_outputs(6660));
    outputs(9260) <= not(layer2_outputs(5520));
    outputs(9261) <= layer2_outputs(4597);
    outputs(9262) <= not(layer2_outputs(8508));
    outputs(9263) <= not(layer2_outputs(1449));
    outputs(9264) <= layer2_outputs(3462);
    outputs(9265) <= not(layer2_outputs(1236)) or (layer2_outputs(8206));
    outputs(9266) <= not(layer2_outputs(2994));
    outputs(9267) <= not(layer2_outputs(8618));
    outputs(9268) <= not(layer2_outputs(4975));
    outputs(9269) <= layer2_outputs(7258);
    outputs(9270) <= not((layer2_outputs(241)) xor (layer2_outputs(9275)));
    outputs(9271) <= not((layer2_outputs(2276)) xor (layer2_outputs(3480)));
    outputs(9272) <= not(layer2_outputs(3957));
    outputs(9273) <= (layer2_outputs(8006)) xor (layer2_outputs(5175));
    outputs(9274) <= layer2_outputs(4772);
    outputs(9275) <= layer2_outputs(5377);
    outputs(9276) <= not(layer2_outputs(5205));
    outputs(9277) <= (layer2_outputs(9525)) and not (layer2_outputs(9610));
    outputs(9278) <= not((layer2_outputs(5634)) xor (layer2_outputs(1997)));
    outputs(9279) <= not(layer2_outputs(8127));
    outputs(9280) <= not((layer2_outputs(3008)) xor (layer2_outputs(9992)));
    outputs(9281) <= not((layer2_outputs(2124)) xor (layer2_outputs(6325)));
    outputs(9282) <= not(layer2_outputs(699));
    outputs(9283) <= not(layer2_outputs(646));
    outputs(9284) <= layer2_outputs(9397);
    outputs(9285) <= (layer2_outputs(9884)) xor (layer2_outputs(7215));
    outputs(9286) <= (layer2_outputs(925)) xor (layer2_outputs(2204));
    outputs(9287) <= (layer2_outputs(5882)) xor (layer2_outputs(3020));
    outputs(9288) <= not(layer2_outputs(2958));
    outputs(9289) <= not(layer2_outputs(4680));
    outputs(9290) <= layer2_outputs(1620);
    outputs(9291) <= not(layer2_outputs(8703));
    outputs(9292) <= not((layer2_outputs(8256)) and (layer2_outputs(7734)));
    outputs(9293) <= not(layer2_outputs(7468)) or (layer2_outputs(5718));
    outputs(9294) <= not((layer2_outputs(5860)) xor (layer2_outputs(9076)));
    outputs(9295) <= not(layer2_outputs(2590));
    outputs(9296) <= (layer2_outputs(540)) xor (layer2_outputs(671));
    outputs(9297) <= layer2_outputs(6816);
    outputs(9298) <= not((layer2_outputs(3407)) or (layer2_outputs(9389)));
    outputs(9299) <= not((layer2_outputs(3013)) xor (layer2_outputs(5672)));
    outputs(9300) <= layer2_outputs(827);
    outputs(9301) <= (layer2_outputs(3677)) and (layer2_outputs(2026));
    outputs(9302) <= layer2_outputs(659);
    outputs(9303) <= (layer2_outputs(6439)) or (layer2_outputs(7262));
    outputs(9304) <= not(layer2_outputs(2024));
    outputs(9305) <= (layer2_outputs(6414)) xor (layer2_outputs(4898));
    outputs(9306) <= not(layer2_outputs(1170));
    outputs(9307) <= (layer2_outputs(2525)) xor (layer2_outputs(4462));
    outputs(9308) <= not(layer2_outputs(7495));
    outputs(9309) <= not((layer2_outputs(6108)) xor (layer2_outputs(9176)));
    outputs(9310) <= layer2_outputs(6537);
    outputs(9311) <= not(layer2_outputs(6455));
    outputs(9312) <= not(layer2_outputs(5132)) or (layer2_outputs(3542));
    outputs(9313) <= layer2_outputs(5896);
    outputs(9314) <= layer2_outputs(9043);
    outputs(9315) <= (layer2_outputs(514)) and not (layer2_outputs(7003));
    outputs(9316) <= not(layer2_outputs(693));
    outputs(9317) <= layer2_outputs(8398);
    outputs(9318) <= (layer2_outputs(5770)) xor (layer2_outputs(7501));
    outputs(9319) <= not(layer2_outputs(1246));
    outputs(9320) <= layer2_outputs(4465);
    outputs(9321) <= layer2_outputs(6860);
    outputs(9322) <= not(layer2_outputs(1612)) or (layer2_outputs(8962));
    outputs(9323) <= not((layer2_outputs(600)) or (layer2_outputs(7328)));
    outputs(9324) <= layer2_outputs(7095);
    outputs(9325) <= not(layer2_outputs(643));
    outputs(9326) <= (layer2_outputs(1546)) xor (layer2_outputs(9252));
    outputs(9327) <= (layer2_outputs(5033)) xor (layer2_outputs(9226));
    outputs(9328) <= not(layer2_outputs(3038));
    outputs(9329) <= not(layer2_outputs(3404));
    outputs(9330) <= layer2_outputs(1545);
    outputs(9331) <= (layer2_outputs(1164)) xor (layer2_outputs(9395));
    outputs(9332) <= not(layer2_outputs(449));
    outputs(9333) <= layer2_outputs(4481);
    outputs(9334) <= layer2_outputs(1958);
    outputs(9335) <= layer2_outputs(6152);
    outputs(9336) <= layer2_outputs(5369);
    outputs(9337) <= not((layer2_outputs(4476)) xor (layer2_outputs(1411)));
    outputs(9338) <= not(layer2_outputs(6493)) or (layer2_outputs(6483));
    outputs(9339) <= layer2_outputs(5093);
    outputs(9340) <= (layer2_outputs(5150)) xor (layer2_outputs(5749));
    outputs(9341) <= layer2_outputs(10011);
    outputs(9342) <= not((layer2_outputs(4660)) xor (layer2_outputs(5981)));
    outputs(9343) <= layer2_outputs(3183);
    outputs(9344) <= layer2_outputs(1165);
    outputs(9345) <= not(layer2_outputs(354));
    outputs(9346) <= not(layer2_outputs(8640)) or (layer2_outputs(5663));
    outputs(9347) <= not((layer2_outputs(6956)) xor (layer2_outputs(4149)));
    outputs(9348) <= layer2_outputs(6549);
    outputs(9349) <= layer2_outputs(1224);
    outputs(9350) <= layer2_outputs(8022);
    outputs(9351) <= layer2_outputs(9094);
    outputs(9352) <= not(layer2_outputs(5822)) or (layer2_outputs(313));
    outputs(9353) <= (layer2_outputs(8667)) xor (layer2_outputs(7912));
    outputs(9354) <= not(layer2_outputs(1629));
    outputs(9355) <= not(layer2_outputs(2022));
    outputs(9356) <= layer2_outputs(5428);
    outputs(9357) <= not(layer2_outputs(3899));
    outputs(9358) <= not(layer2_outputs(5257));
    outputs(9359) <= layer2_outputs(5967);
    outputs(9360) <= layer2_outputs(7811);
    outputs(9361) <= not(layer2_outputs(9124));
    outputs(9362) <= not(layer2_outputs(8391));
    outputs(9363) <= layer2_outputs(4666);
    outputs(9364) <= layer2_outputs(5367);
    outputs(9365) <= layer2_outputs(7286);
    outputs(9366) <= not(layer2_outputs(3913));
    outputs(9367) <= (layer2_outputs(866)) xor (layer2_outputs(1069));
    outputs(9368) <= not(layer2_outputs(9013));
    outputs(9369) <= layer2_outputs(5232);
    outputs(9370) <= layer2_outputs(3885);
    outputs(9371) <= (layer2_outputs(3782)) and not (layer2_outputs(4285));
    outputs(9372) <= not((layer2_outputs(6294)) or (layer2_outputs(1370)));
    outputs(9373) <= not((layer2_outputs(8126)) xor (layer2_outputs(8186)));
    outputs(9374) <= not(layer2_outputs(831));
    outputs(9375) <= not(layer2_outputs(1242));
    outputs(9376) <= not(layer2_outputs(7078));
    outputs(9377) <= not((layer2_outputs(4901)) and (layer2_outputs(1054)));
    outputs(9378) <= not((layer2_outputs(1707)) xor (layer2_outputs(10058)));
    outputs(9379) <= not((layer2_outputs(141)) xor (layer2_outputs(1860)));
    outputs(9380) <= not(layer2_outputs(719));
    outputs(9381) <= layer2_outputs(8446);
    outputs(9382) <= layer2_outputs(5271);
    outputs(9383) <= layer2_outputs(3584);
    outputs(9384) <= not((layer2_outputs(13)) xor (layer2_outputs(1201)));
    outputs(9385) <= layer2_outputs(4082);
    outputs(9386) <= not(layer2_outputs(1998));
    outputs(9387) <= not((layer2_outputs(9117)) or (layer2_outputs(2551)));
    outputs(9388) <= not(layer2_outputs(9910));
    outputs(9389) <= not(layer2_outputs(7229));
    outputs(9390) <= (layer2_outputs(3350)) and not (layer2_outputs(3569));
    outputs(9391) <= not((layer2_outputs(6728)) or (layer2_outputs(2611)));
    outputs(9392) <= not((layer2_outputs(2620)) or (layer2_outputs(1712)));
    outputs(9393) <= layer2_outputs(5372);
    outputs(9394) <= not((layer2_outputs(5879)) xor (layer2_outputs(9825)));
    outputs(9395) <= layer2_outputs(10171);
    outputs(9396) <= (layer2_outputs(4783)) and (layer2_outputs(9099));
    outputs(9397) <= not((layer2_outputs(3496)) and (layer2_outputs(6186)));
    outputs(9398) <= layer2_outputs(9107);
    outputs(9399) <= layer2_outputs(447);
    outputs(9400) <= layer2_outputs(1034);
    outputs(9401) <= not((layer2_outputs(3285)) xor (layer2_outputs(3477)));
    outputs(9402) <= not(layer2_outputs(6987)) or (layer2_outputs(4563));
    outputs(9403) <= not(layer2_outputs(9259));
    outputs(9404) <= (layer2_outputs(2127)) and not (layer2_outputs(7343));
    outputs(9405) <= not(layer2_outputs(1388));
    outputs(9406) <= layer2_outputs(1136);
    outputs(9407) <= not(layer2_outputs(3031));
    outputs(9408) <= layer2_outputs(4574);
    outputs(9409) <= not(layer2_outputs(2041));
    outputs(9410) <= layer2_outputs(9508);
    outputs(9411) <= not(layer2_outputs(9562));
    outputs(9412) <= not(layer2_outputs(66));
    outputs(9413) <= (layer2_outputs(8348)) xor (layer2_outputs(7758));
    outputs(9414) <= layer2_outputs(4333);
    outputs(9415) <= not(layer2_outputs(7543));
    outputs(9416) <= (layer2_outputs(6284)) and (layer2_outputs(3505));
    outputs(9417) <= not(layer2_outputs(8237));
    outputs(9418) <= layer2_outputs(4666);
    outputs(9419) <= not((layer2_outputs(3218)) xor (layer2_outputs(7159)));
    outputs(9420) <= not(layer2_outputs(9480)) or (layer2_outputs(5532));
    outputs(9421) <= layer2_outputs(8979);
    outputs(9422) <= not(layer2_outputs(8540));
    outputs(9423) <= (layer2_outputs(8126)) and not (layer2_outputs(6379));
    outputs(9424) <= not(layer2_outputs(9700));
    outputs(9425) <= (layer2_outputs(5408)) xor (layer2_outputs(4792));
    outputs(9426) <= layer2_outputs(5572);
    outputs(9427) <= not((layer2_outputs(9698)) xor (layer2_outputs(7859)));
    outputs(9428) <= not(layer2_outputs(1978));
    outputs(9429) <= not(layer2_outputs(1449));
    outputs(9430) <= (layer2_outputs(9909)) and (layer2_outputs(2307));
    outputs(9431) <= layer2_outputs(2808);
    outputs(9432) <= (layer2_outputs(4255)) xor (layer2_outputs(1756));
    outputs(9433) <= not(layer2_outputs(6450));
    outputs(9434) <= not(layer2_outputs(4205));
    outputs(9435) <= not(layer2_outputs(10031));
    outputs(9436) <= not(layer2_outputs(5465));
    outputs(9437) <= layer2_outputs(3660);
    outputs(9438) <= layer2_outputs(6560);
    outputs(9439) <= layer2_outputs(2835);
    outputs(9440) <= not((layer2_outputs(3172)) xor (layer2_outputs(5927)));
    outputs(9441) <= not(layer2_outputs(2144));
    outputs(9442) <= not(layer2_outputs(9582));
    outputs(9443) <= (layer2_outputs(8645)) and (layer2_outputs(633));
    outputs(9444) <= layer2_outputs(9788);
    outputs(9445) <= not(layer2_outputs(6508));
    outputs(9446) <= not(layer2_outputs(5850));
    outputs(9447) <= (layer2_outputs(1989)) xor (layer2_outputs(6072));
    outputs(9448) <= layer2_outputs(8182);
    outputs(9449) <= layer2_outputs(2263);
    outputs(9450) <= not((layer2_outputs(5712)) or (layer2_outputs(4190)));
    outputs(9451) <= not(layer2_outputs(4445));
    outputs(9452) <= not(layer2_outputs(8996));
    outputs(9453) <= layer2_outputs(5387);
    outputs(9454) <= layer2_outputs(3515);
    outputs(9455) <= layer2_outputs(8486);
    outputs(9456) <= (layer2_outputs(504)) xor (layer2_outputs(2813));
    outputs(9457) <= (layer2_outputs(3936)) or (layer2_outputs(2612));
    outputs(9458) <= not(layer2_outputs(8109));
    outputs(9459) <= not(layer2_outputs(3278));
    outputs(9460) <= not(layer2_outputs(6237));
    outputs(9461) <= layer2_outputs(1921);
    outputs(9462) <= not((layer2_outputs(540)) xor (layer2_outputs(7707)));
    outputs(9463) <= layer2_outputs(4512);
    outputs(9464) <= layer2_outputs(6016);
    outputs(9465) <= layer2_outputs(8327);
    outputs(9466) <= not(layer2_outputs(9604)) or (layer2_outputs(10105));
    outputs(9467) <= (layer2_outputs(7992)) or (layer2_outputs(2333));
    outputs(9468) <= (layer2_outputs(6855)) and not (layer2_outputs(2698));
    outputs(9469) <= not(layer2_outputs(1213));
    outputs(9470) <= (layer2_outputs(7688)) and not (layer2_outputs(7700));
    outputs(9471) <= not(layer2_outputs(2978));
    outputs(9472) <= (layer2_outputs(1481)) or (layer2_outputs(9091));
    outputs(9473) <= not(layer2_outputs(4672));
    outputs(9474) <= not(layer2_outputs(5014));
    outputs(9475) <= layer2_outputs(2863);
    outputs(9476) <= layer2_outputs(6471);
    outputs(9477) <= not(layer2_outputs(4746));
    outputs(9478) <= not(layer2_outputs(4094));
    outputs(9479) <= not(layer2_outputs(7661));
    outputs(9480) <= not((layer2_outputs(878)) xor (layer2_outputs(3289)));
    outputs(9481) <= (layer2_outputs(2801)) xor (layer2_outputs(2783));
    outputs(9482) <= (layer2_outputs(9477)) xor (layer2_outputs(8137));
    outputs(9483) <= not(layer2_outputs(2249));
    outputs(9484) <= not(layer2_outputs(6149));
    outputs(9485) <= not((layer2_outputs(4405)) xor (layer2_outputs(2834)));
    outputs(9486) <= layer2_outputs(4302);
    outputs(9487) <= not(layer2_outputs(3907)) or (layer2_outputs(605));
    outputs(9488) <= layer2_outputs(3791);
    outputs(9489) <= not(layer2_outputs(3535));
    outputs(9490) <= layer2_outputs(9041);
    outputs(9491) <= layer2_outputs(181);
    outputs(9492) <= not(layer2_outputs(797));
    outputs(9493) <= not(layer2_outputs(2510));
    outputs(9494) <= not((layer2_outputs(5477)) and (layer2_outputs(8105)));
    outputs(9495) <= (layer2_outputs(2486)) xor (layer2_outputs(10021));
    outputs(9496) <= not((layer2_outputs(5803)) or (layer2_outputs(2953)));
    outputs(9497) <= layer2_outputs(4448);
    outputs(9498) <= not(layer2_outputs(6847));
    outputs(9499) <= not(layer2_outputs(3734));
    outputs(9500) <= not((layer2_outputs(4048)) and (layer2_outputs(6838)));
    outputs(9501) <= not(layer2_outputs(8794));
    outputs(9502) <= layer2_outputs(1631);
    outputs(9503) <= (layer2_outputs(7130)) and (layer2_outputs(6222));
    outputs(9504) <= not(layer2_outputs(8161));
    outputs(9505) <= not(layer2_outputs(4888)) or (layer2_outputs(2152));
    outputs(9506) <= layer2_outputs(8481);
    outputs(9507) <= not(layer2_outputs(7665));
    outputs(9508) <= not((layer2_outputs(4059)) or (layer2_outputs(4668)));
    outputs(9509) <= layer2_outputs(3975);
    outputs(9510) <= not(layer2_outputs(5425));
    outputs(9511) <= layer2_outputs(3649);
    outputs(9512) <= (layer2_outputs(1191)) xor (layer2_outputs(4980));
    outputs(9513) <= not(layer2_outputs(6464));
    outputs(9514) <= layer2_outputs(4440);
    outputs(9515) <= not(layer2_outputs(10092));
    outputs(9516) <= not((layer2_outputs(2423)) xor (layer2_outputs(8705)));
    outputs(9517) <= layer2_outputs(7123);
    outputs(9518) <= (layer2_outputs(1575)) or (layer2_outputs(4465));
    outputs(9519) <= not(layer2_outputs(1507)) or (layer2_outputs(116));
    outputs(9520) <= layer2_outputs(7789);
    outputs(9521) <= (layer2_outputs(8049)) or (layer2_outputs(3411));
    outputs(9522) <= layer2_outputs(5680);
    outputs(9523) <= not(layer2_outputs(5820));
    outputs(9524) <= not(layer2_outputs(3681));
    outputs(9525) <= layer2_outputs(10239);
    outputs(9526) <= layer2_outputs(5857);
    outputs(9527) <= layer2_outputs(9059);
    outputs(9528) <= layer2_outputs(50);
    outputs(9529) <= (layer2_outputs(6858)) or (layer2_outputs(6569));
    outputs(9530) <= layer2_outputs(2929);
    outputs(9531) <= not((layer2_outputs(2709)) xor (layer2_outputs(6376)));
    outputs(9532) <= not(layer2_outputs(702));
    outputs(9533) <= layer2_outputs(7134);
    outputs(9534) <= layer2_outputs(5326);
    outputs(9535) <= not((layer2_outputs(8863)) or (layer2_outputs(1953)));
    outputs(9536) <= not((layer2_outputs(8271)) or (layer2_outputs(7734)));
    outputs(9537) <= (layer2_outputs(8779)) xor (layer2_outputs(1038));
    outputs(9538) <= (layer2_outputs(6657)) and (layer2_outputs(3900));
    outputs(9539) <= (layer2_outputs(3145)) and not (layer2_outputs(2295));
    outputs(9540) <= (layer2_outputs(7420)) xor (layer2_outputs(2504));
    outputs(9541) <= (layer2_outputs(6799)) and not (layer2_outputs(9216));
    outputs(9542) <= layer2_outputs(8515);
    outputs(9543) <= layer2_outputs(1686);
    outputs(9544) <= layer2_outputs(3905);
    outputs(9545) <= layer2_outputs(1605);
    outputs(9546) <= layer2_outputs(6287);
    outputs(9547) <= layer2_outputs(3748);
    outputs(9548) <= not(layer2_outputs(411));
    outputs(9549) <= layer2_outputs(3142);
    outputs(9550) <= (layer2_outputs(6417)) and (layer2_outputs(415));
    outputs(9551) <= not(layer2_outputs(2376));
    outputs(9552) <= layer2_outputs(3745);
    outputs(9553) <= not(layer2_outputs(9816));
    outputs(9554) <= (layer2_outputs(8381)) and not (layer2_outputs(675));
    outputs(9555) <= not(layer2_outputs(8299));
    outputs(9556) <= layer2_outputs(4835);
    outputs(9557) <= (layer2_outputs(5626)) xor (layer2_outputs(4446));
    outputs(9558) <= layer2_outputs(3715);
    outputs(9559) <= not(layer2_outputs(7951));
    outputs(9560) <= layer2_outputs(7290);
    outputs(9561) <= layer2_outputs(9447);
    outputs(9562) <= (layer2_outputs(553)) or (layer2_outputs(6727));
    outputs(9563) <= layer2_outputs(7766);
    outputs(9564) <= (layer2_outputs(7691)) and not (layer2_outputs(1186));
    outputs(9565) <= (layer2_outputs(7644)) xor (layer2_outputs(5865));
    outputs(9566) <= layer2_outputs(5089);
    outputs(9567) <= not(layer2_outputs(1790));
    outputs(9568) <= (layer2_outputs(2001)) xor (layer2_outputs(2420));
    outputs(9569) <= layer2_outputs(4139);
    outputs(9570) <= (layer2_outputs(6683)) xor (layer2_outputs(2007));
    outputs(9571) <= (layer2_outputs(7394)) xor (layer2_outputs(8524));
    outputs(9572) <= (layer2_outputs(6919)) xor (layer2_outputs(6017));
    outputs(9573) <= (layer2_outputs(1004)) and (layer2_outputs(6995));
    outputs(9574) <= not(layer2_outputs(10060)) or (layer2_outputs(6975));
    outputs(9575) <= layer2_outputs(10127);
    outputs(9576) <= layer2_outputs(7223);
    outputs(9577) <= (layer2_outputs(8931)) and (layer2_outputs(809));
    outputs(9578) <= not(layer2_outputs(4001));
    outputs(9579) <= not(layer2_outputs(1107));
    outputs(9580) <= not((layer2_outputs(6184)) xor (layer2_outputs(7632)));
    outputs(9581) <= (layer2_outputs(9296)) xor (layer2_outputs(6445));
    outputs(9582) <= layer2_outputs(5853);
    outputs(9583) <= not(layer2_outputs(7655));
    outputs(9584) <= (layer2_outputs(8092)) xor (layer2_outputs(4517));
    outputs(9585) <= (layer2_outputs(607)) and (layer2_outputs(653));
    outputs(9586) <= layer2_outputs(9031);
    outputs(9587) <= layer2_outputs(5336);
    outputs(9588) <= layer2_outputs(1353);
    outputs(9589) <= not(layer2_outputs(9274));
    outputs(9590) <= layer2_outputs(9349);
    outputs(9591) <= layer2_outputs(3315);
    outputs(9592) <= not(layer2_outputs(2668));
    outputs(9593) <= (layer2_outputs(8315)) xor (layer2_outputs(4565));
    outputs(9594) <= not((layer2_outputs(2522)) xor (layer2_outputs(9868)));
    outputs(9595) <= (layer2_outputs(1357)) and not (layer2_outputs(7386));
    outputs(9596) <= not(layer2_outputs(3069));
    outputs(9597) <= not(layer2_outputs(9943));
    outputs(9598) <= not(layer2_outputs(7464));
    outputs(9599) <= layer2_outputs(3473);
    outputs(9600) <= layer2_outputs(9354);
    outputs(9601) <= not(layer2_outputs(4821));
    outputs(9602) <= layer2_outputs(3779);
    outputs(9603) <= not((layer2_outputs(5736)) xor (layer2_outputs(6685)));
    outputs(9604) <= not((layer2_outputs(506)) xor (layer2_outputs(9857)));
    outputs(9605) <= not(layer2_outputs(2166));
    outputs(9606) <= layer2_outputs(5136);
    outputs(9607) <= not(layer2_outputs(3999));
    outputs(9608) <= not((layer2_outputs(4875)) xor (layer2_outputs(879)));
    outputs(9609) <= layer2_outputs(5432);
    outputs(9610) <= layer2_outputs(3283);
    outputs(9611) <= not(layer2_outputs(9457));
    outputs(9612) <= layer2_outputs(3230);
    outputs(9613) <= not((layer2_outputs(980)) and (layer2_outputs(4794)));
    outputs(9614) <= not((layer2_outputs(4880)) xor (layer2_outputs(6951)));
    outputs(9615) <= not(layer2_outputs(3955));
    outputs(9616) <= layer2_outputs(2713);
    outputs(9617) <= not(layer2_outputs(3295)) or (layer2_outputs(5897));
    outputs(9618) <= layer2_outputs(1693);
    outputs(9619) <= layer2_outputs(9554);
    outputs(9620) <= layer2_outputs(5075);
    outputs(9621) <= layer2_outputs(3095);
    outputs(9622) <= layer2_outputs(6704);
    outputs(9623) <= not(layer2_outputs(6280));
    outputs(9624) <= (layer2_outputs(2784)) or (layer2_outputs(9607));
    outputs(9625) <= not(layer2_outputs(3482));
    outputs(9626) <= (layer2_outputs(6656)) and not (layer2_outputs(3621));
    outputs(9627) <= not(layer2_outputs(6608));
    outputs(9628) <= not((layer2_outputs(3255)) or (layer2_outputs(7343)));
    outputs(9629) <= (layer2_outputs(8169)) xor (layer2_outputs(4061));
    outputs(9630) <= not((layer2_outputs(2149)) or (layer2_outputs(10187)));
    outputs(9631) <= not((layer2_outputs(3324)) or (layer2_outputs(3962)));
    outputs(9632) <= layer2_outputs(3832);
    outputs(9633) <= not(layer2_outputs(6811));
    outputs(9634) <= not(layer2_outputs(6889)) or (layer2_outputs(6254));
    outputs(9635) <= layer2_outputs(9644);
    outputs(9636) <= layer2_outputs(3989);
    outputs(9637) <= not((layer2_outputs(1044)) xor (layer2_outputs(1430)));
    outputs(9638) <= layer2_outputs(5652);
    outputs(9639) <= not((layer2_outputs(9156)) or (layer2_outputs(1867)));
    outputs(9640) <= layer2_outputs(435);
    outputs(9641) <= layer2_outputs(843);
    outputs(9642) <= not(layer2_outputs(6218));
    outputs(9643) <= layer2_outputs(4732);
    outputs(9644) <= not(layer2_outputs(2852));
    outputs(9645) <= not(layer2_outputs(5127));
    outputs(9646) <= (layer2_outputs(19)) xor (layer2_outputs(6188));
    outputs(9647) <= layer2_outputs(4766);
    outputs(9648) <= (layer2_outputs(2750)) and not (layer2_outputs(7369));
    outputs(9649) <= layer2_outputs(6804);
    outputs(9650) <= not(layer2_outputs(2303));
    outputs(9651) <= not(layer2_outputs(6886));
    outputs(9652) <= not(layer2_outputs(9300));
    outputs(9653) <= not((layer2_outputs(2600)) and (layer2_outputs(8440)));
    outputs(9654) <= layer2_outputs(5955);
    outputs(9655) <= not((layer2_outputs(5335)) and (layer2_outputs(8381)));
    outputs(9656) <= not((layer2_outputs(1590)) xor (layer2_outputs(4207)));
    outputs(9657) <= not(layer2_outputs(3271));
    outputs(9658) <= not((layer2_outputs(9046)) xor (layer2_outputs(1848)));
    outputs(9659) <= (layer2_outputs(9639)) or (layer2_outputs(8057));
    outputs(9660) <= not(layer2_outputs(7464));
    outputs(9661) <= not((layer2_outputs(6809)) xor (layer2_outputs(5277)));
    outputs(9662) <= (layer2_outputs(7039)) and (layer2_outputs(9375));
    outputs(9663) <= (layer2_outputs(6422)) and not (layer2_outputs(2906));
    outputs(9664) <= not((layer2_outputs(6679)) xor (layer2_outputs(6839)));
    outputs(9665) <= not(layer2_outputs(557));
    outputs(9666) <= not((layer2_outputs(4235)) xor (layer2_outputs(16)));
    outputs(9667) <= not((layer2_outputs(1685)) or (layer2_outputs(9732)));
    outputs(9668) <= not(layer2_outputs(7903));
    outputs(9669) <= (layer2_outputs(1675)) xor (layer2_outputs(8112));
    outputs(9670) <= (layer2_outputs(5902)) xor (layer2_outputs(6514));
    outputs(9671) <= layer2_outputs(7298);
    outputs(9672) <= layer2_outputs(8914);
    outputs(9673) <= layer2_outputs(8310);
    outputs(9674) <= (layer2_outputs(5689)) and not (layer2_outputs(10226));
    outputs(9675) <= (layer2_outputs(707)) xor (layer2_outputs(697));
    outputs(9676) <= not((layer2_outputs(2813)) and (layer2_outputs(1538)));
    outputs(9677) <= not((layer2_outputs(5455)) xor (layer2_outputs(7900)));
    outputs(9678) <= not(layer2_outputs(4253));
    outputs(9679) <= layer2_outputs(6063);
    outputs(9680) <= not(layer2_outputs(3592));
    outputs(9681) <= not(layer2_outputs(9941));
    outputs(9682) <= not(layer2_outputs(6570));
    outputs(9683) <= layer2_outputs(4264);
    outputs(9684) <= not(layer2_outputs(8440));
    outputs(9685) <= layer2_outputs(7020);
    outputs(9686) <= layer2_outputs(3670);
    outputs(9687) <= layer2_outputs(3625);
    outputs(9688) <= (layer2_outputs(4497)) xor (layer2_outputs(7263));
    outputs(9689) <= layer2_outputs(6704);
    outputs(9690) <= layer2_outputs(4157);
    outputs(9691) <= not(layer2_outputs(7057));
    outputs(9692) <= layer2_outputs(6883);
    outputs(9693) <= layer2_outputs(9622);
    outputs(9694) <= not((layer2_outputs(9934)) xor (layer2_outputs(7922)));
    outputs(9695) <= (layer2_outputs(5607)) and not (layer2_outputs(5431));
    outputs(9696) <= layer2_outputs(4973);
    outputs(9697) <= layer2_outputs(1294);
    outputs(9698) <= not(layer2_outputs(1052));
    outputs(9699) <= not(layer2_outputs(8727));
    outputs(9700) <= not((layer2_outputs(2366)) xor (layer2_outputs(10180)));
    outputs(9701) <= not(layer2_outputs(8321));
    outputs(9702) <= layer2_outputs(9960);
    outputs(9703) <= not(layer2_outputs(1371));
    outputs(9704) <= layer2_outputs(5529);
    outputs(9705) <= not(layer2_outputs(4765));
    outputs(9706) <= not(layer2_outputs(9369));
    outputs(9707) <= layer2_outputs(9355);
    outputs(9708) <= not(layer2_outputs(9743));
    outputs(9709) <= not((layer2_outputs(8664)) xor (layer2_outputs(9579)));
    outputs(9710) <= (layer2_outputs(10021)) and not (layer2_outputs(410));
    outputs(9711) <= (layer2_outputs(9768)) xor (layer2_outputs(7952));
    outputs(9712) <= layer2_outputs(9327);
    outputs(9713) <= (layer2_outputs(9817)) xor (layer2_outputs(553));
    outputs(9714) <= not(layer2_outputs(7410)) or (layer2_outputs(1305));
    outputs(9715) <= (layer2_outputs(8964)) xor (layer2_outputs(7627));
    outputs(9716) <= layer2_outputs(447);
    outputs(9717) <= layer2_outputs(8545);
    outputs(9718) <= layer2_outputs(9783);
    outputs(9719) <= (layer2_outputs(4092)) and (layer2_outputs(2686));
    outputs(9720) <= not(layer2_outputs(1009));
    outputs(9721) <= (layer2_outputs(6687)) and not (layer2_outputs(3778));
    outputs(9722) <= not(layer2_outputs(4979));
    outputs(9723) <= (layer2_outputs(5548)) xor (layer2_outputs(9614));
    outputs(9724) <= not((layer2_outputs(2864)) and (layer2_outputs(3766)));
    outputs(9725) <= not((layer2_outputs(6942)) xor (layer2_outputs(3122)));
    outputs(9726) <= not((layer2_outputs(1544)) xor (layer2_outputs(8357)));
    outputs(9727) <= layer2_outputs(5159);
    outputs(9728) <= (layer2_outputs(6261)) and not (layer2_outputs(5092));
    outputs(9729) <= layer2_outputs(1647);
    outputs(9730) <= layer2_outputs(1644);
    outputs(9731) <= (layer2_outputs(3760)) xor (layer2_outputs(9310));
    outputs(9732) <= layer2_outputs(5830);
    outputs(9733) <= not((layer2_outputs(10137)) xor (layer2_outputs(3312)));
    outputs(9734) <= not((layer2_outputs(5241)) or (layer2_outputs(9690)));
    outputs(9735) <= not(layer2_outputs(3186));
    outputs(9736) <= layer2_outputs(9821);
    outputs(9737) <= not(layer2_outputs(2646));
    outputs(9738) <= (layer2_outputs(1302)) and not (layer2_outputs(4267));
    outputs(9739) <= layer2_outputs(8675);
    outputs(9740) <= layer2_outputs(3193);
    outputs(9741) <= (layer2_outputs(7612)) xor (layer2_outputs(2882));
    outputs(9742) <= not((layer2_outputs(9148)) or (layer2_outputs(8822)));
    outputs(9743) <= (layer2_outputs(5507)) xor (layer2_outputs(6125));
    outputs(9744) <= (layer2_outputs(6797)) or (layer2_outputs(6364));
    outputs(9745) <= not(layer2_outputs(4936));
    outputs(9746) <= not(layer2_outputs(2400));
    outputs(9747) <= (layer2_outputs(9939)) xor (layer2_outputs(4542));
    outputs(9748) <= not(layer2_outputs(9928));
    outputs(9749) <= not(layer2_outputs(5028));
    outputs(9750) <= (layer2_outputs(4630)) xor (layer2_outputs(7686));
    outputs(9751) <= not((layer2_outputs(2674)) or (layer2_outputs(2153)));
    outputs(9752) <= layer2_outputs(5409);
    outputs(9753) <= not(layer2_outputs(988));
    outputs(9754) <= not(layer2_outputs(5361));
    outputs(9755) <= layer2_outputs(3282);
    outputs(9756) <= layer2_outputs(6169);
    outputs(9757) <= not((layer2_outputs(4764)) xor (layer2_outputs(845)));
    outputs(9758) <= (layer2_outputs(961)) or (layer2_outputs(5499));
    outputs(9759) <= not(layer2_outputs(131));
    outputs(9760) <= layer2_outputs(5023);
    outputs(9761) <= not(layer2_outputs(5022));
    outputs(9762) <= layer2_outputs(5570);
    outputs(9763) <= not((layer2_outputs(7060)) xor (layer2_outputs(807)));
    outputs(9764) <= layer2_outputs(3945);
    outputs(9765) <= not(layer2_outputs(7645));
    outputs(9766) <= (layer2_outputs(359)) xor (layer2_outputs(1730));
    outputs(9767) <= layer2_outputs(2830);
    outputs(9768) <= not(layer2_outputs(475));
    outputs(9769) <= layer2_outputs(647);
    outputs(9770) <= not(layer2_outputs(5281)) or (layer2_outputs(2681));
    outputs(9771) <= not((layer2_outputs(7477)) xor (layer2_outputs(336)));
    outputs(9772) <= not(layer2_outputs(2268));
    outputs(9773) <= (layer2_outputs(3500)) and not (layer2_outputs(2085));
    outputs(9774) <= layer2_outputs(2408);
    outputs(9775) <= not(layer2_outputs(1678));
    outputs(9776) <= not((layer2_outputs(9117)) and (layer2_outputs(7478)));
    outputs(9777) <= not(layer2_outputs(4695));
    outputs(9778) <= layer2_outputs(7309);
    outputs(9779) <= layer2_outputs(2748);
    outputs(9780) <= layer2_outputs(684);
    outputs(9781) <= layer2_outputs(2734);
    outputs(9782) <= not(layer2_outputs(3196));
    outputs(9783) <= not(layer2_outputs(642));
    outputs(9784) <= not(layer2_outputs(3788));
    outputs(9785) <= (layer2_outputs(1823)) xor (layer2_outputs(10114));
    outputs(9786) <= not(layer2_outputs(6459));
    outputs(9787) <= not(layer2_outputs(9881));
    outputs(9788) <= (layer2_outputs(1574)) and not (layer2_outputs(4509));
    outputs(9789) <= layer2_outputs(8704);
    outputs(9790) <= layer2_outputs(4043);
    outputs(9791) <= not(layer2_outputs(8017));
    outputs(9792) <= not(layer2_outputs(5632));
    outputs(9793) <= layer2_outputs(5406);
    outputs(9794) <= layer2_outputs(9448);
    outputs(9795) <= (layer2_outputs(8565)) xor (layer2_outputs(3262));
    outputs(9796) <= not(layer2_outputs(6684));
    outputs(9797) <= layer2_outputs(1367);
    outputs(9798) <= not((layer2_outputs(7596)) xor (layer2_outputs(6610)));
    outputs(9799) <= (layer2_outputs(1773)) xor (layer2_outputs(6102));
    outputs(9800) <= not((layer2_outputs(5162)) or (layer2_outputs(237)));
    outputs(9801) <= not(layer2_outputs(1099));
    outputs(9802) <= not((layer2_outputs(155)) and (layer2_outputs(1009)));
    outputs(9803) <= not(layer2_outputs(480));
    outputs(9804) <= layer2_outputs(2538);
    outputs(9805) <= layer2_outputs(5038);
    outputs(9806) <= layer2_outputs(1276);
    outputs(9807) <= (layer2_outputs(4594)) xor (layer2_outputs(2441));
    outputs(9808) <= (layer2_outputs(3393)) xor (layer2_outputs(2437));
    outputs(9809) <= layer2_outputs(247);
    outputs(9810) <= (layer2_outputs(2750)) xor (layer2_outputs(7795));
    outputs(9811) <= not(layer2_outputs(6027));
    outputs(9812) <= (layer2_outputs(156)) xor (layer2_outputs(8169));
    outputs(9813) <= layer2_outputs(8656);
    outputs(9814) <= layer2_outputs(6840);
    outputs(9815) <= not(layer2_outputs(555));
    outputs(9816) <= layer2_outputs(1993);
    outputs(9817) <= (layer2_outputs(2048)) or (layer2_outputs(1895));
    outputs(9818) <= (layer2_outputs(6781)) xor (layer2_outputs(10221));
    outputs(9819) <= layer2_outputs(1529);
    outputs(9820) <= layer2_outputs(6984);
    outputs(9821) <= layer2_outputs(3648);
    outputs(9822) <= not((layer2_outputs(836)) xor (layer2_outputs(10096)));
    outputs(9823) <= not(layer2_outputs(6319));
    outputs(9824) <= not(layer2_outputs(3571)) or (layer2_outputs(6600));
    outputs(9825) <= not(layer2_outputs(2566));
    outputs(9826) <= not((layer2_outputs(7669)) xor (layer2_outputs(7740)));
    outputs(9827) <= not(layer2_outputs(6134)) or (layer2_outputs(7348));
    outputs(9828) <= layer2_outputs(4010);
    outputs(9829) <= (layer2_outputs(8892)) xor (layer2_outputs(7166));
    outputs(9830) <= not(layer2_outputs(10108)) or (layer2_outputs(827));
    outputs(9831) <= layer2_outputs(8330);
    outputs(9832) <= not(layer2_outputs(10066));
    outputs(9833) <= layer2_outputs(7151);
    outputs(9834) <= layer2_outputs(4170);
    outputs(9835) <= layer2_outputs(9263);
    outputs(9836) <= not(layer2_outputs(6049));
    outputs(9837) <= not((layer2_outputs(6166)) xor (layer2_outputs(4019)));
    outputs(9838) <= not(layer2_outputs(5063));
    outputs(9839) <= not(layer2_outputs(4750));
    outputs(9840) <= not((layer2_outputs(6469)) or (layer2_outputs(6986)));
    outputs(9841) <= not((layer2_outputs(9311)) and (layer2_outputs(5686)));
    outputs(9842) <= not((layer2_outputs(9937)) xor (layer2_outputs(4219)));
    outputs(9843) <= (layer2_outputs(2211)) xor (layer2_outputs(6328));
    outputs(9844) <= layer2_outputs(951);
    outputs(9845) <= layer2_outputs(8708);
    outputs(9846) <= (layer2_outputs(7411)) and not (layer2_outputs(5495));
    outputs(9847) <= not(layer2_outputs(835));
    outputs(9848) <= layer2_outputs(5388);
    outputs(9849) <= layer2_outputs(8028);
    outputs(9850) <= (layer2_outputs(9974)) and (layer2_outputs(8439));
    outputs(9851) <= not(layer2_outputs(10228));
    outputs(9852) <= layer2_outputs(3625);
    outputs(9853) <= layer2_outputs(3821);
    outputs(9854) <= (layer2_outputs(4919)) and (layer2_outputs(5763));
    outputs(9855) <= not(layer2_outputs(5933));
    outputs(9856) <= not(layer2_outputs(5482));
    outputs(9857) <= layer2_outputs(10208);
    outputs(9858) <= not(layer2_outputs(7034));
    outputs(9859) <= layer2_outputs(8225);
    outputs(9860) <= not((layer2_outputs(6133)) or (layer2_outputs(2176)));
    outputs(9861) <= (layer2_outputs(5425)) xor (layer2_outputs(4220));
    outputs(9862) <= not(layer2_outputs(4933));
    outputs(9863) <= layer2_outputs(5269);
    outputs(9864) <= layer2_outputs(9354);
    outputs(9865) <= layer2_outputs(2086);
    outputs(9866) <= layer2_outputs(8051);
    outputs(9867) <= not((layer2_outputs(8873)) or (layer2_outputs(465)));
    outputs(9868) <= not(layer2_outputs(9116));
    outputs(9869) <= not(layer2_outputs(5355));
    outputs(9870) <= (layer2_outputs(7583)) xor (layer2_outputs(9964));
    outputs(9871) <= not((layer2_outputs(4756)) xor (layer2_outputs(5963)));
    outputs(9872) <= (layer2_outputs(4093)) xor (layer2_outputs(3098));
    outputs(9873) <= not(layer2_outputs(2410));
    outputs(9874) <= not(layer2_outputs(2399));
    outputs(9875) <= layer2_outputs(1117);
    outputs(9876) <= not(layer2_outputs(7710));
    outputs(9877) <= not((layer2_outputs(8740)) or (layer2_outputs(4965)));
    outputs(9878) <= (layer2_outputs(919)) and (layer2_outputs(9071));
    outputs(9879) <= layer2_outputs(8269);
    outputs(9880) <= not(layer2_outputs(7595));
    outputs(9881) <= (layer2_outputs(6291)) xor (layer2_outputs(4035));
    outputs(9882) <= (layer2_outputs(5155)) xor (layer2_outputs(3465));
    outputs(9883) <= not(layer2_outputs(5495));
    outputs(9884) <= not(layer2_outputs(3007));
    outputs(9885) <= not(layer2_outputs(5813));
    outputs(9886) <= (layer2_outputs(7751)) xor (layer2_outputs(10096));
    outputs(9887) <= (layer2_outputs(3744)) and (layer2_outputs(1509));
    outputs(9888) <= (layer2_outputs(7861)) and not (layer2_outputs(375));
    outputs(9889) <= layer2_outputs(1523);
    outputs(9890) <= not((layer2_outputs(8828)) or (layer2_outputs(4160)));
    outputs(9891) <= layer2_outputs(1056);
    outputs(9892) <= not(layer2_outputs(2873));
    outputs(9893) <= not(layer2_outputs(4752));
    outputs(9894) <= layer2_outputs(4596);
    outputs(9895) <= (layer2_outputs(6069)) or (layer2_outputs(6829));
    outputs(9896) <= layer2_outputs(4595);
    outputs(9897) <= layer2_outputs(503);
    outputs(9898) <= layer2_outputs(1306);
    outputs(9899) <= not((layer2_outputs(4724)) xor (layer2_outputs(1778)));
    outputs(9900) <= layer2_outputs(4890);
    outputs(9901) <= layer2_outputs(5858);
    outputs(9902) <= layer2_outputs(5202);
    outputs(9903) <= not(layer2_outputs(7014));
    outputs(9904) <= layer2_outputs(8809);
    outputs(9905) <= (layer2_outputs(527)) or (layer2_outputs(1675));
    outputs(9906) <= not(layer2_outputs(7830));
    outputs(9907) <= layer2_outputs(122);
    outputs(9908) <= not(layer2_outputs(5454));
    outputs(9909) <= not((layer2_outputs(6095)) or (layer2_outputs(1202)));
    outputs(9910) <= not((layer2_outputs(524)) xor (layer2_outputs(728)));
    outputs(9911) <= not(layer2_outputs(1801));
    outputs(9912) <= not(layer2_outputs(9583));
    outputs(9913) <= layer2_outputs(6540);
    outputs(9914) <= not(layer2_outputs(9584));
    outputs(9915) <= layer2_outputs(5999);
    outputs(9916) <= not(layer2_outputs(4276));
    outputs(9917) <= not((layer2_outputs(9276)) and (layer2_outputs(2107)));
    outputs(9918) <= layer2_outputs(2748);
    outputs(9919) <= layer2_outputs(5186);
    outputs(9920) <= not(layer2_outputs(4117));
    outputs(9921) <= layer2_outputs(2516);
    outputs(9922) <= layer2_outputs(8475);
    outputs(9923) <= layer2_outputs(9359);
    outputs(9924) <= not(layer2_outputs(5201));
    outputs(9925) <= layer2_outputs(5755);
    outputs(9926) <= not(layer2_outputs(5265));
    outputs(9927) <= not(layer2_outputs(2014));
    outputs(9928) <= not(layer2_outputs(4729));
    outputs(9929) <= (layer2_outputs(4290)) and not (layer2_outputs(1110));
    outputs(9930) <= not((layer2_outputs(3168)) and (layer2_outputs(10094)));
    outputs(9931) <= not(layer2_outputs(2977));
    outputs(9932) <= (layer2_outputs(9870)) xor (layer2_outputs(6140));
    outputs(9933) <= (layer2_outputs(3204)) xor (layer2_outputs(2404));
    outputs(9934) <= not(layer2_outputs(3771));
    outputs(9935) <= not(layer2_outputs(406));
    outputs(9936) <= not(layer2_outputs(6655));
    outputs(9937) <= (layer2_outputs(5255)) xor (layer2_outputs(867));
    outputs(9938) <= not(layer2_outputs(4782));
    outputs(9939) <= layer2_outputs(4758);
    outputs(9940) <= not(layer2_outputs(5162));
    outputs(9941) <= not(layer2_outputs(8856));
    outputs(9942) <= (layer2_outputs(4127)) xor (layer2_outputs(8677));
    outputs(9943) <= layer2_outputs(6330);
    outputs(9944) <= layer2_outputs(5110);
    outputs(9945) <= layer2_outputs(9966);
    outputs(9946) <= not(layer2_outputs(6790));
    outputs(9947) <= not(layer2_outputs(8308));
    outputs(9948) <= not(layer2_outputs(6275));
    outputs(9949) <= layer2_outputs(9976);
    outputs(9950) <= layer2_outputs(4114);
    outputs(9951) <= layer2_outputs(5339);
    outputs(9952) <= layer2_outputs(8320);
    outputs(9953) <= layer2_outputs(2830);
    outputs(9954) <= layer2_outputs(7024);
    outputs(9955) <= layer2_outputs(7757);
    outputs(9956) <= layer2_outputs(5227);
    outputs(9957) <= (layer2_outputs(7806)) xor (layer2_outputs(5478));
    outputs(9958) <= not(layer2_outputs(5781));
    outputs(9959) <= not((layer2_outputs(178)) or (layer2_outputs(8928)));
    outputs(9960) <= layer2_outputs(4870);
    outputs(9961) <= layer2_outputs(5694);
    outputs(9962) <= not(layer2_outputs(4905));
    outputs(9963) <= not(layer2_outputs(6002));
    outputs(9964) <= not(layer2_outputs(9133));
    outputs(9965) <= layer2_outputs(4684);
    outputs(9966) <= layer2_outputs(4004);
    outputs(9967) <= not((layer2_outputs(3134)) xor (layer2_outputs(396)));
    outputs(9968) <= not(layer2_outputs(7181));
    outputs(9969) <= layer2_outputs(804);
    outputs(9970) <= not(layer2_outputs(10167));
    outputs(9971) <= layer2_outputs(598);
    outputs(9972) <= layer2_outputs(8748);
    outputs(9973) <= not((layer2_outputs(9285)) xor (layer2_outputs(3794)));
    outputs(9974) <= layer2_outputs(7899);
    outputs(9975) <= not(layer2_outputs(4016));
    outputs(9976) <= not(layer2_outputs(8111));
    outputs(9977) <= not((layer2_outputs(8535)) xor (layer2_outputs(3149)));
    outputs(9978) <= not(layer2_outputs(726));
    outputs(9979) <= not(layer2_outputs(2590));
    outputs(9980) <= layer2_outputs(10139);
    outputs(9981) <= not((layer2_outputs(6583)) xor (layer2_outputs(5258)));
    outputs(9982) <= layer2_outputs(3735);
    outputs(9983) <= layer2_outputs(2155);
    outputs(9984) <= layer2_outputs(4261);
    outputs(9985) <= (layer2_outputs(1976)) xor (layer2_outputs(8177));
    outputs(9986) <= not(layer2_outputs(3184));
    outputs(9987) <= (layer2_outputs(3348)) xor (layer2_outputs(5584));
    outputs(9988) <= layer2_outputs(5611);
    outputs(9989) <= layer2_outputs(4891);
    outputs(9990) <= layer2_outputs(1741);
    outputs(9991) <= layer2_outputs(8046);
    outputs(9992) <= (layer2_outputs(7531)) xor (layer2_outputs(8975));
    outputs(9993) <= not((layer2_outputs(6581)) xor (layer2_outputs(8599)));
    outputs(9994) <= (layer2_outputs(6637)) or (layer2_outputs(8067));
    outputs(9995) <= layer2_outputs(8951);
    outputs(9996) <= (layer2_outputs(8208)) xor (layer2_outputs(1068));
    outputs(9997) <= (layer2_outputs(4088)) and (layer2_outputs(1694));
    outputs(9998) <= not((layer2_outputs(8162)) xor (layer2_outputs(9126)));
    outputs(9999) <= not(layer2_outputs(2601));
    outputs(10000) <= not(layer2_outputs(6452)) or (layer2_outputs(9107));
    outputs(10001) <= (layer2_outputs(5612)) and (layer2_outputs(7206));
    outputs(10002) <= not((layer2_outputs(1032)) xor (layer2_outputs(3953)));
    outputs(10003) <= not(layer2_outputs(394));
    outputs(10004) <= not(layer2_outputs(3740));
    outputs(10005) <= (layer2_outputs(6749)) and not (layer2_outputs(9367));
    outputs(10006) <= layer2_outputs(3350);
    outputs(10007) <= not(layer2_outputs(10152));
    outputs(10008) <= layer2_outputs(8261);
    outputs(10009) <= layer2_outputs(4856);
    outputs(10010) <= (layer2_outputs(9146)) and not (layer2_outputs(1874));
    outputs(10011) <= layer2_outputs(277);
    outputs(10012) <= not((layer2_outputs(6070)) xor (layer2_outputs(3641)));
    outputs(10013) <= not((layer2_outputs(6904)) xor (layer2_outputs(9376)));
    outputs(10014) <= not(layer2_outputs(5168));
    outputs(10015) <= layer2_outputs(1348);
    outputs(10016) <= layer2_outputs(1863);
    outputs(10017) <= layer2_outputs(706);
    outputs(10018) <= (layer2_outputs(2310)) xor (layer2_outputs(221));
    outputs(10019) <= not((layer2_outputs(2616)) and (layer2_outputs(386)));
    outputs(10020) <= layer2_outputs(7018);
    outputs(10021) <= not(layer2_outputs(7339));
    outputs(10022) <= not(layer2_outputs(9430));
    outputs(10023) <= not(layer2_outputs(7234));
    outputs(10024) <= not(layer2_outputs(8333));
    outputs(10025) <= layer2_outputs(864);
    outputs(10026) <= layer2_outputs(2524);
    outputs(10027) <= not((layer2_outputs(5655)) xor (layer2_outputs(1478)));
    outputs(10028) <= layer2_outputs(8720);
    outputs(10029) <= not(layer2_outputs(4276));
    outputs(10030) <= layer2_outputs(3287);
    outputs(10031) <= layer2_outputs(7458);
    outputs(10032) <= layer2_outputs(8148);
    outputs(10033) <= layer2_outputs(2626);
    outputs(10034) <= not((layer2_outputs(8172)) xor (layer2_outputs(4893)));
    outputs(10035) <= not((layer2_outputs(5005)) xor (layer2_outputs(8041)));
    outputs(10036) <= layer2_outputs(9316);
    outputs(10037) <= not(layer2_outputs(6899));
    outputs(10038) <= not(layer2_outputs(6998)) or (layer2_outputs(4708));
    outputs(10039) <= not(layer2_outputs(10181));
    outputs(10040) <= not((layer2_outputs(6884)) xor (layer2_outputs(3730)));
    outputs(10041) <= not(layer2_outputs(6866));
    outputs(10042) <= layer2_outputs(4155);
    outputs(10043) <= layer2_outputs(6542);
    outputs(10044) <= not(layer2_outputs(2430));
    outputs(10045) <= not((layer2_outputs(2107)) xor (layer2_outputs(3544)));
    outputs(10046) <= not((layer2_outputs(8923)) xor (layer2_outputs(289)));
    outputs(10047) <= not(layer2_outputs(7815));
    outputs(10048) <= not(layer2_outputs(1508));
    outputs(10049) <= not(layer2_outputs(6947));
    outputs(10050) <= not(layer2_outputs(8776));
    outputs(10051) <= layer2_outputs(559);
    outputs(10052) <= not(layer2_outputs(6093)) or (layer2_outputs(7534));
    outputs(10053) <= not(layer2_outputs(2259));
    outputs(10054) <= not(layer2_outputs(3778));
    outputs(10055) <= not(layer2_outputs(7801));
    outputs(10056) <= (layer2_outputs(6629)) xor (layer2_outputs(4270));
    outputs(10057) <= not(layer2_outputs(9101));
    outputs(10058) <= layer2_outputs(8771);
    outputs(10059) <= not((layer2_outputs(3894)) xor (layer2_outputs(3510)));
    outputs(10060) <= not(layer2_outputs(1203));
    outputs(10061) <= (layer2_outputs(3699)) xor (layer2_outputs(6005));
    outputs(10062) <= not((layer2_outputs(5493)) and (layer2_outputs(7004)));
    outputs(10063) <= layer2_outputs(9952);
    outputs(10064) <= not(layer2_outputs(6446));
    outputs(10065) <= layer2_outputs(251);
    outputs(10066) <= layer2_outputs(4145);
    outputs(10067) <= not(layer2_outputs(1926));
    outputs(10068) <= not(layer2_outputs(7848));
    outputs(10069) <= layer2_outputs(4260);
    outputs(10070) <= not(layer2_outputs(1837));
    outputs(10071) <= layer2_outputs(6712);
    outputs(10072) <= layer2_outputs(250);
    outputs(10073) <= (layer2_outputs(422)) or (layer2_outputs(1469));
    outputs(10074) <= not(layer2_outputs(8429));
    outputs(10075) <= layer2_outputs(8456);
    outputs(10076) <= layer2_outputs(2496);
    outputs(10077) <= (layer2_outputs(3525)) xor (layer2_outputs(1740));
    outputs(10078) <= not(layer2_outputs(9834));
    outputs(10079) <= not(layer2_outputs(7571));
    outputs(10080) <= layer2_outputs(997);
    outputs(10081) <= layer2_outputs(9082);
    outputs(10082) <= not((layer2_outputs(4050)) and (layer2_outputs(765)));
    outputs(10083) <= not(layer2_outputs(1761)) or (layer2_outputs(97));
    outputs(10084) <= not(layer2_outputs(9823));
    outputs(10085) <= not(layer2_outputs(4701));
    outputs(10086) <= layer2_outputs(3389);
    outputs(10087) <= not(layer2_outputs(1423));
    outputs(10088) <= (layer2_outputs(704)) and not (layer2_outputs(7454));
    outputs(10089) <= not(layer2_outputs(3382));
    outputs(10090) <= not(layer2_outputs(1135));
    outputs(10091) <= (layer2_outputs(3632)) and not (layer2_outputs(4051));
    outputs(10092) <= not(layer2_outputs(3033));
    outputs(10093) <= layer2_outputs(6492);
    outputs(10094) <= (layer2_outputs(5929)) or (layer2_outputs(5074));
    outputs(10095) <= (layer2_outputs(1696)) and not (layer2_outputs(2828));
    outputs(10096) <= layer2_outputs(1884);
    outputs(10097) <= not(layer2_outputs(986));
    outputs(10098) <= not((layer2_outputs(5988)) xor (layer2_outputs(5194)));
    outputs(10099) <= not(layer2_outputs(9093));
    outputs(10100) <= not(layer2_outputs(2294));
    outputs(10101) <= (layer2_outputs(7453)) and not (layer2_outputs(853));
    outputs(10102) <= not((layer2_outputs(6698)) xor (layer2_outputs(6628)));
    outputs(10103) <= layer2_outputs(1367);
    outputs(10104) <= layer2_outputs(4100);
    outputs(10105) <= not((layer2_outputs(1146)) xor (layer2_outputs(1296)));
    outputs(10106) <= (layer2_outputs(443)) and not (layer2_outputs(3519));
    outputs(10107) <= layer2_outputs(8987);
    outputs(10108) <= (layer2_outputs(1877)) and not (layer2_outputs(5867));
    outputs(10109) <= (layer2_outputs(1179)) and (layer2_outputs(3534));
    outputs(10110) <= layer2_outputs(4993);
    outputs(10111) <= layer2_outputs(2916);
    outputs(10112) <= not(layer2_outputs(5618));
    outputs(10113) <= not(layer2_outputs(7544));
    outputs(10114) <= layer2_outputs(6399);
    outputs(10115) <= (layer2_outputs(6142)) xor (layer2_outputs(9773));
    outputs(10116) <= not((layer2_outputs(3463)) xor (layer2_outputs(431)));
    outputs(10117) <= (layer2_outputs(3836)) xor (layer2_outputs(1420));
    outputs(10118) <= not((layer2_outputs(1930)) or (layer2_outputs(3793)));
    outputs(10119) <= (layer2_outputs(3480)) xor (layer2_outputs(3095));
    outputs(10120) <= (layer2_outputs(7469)) and (layer2_outputs(5439));
    outputs(10121) <= (layer2_outputs(8812)) xor (layer2_outputs(2785));
    outputs(10122) <= not(layer2_outputs(3236));
    outputs(10123) <= layer2_outputs(2654);
    outputs(10124) <= layer2_outputs(9639);
    outputs(10125) <= layer2_outputs(2826);
    outputs(10126) <= not(layer2_outputs(4671));
    outputs(10127) <= not(layer2_outputs(4445));
    outputs(10128) <= layer2_outputs(4372);
    outputs(10129) <= not(layer2_outputs(2690));
    outputs(10130) <= '1';
    outputs(10131) <= not(layer2_outputs(4422)) or (layer2_outputs(4274));
    outputs(10132) <= layer2_outputs(7518);
    outputs(10133) <= (layer2_outputs(5619)) and (layer2_outputs(1119));
    outputs(10134) <= not(layer2_outputs(8447));
    outputs(10135) <= layer2_outputs(142);
    outputs(10136) <= layer2_outputs(2724);
    outputs(10137) <= not(layer2_outputs(8025));
    outputs(10138) <= not(layer2_outputs(3755));
    outputs(10139) <= (layer2_outputs(4428)) xor (layer2_outputs(10112));
    outputs(10140) <= not(layer2_outputs(2792)) or (layer2_outputs(111));
    outputs(10141) <= not(layer2_outputs(565));
    outputs(10142) <= layer2_outputs(167);
    outputs(10143) <= not(layer2_outputs(786));
    outputs(10144) <= (layer2_outputs(1259)) and not (layer2_outputs(9950));
    outputs(10145) <= not((layer2_outputs(9189)) xor (layer2_outputs(6949)));
    outputs(10146) <= not(layer2_outputs(2758)) or (layer2_outputs(5940));
    outputs(10147) <= not((layer2_outputs(4314)) or (layer2_outputs(2021)));
    outputs(10148) <= layer2_outputs(380);
    outputs(10149) <= not(layer2_outputs(7115));
    outputs(10150) <= layer2_outputs(8513);
    outputs(10151) <= layer2_outputs(4616);
    outputs(10152) <= layer2_outputs(3427);
    outputs(10153) <= not(layer2_outputs(4838));
    outputs(10154) <= not(layer2_outputs(6035));
    outputs(10155) <= layer2_outputs(7591);
    outputs(10156) <= not(layer2_outputs(1660));
    outputs(10157) <= not(layer2_outputs(7122));
    outputs(10158) <= (layer2_outputs(4620)) xor (layer2_outputs(4548));
    outputs(10159) <= not((layer2_outputs(2891)) xor (layer2_outputs(1276)));
    outputs(10160) <= not(layer2_outputs(10019));
    outputs(10161) <= not(layer2_outputs(7889));
    outputs(10162) <= layer2_outputs(5367);
    outputs(10163) <= (layer2_outputs(8585)) and (layer2_outputs(6302));
    outputs(10164) <= not(layer2_outputs(7790));
    outputs(10165) <= (layer2_outputs(2862)) xor (layer2_outputs(2251));
    outputs(10166) <= not(layer2_outputs(7196));
    outputs(10167) <= layer2_outputs(9151);
    outputs(10168) <= (layer2_outputs(6015)) and not (layer2_outputs(9687));
    outputs(10169) <= not(layer2_outputs(1251));
    outputs(10170) <= layer2_outputs(2840);
    outputs(10171) <= not((layer2_outputs(1142)) xor (layer2_outputs(2394)));
    outputs(10172) <= not(layer2_outputs(3817));
    outputs(10173) <= not((layer2_outputs(9942)) xor (layer2_outputs(7972)));
    outputs(10174) <= layer2_outputs(672);
    outputs(10175) <= not(layer2_outputs(2992));
    outputs(10176) <= not((layer2_outputs(1284)) and (layer2_outputs(1366)));
    outputs(10177) <= layer2_outputs(8433);
    outputs(10178) <= not(layer2_outputs(4913));
    outputs(10179) <= not(layer2_outputs(6912));
    outputs(10180) <= not(layer2_outputs(1054));
    outputs(10181) <= (layer2_outputs(8428)) and (layer2_outputs(5531));
    outputs(10182) <= not((layer2_outputs(5891)) or (layer2_outputs(105)));
    outputs(10183) <= not(layer2_outputs(2523));
    outputs(10184) <= not(layer2_outputs(5188));
    outputs(10185) <= layer2_outputs(7092);
    outputs(10186) <= not((layer2_outputs(5605)) xor (layer2_outputs(5178)));
    outputs(10187) <= layer2_outputs(9017);
    outputs(10188) <= not(layer2_outputs(2116));
    outputs(10189) <= not(layer2_outputs(4823));
    outputs(10190) <= not(layer2_outputs(1169));
    outputs(10191) <= layer2_outputs(3643);
    outputs(10192) <= not(layer2_outputs(2774));
    outputs(10193) <= not(layer2_outputs(4154)) or (layer2_outputs(7660));
    outputs(10194) <= layer2_outputs(697);
    outputs(10195) <= (layer2_outputs(8236)) xor (layer2_outputs(2771));
    outputs(10196) <= (layer2_outputs(5468)) xor (layer2_outputs(8534));
    outputs(10197) <= layer2_outputs(8915);
    outputs(10198) <= (layer2_outputs(9575)) xor (layer2_outputs(6876));
    outputs(10199) <= not(layer2_outputs(4420));
    outputs(10200) <= layer2_outputs(6142);
    outputs(10201) <= (layer2_outputs(2496)) and (layer2_outputs(4427));
    outputs(10202) <= not(layer2_outputs(7072));
    outputs(10203) <= not((layer2_outputs(8796)) and (layer2_outputs(9502)));
    outputs(10204) <= layer2_outputs(5029);
    outputs(10205) <= layer2_outputs(2464);
    outputs(10206) <= layer2_outputs(5412);
    outputs(10207) <= (layer2_outputs(7013)) or (layer2_outputs(10069));
    outputs(10208) <= layer2_outputs(4954);
    outputs(10209) <= layer2_outputs(6852);
    outputs(10210) <= not(layer2_outputs(9834));
    outputs(10211) <= not(layer2_outputs(4259));
    outputs(10212) <= not(layer2_outputs(5374));
    outputs(10213) <= (layer2_outputs(5121)) xor (layer2_outputs(5944));
    outputs(10214) <= (layer2_outputs(7563)) and not (layer2_outputs(10093));
    outputs(10215) <= not((layer2_outputs(9685)) xor (layer2_outputs(3923)));
    outputs(10216) <= not((layer2_outputs(4669)) and (layer2_outputs(7572)));
    outputs(10217) <= layer2_outputs(8810);
    outputs(10218) <= not(layer2_outputs(3580));
    outputs(10219) <= not(layer2_outputs(3594));
    outputs(10220) <= not(layer2_outputs(2651));
    outputs(10221) <= not((layer2_outputs(7178)) or (layer2_outputs(5823)));
    outputs(10222) <= not(layer2_outputs(5504)) or (layer2_outputs(4459));
    outputs(10223) <= (layer2_outputs(968)) xor (layer2_outputs(7005));
    outputs(10224) <= (layer2_outputs(1028)) xor (layer2_outputs(8533));
    outputs(10225) <= layer2_outputs(7789);
    outputs(10226) <= layer2_outputs(7482);
    outputs(10227) <= layer2_outputs(10040);
    outputs(10228) <= not((layer2_outputs(1861)) xor (layer2_outputs(3445)));
    outputs(10229) <= not(layer2_outputs(300));
    outputs(10230) <= layer2_outputs(1982);
    outputs(10231) <= layer2_outputs(3512);
    outputs(10232) <= (layer2_outputs(652)) xor (layer2_outputs(66));
    outputs(10233) <= not(layer2_outputs(2226));
    outputs(10234) <= (layer2_outputs(1910)) xor (layer2_outputs(5569));
    outputs(10235) <= not(layer2_outputs(882));
    outputs(10236) <= (layer2_outputs(4443)) and (layer2_outputs(6865));
    outputs(10237) <= layer2_outputs(5904);
    outputs(10238) <= layer2_outputs(9327);
    outputs(10239) <= layer2_outputs(7717);

end Behavioral;
