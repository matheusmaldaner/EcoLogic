module logic_network(
    input wire [255:0] inputs,
    output wire [9:0] outputs
);

    wire [5119:0] layer0_outputs;

    assign layer0_outputs[0] = (inputs[68]) & ~(inputs[17]);
    assign layer0_outputs[1] = (inputs[232]) ^ (inputs[239]);
    assign layer0_outputs[2] = ~(inputs[243]);
    assign layer0_outputs[3] = ~(inputs[41]);
    assign layer0_outputs[4] = ~(inputs[78]) | (inputs[142]);
    assign layer0_outputs[5] = ~(inputs[19]);
    assign layer0_outputs[6] = ~(inputs[90]) | (inputs[47]);
    assign layer0_outputs[7] = ~((inputs[233]) | (inputs[90]));
    assign layer0_outputs[8] = (inputs[197]) ^ (inputs[51]);
    assign layer0_outputs[9] = ~((inputs[101]) ^ (inputs[8]));
    assign layer0_outputs[10] = (inputs[92]) & ~(inputs[51]);
    assign layer0_outputs[11] = (inputs[196]) | (inputs[99]);
    assign layer0_outputs[12] = ~((inputs[8]) ^ (inputs[131]));
    assign layer0_outputs[13] = (inputs[201]) | (inputs[37]);
    assign layer0_outputs[14] = (inputs[252]) ^ (inputs[22]);
    assign layer0_outputs[15] = inputs[237];
    assign layer0_outputs[16] = (inputs[161]) & (inputs[59]);
    assign layer0_outputs[17] = inputs[67];
    assign layer0_outputs[18] = (inputs[157]) & ~(inputs[35]);
    assign layer0_outputs[19] = ~(inputs[69]) | (inputs[209]);
    assign layer0_outputs[20] = (inputs[50]) ^ (inputs[177]);
    assign layer0_outputs[21] = inputs[246];
    assign layer0_outputs[22] = (inputs[160]) & ~(inputs[1]);
    assign layer0_outputs[23] = ~(inputs[37]);
    assign layer0_outputs[24] = (inputs[158]) | (inputs[141]);
    assign layer0_outputs[25] = ~(inputs[100]);
    assign layer0_outputs[26] = inputs[157];
    assign layer0_outputs[27] = 1'b0;
    assign layer0_outputs[28] = inputs[69];
    assign layer0_outputs[29] = ~((inputs[247]) ^ (inputs[218]));
    assign layer0_outputs[30] = ~((inputs[149]) ^ (inputs[19]));
    assign layer0_outputs[31] = inputs[72];
    assign layer0_outputs[32] = ~(inputs[27]) | (inputs[209]);
    assign layer0_outputs[33] = ~(inputs[174]) | (inputs[47]);
    assign layer0_outputs[34] = ~(inputs[235]);
    assign layer0_outputs[35] = ~((inputs[184]) | (inputs[250]));
    assign layer0_outputs[36] = inputs[20];
    assign layer0_outputs[37] = 1'b1;
    assign layer0_outputs[38] = inputs[221];
    assign layer0_outputs[39] = ~((inputs[124]) | (inputs[189]));
    assign layer0_outputs[40] = ~((inputs[166]) ^ (inputs[4]));
    assign layer0_outputs[41] = ~((inputs[100]) | (inputs[12]));
    assign layer0_outputs[42] = ~(inputs[232]) | (inputs[171]);
    assign layer0_outputs[43] = ~(inputs[68]);
    assign layer0_outputs[44] = ~((inputs[250]) | (inputs[215]));
    assign layer0_outputs[45] = (inputs[157]) | (inputs[194]);
    assign layer0_outputs[46] = (inputs[140]) ^ (inputs[14]);
    assign layer0_outputs[47] = ~((inputs[202]) | (inputs[189]));
    assign layer0_outputs[48] = (inputs[219]) | (inputs[84]);
    assign layer0_outputs[49] = (inputs[178]) | (inputs[65]);
    assign layer0_outputs[50] = (inputs[217]) & ~(inputs[208]);
    assign layer0_outputs[51] = (inputs[106]) | (inputs[5]);
    assign layer0_outputs[52] = (inputs[92]) | (inputs[122]);
    assign layer0_outputs[53] = ~((inputs[59]) | (inputs[162]));
    assign layer0_outputs[54] = ~((inputs[40]) | (inputs[174]));
    assign layer0_outputs[55] = ~((inputs[227]) ^ (inputs[243]));
    assign layer0_outputs[56] = ~(inputs[92]);
    assign layer0_outputs[57] = ~((inputs[44]) | (inputs[99]));
    assign layer0_outputs[58] = (inputs[70]) | (inputs[251]);
    assign layer0_outputs[59] = ~(inputs[185]) | (inputs[240]);
    assign layer0_outputs[60] = ~((inputs[7]) | (inputs[234]));
    assign layer0_outputs[61] = (inputs[143]) & ~(inputs[178]);
    assign layer0_outputs[62] = 1'b0;
    assign layer0_outputs[63] = (inputs[186]) ^ (inputs[52]);
    assign layer0_outputs[64] = (inputs[23]) ^ (inputs[29]);
    assign layer0_outputs[65] = inputs[143];
    assign layer0_outputs[66] = ~(inputs[21]);
    assign layer0_outputs[67] = ~(inputs[152]) | (inputs[73]);
    assign layer0_outputs[68] = (inputs[48]) & (inputs[223]);
    assign layer0_outputs[69] = inputs[202];
    assign layer0_outputs[70] = inputs[229];
    assign layer0_outputs[71] = (inputs[237]) | (inputs[56]);
    assign layer0_outputs[72] = (inputs[193]) & ~(inputs[31]);
    assign layer0_outputs[73] = ~(inputs[111]) | (inputs[235]);
    assign layer0_outputs[74] = ~((inputs[47]) | (inputs[253]));
    assign layer0_outputs[75] = (inputs[97]) & (inputs[89]);
    assign layer0_outputs[76] = (inputs[178]) & (inputs[244]);
    assign layer0_outputs[77] = 1'b0;
    assign layer0_outputs[78] = (inputs[181]) | (inputs[59]);
    assign layer0_outputs[79] = ~((inputs[2]) & (inputs[20]));
    assign layer0_outputs[80] = ~((inputs[135]) | (inputs[197]));
    assign layer0_outputs[81] = (inputs[240]) & ~(inputs[101]);
    assign layer0_outputs[82] = ~(inputs[103]);
    assign layer0_outputs[83] = (inputs[234]) ^ (inputs[82]);
    assign layer0_outputs[84] = (inputs[153]) | (inputs[132]);
    assign layer0_outputs[85] = (inputs[47]) | (inputs[84]);
    assign layer0_outputs[86] = (inputs[206]) ^ (inputs[102]);
    assign layer0_outputs[87] = (inputs[70]) & ~(inputs[242]);
    assign layer0_outputs[88] = (inputs[83]) ^ (inputs[174]);
    assign layer0_outputs[89] = ~((inputs[39]) | (inputs[40]));
    assign layer0_outputs[90] = ~((inputs[7]) ^ (inputs[181]));
    assign layer0_outputs[91] = (inputs[98]) | (inputs[166]);
    assign layer0_outputs[92] = (inputs[225]) & ~(inputs[248]);
    assign layer0_outputs[93] = ~((inputs[58]) | (inputs[150]));
    assign layer0_outputs[94] = ~((inputs[243]) ^ (inputs[242]));
    assign layer0_outputs[95] = (inputs[114]) ^ (inputs[174]);
    assign layer0_outputs[96] = ~((inputs[237]) | (inputs[236]));
    assign layer0_outputs[97] = inputs[199];
    assign layer0_outputs[98] = (inputs[236]) ^ (inputs[185]);
    assign layer0_outputs[99] = ~(inputs[20]);
    assign layer0_outputs[100] = (inputs[104]) & ~(inputs[224]);
    assign layer0_outputs[101] = ~((inputs[180]) | (inputs[60]));
    assign layer0_outputs[102] = ~((inputs[247]) ^ (inputs[218]));
    assign layer0_outputs[103] = inputs[69];
    assign layer0_outputs[104] = ~(inputs[95]);
    assign layer0_outputs[105] = ~((inputs[62]) ^ (inputs[16]));
    assign layer0_outputs[106] = ~(inputs[104]) | (inputs[137]);
    assign layer0_outputs[107] = (inputs[153]) & ~(inputs[11]);
    assign layer0_outputs[108] = (inputs[101]) | (inputs[86]);
    assign layer0_outputs[109] = ~((inputs[227]) & (inputs[248]));
    assign layer0_outputs[110] = (inputs[163]) ^ (inputs[191]);
    assign layer0_outputs[111] = inputs[228];
    assign layer0_outputs[112] = ~((inputs[199]) | (inputs[15]));
    assign layer0_outputs[113] = 1'b1;
    assign layer0_outputs[114] = (inputs[159]) | (inputs[107]);
    assign layer0_outputs[115] = ~((inputs[102]) ^ (inputs[167]));
    assign layer0_outputs[116] = ~((inputs[170]) | (inputs[236]));
    assign layer0_outputs[117] = (inputs[4]) & ~(inputs[21]);
    assign layer0_outputs[118] = (inputs[168]) ^ (inputs[239]);
    assign layer0_outputs[119] = ~(inputs[106]);
    assign layer0_outputs[120] = ~(inputs[102]);
    assign layer0_outputs[121] = (inputs[234]) & ~(inputs[141]);
    assign layer0_outputs[122] = (inputs[28]) & (inputs[65]);
    assign layer0_outputs[123] = (inputs[161]) ^ (inputs[6]);
    assign layer0_outputs[124] = ~(inputs[121]) | (inputs[69]);
    assign layer0_outputs[125] = inputs[151];
    assign layer0_outputs[126] = (inputs[222]) | (inputs[58]);
    assign layer0_outputs[127] = ~(inputs[88]) | (inputs[82]);
    assign layer0_outputs[128] = (inputs[122]) | (inputs[0]);
    assign layer0_outputs[129] = ~((inputs[253]) ^ (inputs[123]));
    assign layer0_outputs[130] = inputs[77];
    assign layer0_outputs[131] = ~((inputs[147]) | (inputs[164]));
    assign layer0_outputs[132] = ~(inputs[200]);
    assign layer0_outputs[133] = ~(inputs[198]);
    assign layer0_outputs[134] = ~((inputs[188]) | (inputs[59]));
    assign layer0_outputs[135] = ~((inputs[247]) ^ (inputs[181]));
    assign layer0_outputs[136] = inputs[25];
    assign layer0_outputs[137] = 1'b1;
    assign layer0_outputs[138] = (inputs[102]) & ~(inputs[28]);
    assign layer0_outputs[139] = ~(inputs[102]) | (inputs[161]);
    assign layer0_outputs[140] = ~(inputs[202]) | (inputs[29]);
    assign layer0_outputs[141] = ~(inputs[173]);
    assign layer0_outputs[142] = ~(inputs[131]) | (inputs[24]);
    assign layer0_outputs[143] = 1'b1;
    assign layer0_outputs[144] = (inputs[33]) & ~(inputs[218]);
    assign layer0_outputs[145] = (inputs[14]) | (inputs[139]);
    assign layer0_outputs[146] = (inputs[196]) & ~(inputs[114]);
    assign layer0_outputs[147] = (inputs[57]) | (inputs[77]);
    assign layer0_outputs[148] = inputs[122];
    assign layer0_outputs[149] = inputs[183];
    assign layer0_outputs[150] = ~((inputs[39]) ^ (inputs[81]));
    assign layer0_outputs[151] = (inputs[53]) & ~(inputs[38]);
    assign layer0_outputs[152] = ~(inputs[193]);
    assign layer0_outputs[153] = ~(inputs[85]);
    assign layer0_outputs[154] = (inputs[71]) | (inputs[95]);
    assign layer0_outputs[155] = ~(inputs[87]) | (inputs[205]);
    assign layer0_outputs[156] = ~(inputs[190]) | (inputs[30]);
    assign layer0_outputs[157] = inputs[56];
    assign layer0_outputs[158] = (inputs[48]) ^ (inputs[210]);
    assign layer0_outputs[159] = ~(inputs[21]) | (inputs[82]);
    assign layer0_outputs[160] = (inputs[199]) & ~(inputs[177]);
    assign layer0_outputs[161] = (inputs[10]) & ~(inputs[128]);
    assign layer0_outputs[162] = ~(inputs[151]) | (inputs[248]);
    assign layer0_outputs[163] = ~((inputs[93]) | (inputs[197]));
    assign layer0_outputs[164] = (inputs[225]) ^ (inputs[166]);
    assign layer0_outputs[165] = (inputs[29]) & ~(inputs[4]);
    assign layer0_outputs[166] = ~(inputs[181]) | (inputs[29]);
    assign layer0_outputs[167] = ~((inputs[205]) ^ (inputs[231]));
    assign layer0_outputs[168] = ~((inputs[251]) | (inputs[101]));
    assign layer0_outputs[169] = ~(inputs[181]);
    assign layer0_outputs[170] = (inputs[96]) ^ (inputs[58]);
    assign layer0_outputs[171] = ~((inputs[37]) | (inputs[158]));
    assign layer0_outputs[172] = ~(inputs[215]);
    assign layer0_outputs[173] = (inputs[153]) & ~(inputs[116]);
    assign layer0_outputs[174] = (inputs[41]) ^ (inputs[254]);
    assign layer0_outputs[175] = (inputs[118]) & ~(inputs[240]);
    assign layer0_outputs[176] = ~((inputs[218]) | (inputs[204]));
    assign layer0_outputs[177] = (inputs[237]) & (inputs[241]);
    assign layer0_outputs[178] = (inputs[33]) ^ (inputs[251]);
    assign layer0_outputs[179] = inputs[66];
    assign layer0_outputs[180] = ~((inputs[251]) | (inputs[242]));
    assign layer0_outputs[181] = inputs[10];
    assign layer0_outputs[182] = (inputs[181]) & ~(inputs[78]);
    assign layer0_outputs[183] = inputs[121];
    assign layer0_outputs[184] = (inputs[52]) | (inputs[8]);
    assign layer0_outputs[185] = (inputs[104]) & ~(inputs[186]);
    assign layer0_outputs[186] = (inputs[2]) & ~(inputs[124]);
    assign layer0_outputs[187] = ~(inputs[108]);
    assign layer0_outputs[188] = (inputs[126]) & ~(inputs[19]);
    assign layer0_outputs[189] = (inputs[16]) ^ (inputs[229]);
    assign layer0_outputs[190] = inputs[179];
    assign layer0_outputs[191] = ~(inputs[118]) | (inputs[18]);
    assign layer0_outputs[192] = ~((inputs[156]) ^ (inputs[127]));
    assign layer0_outputs[193] = ~(inputs[220]);
    assign layer0_outputs[194] = (inputs[240]) | (inputs[159]);
    assign layer0_outputs[195] = (inputs[62]) | (inputs[78]);
    assign layer0_outputs[196] = ~(inputs[136]);
    assign layer0_outputs[197] = ~(inputs[64]) | (inputs[11]);
    assign layer0_outputs[198] = (inputs[255]) & (inputs[32]);
    assign layer0_outputs[199] = (inputs[43]) ^ (inputs[34]);
    assign layer0_outputs[200] = ~(inputs[183]);
    assign layer0_outputs[201] = (inputs[213]) & ~(inputs[13]);
    assign layer0_outputs[202] = ~(inputs[214]) | (inputs[211]);
    assign layer0_outputs[203] = ~(inputs[66]);
    assign layer0_outputs[204] = ~(inputs[220]) | (inputs[226]);
    assign layer0_outputs[205] = ~(inputs[151]);
    assign layer0_outputs[206] = ~(inputs[132]) | (inputs[79]);
    assign layer0_outputs[207] = (inputs[203]) & ~(inputs[10]);
    assign layer0_outputs[208] = (inputs[101]) | (inputs[225]);
    assign layer0_outputs[209] = inputs[198];
    assign layer0_outputs[210] = ~((inputs[102]) | (inputs[141]));
    assign layer0_outputs[211] = (inputs[27]) | (inputs[200]);
    assign layer0_outputs[212] = ~(inputs[37]) | (inputs[125]);
    assign layer0_outputs[213] = ~((inputs[194]) | (inputs[170]));
    assign layer0_outputs[214] = ~(inputs[237]);
    assign layer0_outputs[215] = inputs[165];
    assign layer0_outputs[216] = ~((inputs[165]) | (inputs[97]));
    assign layer0_outputs[217] = inputs[119];
    assign layer0_outputs[218] = inputs[230];
    assign layer0_outputs[219] = inputs[56];
    assign layer0_outputs[220] = ~(inputs[66]);
    assign layer0_outputs[221] = ~((inputs[151]) | (inputs[228]));
    assign layer0_outputs[222] = (inputs[61]) | (inputs[139]);
    assign layer0_outputs[223] = ~((inputs[174]) | (inputs[247]));
    assign layer0_outputs[224] = ~(inputs[88]) | (inputs[16]);
    assign layer0_outputs[225] = inputs[246];
    assign layer0_outputs[226] = inputs[118];
    assign layer0_outputs[227] = ~(inputs[180]) | (inputs[127]);
    assign layer0_outputs[228] = (inputs[166]) & ~(inputs[94]);
    assign layer0_outputs[229] = (inputs[41]) ^ (inputs[73]);
    assign layer0_outputs[230] = ~((inputs[82]) | (inputs[150]));
    assign layer0_outputs[231] = ~(inputs[82]);
    assign layer0_outputs[232] = ~(inputs[197]);
    assign layer0_outputs[233] = ~(inputs[27]);
    assign layer0_outputs[234] = 1'b1;
    assign layer0_outputs[235] = (inputs[14]) ^ (inputs[135]);
    assign layer0_outputs[236] = ~((inputs[220]) ^ (inputs[31]));
    assign layer0_outputs[237] = inputs[153];
    assign layer0_outputs[238] = ~(inputs[184]) | (inputs[231]);
    assign layer0_outputs[239] = (inputs[64]) | (inputs[153]);
    assign layer0_outputs[240] = ~(inputs[166]) | (inputs[249]);
    assign layer0_outputs[241] = ~(inputs[99]) | (inputs[66]);
    assign layer0_outputs[242] = ~(inputs[99]) | (inputs[253]);
    assign layer0_outputs[243] = (inputs[244]) | (inputs[225]);
    assign layer0_outputs[244] = inputs[218];
    assign layer0_outputs[245] = ~(inputs[7]) | (inputs[238]);
    assign layer0_outputs[246] = ~(inputs[150]) | (inputs[66]);
    assign layer0_outputs[247] = ~((inputs[218]) | (inputs[190]));
    assign layer0_outputs[248] = inputs[38];
    assign layer0_outputs[249] = ~(inputs[204]);
    assign layer0_outputs[250] = (inputs[187]) & ~(inputs[114]);
    assign layer0_outputs[251] = ~(inputs[173]);
    assign layer0_outputs[252] = (inputs[57]) | (inputs[147]);
    assign layer0_outputs[253] = ~(inputs[203]) | (inputs[19]);
    assign layer0_outputs[254] = ~(inputs[70]);
    assign layer0_outputs[255] = ~((inputs[51]) | (inputs[220]));
    assign layer0_outputs[256] = ~(inputs[157]);
    assign layer0_outputs[257] = ~(inputs[232]) | (inputs[69]);
    assign layer0_outputs[258] = ~((inputs[139]) | (inputs[39]));
    assign layer0_outputs[259] = ~(inputs[88]);
    assign layer0_outputs[260] = inputs[131];
    assign layer0_outputs[261] = ~((inputs[118]) ^ (inputs[174]));
    assign layer0_outputs[262] = ~(inputs[126]);
    assign layer0_outputs[263] = inputs[12];
    assign layer0_outputs[264] = ~((inputs[93]) | (inputs[222]));
    assign layer0_outputs[265] = ~((inputs[214]) & (inputs[234]));
    assign layer0_outputs[266] = ~((inputs[42]) | (inputs[38]));
    assign layer0_outputs[267] = ~(inputs[207]);
    assign layer0_outputs[268] = (inputs[28]) & (inputs[5]);
    assign layer0_outputs[269] = (inputs[196]) ^ (inputs[26]);
    assign layer0_outputs[270] = ~(inputs[150]);
    assign layer0_outputs[271] = (inputs[210]) ^ (inputs[178]);
    assign layer0_outputs[272] = ~(inputs[28]);
    assign layer0_outputs[273] = ~(inputs[163]);
    assign layer0_outputs[274] = ~(inputs[126]);
    assign layer0_outputs[275] = (inputs[89]) & ~(inputs[233]);
    assign layer0_outputs[276] = (inputs[94]) | (inputs[96]);
    assign layer0_outputs[277] = ~((inputs[27]) | (inputs[103]));
    assign layer0_outputs[278] = inputs[1];
    assign layer0_outputs[279] = (inputs[34]) | (inputs[68]);
    assign layer0_outputs[280] = ~((inputs[117]) | (inputs[45]));
    assign layer0_outputs[281] = ~(inputs[194]) | (inputs[205]);
    assign layer0_outputs[282] = ~(inputs[175]);
    assign layer0_outputs[283] = ~(inputs[165]);
    assign layer0_outputs[284] = ~((inputs[157]) | (inputs[169]));
    assign layer0_outputs[285] = ~(inputs[68]) | (inputs[158]);
    assign layer0_outputs[286] = ~((inputs[92]) | (inputs[235]));
    assign layer0_outputs[287] = ~((inputs[100]) ^ (inputs[57]));
    assign layer0_outputs[288] = inputs[121];
    assign layer0_outputs[289] = inputs[150];
    assign layer0_outputs[290] = 1'b1;
    assign layer0_outputs[291] = ~((inputs[240]) ^ (inputs[174]));
    assign layer0_outputs[292] = ~(inputs[137]) | (inputs[95]);
    assign layer0_outputs[293] = (inputs[221]) | (inputs[147]);
    assign layer0_outputs[294] = ~(inputs[199]) | (inputs[137]);
    assign layer0_outputs[295] = (inputs[197]) | (inputs[198]);
    assign layer0_outputs[296] = ~(inputs[38]);
    assign layer0_outputs[297] = inputs[151];
    assign layer0_outputs[298] = ~(inputs[172]) | (inputs[98]);
    assign layer0_outputs[299] = ~(inputs[93]);
    assign layer0_outputs[300] = ~((inputs[61]) | (inputs[115]));
    assign layer0_outputs[301] = (inputs[75]) & ~(inputs[80]);
    assign layer0_outputs[302] = ~((inputs[207]) | (inputs[92]));
    assign layer0_outputs[303] = (inputs[16]) ^ (inputs[157]);
    assign layer0_outputs[304] = ~(inputs[229]) | (inputs[220]);
    assign layer0_outputs[305] = ~(inputs[166]);
    assign layer0_outputs[306] = (inputs[170]) & (inputs[88]);
    assign layer0_outputs[307] = inputs[130];
    assign layer0_outputs[308] = (inputs[211]) | (inputs[214]);
    assign layer0_outputs[309] = ~((inputs[148]) | (inputs[134]));
    assign layer0_outputs[310] = ~((inputs[132]) | (inputs[76]));
    assign layer0_outputs[311] = inputs[124];
    assign layer0_outputs[312] = (inputs[233]) | (inputs[97]);
    assign layer0_outputs[313] = ~((inputs[177]) | (inputs[73]));
    assign layer0_outputs[314] = (inputs[133]) & ~(inputs[239]);
    assign layer0_outputs[315] = inputs[91];
    assign layer0_outputs[316] = (inputs[201]) ^ (inputs[252]);
    assign layer0_outputs[317] = ~((inputs[6]) | (inputs[84]));
    assign layer0_outputs[318] = ~((inputs[171]) ^ (inputs[10]));
    assign layer0_outputs[319] = (inputs[246]) | (inputs[107]);
    assign layer0_outputs[320] = (inputs[160]) & ~(inputs[105]);
    assign layer0_outputs[321] = inputs[152];
    assign layer0_outputs[322] = ~((inputs[234]) | (inputs[70]));
    assign layer0_outputs[323] = ~(inputs[90]) | (inputs[45]);
    assign layer0_outputs[324] = ~((inputs[223]) | (inputs[56]));
    assign layer0_outputs[325] = ~((inputs[150]) | (inputs[39]));
    assign layer0_outputs[326] = ~(inputs[216]);
    assign layer0_outputs[327] = 1'b1;
    assign layer0_outputs[328] = (inputs[153]) | (inputs[68]);
    assign layer0_outputs[329] = (inputs[180]) ^ (inputs[9]);
    assign layer0_outputs[330] = (inputs[138]) & ~(inputs[45]);
    assign layer0_outputs[331] = inputs[58];
    assign layer0_outputs[332] = ~(inputs[232]);
    assign layer0_outputs[333] = inputs[180];
    assign layer0_outputs[334] = (inputs[179]) | (inputs[203]);
    assign layer0_outputs[335] = (inputs[245]) & ~(inputs[129]);
    assign layer0_outputs[336] = (inputs[180]) & ~(inputs[214]);
    assign layer0_outputs[337] = 1'b0;
    assign layer0_outputs[338] = ~(inputs[136]) | (inputs[31]);
    assign layer0_outputs[339] = (inputs[211]) & ~(inputs[49]);
    assign layer0_outputs[340] = (inputs[153]) | (inputs[203]);
    assign layer0_outputs[341] = ~(inputs[142]);
    assign layer0_outputs[342] = ~(inputs[236]);
    assign layer0_outputs[343] = (inputs[7]) | (inputs[207]);
    assign layer0_outputs[344] = ~(inputs[150]) | (inputs[222]);
    assign layer0_outputs[345] = (inputs[32]) & (inputs[169]);
    assign layer0_outputs[346] = (inputs[34]) ^ (inputs[191]);
    assign layer0_outputs[347] = inputs[252];
    assign layer0_outputs[348] = (inputs[235]) & ~(inputs[227]);
    assign layer0_outputs[349] = (inputs[97]) | (inputs[107]);
    assign layer0_outputs[350] = (inputs[116]) & ~(inputs[234]);
    assign layer0_outputs[351] = ~(inputs[139]) | (inputs[76]);
    assign layer0_outputs[352] = ~((inputs[94]) | (inputs[199]));
    assign layer0_outputs[353] = (inputs[155]) & ~(inputs[22]);
    assign layer0_outputs[354] = ~((inputs[208]) | (inputs[170]));
    assign layer0_outputs[355] = ~((inputs[24]) | (inputs[190]));
    assign layer0_outputs[356] = (inputs[72]) & (inputs[212]);
    assign layer0_outputs[357] = ~((inputs[143]) & (inputs[54]));
    assign layer0_outputs[358] = ~((inputs[64]) ^ (inputs[106]));
    assign layer0_outputs[359] = (inputs[13]) | (inputs[75]);
    assign layer0_outputs[360] = ~(inputs[102]);
    assign layer0_outputs[361] = ~((inputs[236]) | (inputs[218]));
    assign layer0_outputs[362] = ~(inputs[178]);
    assign layer0_outputs[363] = (inputs[221]) & ~(inputs[226]);
    assign layer0_outputs[364] = (inputs[102]) & ~(inputs[244]);
    assign layer0_outputs[365] = ~(inputs[141]) | (inputs[205]);
    assign layer0_outputs[366] = ~(inputs[162]);
    assign layer0_outputs[367] = inputs[135];
    assign layer0_outputs[368] = ~((inputs[138]) | (inputs[250]));
    assign layer0_outputs[369] = ~(inputs[135]);
    assign layer0_outputs[370] = ~((inputs[61]) & (inputs[171]));
    assign layer0_outputs[371] = ~((inputs[7]) ^ (inputs[233]));
    assign layer0_outputs[372] = ~(inputs[3]) | (inputs[241]);
    assign layer0_outputs[373] = ~((inputs[202]) | (inputs[218]));
    assign layer0_outputs[374] = ~((inputs[147]) ^ (inputs[252]));
    assign layer0_outputs[375] = ~(inputs[84]) | (inputs[221]);
    assign layer0_outputs[376] = ~(inputs[90]) | (inputs[204]);
    assign layer0_outputs[377] = 1'b0;
    assign layer0_outputs[378] = inputs[102];
    assign layer0_outputs[379] = ~((inputs[114]) ^ (inputs[147]));
    assign layer0_outputs[380] = ~(inputs[167]);
    assign layer0_outputs[381] = (inputs[77]) | (inputs[63]);
    assign layer0_outputs[382] = ~((inputs[58]) ^ (inputs[141]));
    assign layer0_outputs[383] = (inputs[54]) ^ (inputs[236]);
    assign layer0_outputs[384] = ~(inputs[118]);
    assign layer0_outputs[385] = ~((inputs[228]) | (inputs[223]));
    assign layer0_outputs[386] = (inputs[0]) ^ (inputs[219]);
    assign layer0_outputs[387] = (inputs[65]) & ~(inputs[37]);
    assign layer0_outputs[388] = ~((inputs[93]) | (inputs[253]));
    assign layer0_outputs[389] = (inputs[155]) & ~(inputs[114]);
    assign layer0_outputs[390] = ~((inputs[152]) & (inputs[152]));
    assign layer0_outputs[391] = ~(inputs[101]) | (inputs[64]);
    assign layer0_outputs[392] = (inputs[27]) ^ (inputs[20]);
    assign layer0_outputs[393] = inputs[130];
    assign layer0_outputs[394] = (inputs[211]) | (inputs[51]);
    assign layer0_outputs[395] = ~(inputs[164]);
    assign layer0_outputs[396] = ~(inputs[91]) | (inputs[128]);
    assign layer0_outputs[397] = (inputs[246]) | (inputs[251]);
    assign layer0_outputs[398] = (inputs[160]) & ~(inputs[62]);
    assign layer0_outputs[399] = (inputs[23]) | (inputs[170]);
    assign layer0_outputs[400] = (inputs[185]) & ~(inputs[234]);
    assign layer0_outputs[401] = ~(inputs[152]);
    assign layer0_outputs[402] = (inputs[237]) & (inputs[8]);
    assign layer0_outputs[403] = ~(inputs[235]) | (inputs[213]);
    assign layer0_outputs[404] = inputs[228];
    assign layer0_outputs[405] = (inputs[168]) & ~(inputs[92]);
    assign layer0_outputs[406] = ~(inputs[253]) | (inputs[209]);
    assign layer0_outputs[407] = (inputs[20]) & ~(inputs[165]);
    assign layer0_outputs[408] = (inputs[127]) ^ (inputs[55]);
    assign layer0_outputs[409] = (inputs[168]) & ~(inputs[13]);
    assign layer0_outputs[410] = ~(inputs[200]) | (inputs[53]);
    assign layer0_outputs[411] = (inputs[52]) ^ (inputs[193]);
    assign layer0_outputs[412] = inputs[182];
    assign layer0_outputs[413] = (inputs[123]) & ~(inputs[94]);
    assign layer0_outputs[414] = ~(inputs[51]) | (inputs[133]);
    assign layer0_outputs[415] = inputs[120];
    assign layer0_outputs[416] = ~((inputs[81]) | (inputs[136]));
    assign layer0_outputs[417] = ~((inputs[2]) | (inputs[172]));
    assign layer0_outputs[418] = inputs[92];
    assign layer0_outputs[419] = (inputs[147]) & ~(inputs[189]);
    assign layer0_outputs[420] = inputs[89];
    assign layer0_outputs[421] = (inputs[119]) & ~(inputs[221]);
    assign layer0_outputs[422] = inputs[249];
    assign layer0_outputs[423] = (inputs[157]) | (inputs[23]);
    assign layer0_outputs[424] = ~((inputs[81]) ^ (inputs[46]));
    assign layer0_outputs[425] = ~((inputs[62]) | (inputs[109]));
    assign layer0_outputs[426] = (inputs[94]) ^ (inputs[113]);
    assign layer0_outputs[427] = ~((inputs[124]) | (inputs[26]));
    assign layer0_outputs[428] = inputs[165];
    assign layer0_outputs[429] = ~((inputs[4]) | (inputs[37]));
    assign layer0_outputs[430] = (inputs[200]) & (inputs[171]);
    assign layer0_outputs[431] = (inputs[142]) ^ (inputs[201]);
    assign layer0_outputs[432] = (inputs[94]) | (inputs[181]);
    assign layer0_outputs[433] = (inputs[22]) | (inputs[162]);
    assign layer0_outputs[434] = (inputs[227]) & ~(inputs[115]);
    assign layer0_outputs[435] = ~(inputs[41]) | (inputs[4]);
    assign layer0_outputs[436] = ~((inputs[194]) ^ (inputs[205]));
    assign layer0_outputs[437] = (inputs[136]) & ~(inputs[213]);
    assign layer0_outputs[438] = (inputs[76]) & ~(inputs[202]);
    assign layer0_outputs[439] = ~((inputs[201]) ^ (inputs[11]));
    assign layer0_outputs[440] = ~(inputs[56]);
    assign layer0_outputs[441] = (inputs[191]) | (inputs[82]);
    assign layer0_outputs[442] = inputs[60];
    assign layer0_outputs[443] = (inputs[200]) ^ (inputs[63]);
    assign layer0_outputs[444] = (inputs[123]) & (inputs[252]);
    assign layer0_outputs[445] = ~(inputs[87]);
    assign layer0_outputs[446] = (inputs[55]) ^ (inputs[7]);
    assign layer0_outputs[447] = (inputs[101]) ^ (inputs[131]);
    assign layer0_outputs[448] = ~((inputs[27]) | (inputs[43]));
    assign layer0_outputs[449] = ~((inputs[104]) | (inputs[63]));
    assign layer0_outputs[450] = ~(inputs[54]) | (inputs[249]);
    assign layer0_outputs[451] = (inputs[107]) & ~(inputs[61]);
    assign layer0_outputs[452] = (inputs[173]) | (inputs[78]);
    assign layer0_outputs[453] = ~((inputs[199]) | (inputs[131]));
    assign layer0_outputs[454] = (inputs[137]) ^ (inputs[170]);
    assign layer0_outputs[455] = (inputs[178]) & ~(inputs[112]);
    assign layer0_outputs[456] = ~((inputs[96]) ^ (inputs[200]));
    assign layer0_outputs[457] = ~(inputs[137]) | (inputs[250]);
    assign layer0_outputs[458] = (inputs[72]) & ~(inputs[167]);
    assign layer0_outputs[459] = ~((inputs[44]) | (inputs[127]));
    assign layer0_outputs[460] = ~((inputs[164]) | (inputs[50]));
    assign layer0_outputs[461] = ~((inputs[218]) | (inputs[188]));
    assign layer0_outputs[462] = (inputs[127]) & ~(inputs[238]);
    assign layer0_outputs[463] = (inputs[125]) | (inputs[109]);
    assign layer0_outputs[464] = (inputs[33]) & (inputs[145]);
    assign layer0_outputs[465] = (inputs[24]) & (inputs[129]);
    assign layer0_outputs[466] = inputs[251];
    assign layer0_outputs[467] = ~(inputs[102]) | (inputs[53]);
    assign layer0_outputs[468] = (inputs[228]) | (inputs[149]);
    assign layer0_outputs[469] = (inputs[224]) ^ (inputs[212]);
    assign layer0_outputs[470] = ~(inputs[57]) | (inputs[172]);
    assign layer0_outputs[471] = 1'b1;
    assign layer0_outputs[472] = inputs[215];
    assign layer0_outputs[473] = ~(inputs[91]);
    assign layer0_outputs[474] = (inputs[240]) & (inputs[193]);
    assign layer0_outputs[475] = (inputs[98]) ^ (inputs[117]);
    assign layer0_outputs[476] = (inputs[92]) ^ (inputs[90]);
    assign layer0_outputs[477] = (inputs[200]) | (inputs[163]);
    assign layer0_outputs[478] = 1'b0;
    assign layer0_outputs[479] = ~(inputs[122]);
    assign layer0_outputs[480] = ~((inputs[18]) | (inputs[144]));
    assign layer0_outputs[481] = ~((inputs[33]) | (inputs[120]));
    assign layer0_outputs[482] = (inputs[251]) & (inputs[79]);
    assign layer0_outputs[483] = ~(inputs[215]) | (inputs[61]);
    assign layer0_outputs[484] = (inputs[250]) & (inputs[168]);
    assign layer0_outputs[485] = ~(inputs[97]);
    assign layer0_outputs[486] = (inputs[214]) & ~(inputs[147]);
    assign layer0_outputs[487] = ~((inputs[23]) | (inputs[109]));
    assign layer0_outputs[488] = ~((inputs[89]) | (inputs[189]));
    assign layer0_outputs[489] = (inputs[123]) & ~(inputs[82]);
    assign layer0_outputs[490] = (inputs[183]) & ~(inputs[114]);
    assign layer0_outputs[491] = ~(inputs[155]) | (inputs[13]);
    assign layer0_outputs[492] = ~(inputs[39]) | (inputs[13]);
    assign layer0_outputs[493] = ~(inputs[40]) | (inputs[48]);
    assign layer0_outputs[494] = inputs[59];
    assign layer0_outputs[495] = ~((inputs[249]) | (inputs[233]));
    assign layer0_outputs[496] = ~(inputs[155]) | (inputs[49]);
    assign layer0_outputs[497] = inputs[80];
    assign layer0_outputs[498] = (inputs[187]) & ~(inputs[95]);
    assign layer0_outputs[499] = (inputs[235]) ^ (inputs[230]);
    assign layer0_outputs[500] = (inputs[32]) | (inputs[23]);
    assign layer0_outputs[501] = ~(inputs[120]) | (inputs[12]);
    assign layer0_outputs[502] = inputs[122];
    assign layer0_outputs[503] = inputs[221];
    assign layer0_outputs[504] = inputs[189];
    assign layer0_outputs[505] = (inputs[156]) & ~(inputs[98]);
    assign layer0_outputs[506] = (inputs[160]) ^ (inputs[248]);
    assign layer0_outputs[507] = inputs[120];
    assign layer0_outputs[508] = (inputs[99]) & ~(inputs[59]);
    assign layer0_outputs[509] = ~(inputs[76]);
    assign layer0_outputs[510] = ~(inputs[39]) | (inputs[228]);
    assign layer0_outputs[511] = (inputs[128]) | (inputs[114]);
    assign layer0_outputs[512] = ~((inputs[159]) ^ (inputs[217]));
    assign layer0_outputs[513] = ~(inputs[106]) | (inputs[13]);
    assign layer0_outputs[514] = ~((inputs[176]) & (inputs[17]));
    assign layer0_outputs[515] = ~((inputs[205]) | (inputs[189]));
    assign layer0_outputs[516] = ~(inputs[231]);
    assign layer0_outputs[517] = ~((inputs[230]) & (inputs[1]));
    assign layer0_outputs[518] = ~((inputs[49]) ^ (inputs[105]));
    assign layer0_outputs[519] = inputs[153];
    assign layer0_outputs[520] = inputs[92];
    assign layer0_outputs[521] = (inputs[196]) & ~(inputs[246]);
    assign layer0_outputs[522] = 1'b1;
    assign layer0_outputs[523] = inputs[107];
    assign layer0_outputs[524] = (inputs[102]) & ~(inputs[254]);
    assign layer0_outputs[525] = (inputs[71]) | (inputs[242]);
    assign layer0_outputs[526] = (inputs[130]) ^ (inputs[195]);
    assign layer0_outputs[527] = ~((inputs[79]) ^ (inputs[120]));
    assign layer0_outputs[528] = ~(inputs[27]) | (inputs[18]);
    assign layer0_outputs[529] = ~(inputs[105]);
    assign layer0_outputs[530] = (inputs[148]) ^ (inputs[224]);
    assign layer0_outputs[531] = ~((inputs[153]) | (inputs[34]));
    assign layer0_outputs[532] = ~((inputs[46]) & (inputs[163]));
    assign layer0_outputs[533] = (inputs[238]) & (inputs[216]);
    assign layer0_outputs[534] = ~(inputs[130]) | (inputs[74]);
    assign layer0_outputs[535] = (inputs[14]) & (inputs[33]);
    assign layer0_outputs[536] = (inputs[115]) | (inputs[138]);
    assign layer0_outputs[537] = ~(inputs[154]);
    assign layer0_outputs[538] = ~((inputs[151]) | (inputs[233]));
    assign layer0_outputs[539] = ~((inputs[165]) | (inputs[37]));
    assign layer0_outputs[540] = ~(inputs[107]);
    assign layer0_outputs[541] = inputs[40];
    assign layer0_outputs[542] = inputs[240];
    assign layer0_outputs[543] = (inputs[48]) | (inputs[157]);
    assign layer0_outputs[544] = ~((inputs[3]) | (inputs[148]));
    assign layer0_outputs[545] = inputs[173];
    assign layer0_outputs[546] = inputs[56];
    assign layer0_outputs[547] = (inputs[29]) ^ (inputs[67]);
    assign layer0_outputs[548] = ~((inputs[249]) | (inputs[135]));
    assign layer0_outputs[549] = (inputs[114]) ^ (inputs[67]);
    assign layer0_outputs[550] = ~(inputs[112]);
    assign layer0_outputs[551] = ~(inputs[70]);
    assign layer0_outputs[552] = (inputs[3]) | (inputs[122]);
    assign layer0_outputs[553] = (inputs[194]) ^ (inputs[230]);
    assign layer0_outputs[554] = (inputs[149]) & ~(inputs[211]);
    assign layer0_outputs[555] = (inputs[235]) & ~(inputs[17]);
    assign layer0_outputs[556] = inputs[124];
    assign layer0_outputs[557] = (inputs[163]) & ~(inputs[247]);
    assign layer0_outputs[558] = (inputs[156]) | (inputs[232]);
    assign layer0_outputs[559] = ~(inputs[165]);
    assign layer0_outputs[560] = (inputs[234]) ^ (inputs[116]);
    assign layer0_outputs[561] = (inputs[231]) & ~(inputs[196]);
    assign layer0_outputs[562] = ~((inputs[74]) ^ (inputs[11]));
    assign layer0_outputs[563] = (inputs[32]) | (inputs[16]);
    assign layer0_outputs[564] = (inputs[214]) | (inputs[222]);
    assign layer0_outputs[565] = ~((inputs[139]) ^ (inputs[134]));
    assign layer0_outputs[566] = (inputs[175]) ^ (inputs[226]);
    assign layer0_outputs[567] = ~(inputs[39]);
    assign layer0_outputs[568] = ~((inputs[109]) ^ (inputs[87]));
    assign layer0_outputs[569] = (inputs[190]) | (inputs[75]);
    assign layer0_outputs[570] = (inputs[220]) | (inputs[201]);
    assign layer0_outputs[571] = (inputs[69]) | (inputs[172]);
    assign layer0_outputs[572] = ~(inputs[250]) | (inputs[154]);
    assign layer0_outputs[573] = ~((inputs[72]) | (inputs[2]));
    assign layer0_outputs[574] = ~((inputs[88]) | (inputs[13]));
    assign layer0_outputs[575] = ~((inputs[133]) | (inputs[220]));
    assign layer0_outputs[576] = ~(inputs[77]) | (inputs[246]);
    assign layer0_outputs[577] = ~(inputs[121]) | (inputs[13]);
    assign layer0_outputs[578] = (inputs[29]) | (inputs[152]);
    assign layer0_outputs[579] = ~(inputs[130]) | (inputs[145]);
    assign layer0_outputs[580] = (inputs[72]) & ~(inputs[11]);
    assign layer0_outputs[581] = (inputs[102]) & ~(inputs[32]);
    assign layer0_outputs[582] = ~((inputs[91]) | (inputs[237]));
    assign layer0_outputs[583] = ~(inputs[125]) | (inputs[20]);
    assign layer0_outputs[584] = (inputs[119]) | (inputs[250]);
    assign layer0_outputs[585] = ~((inputs[143]) & (inputs[30]));
    assign layer0_outputs[586] = ~(inputs[76]);
    assign layer0_outputs[587] = (inputs[54]) ^ (inputs[30]);
    assign layer0_outputs[588] = (inputs[89]) | (inputs[111]);
    assign layer0_outputs[589] = (inputs[246]) ^ (inputs[1]);
    assign layer0_outputs[590] = 1'b0;
    assign layer0_outputs[591] = ~((inputs[77]) ^ (inputs[44]));
    assign layer0_outputs[592] = ~(inputs[185]) | (inputs[117]);
    assign layer0_outputs[593] = ~(inputs[50]);
    assign layer0_outputs[594] = ~(inputs[216]) | (inputs[146]);
    assign layer0_outputs[595] = (inputs[173]) ^ (inputs[140]);
    assign layer0_outputs[596] = (inputs[135]) | (inputs[79]);
    assign layer0_outputs[597] = ~(inputs[204]);
    assign layer0_outputs[598] = (inputs[30]) | (inputs[147]);
    assign layer0_outputs[599] = (inputs[5]) | (inputs[178]);
    assign layer0_outputs[600] = (inputs[26]) & ~(inputs[7]);
    assign layer0_outputs[601] = ~((inputs[132]) ^ (inputs[241]));
    assign layer0_outputs[602] = (inputs[19]) & (inputs[50]);
    assign layer0_outputs[603] = ~((inputs[70]) | (inputs[147]));
    assign layer0_outputs[604] = 1'b1;
    assign layer0_outputs[605] = ~(inputs[101]);
    assign layer0_outputs[606] = ~(inputs[167]) | (inputs[10]);
    assign layer0_outputs[607] = (inputs[251]) | (inputs[21]);
    assign layer0_outputs[608] = ~(inputs[115]);
    assign layer0_outputs[609] = (inputs[106]) | (inputs[6]);
    assign layer0_outputs[610] = (inputs[112]) | (inputs[54]);
    assign layer0_outputs[611] = ~(inputs[170]);
    assign layer0_outputs[612] = (inputs[205]) | (inputs[101]);
    assign layer0_outputs[613] = (inputs[192]) | (inputs[207]);
    assign layer0_outputs[614] = ~(inputs[134]) | (inputs[245]);
    assign layer0_outputs[615] = inputs[94];
    assign layer0_outputs[616] = (inputs[53]) ^ (inputs[112]);
    assign layer0_outputs[617] = ~((inputs[190]) | (inputs[178]));
    assign layer0_outputs[618] = ~(inputs[105]);
    assign layer0_outputs[619] = ~((inputs[202]) & (inputs[113]));
    assign layer0_outputs[620] = inputs[101];
    assign layer0_outputs[621] = (inputs[38]) | (inputs[183]);
    assign layer0_outputs[622] = ~(inputs[119]) | (inputs[149]);
    assign layer0_outputs[623] = (inputs[184]) | (inputs[211]);
    assign layer0_outputs[624] = (inputs[223]) | (inputs[165]);
    assign layer0_outputs[625] = 1'b0;
    assign layer0_outputs[626] = (inputs[19]) & ~(inputs[163]);
    assign layer0_outputs[627] = (inputs[98]) | (inputs[233]);
    assign layer0_outputs[628] = (inputs[222]) | (inputs[126]);
    assign layer0_outputs[629] = (inputs[155]) & ~(inputs[235]);
    assign layer0_outputs[630] = inputs[51];
    assign layer0_outputs[631] = ~(inputs[104]);
    assign layer0_outputs[632] = (inputs[231]) ^ (inputs[227]);
    assign layer0_outputs[633] = (inputs[21]) | (inputs[187]);
    assign layer0_outputs[634] = ~((inputs[164]) ^ (inputs[186]));
    assign layer0_outputs[635] = ~((inputs[253]) ^ (inputs[193]));
    assign layer0_outputs[636] = (inputs[150]) & (inputs[237]);
    assign layer0_outputs[637] = (inputs[230]) & ~(inputs[202]);
    assign layer0_outputs[638] = ~(inputs[201]) | (inputs[32]);
    assign layer0_outputs[639] = ~(inputs[152]);
    assign layer0_outputs[640] = ~(inputs[85]) | (inputs[24]);
    assign layer0_outputs[641] = inputs[233];
    assign layer0_outputs[642] = ~(inputs[210]);
    assign layer0_outputs[643] = ~(inputs[229]) | (inputs[176]);
    assign layer0_outputs[644] = (inputs[98]) | (inputs[122]);
    assign layer0_outputs[645] = ~(inputs[158]);
    assign layer0_outputs[646] = ~(inputs[76]);
    assign layer0_outputs[647] = ~((inputs[101]) | (inputs[70]));
    assign layer0_outputs[648] = (inputs[252]) & (inputs[17]);
    assign layer0_outputs[649] = 1'b1;
    assign layer0_outputs[650] = ~(inputs[43]) | (inputs[6]);
    assign layer0_outputs[651] = ~(inputs[58]);
    assign layer0_outputs[652] = ~((inputs[28]) & (inputs[161]));
    assign layer0_outputs[653] = (inputs[64]) | (inputs[99]);
    assign layer0_outputs[654] = (inputs[132]) & ~(inputs[112]);
    assign layer0_outputs[655] = ~(inputs[79]) | (inputs[25]);
    assign layer0_outputs[656] = ~(inputs[195]) | (inputs[177]);
    assign layer0_outputs[657] = ~(inputs[90]) | (inputs[0]);
    assign layer0_outputs[658] = (inputs[209]) | (inputs[171]);
    assign layer0_outputs[659] = ~(inputs[227]) | (inputs[6]);
    assign layer0_outputs[660] = (inputs[245]) & ~(inputs[175]);
    assign layer0_outputs[661] = (inputs[31]) | (inputs[7]);
    assign layer0_outputs[662] = (inputs[201]) & ~(inputs[131]);
    assign layer0_outputs[663] = (inputs[211]) & (inputs[143]);
    assign layer0_outputs[664] = inputs[188];
    assign layer0_outputs[665] = (inputs[86]) & ~(inputs[43]);
    assign layer0_outputs[666] = ~((inputs[232]) | (inputs[66]));
    assign layer0_outputs[667] = inputs[107];
    assign layer0_outputs[668] = (inputs[71]) & ~(inputs[30]);
    assign layer0_outputs[669] = ~((inputs[196]) | (inputs[218]));
    assign layer0_outputs[670] = (inputs[213]) ^ (inputs[244]);
    assign layer0_outputs[671] = (inputs[44]) ^ (inputs[219]);
    assign layer0_outputs[672] = ~(inputs[103]) | (inputs[220]);
    assign layer0_outputs[673] = inputs[61];
    assign layer0_outputs[674] = ~(inputs[178]) | (inputs[26]);
    assign layer0_outputs[675] = ~(inputs[49]);
    assign layer0_outputs[676] = (inputs[210]) & (inputs[250]);
    assign layer0_outputs[677] = ~(inputs[134]);
    assign layer0_outputs[678] = ~((inputs[92]) & (inputs[74]));
    assign layer0_outputs[679] = ~(inputs[112]) | (inputs[20]);
    assign layer0_outputs[680] = ~((inputs[249]) | (inputs[45]));
    assign layer0_outputs[681] = ~((inputs[20]) ^ (inputs[238]));
    assign layer0_outputs[682] = ~((inputs[87]) ^ (inputs[224]));
    assign layer0_outputs[683] = ~(inputs[149]);
    assign layer0_outputs[684] = ~(inputs[112]);
    assign layer0_outputs[685] = ~(inputs[119]);
    assign layer0_outputs[686] = ~((inputs[50]) ^ (inputs[0]));
    assign layer0_outputs[687] = ~((inputs[96]) ^ (inputs[67]));
    assign layer0_outputs[688] = (inputs[67]) & ~(inputs[1]);
    assign layer0_outputs[689] = inputs[104];
    assign layer0_outputs[690] = ~(inputs[72]);
    assign layer0_outputs[691] = ~((inputs[188]) ^ (inputs[225]));
    assign layer0_outputs[692] = ~(inputs[180]);
    assign layer0_outputs[693] = ~(inputs[88]);
    assign layer0_outputs[694] = (inputs[127]) | (inputs[1]);
    assign layer0_outputs[695] = ~((inputs[113]) ^ (inputs[67]));
    assign layer0_outputs[696] = inputs[182];
    assign layer0_outputs[697] = inputs[227];
    assign layer0_outputs[698] = ~((inputs[224]) | (inputs[149]));
    assign layer0_outputs[699] = inputs[202];
    assign layer0_outputs[700] = (inputs[229]) & ~(inputs[11]);
    assign layer0_outputs[701] = (inputs[238]) | (inputs[195]);
    assign layer0_outputs[702] = ~(inputs[137]);
    assign layer0_outputs[703] = (inputs[177]) & (inputs[42]);
    assign layer0_outputs[704] = ~(inputs[171]) | (inputs[27]);
    assign layer0_outputs[705] = (inputs[147]) & (inputs[127]);
    assign layer0_outputs[706] = ~(inputs[162]);
    assign layer0_outputs[707] = (inputs[230]) & ~(inputs[16]);
    assign layer0_outputs[708] = ~(inputs[159]);
    assign layer0_outputs[709] = ~((inputs[239]) | (inputs[56]));
    assign layer0_outputs[710] = (inputs[39]) ^ (inputs[139]);
    assign layer0_outputs[711] = ~(inputs[134]) | (inputs[214]);
    assign layer0_outputs[712] = (inputs[118]) & ~(inputs[161]);
    assign layer0_outputs[713] = ~((inputs[181]) & (inputs[179]));
    assign layer0_outputs[714] = 1'b1;
    assign layer0_outputs[715] = (inputs[33]) ^ (inputs[3]);
    assign layer0_outputs[716] = 1'b1;
    assign layer0_outputs[717] = (inputs[58]) & (inputs[154]);
    assign layer0_outputs[718] = ~(inputs[200]) | (inputs[78]);
    assign layer0_outputs[719] = ~((inputs[190]) & (inputs[251]));
    assign layer0_outputs[720] = ~(inputs[104]);
    assign layer0_outputs[721] = ~((inputs[61]) ^ (inputs[158]));
    assign layer0_outputs[722] = (inputs[51]) & ~(inputs[241]);
    assign layer0_outputs[723] = 1'b0;
    assign layer0_outputs[724] = ~(inputs[201]) | (inputs[20]);
    assign layer0_outputs[725] = inputs[74];
    assign layer0_outputs[726] = (inputs[155]) | (inputs[207]);
    assign layer0_outputs[727] = (inputs[5]) | (inputs[137]);
    assign layer0_outputs[728] = inputs[8];
    assign layer0_outputs[729] = (inputs[144]) | (inputs[201]);
    assign layer0_outputs[730] = inputs[96];
    assign layer0_outputs[731] = (inputs[230]) | (inputs[105]);
    assign layer0_outputs[732] = ~(inputs[188]) | (inputs[108]);
    assign layer0_outputs[733] = inputs[219];
    assign layer0_outputs[734] = ~(inputs[129]);
    assign layer0_outputs[735] = ~((inputs[171]) ^ (inputs[52]));
    assign layer0_outputs[736] = 1'b1;
    assign layer0_outputs[737] = ~((inputs[251]) | (inputs[90]));
    assign layer0_outputs[738] = ~(inputs[119]);
    assign layer0_outputs[739] = (inputs[47]) & ~(inputs[226]);
    assign layer0_outputs[740] = (inputs[130]) & (inputs[21]);
    assign layer0_outputs[741] = ~(inputs[196]);
    assign layer0_outputs[742] = (inputs[10]) & ~(inputs[26]);
    assign layer0_outputs[743] = ~((inputs[207]) ^ (inputs[171]));
    assign layer0_outputs[744] = ~((inputs[42]) | (inputs[181]));
    assign layer0_outputs[745] = ~(inputs[242]) | (inputs[190]);
    assign layer0_outputs[746] = (inputs[179]) & ~(inputs[13]);
    assign layer0_outputs[747] = ~(inputs[116]) | (inputs[228]);
    assign layer0_outputs[748] = inputs[168];
    assign layer0_outputs[749] = ~((inputs[232]) ^ (inputs[6]));
    assign layer0_outputs[750] = inputs[57];
    assign layer0_outputs[751] = (inputs[13]) | (inputs[18]);
    assign layer0_outputs[752] = ~((inputs[35]) | (inputs[215]));
    assign layer0_outputs[753] = (inputs[31]) | (inputs[103]);
    assign layer0_outputs[754] = (inputs[254]) | (inputs[50]);
    assign layer0_outputs[755] = ~((inputs[10]) ^ (inputs[132]));
    assign layer0_outputs[756] = (inputs[44]) ^ (inputs[9]);
    assign layer0_outputs[757] = ~(inputs[0]) | (inputs[11]);
    assign layer0_outputs[758] = (inputs[248]) & (inputs[185]);
    assign layer0_outputs[759] = (inputs[20]) | (inputs[20]);
    assign layer0_outputs[760] = ~((inputs[249]) | (inputs[218]));
    assign layer0_outputs[761] = inputs[105];
    assign layer0_outputs[762] = (inputs[77]) | (inputs[138]);
    assign layer0_outputs[763] = 1'b0;
    assign layer0_outputs[764] = ~(inputs[143]) | (inputs[242]);
    assign layer0_outputs[765] = ~((inputs[238]) ^ (inputs[102]));
    assign layer0_outputs[766] = ~((inputs[218]) ^ (inputs[45]));
    assign layer0_outputs[767] = (inputs[216]) | (inputs[30]);
    assign layer0_outputs[768] = ~((inputs[145]) ^ (inputs[190]));
    assign layer0_outputs[769] = ~(inputs[216]) | (inputs[18]);
    assign layer0_outputs[770] = inputs[140];
    assign layer0_outputs[771] = ~((inputs[181]) | (inputs[128]));
    assign layer0_outputs[772] = 1'b0;
    assign layer0_outputs[773] = (inputs[180]) ^ (inputs[115]);
    assign layer0_outputs[774] = inputs[135];
    assign layer0_outputs[775] = inputs[61];
    assign layer0_outputs[776] = 1'b1;
    assign layer0_outputs[777] = ~((inputs[128]) ^ (inputs[78]));
    assign layer0_outputs[778] = ~((inputs[129]) | (inputs[137]));
    assign layer0_outputs[779] = ~((inputs[166]) | (inputs[194]));
    assign layer0_outputs[780] = inputs[43];
    assign layer0_outputs[781] = (inputs[116]) | (inputs[0]);
    assign layer0_outputs[782] = ~((inputs[81]) ^ (inputs[60]));
    assign layer0_outputs[783] = ~(inputs[118]);
    assign layer0_outputs[784] = (inputs[95]) & ~(inputs[247]);
    assign layer0_outputs[785] = (inputs[63]) ^ (inputs[56]);
    assign layer0_outputs[786] = ~((inputs[206]) | (inputs[77]));
    assign layer0_outputs[787] = (inputs[168]) & ~(inputs[201]);
    assign layer0_outputs[788] = inputs[68];
    assign layer0_outputs[789] = ~((inputs[156]) ^ (inputs[223]));
    assign layer0_outputs[790] = ~(inputs[24]);
    assign layer0_outputs[791] = (inputs[119]) | (inputs[146]);
    assign layer0_outputs[792] = (inputs[4]) ^ (inputs[17]);
    assign layer0_outputs[793] = (inputs[230]) | (inputs[229]);
    assign layer0_outputs[794] = (inputs[154]) & ~(inputs[3]);
    assign layer0_outputs[795] = ~((inputs[239]) ^ (inputs[163]));
    assign layer0_outputs[796] = ~((inputs[194]) | (inputs[235]));
    assign layer0_outputs[797] = ~(inputs[34]);
    assign layer0_outputs[798] = ~(inputs[155]);
    assign layer0_outputs[799] = (inputs[173]) & ~(inputs[31]);
    assign layer0_outputs[800] = ~((inputs[119]) | (inputs[132]));
    assign layer0_outputs[801] = ~(inputs[55]);
    assign layer0_outputs[802] = (inputs[1]) ^ (inputs[100]);
    assign layer0_outputs[803] = (inputs[232]) & ~(inputs[188]);
    assign layer0_outputs[804] = ~(inputs[28]) | (inputs[109]);
    assign layer0_outputs[805] = inputs[118];
    assign layer0_outputs[806] = (inputs[61]) | (inputs[68]);
    assign layer0_outputs[807] = (inputs[60]) ^ (inputs[93]);
    assign layer0_outputs[808] = (inputs[74]) & ~(inputs[23]);
    assign layer0_outputs[809] = ~(inputs[145]) | (inputs[208]);
    assign layer0_outputs[810] = (inputs[183]) & ~(inputs[189]);
    assign layer0_outputs[811] = ~(inputs[0]) | (inputs[185]);
    assign layer0_outputs[812] = (inputs[27]) ^ (inputs[12]);
    assign layer0_outputs[813] = ~((inputs[232]) ^ (inputs[22]));
    assign layer0_outputs[814] = ~((inputs[219]) ^ (inputs[199]));
    assign layer0_outputs[815] = (inputs[184]) | (inputs[162]);
    assign layer0_outputs[816] = inputs[39];
    assign layer0_outputs[817] = ~(inputs[79]) | (inputs[5]);
    assign layer0_outputs[818] = ~(inputs[106]);
    assign layer0_outputs[819] = inputs[119];
    assign layer0_outputs[820] = inputs[229];
    assign layer0_outputs[821] = ~((inputs[255]) | (inputs[36]));
    assign layer0_outputs[822] = (inputs[162]) ^ (inputs[84]);
    assign layer0_outputs[823] = 1'b0;
    assign layer0_outputs[824] = (inputs[12]) | (inputs[221]);
    assign layer0_outputs[825] = ~(inputs[250]) | (inputs[50]);
    assign layer0_outputs[826] = ~(inputs[11]) | (inputs[17]);
    assign layer0_outputs[827] = ~((inputs[96]) ^ (inputs[80]));
    assign layer0_outputs[828] = (inputs[201]) & ~(inputs[162]);
    assign layer0_outputs[829] = ~(inputs[46]) | (inputs[190]);
    assign layer0_outputs[830] = ~(inputs[136]) | (inputs[21]);
    assign layer0_outputs[831] = ~((inputs[255]) ^ (inputs[52]));
    assign layer0_outputs[832] = ~((inputs[218]) ^ (inputs[32]));
    assign layer0_outputs[833] = ~(inputs[156]) | (inputs[66]);
    assign layer0_outputs[834] = ~((inputs[48]) ^ (inputs[152]));
    assign layer0_outputs[835] = (inputs[205]) | (inputs[26]);
    assign layer0_outputs[836] = ~(inputs[121]);
    assign layer0_outputs[837] = (inputs[81]) ^ (inputs[140]);
    assign layer0_outputs[838] = inputs[115];
    assign layer0_outputs[839] = (inputs[153]) & ~(inputs[40]);
    assign layer0_outputs[840] = (inputs[64]) | (inputs[251]);
    assign layer0_outputs[841] = ~(inputs[245]);
    assign layer0_outputs[842] = (inputs[141]) | (inputs[237]);
    assign layer0_outputs[843] = 1'b1;
    assign layer0_outputs[844] = ~((inputs[168]) ^ (inputs[60]));
    assign layer0_outputs[845] = ~(inputs[212]);
    assign layer0_outputs[846] = (inputs[185]) | (inputs[206]);
    assign layer0_outputs[847] = (inputs[208]) & ~(inputs[47]);
    assign layer0_outputs[848] = ~(inputs[100]);
    assign layer0_outputs[849] = ~((inputs[11]) ^ (inputs[108]));
    assign layer0_outputs[850] = (inputs[23]) & (inputs[241]);
    assign layer0_outputs[851] = ~((inputs[168]) ^ (inputs[215]));
    assign layer0_outputs[852] = (inputs[98]) & (inputs[53]);
    assign layer0_outputs[853] = ~(inputs[101]);
    assign layer0_outputs[854] = ~(inputs[220]) | (inputs[160]);
    assign layer0_outputs[855] = 1'b0;
    assign layer0_outputs[856] = ~(inputs[153]) | (inputs[180]);
    assign layer0_outputs[857] = (inputs[3]) & ~(inputs[163]);
    assign layer0_outputs[858] = (inputs[215]) & ~(inputs[44]);
    assign layer0_outputs[859] = 1'b1;
    assign layer0_outputs[860] = inputs[154];
    assign layer0_outputs[861] = inputs[251];
    assign layer0_outputs[862] = ~((inputs[106]) | (inputs[153]));
    assign layer0_outputs[863] = (inputs[36]) & (inputs[252]);
    assign layer0_outputs[864] = (inputs[228]) ^ (inputs[161]);
    assign layer0_outputs[865] = (inputs[246]) & ~(inputs[243]);
    assign layer0_outputs[866] = ~(inputs[14]) | (inputs[114]);
    assign layer0_outputs[867] = ~(inputs[220]);
    assign layer0_outputs[868] = (inputs[166]) | (inputs[141]);
    assign layer0_outputs[869] = ~((inputs[249]) & (inputs[111]));
    assign layer0_outputs[870] = ~((inputs[99]) | (inputs[106]));
    assign layer0_outputs[871] = (inputs[88]) & ~(inputs[134]);
    assign layer0_outputs[872] = (inputs[167]) & ~(inputs[244]);
    assign layer0_outputs[873] = ~((inputs[160]) | (inputs[166]));
    assign layer0_outputs[874] = ~((inputs[162]) | (inputs[164]));
    assign layer0_outputs[875] = inputs[155];
    assign layer0_outputs[876] = (inputs[132]) & ~(inputs[193]);
    assign layer0_outputs[877] = (inputs[73]) & ~(inputs[127]);
    assign layer0_outputs[878] = ~(inputs[204]);
    assign layer0_outputs[879] = inputs[25];
    assign layer0_outputs[880] = ~((inputs[205]) | (inputs[249]));
    assign layer0_outputs[881] = 1'b1;
    assign layer0_outputs[882] = inputs[132];
    assign layer0_outputs[883] = (inputs[192]) & ~(inputs[160]);
    assign layer0_outputs[884] = ~((inputs[60]) ^ (inputs[236]));
    assign layer0_outputs[885] = ~(inputs[102]) | (inputs[195]);
    assign layer0_outputs[886] = (inputs[115]) & ~(inputs[22]);
    assign layer0_outputs[887] = 1'b0;
    assign layer0_outputs[888] = inputs[39];
    assign layer0_outputs[889] = ~((inputs[128]) | (inputs[208]));
    assign layer0_outputs[890] = inputs[65];
    assign layer0_outputs[891] = ~((inputs[90]) | (inputs[229]));
    assign layer0_outputs[892] = ~(inputs[36]);
    assign layer0_outputs[893] = ~((inputs[58]) & (inputs[223]));
    assign layer0_outputs[894] = ~(inputs[124]);
    assign layer0_outputs[895] = ~((inputs[234]) | (inputs[54]));
    assign layer0_outputs[896] = ~((inputs[60]) | (inputs[220]));
    assign layer0_outputs[897] = inputs[12];
    assign layer0_outputs[898] = ~((inputs[70]) | (inputs[75]));
    assign layer0_outputs[899] = inputs[47];
    assign layer0_outputs[900] = (inputs[199]) & ~(inputs[215]);
    assign layer0_outputs[901] = ~((inputs[85]) ^ (inputs[159]));
    assign layer0_outputs[902] = (inputs[206]) ^ (inputs[59]);
    assign layer0_outputs[903] = 1'b0;
    assign layer0_outputs[904] = (inputs[28]) & ~(inputs[247]);
    assign layer0_outputs[905] = (inputs[230]) ^ (inputs[29]);
    assign layer0_outputs[906] = ~((inputs[232]) ^ (inputs[168]));
    assign layer0_outputs[907] = (inputs[60]) | (inputs[8]);
    assign layer0_outputs[908] = inputs[155];
    assign layer0_outputs[909] = ~((inputs[192]) ^ (inputs[68]));
    assign layer0_outputs[910] = ~(inputs[152]) | (inputs[52]);
    assign layer0_outputs[911] = ~(inputs[196]);
    assign layer0_outputs[912] = (inputs[25]) ^ (inputs[219]);
    assign layer0_outputs[913] = ~((inputs[226]) ^ (inputs[84]));
    assign layer0_outputs[914] = ~(inputs[101]);
    assign layer0_outputs[915] = (inputs[125]) & ~(inputs[13]);
    assign layer0_outputs[916] = (inputs[72]) & ~(inputs[103]);
    assign layer0_outputs[917] = ~(inputs[26]) | (inputs[250]);
    assign layer0_outputs[918] = ~((inputs[255]) | (inputs[159]));
    assign layer0_outputs[919] = ~(inputs[121]) | (inputs[204]);
    assign layer0_outputs[920] = ~((inputs[113]) | (inputs[246]));
    assign layer0_outputs[921] = 1'b1;
    assign layer0_outputs[922] = ~((inputs[104]) | (inputs[255]));
    assign layer0_outputs[923] = (inputs[49]) | (inputs[121]);
    assign layer0_outputs[924] = ~((inputs[255]) | (inputs[183]));
    assign layer0_outputs[925] = inputs[67];
    assign layer0_outputs[926] = inputs[56];
    assign layer0_outputs[927] = (inputs[42]) | (inputs[197]);
    assign layer0_outputs[928] = ~((inputs[164]) | (inputs[185]));
    assign layer0_outputs[929] = inputs[197];
    assign layer0_outputs[930] = ~((inputs[197]) | (inputs[76]));
    assign layer0_outputs[931] = (inputs[155]) & ~(inputs[75]);
    assign layer0_outputs[932] = (inputs[23]) | (inputs[7]);
    assign layer0_outputs[933] = ~((inputs[149]) ^ (inputs[112]));
    assign layer0_outputs[934] = (inputs[183]) & ~(inputs[241]);
    assign layer0_outputs[935] = ~(inputs[101]) | (inputs[244]);
    assign layer0_outputs[936] = (inputs[39]) & (inputs[185]);
    assign layer0_outputs[937] = (inputs[250]) & ~(inputs[242]);
    assign layer0_outputs[938] = ~(inputs[243]);
    assign layer0_outputs[939] = (inputs[243]) & ~(inputs[53]);
    assign layer0_outputs[940] = (inputs[87]) | (inputs[235]);
    assign layer0_outputs[941] = ~((inputs[217]) ^ (inputs[168]));
    assign layer0_outputs[942] = ~(inputs[168]);
    assign layer0_outputs[943] = ~((inputs[37]) & (inputs[227]));
    assign layer0_outputs[944] = inputs[118];
    assign layer0_outputs[945] = inputs[7];
    assign layer0_outputs[946] = inputs[106];
    assign layer0_outputs[947] = ~(inputs[248]) | (inputs[36]);
    assign layer0_outputs[948] = ~(inputs[60]) | (inputs[119]);
    assign layer0_outputs[949] = ~(inputs[207]) | (inputs[207]);
    assign layer0_outputs[950] = (inputs[113]) ^ (inputs[30]);
    assign layer0_outputs[951] = ~((inputs[65]) ^ (inputs[221]));
    assign layer0_outputs[952] = (inputs[103]) | (inputs[139]);
    assign layer0_outputs[953] = 1'b0;
    assign layer0_outputs[954] = ~(inputs[85]);
    assign layer0_outputs[955] = (inputs[222]) | (inputs[42]);
    assign layer0_outputs[956] = inputs[149];
    assign layer0_outputs[957] = (inputs[254]) | (inputs[240]);
    assign layer0_outputs[958] = (inputs[148]) & ~(inputs[254]);
    assign layer0_outputs[959] = (inputs[156]) & ~(inputs[161]);
    assign layer0_outputs[960] = ~(inputs[109]) | (inputs[227]);
    assign layer0_outputs[961] = (inputs[181]) & ~(inputs[8]);
    assign layer0_outputs[962] = inputs[71];
    assign layer0_outputs[963] = ~((inputs[217]) | (inputs[228]));
    assign layer0_outputs[964] = ~(inputs[39]);
    assign layer0_outputs[965] = ~(inputs[102]) | (inputs[65]);
    assign layer0_outputs[966] = ~((inputs[141]) | (inputs[96]));
    assign layer0_outputs[967] = inputs[202];
    assign layer0_outputs[968] = (inputs[123]) & ~(inputs[66]);
    assign layer0_outputs[969] = (inputs[219]) & (inputs[33]);
    assign layer0_outputs[970] = ~(inputs[13]) | (inputs[37]);
    assign layer0_outputs[971] = 1'b1;
    assign layer0_outputs[972] = (inputs[79]) ^ (inputs[165]);
    assign layer0_outputs[973] = (inputs[128]) & ~(inputs[94]);
    assign layer0_outputs[974] = (inputs[161]) & ~(inputs[231]);
    assign layer0_outputs[975] = inputs[164];
    assign layer0_outputs[976] = (inputs[141]) & ~(inputs[251]);
    assign layer0_outputs[977] = ~(inputs[71]);
    assign layer0_outputs[978] = ~(inputs[137]) | (inputs[158]);
    assign layer0_outputs[979] = ~((inputs[104]) ^ (inputs[20]));
    assign layer0_outputs[980] = ~(inputs[58]) | (inputs[114]);
    assign layer0_outputs[981] = ~((inputs[84]) | (inputs[110]));
    assign layer0_outputs[982] = (inputs[142]) & (inputs[112]);
    assign layer0_outputs[983] = ~(inputs[117]) | (inputs[249]);
    assign layer0_outputs[984] = ~(inputs[58]);
    assign layer0_outputs[985] = inputs[41];
    assign layer0_outputs[986] = inputs[215];
    assign layer0_outputs[987] = (inputs[83]) | (inputs[105]);
    assign layer0_outputs[988] = inputs[107];
    assign layer0_outputs[989] = (inputs[246]) & (inputs[31]);
    assign layer0_outputs[990] = ~(inputs[46]);
    assign layer0_outputs[991] = ~((inputs[60]) | (inputs[76]));
    assign layer0_outputs[992] = ~((inputs[210]) | (inputs[142]));
    assign layer0_outputs[993] = ~((inputs[39]) | (inputs[158]));
    assign layer0_outputs[994] = (inputs[55]) & ~(inputs[244]);
    assign layer0_outputs[995] = (inputs[214]) ^ (inputs[32]);
    assign layer0_outputs[996] = ~((inputs[128]) ^ (inputs[135]));
    assign layer0_outputs[997] = (inputs[146]) & ~(inputs[252]);
    assign layer0_outputs[998] = ~(inputs[153]) | (inputs[245]);
    assign layer0_outputs[999] = (inputs[238]) & ~(inputs[71]);
    assign layer0_outputs[1000] = inputs[118];
    assign layer0_outputs[1001] = ~((inputs[138]) ^ (inputs[209]));
    assign layer0_outputs[1002] = inputs[137];
    assign layer0_outputs[1003] = (inputs[96]) ^ (inputs[216]);
    assign layer0_outputs[1004] = ~(inputs[198]);
    assign layer0_outputs[1005] = inputs[55];
    assign layer0_outputs[1006] = inputs[89];
    assign layer0_outputs[1007] = ~((inputs[103]) | (inputs[94]));
    assign layer0_outputs[1008] = ~(inputs[127]) | (inputs[8]);
    assign layer0_outputs[1009] = ~((inputs[31]) | (inputs[240]));
    assign layer0_outputs[1010] = ~((inputs[190]) ^ (inputs[178]));
    assign layer0_outputs[1011] = (inputs[72]) | (inputs[67]);
    assign layer0_outputs[1012] = ~(inputs[243]);
    assign layer0_outputs[1013] = (inputs[197]) & ~(inputs[210]);
    assign layer0_outputs[1014] = ~(inputs[66]);
    assign layer0_outputs[1015] = ~(inputs[145]);
    assign layer0_outputs[1016] = 1'b0;
    assign layer0_outputs[1017] = ~(inputs[27]);
    assign layer0_outputs[1018] = ~((inputs[120]) ^ (inputs[129]));
    assign layer0_outputs[1019] = ~(inputs[103]) | (inputs[29]);
    assign layer0_outputs[1020] = ~(inputs[55]) | (inputs[167]);
    assign layer0_outputs[1021] = (inputs[77]) | (inputs[40]);
    assign layer0_outputs[1022] = (inputs[58]) ^ (inputs[11]);
    assign layer0_outputs[1023] = 1'b1;
    assign layer0_outputs[1024] = inputs[106];
    assign layer0_outputs[1025] = inputs[100];
    assign layer0_outputs[1026] = inputs[140];
    assign layer0_outputs[1027] = ~(inputs[93]) | (inputs[194]);
    assign layer0_outputs[1028] = inputs[119];
    assign layer0_outputs[1029] = ~((inputs[154]) | (inputs[8]));
    assign layer0_outputs[1030] = ~(inputs[150]) | (inputs[215]);
    assign layer0_outputs[1031] = (inputs[84]) & ~(inputs[208]);
    assign layer0_outputs[1032] = (inputs[84]) | (inputs[180]);
    assign layer0_outputs[1033] = ~((inputs[49]) ^ (inputs[171]));
    assign layer0_outputs[1034] = ~(inputs[119]);
    assign layer0_outputs[1035] = (inputs[152]) & ~(inputs[27]);
    assign layer0_outputs[1036] = (inputs[55]) | (inputs[54]);
    assign layer0_outputs[1037] = ~(inputs[39]);
    assign layer0_outputs[1038] = inputs[172];
    assign layer0_outputs[1039] = ~((inputs[228]) | (inputs[154]));
    assign layer0_outputs[1040] = (inputs[151]) ^ (inputs[95]);
    assign layer0_outputs[1041] = (inputs[248]) ^ (inputs[250]);
    assign layer0_outputs[1042] = (inputs[15]) ^ (inputs[198]);
    assign layer0_outputs[1043] = ~(inputs[73]) | (inputs[27]);
    assign layer0_outputs[1044] = (inputs[8]) ^ (inputs[120]);
    assign layer0_outputs[1045] = 1'b0;
    assign layer0_outputs[1046] = ~(inputs[136]) | (inputs[171]);
    assign layer0_outputs[1047] = ~((inputs[179]) ^ (inputs[24]));
    assign layer0_outputs[1048] = ~(inputs[221]);
    assign layer0_outputs[1049] = ~((inputs[153]) ^ (inputs[19]));
    assign layer0_outputs[1050] = (inputs[141]) ^ (inputs[206]);
    assign layer0_outputs[1051] = (inputs[115]) & ~(inputs[242]);
    assign layer0_outputs[1052] = 1'b1;
    assign layer0_outputs[1053] = (inputs[125]) & ~(inputs[210]);
    assign layer0_outputs[1054] = inputs[47];
    assign layer0_outputs[1055] = ~((inputs[141]) | (inputs[147]));
    assign layer0_outputs[1056] = ~(inputs[106]) | (inputs[195]);
    assign layer0_outputs[1057] = ~(inputs[69]) | (inputs[8]);
    assign layer0_outputs[1058] = ~((inputs[39]) | (inputs[123]));
    assign layer0_outputs[1059] = ~((inputs[254]) | (inputs[163]));
    assign layer0_outputs[1060] = (inputs[106]) & ~(inputs[177]);
    assign layer0_outputs[1061] = inputs[112];
    assign layer0_outputs[1062] = (inputs[158]) & ~(inputs[177]);
    assign layer0_outputs[1063] = inputs[121];
    assign layer0_outputs[1064] = ~((inputs[78]) ^ (inputs[164]));
    assign layer0_outputs[1065] = ~(inputs[120]) | (inputs[202]);
    assign layer0_outputs[1066] = (inputs[67]) & ~(inputs[191]);
    assign layer0_outputs[1067] = (inputs[73]) | (inputs[144]);
    assign layer0_outputs[1068] = inputs[112];
    assign layer0_outputs[1069] = (inputs[165]) | (inputs[223]);
    assign layer0_outputs[1070] = ~((inputs[195]) | (inputs[191]));
    assign layer0_outputs[1071] = inputs[49];
    assign layer0_outputs[1072] = ~(inputs[119]) | (inputs[7]);
    assign layer0_outputs[1073] = ~(inputs[197]);
    assign layer0_outputs[1074] = inputs[249];
    assign layer0_outputs[1075] = ~((inputs[65]) & (inputs[61]));
    assign layer0_outputs[1076] = ~(inputs[112]) | (inputs[210]);
    assign layer0_outputs[1077] = inputs[200];
    assign layer0_outputs[1078] = ~(inputs[100]);
    assign layer0_outputs[1079] = (inputs[139]) & ~(inputs[194]);
    assign layer0_outputs[1080] = inputs[104];
    assign layer0_outputs[1081] = (inputs[109]) | (inputs[109]);
    assign layer0_outputs[1082] = (inputs[3]) | (inputs[237]);
    assign layer0_outputs[1083] = ~(inputs[210]) | (inputs[66]);
    assign layer0_outputs[1084] = (inputs[9]) | (inputs[63]);
    assign layer0_outputs[1085] = (inputs[152]) ^ (inputs[248]);
    assign layer0_outputs[1086] = (inputs[158]) & (inputs[104]);
    assign layer0_outputs[1087] = (inputs[9]) ^ (inputs[186]);
    assign layer0_outputs[1088] = ~((inputs[32]) ^ (inputs[214]));
    assign layer0_outputs[1089] = (inputs[229]) & ~(inputs[84]);
    assign layer0_outputs[1090] = ~(inputs[53]);
    assign layer0_outputs[1091] = (inputs[103]) | (inputs[118]);
    assign layer0_outputs[1092] = (inputs[222]) ^ (inputs[91]);
    assign layer0_outputs[1093] = (inputs[52]) | (inputs[199]);
    assign layer0_outputs[1094] = 1'b1;
    assign layer0_outputs[1095] = (inputs[237]) ^ (inputs[166]);
    assign layer0_outputs[1096] = ~((inputs[90]) | (inputs[228]));
    assign layer0_outputs[1097] = inputs[103];
    assign layer0_outputs[1098] = ~(inputs[187]);
    assign layer0_outputs[1099] = inputs[96];
    assign layer0_outputs[1100] = inputs[241];
    assign layer0_outputs[1101] = ~((inputs[60]) ^ (inputs[78]));
    assign layer0_outputs[1102] = ~(inputs[238]) | (inputs[14]);
    assign layer0_outputs[1103] = (inputs[18]) ^ (inputs[163]);
    assign layer0_outputs[1104] = (inputs[96]) | (inputs[212]);
    assign layer0_outputs[1105] = (inputs[196]) & (inputs[42]);
    assign layer0_outputs[1106] = (inputs[117]) & ~(inputs[52]);
    assign layer0_outputs[1107] = (inputs[30]) ^ (inputs[148]);
    assign layer0_outputs[1108] = ~(inputs[74]);
    assign layer0_outputs[1109] = (inputs[63]) & ~(inputs[110]);
    assign layer0_outputs[1110] = ~(inputs[236]);
    assign layer0_outputs[1111] = (inputs[21]) | (inputs[5]);
    assign layer0_outputs[1112] = (inputs[94]) | (inputs[140]);
    assign layer0_outputs[1113] = ~((inputs[243]) | (inputs[110]));
    assign layer0_outputs[1114] = ~((inputs[17]) ^ (inputs[159]));
    assign layer0_outputs[1115] = inputs[186];
    assign layer0_outputs[1116] = (inputs[98]) | (inputs[59]);
    assign layer0_outputs[1117] = ~((inputs[40]) ^ (inputs[8]));
    assign layer0_outputs[1118] = inputs[59];
    assign layer0_outputs[1119] = ~(inputs[226]);
    assign layer0_outputs[1120] = (inputs[243]) & ~(inputs[53]);
    assign layer0_outputs[1121] = ~((inputs[211]) | (inputs[114]));
    assign layer0_outputs[1122] = ~((inputs[48]) | (inputs[140]));
    assign layer0_outputs[1123] = ~((inputs[144]) & (inputs[110]));
    assign layer0_outputs[1124] = 1'b1;
    assign layer0_outputs[1125] = (inputs[238]) | (inputs[40]);
    assign layer0_outputs[1126] = inputs[111];
    assign layer0_outputs[1127] = 1'b0;
    assign layer0_outputs[1128] = inputs[90];
    assign layer0_outputs[1129] = (inputs[153]) | (inputs[119]);
    assign layer0_outputs[1130] = ~((inputs[31]) | (inputs[206]));
    assign layer0_outputs[1131] = inputs[221];
    assign layer0_outputs[1132] = ~((inputs[160]) | (inputs[167]));
    assign layer0_outputs[1133] = ~(inputs[195]) | (inputs[29]);
    assign layer0_outputs[1134] = ~(inputs[121]) | (inputs[50]);
    assign layer0_outputs[1135] = (inputs[11]) & ~(inputs[50]);
    assign layer0_outputs[1136] = inputs[94];
    assign layer0_outputs[1137] = (inputs[160]) | (inputs[90]);
    assign layer0_outputs[1138] = ~((inputs[161]) | (inputs[197]));
    assign layer0_outputs[1139] = 1'b1;
    assign layer0_outputs[1140] = (inputs[23]) & ~(inputs[202]);
    assign layer0_outputs[1141] = ~(inputs[29]) | (inputs[224]);
    assign layer0_outputs[1142] = ~((inputs[172]) & (inputs[132]));
    assign layer0_outputs[1143] = (inputs[119]) & ~(inputs[235]);
    assign layer0_outputs[1144] = ~(inputs[111]);
    assign layer0_outputs[1145] = ~((inputs[188]) | (inputs[6]));
    assign layer0_outputs[1146] = inputs[160];
    assign layer0_outputs[1147] = inputs[94];
    assign layer0_outputs[1148] = (inputs[180]) & ~(inputs[226]);
    assign layer0_outputs[1149] = ~((inputs[226]) ^ (inputs[158]));
    assign layer0_outputs[1150] = 1'b1;
    assign layer0_outputs[1151] = ~((inputs[14]) | (inputs[51]));
    assign layer0_outputs[1152] = ~((inputs[172]) | (inputs[171]));
    assign layer0_outputs[1153] = (inputs[110]) ^ (inputs[193]);
    assign layer0_outputs[1154] = inputs[209];
    assign layer0_outputs[1155] = inputs[136];
    assign layer0_outputs[1156] = (inputs[176]) & ~(inputs[245]);
    assign layer0_outputs[1157] = (inputs[204]) | (inputs[194]);
    assign layer0_outputs[1158] = ~(inputs[117]);
    assign layer0_outputs[1159] = 1'b0;
    assign layer0_outputs[1160] = (inputs[214]) | (inputs[13]);
    assign layer0_outputs[1161] = ~(inputs[63]) | (inputs[43]);
    assign layer0_outputs[1162] = ~(inputs[148]);
    assign layer0_outputs[1163] = (inputs[136]) & ~(inputs[50]);
    assign layer0_outputs[1164] = inputs[88];
    assign layer0_outputs[1165] = ~(inputs[187]) | (inputs[169]);
    assign layer0_outputs[1166] = ~((inputs[27]) ^ (inputs[247]));
    assign layer0_outputs[1167] = inputs[158];
    assign layer0_outputs[1168] = (inputs[115]) | (inputs[124]);
    assign layer0_outputs[1169] = inputs[254];
    assign layer0_outputs[1170] = 1'b1;
    assign layer0_outputs[1171] = ~((inputs[143]) & (inputs[43]));
    assign layer0_outputs[1172] = inputs[77];
    assign layer0_outputs[1173] = ~(inputs[18]) | (inputs[97]);
    assign layer0_outputs[1174] = (inputs[147]) ^ (inputs[32]);
    assign layer0_outputs[1175] = ~((inputs[243]) ^ (inputs[115]));
    assign layer0_outputs[1176] = (inputs[239]) | (inputs[205]);
    assign layer0_outputs[1177] = ~(inputs[158]);
    assign layer0_outputs[1178] = (inputs[241]) ^ (inputs[217]);
    assign layer0_outputs[1179] = (inputs[241]) ^ (inputs[69]);
    assign layer0_outputs[1180] = (inputs[199]) & ~(inputs[189]);
    assign layer0_outputs[1181] = ~((inputs[201]) | (inputs[128]));
    assign layer0_outputs[1182] = ~(inputs[44]) | (inputs[110]);
    assign layer0_outputs[1183] = (inputs[127]) & ~(inputs[52]);
    assign layer0_outputs[1184] = ~(inputs[69]);
    assign layer0_outputs[1185] = (inputs[189]) | (inputs[36]);
    assign layer0_outputs[1186] = (inputs[198]) & ~(inputs[43]);
    assign layer0_outputs[1187] = ~(inputs[162]);
    assign layer0_outputs[1188] = ~((inputs[44]) ^ (inputs[190]));
    assign layer0_outputs[1189] = ~((inputs[38]) | (inputs[118]));
    assign layer0_outputs[1190] = ~(inputs[137]);
    assign layer0_outputs[1191] = ~((inputs[166]) ^ (inputs[97]));
    assign layer0_outputs[1192] = (inputs[117]) & ~(inputs[65]);
    assign layer0_outputs[1193] = ~(inputs[79]) | (inputs[238]);
    assign layer0_outputs[1194] = ~(inputs[153]);
    assign layer0_outputs[1195] = inputs[70];
    assign layer0_outputs[1196] = inputs[141];
    assign layer0_outputs[1197] = inputs[42];
    assign layer0_outputs[1198] = ~(inputs[87]);
    assign layer0_outputs[1199] = (inputs[82]) & ~(inputs[62]);
    assign layer0_outputs[1200] = (inputs[250]) ^ (inputs[68]);
    assign layer0_outputs[1201] = ~(inputs[166]) | (inputs[209]);
    assign layer0_outputs[1202] = 1'b0;
    assign layer0_outputs[1203] = ~(inputs[42]);
    assign layer0_outputs[1204] = ~((inputs[158]) ^ (inputs[81]));
    assign layer0_outputs[1205] = (inputs[146]) | (inputs[94]);
    assign layer0_outputs[1206] = (inputs[153]) & ~(inputs[103]);
    assign layer0_outputs[1207] = ~(inputs[117]);
    assign layer0_outputs[1208] = ~(inputs[168]) | (inputs[79]);
    assign layer0_outputs[1209] = ~(inputs[202]);
    assign layer0_outputs[1210] = ~(inputs[154]);
    assign layer0_outputs[1211] = (inputs[159]) | (inputs[151]);
    assign layer0_outputs[1212] = (inputs[182]) ^ (inputs[195]);
    assign layer0_outputs[1213] = 1'b1;
    assign layer0_outputs[1214] = (inputs[90]) & ~(inputs[26]);
    assign layer0_outputs[1215] = ~(inputs[187]) | (inputs[146]);
    assign layer0_outputs[1216] = (inputs[240]) ^ (inputs[237]);
    assign layer0_outputs[1217] = inputs[72];
    assign layer0_outputs[1218] = (inputs[183]) ^ (inputs[89]);
    assign layer0_outputs[1219] = ~(inputs[247]);
    assign layer0_outputs[1220] = (inputs[7]) & ~(inputs[239]);
    assign layer0_outputs[1221] = inputs[156];
    assign layer0_outputs[1222] = (inputs[137]) & ~(inputs[188]);
    assign layer0_outputs[1223] = inputs[103];
    assign layer0_outputs[1224] = ~(inputs[59]) | (inputs[210]);
    assign layer0_outputs[1225] = ~(inputs[77]) | (inputs[248]);
    assign layer0_outputs[1226] = ~(inputs[245]) | (inputs[95]);
    assign layer0_outputs[1227] = 1'b0;
    assign layer0_outputs[1228] = ~(inputs[56]);
    assign layer0_outputs[1229] = inputs[17];
    assign layer0_outputs[1230] = (inputs[73]) & ~(inputs[11]);
    assign layer0_outputs[1231] = ~(inputs[237]) | (inputs[67]);
    assign layer0_outputs[1232] = 1'b0;
    assign layer0_outputs[1233] = ~((inputs[44]) | (inputs[20]));
    assign layer0_outputs[1234] = (inputs[70]) | (inputs[208]);
    assign layer0_outputs[1235] = ~(inputs[26]) | (inputs[243]);
    assign layer0_outputs[1236] = ~((inputs[90]) ^ (inputs[253]));
    assign layer0_outputs[1237] = ~((inputs[234]) | (inputs[109]));
    assign layer0_outputs[1238] = ~((inputs[25]) ^ (inputs[122]));
    assign layer0_outputs[1239] = ~((inputs[31]) | (inputs[24]));
    assign layer0_outputs[1240] = ~(inputs[229]);
    assign layer0_outputs[1241] = (inputs[7]) & ~(inputs[145]);
    assign layer0_outputs[1242] = inputs[159];
    assign layer0_outputs[1243] = ~((inputs[201]) ^ (inputs[222]));
    assign layer0_outputs[1244] = ~((inputs[251]) ^ (inputs[25]));
    assign layer0_outputs[1245] = inputs[149];
    assign layer0_outputs[1246] = (inputs[197]) | (inputs[189]);
    assign layer0_outputs[1247] = (inputs[26]) & ~(inputs[245]);
    assign layer0_outputs[1248] = (inputs[113]) & ~(inputs[240]);
    assign layer0_outputs[1249] = inputs[82];
    assign layer0_outputs[1250] = inputs[253];
    assign layer0_outputs[1251] = inputs[167];
    assign layer0_outputs[1252] = ~(inputs[90]);
    assign layer0_outputs[1253] = ~(inputs[136]);
    assign layer0_outputs[1254] = inputs[121];
    assign layer0_outputs[1255] = inputs[144];
    assign layer0_outputs[1256] = ~((inputs[144]) ^ (inputs[53]));
    assign layer0_outputs[1257] = ~((inputs[36]) ^ (inputs[162]));
    assign layer0_outputs[1258] = ~(inputs[181]);
    assign layer0_outputs[1259] = ~(inputs[150]);
    assign layer0_outputs[1260] = inputs[87];
    assign layer0_outputs[1261] = ~(inputs[88]) | (inputs[148]);
    assign layer0_outputs[1262] = ~((inputs[72]) | (inputs[178]));
    assign layer0_outputs[1263] = (inputs[72]) & ~(inputs[53]);
    assign layer0_outputs[1264] = inputs[222];
    assign layer0_outputs[1265] = ~((inputs[218]) ^ (inputs[94]));
    assign layer0_outputs[1266] = (inputs[110]) | (inputs[58]);
    assign layer0_outputs[1267] = (inputs[63]) & ~(inputs[239]);
    assign layer0_outputs[1268] = ~(inputs[68]);
    assign layer0_outputs[1269] = 1'b0;
    assign layer0_outputs[1270] = (inputs[238]) & ~(inputs[177]);
    assign layer0_outputs[1271] = 1'b1;
    assign layer0_outputs[1272] = (inputs[11]) ^ (inputs[253]);
    assign layer0_outputs[1273] = (inputs[153]) & ~(inputs[119]);
    assign layer0_outputs[1274] = (inputs[34]) & ~(inputs[118]);
    assign layer0_outputs[1275] = ~((inputs[187]) | (inputs[215]));
    assign layer0_outputs[1276] = (inputs[154]) | (inputs[36]);
    assign layer0_outputs[1277] = ~(inputs[119]) | (inputs[131]);
    assign layer0_outputs[1278] = ~(inputs[113]);
    assign layer0_outputs[1279] = ~((inputs[224]) ^ (inputs[102]));
    assign layer0_outputs[1280] = ~(inputs[128]);
    assign layer0_outputs[1281] = inputs[182];
    assign layer0_outputs[1282] = ~(inputs[136]) | (inputs[29]);
    assign layer0_outputs[1283] = ~((inputs[144]) ^ (inputs[188]));
    assign layer0_outputs[1284] = (inputs[99]) | (inputs[217]);
    assign layer0_outputs[1285] = ~((inputs[82]) | (inputs[104]));
    assign layer0_outputs[1286] = ~(inputs[165]);
    assign layer0_outputs[1287] = (inputs[108]) | (inputs[25]);
    assign layer0_outputs[1288] = inputs[244];
    assign layer0_outputs[1289] = ~(inputs[159]);
    assign layer0_outputs[1290] = ~((inputs[72]) & (inputs[67]));
    assign layer0_outputs[1291] = ~((inputs[246]) ^ (inputs[74]));
    assign layer0_outputs[1292] = (inputs[217]) & (inputs[251]);
    assign layer0_outputs[1293] = (inputs[122]) & ~(inputs[251]);
    assign layer0_outputs[1294] = ~(inputs[133]);
    assign layer0_outputs[1295] = (inputs[38]) & ~(inputs[204]);
    assign layer0_outputs[1296] = ~(inputs[171]);
    assign layer0_outputs[1297] = ~((inputs[188]) | (inputs[194]));
    assign layer0_outputs[1298] = ~(inputs[224]) | (inputs[191]);
    assign layer0_outputs[1299] = (inputs[131]) & ~(inputs[49]);
    assign layer0_outputs[1300] = (inputs[153]) | (inputs[116]);
    assign layer0_outputs[1301] = ~((inputs[169]) ^ (inputs[128]));
    assign layer0_outputs[1302] = inputs[230];
    assign layer0_outputs[1303] = ~(inputs[198]) | (inputs[45]);
    assign layer0_outputs[1304] = (inputs[124]) & ~(inputs[145]);
    assign layer0_outputs[1305] = ~(inputs[91]);
    assign layer0_outputs[1306] = (inputs[231]) ^ (inputs[241]);
    assign layer0_outputs[1307] = ~(inputs[101]) | (inputs[126]);
    assign layer0_outputs[1308] = inputs[71];
    assign layer0_outputs[1309] = ~(inputs[194]);
    assign layer0_outputs[1310] = (inputs[43]) & ~(inputs[35]);
    assign layer0_outputs[1311] = ~((inputs[129]) ^ (inputs[106]));
    assign layer0_outputs[1312] = (inputs[166]) | (inputs[193]);
    assign layer0_outputs[1313] = ~(inputs[209]);
    assign layer0_outputs[1314] = inputs[90];
    assign layer0_outputs[1315] = ~(inputs[216]);
    assign layer0_outputs[1316] = ~((inputs[80]) & (inputs[13]));
    assign layer0_outputs[1317] = (inputs[210]) | (inputs[212]);
    assign layer0_outputs[1318] = (inputs[0]) & ~(inputs[111]);
    assign layer0_outputs[1319] = ~(inputs[197]) | (inputs[208]);
    assign layer0_outputs[1320] = ~((inputs[99]) ^ (inputs[241]));
    assign layer0_outputs[1321] = inputs[59];
    assign layer0_outputs[1322] = ~((inputs[97]) | (inputs[168]));
    assign layer0_outputs[1323] = ~(inputs[122]);
    assign layer0_outputs[1324] = inputs[152];
    assign layer0_outputs[1325] = ~(inputs[167]) | (inputs[108]);
    assign layer0_outputs[1326] = (inputs[60]) & ~(inputs[14]);
    assign layer0_outputs[1327] = 1'b1;
    assign layer0_outputs[1328] = ~((inputs[87]) ^ (inputs[85]));
    assign layer0_outputs[1329] = ~((inputs[147]) | (inputs[80]));
    assign layer0_outputs[1330] = (inputs[169]) & ~(inputs[78]);
    assign layer0_outputs[1331] = ~(inputs[251]) | (inputs[145]);
    assign layer0_outputs[1332] = inputs[151];
    assign layer0_outputs[1333] = (inputs[118]) & ~(inputs[163]);
    assign layer0_outputs[1334] = inputs[165];
    assign layer0_outputs[1335] = (inputs[189]) & ~(inputs[22]);
    assign layer0_outputs[1336] = (inputs[52]) | (inputs[4]);
    assign layer0_outputs[1337] = (inputs[81]) & (inputs[176]);
    assign layer0_outputs[1338] = inputs[197];
    assign layer0_outputs[1339] = ~((inputs[239]) | (inputs[34]));
    assign layer0_outputs[1340] = inputs[113];
    assign layer0_outputs[1341] = ~(inputs[149]);
    assign layer0_outputs[1342] = (inputs[205]) & ~(inputs[66]);
    assign layer0_outputs[1343] = inputs[159];
    assign layer0_outputs[1344] = ~(inputs[160]);
    assign layer0_outputs[1345] = (inputs[165]) & ~(inputs[238]);
    assign layer0_outputs[1346] = inputs[69];
    assign layer0_outputs[1347] = ~(inputs[101]);
    assign layer0_outputs[1348] = ~(inputs[104]);
    assign layer0_outputs[1349] = inputs[166];
    assign layer0_outputs[1350] = ~((inputs[21]) & (inputs[10]));
    assign layer0_outputs[1351] = 1'b1;
    assign layer0_outputs[1352] = ~(inputs[165]) | (inputs[234]);
    assign layer0_outputs[1353] = ~((inputs[137]) ^ (inputs[63]));
    assign layer0_outputs[1354] = (inputs[75]) ^ (inputs[242]);
    assign layer0_outputs[1355] = ~((inputs[4]) | (inputs[147]));
    assign layer0_outputs[1356] = ~(inputs[99]);
    assign layer0_outputs[1357] = (inputs[234]) & ~(inputs[48]);
    assign layer0_outputs[1358] = (inputs[131]) | (inputs[136]);
    assign layer0_outputs[1359] = ~((inputs[130]) ^ (inputs[81]));
    assign layer0_outputs[1360] = ~(inputs[110]) | (inputs[7]);
    assign layer0_outputs[1361] = ~((inputs[44]) ^ (inputs[181]));
    assign layer0_outputs[1362] = ~((inputs[221]) ^ (inputs[154]));
    assign layer0_outputs[1363] = ~((inputs[54]) | (inputs[172]));
    assign layer0_outputs[1364] = ~(inputs[7]) | (inputs[212]);
    assign layer0_outputs[1365] = inputs[39];
    assign layer0_outputs[1366] = (inputs[221]) & ~(inputs[85]);
    assign layer0_outputs[1367] = ~(inputs[73]) | (inputs[4]);
    assign layer0_outputs[1368] = (inputs[100]) & ~(inputs[194]);
    assign layer0_outputs[1369] = (inputs[149]) ^ (inputs[175]);
    assign layer0_outputs[1370] = (inputs[15]) & ~(inputs[234]);
    assign layer0_outputs[1371] = ~((inputs[39]) | (inputs[162]));
    assign layer0_outputs[1372] = (inputs[19]) | (inputs[123]);
    assign layer0_outputs[1373] = ~(inputs[125]) | (inputs[245]);
    assign layer0_outputs[1374] = ~((inputs[24]) | (inputs[210]));
    assign layer0_outputs[1375] = inputs[81];
    assign layer0_outputs[1376] = (inputs[44]) & (inputs[118]);
    assign layer0_outputs[1377] = ~((inputs[179]) ^ (inputs[238]));
    assign layer0_outputs[1378] = (inputs[108]) ^ (inputs[205]);
    assign layer0_outputs[1379] = 1'b1;
    assign layer0_outputs[1380] = (inputs[154]) ^ (inputs[106]);
    assign layer0_outputs[1381] = ~(inputs[51]) | (inputs[220]);
    assign layer0_outputs[1382] = ~((inputs[158]) ^ (inputs[249]));
    assign layer0_outputs[1383] = (inputs[126]) & ~(inputs[167]);
    assign layer0_outputs[1384] = (inputs[218]) | (inputs[79]);
    assign layer0_outputs[1385] = ~(inputs[254]);
    assign layer0_outputs[1386] = ~(inputs[211]) | (inputs[46]);
    assign layer0_outputs[1387] = (inputs[52]) ^ (inputs[149]);
    assign layer0_outputs[1388] = inputs[34];
    assign layer0_outputs[1389] = ~(inputs[213]) | (inputs[125]);
    assign layer0_outputs[1390] = ~(inputs[19]);
    assign layer0_outputs[1391] = ~((inputs[194]) | (inputs[15]));
    assign layer0_outputs[1392] = ~((inputs[21]) | (inputs[131]));
    assign layer0_outputs[1393] = inputs[137];
    assign layer0_outputs[1394] = ~(inputs[231]) | (inputs[163]);
    assign layer0_outputs[1395] = ~(inputs[21]);
    assign layer0_outputs[1396] = (inputs[247]) & (inputs[175]);
    assign layer0_outputs[1397] = ~((inputs[252]) | (inputs[225]));
    assign layer0_outputs[1398] = ~((inputs[248]) ^ (inputs[57]));
    assign layer0_outputs[1399] = ~((inputs[56]) | (inputs[231]));
    assign layer0_outputs[1400] = inputs[179];
    assign layer0_outputs[1401] = ~(inputs[152]);
    assign layer0_outputs[1402] = inputs[189];
    assign layer0_outputs[1403] = 1'b1;
    assign layer0_outputs[1404] = (inputs[253]) | (inputs[91]);
    assign layer0_outputs[1405] = (inputs[16]) & (inputs[130]);
    assign layer0_outputs[1406] = ~((inputs[246]) ^ (inputs[41]));
    assign layer0_outputs[1407] = (inputs[82]) & ~(inputs[115]);
    assign layer0_outputs[1408] = (inputs[28]) & ~(inputs[112]);
    assign layer0_outputs[1409] = (inputs[193]) ^ (inputs[208]);
    assign layer0_outputs[1410] = inputs[182];
    assign layer0_outputs[1411] = ~((inputs[92]) | (inputs[126]));
    assign layer0_outputs[1412] = ~((inputs[2]) | (inputs[59]));
    assign layer0_outputs[1413] = 1'b1;
    assign layer0_outputs[1414] = (inputs[216]) | (inputs[128]);
    assign layer0_outputs[1415] = inputs[186];
    assign layer0_outputs[1416] = 1'b1;
    assign layer0_outputs[1417] = ~((inputs[71]) ^ (inputs[95]));
    assign layer0_outputs[1418] = (inputs[174]) & ~(inputs[244]);
    assign layer0_outputs[1419] = (inputs[172]) & ~(inputs[14]);
    assign layer0_outputs[1420] = (inputs[198]) | (inputs[213]);
    assign layer0_outputs[1421] = (inputs[186]) | (inputs[243]);
    assign layer0_outputs[1422] = ~((inputs[229]) ^ (inputs[210]));
    assign layer0_outputs[1423] = ~(inputs[129]);
    assign layer0_outputs[1424] = ~(inputs[42]);
    assign layer0_outputs[1425] = ~(inputs[198]);
    assign layer0_outputs[1426] = ~((inputs[247]) | (inputs[182]));
    assign layer0_outputs[1427] = ~(inputs[216]) | (inputs[26]);
    assign layer0_outputs[1428] = (inputs[89]) & ~(inputs[9]);
    assign layer0_outputs[1429] = (inputs[87]) & ~(inputs[236]);
    assign layer0_outputs[1430] = inputs[54];
    assign layer0_outputs[1431] = ~(inputs[132]);
    assign layer0_outputs[1432] = inputs[203];
    assign layer0_outputs[1433] = (inputs[120]) & ~(inputs[82]);
    assign layer0_outputs[1434] = (inputs[141]) & ~(inputs[6]);
    assign layer0_outputs[1435] = ~(inputs[102]) | (inputs[210]);
    assign layer0_outputs[1436] = ~((inputs[126]) ^ (inputs[176]));
    assign layer0_outputs[1437] = (inputs[75]) & (inputs[16]);
    assign layer0_outputs[1438] = ~((inputs[110]) | (inputs[237]));
    assign layer0_outputs[1439] = (inputs[138]) | (inputs[122]);
    assign layer0_outputs[1440] = (inputs[104]) | (inputs[234]);
    assign layer0_outputs[1441] = inputs[10];
    assign layer0_outputs[1442] = ~((inputs[117]) ^ (inputs[236]));
    assign layer0_outputs[1443] = ~(inputs[131]);
    assign layer0_outputs[1444] = (inputs[145]) | (inputs[8]);
    assign layer0_outputs[1445] = ~((inputs[169]) & (inputs[172]));
    assign layer0_outputs[1446] = (inputs[42]) | (inputs[206]);
    assign layer0_outputs[1447] = inputs[182];
    assign layer0_outputs[1448] = inputs[72];
    assign layer0_outputs[1449] = 1'b0;
    assign layer0_outputs[1450] = (inputs[133]) & ~(inputs[16]);
    assign layer0_outputs[1451] = (inputs[192]) ^ (inputs[74]);
    assign layer0_outputs[1452] = inputs[33];
    assign layer0_outputs[1453] = (inputs[4]) | (inputs[44]);
    assign layer0_outputs[1454] = 1'b0;
    assign layer0_outputs[1455] = (inputs[191]) | (inputs[52]);
    assign layer0_outputs[1456] = ~((inputs[162]) ^ (inputs[168]));
    assign layer0_outputs[1457] = ~(inputs[223]);
    assign layer0_outputs[1458] = (inputs[196]) | (inputs[188]);
    assign layer0_outputs[1459] = ~(inputs[47]) | (inputs[234]);
    assign layer0_outputs[1460] = inputs[82];
    assign layer0_outputs[1461] = (inputs[131]) ^ (inputs[68]);
    assign layer0_outputs[1462] = (inputs[247]) ^ (inputs[83]);
    assign layer0_outputs[1463] = (inputs[230]) & ~(inputs[93]);
    assign layer0_outputs[1464] = ~((inputs[215]) | (inputs[73]));
    assign layer0_outputs[1465] = (inputs[214]) & ~(inputs[147]);
    assign layer0_outputs[1466] = (inputs[209]) ^ (inputs[26]);
    assign layer0_outputs[1467] = (inputs[172]) | (inputs[69]);
    assign layer0_outputs[1468] = 1'b1;
    assign layer0_outputs[1469] = (inputs[195]) & ~(inputs[81]);
    assign layer0_outputs[1470] = ~(inputs[54]);
    assign layer0_outputs[1471] = (inputs[180]) | (inputs[125]);
    assign layer0_outputs[1472] = inputs[124];
    assign layer0_outputs[1473] = (inputs[145]) ^ (inputs[109]);
    assign layer0_outputs[1474] = (inputs[7]) ^ (inputs[116]);
    assign layer0_outputs[1475] = (inputs[79]) | (inputs[71]);
    assign layer0_outputs[1476] = inputs[138];
    assign layer0_outputs[1477] = (inputs[236]) & ~(inputs[206]);
    assign layer0_outputs[1478] = ~(inputs[124]);
    assign layer0_outputs[1479] = (inputs[229]) | (inputs[53]);
    assign layer0_outputs[1480] = inputs[135];
    assign layer0_outputs[1481] = ~((inputs[222]) ^ (inputs[126]));
    assign layer0_outputs[1482] = (inputs[9]) | (inputs[166]);
    assign layer0_outputs[1483] = (inputs[124]) | (inputs[135]);
    assign layer0_outputs[1484] = (inputs[96]) ^ (inputs[118]);
    assign layer0_outputs[1485] = ~(inputs[108]);
    assign layer0_outputs[1486] = (inputs[186]) | (inputs[186]);
    assign layer0_outputs[1487] = (inputs[114]) | (inputs[250]);
    assign layer0_outputs[1488] = (inputs[131]) & ~(inputs[31]);
    assign layer0_outputs[1489] = ~((inputs[170]) | (inputs[228]));
    assign layer0_outputs[1490] = ~((inputs[40]) | (inputs[57]));
    assign layer0_outputs[1491] = ~(inputs[202]) | (inputs[225]);
    assign layer0_outputs[1492] = inputs[138];
    assign layer0_outputs[1493] = inputs[246];
    assign layer0_outputs[1494] = (inputs[177]) & (inputs[209]);
    assign layer0_outputs[1495] = ~(inputs[220]) | (inputs[135]);
    assign layer0_outputs[1496] = (inputs[142]) | (inputs[91]);
    assign layer0_outputs[1497] = inputs[120];
    assign layer0_outputs[1498] = ~(inputs[136]) | (inputs[44]);
    assign layer0_outputs[1499] = ~(inputs[87]) | (inputs[29]);
    assign layer0_outputs[1500] = (inputs[147]) ^ (inputs[9]);
    assign layer0_outputs[1501] = ~(inputs[216]) | (inputs[225]);
    assign layer0_outputs[1502] = ~((inputs[72]) ^ (inputs[211]));
    assign layer0_outputs[1503] = (inputs[129]) ^ (inputs[187]);
    assign layer0_outputs[1504] = inputs[215];
    assign layer0_outputs[1505] = inputs[99];
    assign layer0_outputs[1506] = (inputs[5]) & ~(inputs[72]);
    assign layer0_outputs[1507] = ~(inputs[151]);
    assign layer0_outputs[1508] = ~(inputs[105]);
    assign layer0_outputs[1509] = inputs[50];
    assign layer0_outputs[1510] = ~((inputs[174]) | (inputs[164]));
    assign layer0_outputs[1511] = inputs[118];
    assign layer0_outputs[1512] = (inputs[47]) & ~(inputs[216]);
    assign layer0_outputs[1513] = ~((inputs[177]) ^ (inputs[231]));
    assign layer0_outputs[1514] = ~(inputs[59]) | (inputs[255]);
    assign layer0_outputs[1515] = ~((inputs[89]) ^ (inputs[31]));
    assign layer0_outputs[1516] = 1'b0;
    assign layer0_outputs[1517] = inputs[100];
    assign layer0_outputs[1518] = ~(inputs[143]);
    assign layer0_outputs[1519] = ~((inputs[6]) ^ (inputs[71]));
    assign layer0_outputs[1520] = inputs[119];
    assign layer0_outputs[1521] = ~((inputs[239]) ^ (inputs[11]));
    assign layer0_outputs[1522] = ~(inputs[181]) | (inputs[33]);
    assign layer0_outputs[1523] = ~(inputs[148]) | (inputs[223]);
    assign layer0_outputs[1524] = ~(inputs[116]);
    assign layer0_outputs[1525] = 1'b1;
    assign layer0_outputs[1526] = (inputs[86]) & (inputs[201]);
    assign layer0_outputs[1527] = ~(inputs[22]);
    assign layer0_outputs[1528] = (inputs[31]) ^ (inputs[96]);
    assign layer0_outputs[1529] = ~((inputs[85]) & (inputs[143]));
    assign layer0_outputs[1530] = inputs[107];
    assign layer0_outputs[1531] = ~(inputs[53]) | (inputs[157]);
    assign layer0_outputs[1532] = inputs[90];
    assign layer0_outputs[1533] = ~(inputs[155]) | (inputs[179]);
    assign layer0_outputs[1534] = 1'b0;
    assign layer0_outputs[1535] = (inputs[174]) & ~(inputs[100]);
    assign layer0_outputs[1536] = (inputs[143]) ^ (inputs[25]);
    assign layer0_outputs[1537] = inputs[172];
    assign layer0_outputs[1538] = ~(inputs[20]);
    assign layer0_outputs[1539] = ~(inputs[190]);
    assign layer0_outputs[1540] = ~((inputs[171]) ^ (inputs[62]));
    assign layer0_outputs[1541] = ~((inputs[114]) | (inputs[232]));
    assign layer0_outputs[1542] = (inputs[102]) & ~(inputs[146]);
    assign layer0_outputs[1543] = ~((inputs[129]) | (inputs[103]));
    assign layer0_outputs[1544] = ~(inputs[100]) | (inputs[141]);
    assign layer0_outputs[1545] = (inputs[191]) ^ (inputs[70]);
    assign layer0_outputs[1546] = ~((inputs[128]) | (inputs[109]));
    assign layer0_outputs[1547] = ~(inputs[27]);
    assign layer0_outputs[1548] = (inputs[105]) & ~(inputs[9]);
    assign layer0_outputs[1549] = ~((inputs[216]) | (inputs[185]));
    assign layer0_outputs[1550] = ~((inputs[183]) ^ (inputs[214]));
    assign layer0_outputs[1551] = ~(inputs[104]);
    assign layer0_outputs[1552] = (inputs[207]) ^ (inputs[143]);
    assign layer0_outputs[1553] = ~(inputs[82]);
    assign layer0_outputs[1554] = ~((inputs[25]) | (inputs[53]));
    assign layer0_outputs[1555] = ~(inputs[102]);
    assign layer0_outputs[1556] = ~((inputs[96]) | (inputs[50]));
    assign layer0_outputs[1557] = ~((inputs[161]) ^ (inputs[124]));
    assign layer0_outputs[1558] = ~((inputs[48]) ^ (inputs[115]));
    assign layer0_outputs[1559] = ~(inputs[183]);
    assign layer0_outputs[1560] = ~((inputs[144]) & (inputs[5]));
    assign layer0_outputs[1561] = ~((inputs[145]) | (inputs[150]));
    assign layer0_outputs[1562] = inputs[187];
    assign layer0_outputs[1563] = ~(inputs[56]) | (inputs[100]);
    assign layer0_outputs[1564] = ~((inputs[62]) | (inputs[33]));
    assign layer0_outputs[1565] = ~(inputs[183]) | (inputs[134]);
    assign layer0_outputs[1566] = ~((inputs[83]) | (inputs[150]));
    assign layer0_outputs[1567] = (inputs[106]) & ~(inputs[249]);
    assign layer0_outputs[1568] = ~(inputs[211]) | (inputs[114]);
    assign layer0_outputs[1569] = inputs[156];
    assign layer0_outputs[1570] = ~((inputs[179]) | (inputs[6]));
    assign layer0_outputs[1571] = (inputs[162]) | (inputs[229]);
    assign layer0_outputs[1572] = 1'b0;
    assign layer0_outputs[1573] = ~((inputs[222]) & (inputs[43]));
    assign layer0_outputs[1574] = (inputs[177]) ^ (inputs[73]);
    assign layer0_outputs[1575] = (inputs[131]) | (inputs[14]);
    assign layer0_outputs[1576] = (inputs[226]) | (inputs[197]);
    assign layer0_outputs[1577] = inputs[69];
    assign layer0_outputs[1578] = (inputs[197]) | (inputs[195]);
    assign layer0_outputs[1579] = (inputs[167]) & ~(inputs[132]);
    assign layer0_outputs[1580] = ~((inputs[56]) | (inputs[125]));
    assign layer0_outputs[1581] = (inputs[238]) & ~(inputs[144]);
    assign layer0_outputs[1582] = inputs[91];
    assign layer0_outputs[1583] = (inputs[74]) ^ (inputs[126]);
    assign layer0_outputs[1584] = ~(inputs[196]);
    assign layer0_outputs[1585] = (inputs[104]) | (inputs[232]);
    assign layer0_outputs[1586] = 1'b1;
    assign layer0_outputs[1587] = ~((inputs[90]) | (inputs[146]));
    assign layer0_outputs[1588] = ~(inputs[116]) | (inputs[128]);
    assign layer0_outputs[1589] = (inputs[32]) ^ (inputs[40]);
    assign layer0_outputs[1590] = (inputs[120]) & ~(inputs[132]);
    assign layer0_outputs[1591] = (inputs[4]) & ~(inputs[33]);
    assign layer0_outputs[1592] = ~(inputs[169]);
    assign layer0_outputs[1593] = inputs[111];
    assign layer0_outputs[1594] = (inputs[209]) & (inputs[18]);
    assign layer0_outputs[1595] = ~(inputs[41]);
    assign layer0_outputs[1596] = ~((inputs[69]) | (inputs[24]));
    assign layer0_outputs[1597] = (inputs[132]) | (inputs[26]);
    assign layer0_outputs[1598] = 1'b1;
    assign layer0_outputs[1599] = (inputs[249]) & ~(inputs[23]);
    assign layer0_outputs[1600] = ~((inputs[93]) ^ (inputs[16]));
    assign layer0_outputs[1601] = ~((inputs[46]) ^ (inputs[171]));
    assign layer0_outputs[1602] = ~(inputs[182]);
    assign layer0_outputs[1603] = ~(inputs[151]) | (inputs[52]);
    assign layer0_outputs[1604] = (inputs[117]) ^ (inputs[97]);
    assign layer0_outputs[1605] = (inputs[30]) ^ (inputs[74]);
    assign layer0_outputs[1606] = ~((inputs[233]) | (inputs[109]));
    assign layer0_outputs[1607] = ~(inputs[228]);
    assign layer0_outputs[1608] = ~(inputs[149]);
    assign layer0_outputs[1609] = (inputs[178]) & ~(inputs[189]);
    assign layer0_outputs[1610] = ~((inputs[10]) ^ (inputs[63]));
    assign layer0_outputs[1611] = (inputs[117]) & ~(inputs[57]);
    assign layer0_outputs[1612] = (inputs[136]) | (inputs[233]);
    assign layer0_outputs[1613] = (inputs[109]) ^ (inputs[17]);
    assign layer0_outputs[1614] = ~(inputs[165]);
    assign layer0_outputs[1615] = ~(inputs[180]) | (inputs[39]);
    assign layer0_outputs[1616] = ~((inputs[5]) & (inputs[211]));
    assign layer0_outputs[1617] = (inputs[218]) & ~(inputs[171]);
    assign layer0_outputs[1618] = ~((inputs[178]) | (inputs[72]));
    assign layer0_outputs[1619] = inputs[206];
    assign layer0_outputs[1620] = ~((inputs[237]) & (inputs[30]));
    assign layer0_outputs[1621] = ~(inputs[28]) | (inputs[208]);
    assign layer0_outputs[1622] = (inputs[133]) & ~(inputs[58]);
    assign layer0_outputs[1623] = ~(inputs[0]);
    assign layer0_outputs[1624] = (inputs[196]) ^ (inputs[254]);
    assign layer0_outputs[1625] = inputs[53];
    assign layer0_outputs[1626] = ~(inputs[46]);
    assign layer0_outputs[1627] = (inputs[216]) & ~(inputs[208]);
    assign layer0_outputs[1628] = ~((inputs[132]) ^ (inputs[12]));
    assign layer0_outputs[1629] = ~(inputs[213]);
    assign layer0_outputs[1630] = ~(inputs[119]);
    assign layer0_outputs[1631] = (inputs[193]) & (inputs[96]);
    assign layer0_outputs[1632] = (inputs[82]) & ~(inputs[157]);
    assign layer0_outputs[1633] = ~((inputs[78]) | (inputs[229]));
    assign layer0_outputs[1634] = (inputs[131]) & ~(inputs[119]);
    assign layer0_outputs[1635] = (inputs[232]) & ~(inputs[126]);
    assign layer0_outputs[1636] = ~(inputs[132]);
    assign layer0_outputs[1637] = ~(inputs[92]) | (inputs[161]);
    assign layer0_outputs[1638] = (inputs[87]) ^ (inputs[130]);
    assign layer0_outputs[1639] = (inputs[151]) & ~(inputs[229]);
    assign layer0_outputs[1640] = (inputs[194]) ^ (inputs[110]);
    assign layer0_outputs[1641] = (inputs[101]) & ~(inputs[178]);
    assign layer0_outputs[1642] = ~(inputs[180]) | (inputs[159]);
    assign layer0_outputs[1643] = inputs[184];
    assign layer0_outputs[1644] = (inputs[75]) & ~(inputs[153]);
    assign layer0_outputs[1645] = ~(inputs[240]);
    assign layer0_outputs[1646] = ~((inputs[235]) | (inputs[200]));
    assign layer0_outputs[1647] = (inputs[4]) & ~(inputs[37]);
    assign layer0_outputs[1648] = (inputs[141]) & ~(inputs[212]);
    assign layer0_outputs[1649] = (inputs[104]) | (inputs[163]);
    assign layer0_outputs[1650] = ~((inputs[34]) | (inputs[120]));
    assign layer0_outputs[1651] = (inputs[86]) | (inputs[140]);
    assign layer0_outputs[1652] = ~(inputs[248]);
    assign layer0_outputs[1653] = inputs[138];
    assign layer0_outputs[1654] = ~((inputs[39]) ^ (inputs[29]));
    assign layer0_outputs[1655] = (inputs[178]) & ~(inputs[63]);
    assign layer0_outputs[1656] = (inputs[149]) | (inputs[252]);
    assign layer0_outputs[1657] = (inputs[1]) | (inputs[41]);
    assign layer0_outputs[1658] = ~(inputs[205]);
    assign layer0_outputs[1659] = inputs[214];
    assign layer0_outputs[1660] = inputs[130];
    assign layer0_outputs[1661] = ~((inputs[19]) | (inputs[104]));
    assign layer0_outputs[1662] = (inputs[139]) ^ (inputs[44]);
    assign layer0_outputs[1663] = (inputs[131]) & ~(inputs[252]);
    assign layer0_outputs[1664] = inputs[34];
    assign layer0_outputs[1665] = (inputs[124]) | (inputs[74]);
    assign layer0_outputs[1666] = (inputs[164]) | (inputs[44]);
    assign layer0_outputs[1667] = (inputs[209]) & ~(inputs[85]);
    assign layer0_outputs[1668] = ~(inputs[155]) | (inputs[0]);
    assign layer0_outputs[1669] = 1'b1;
    assign layer0_outputs[1670] = (inputs[55]) & ~(inputs[22]);
    assign layer0_outputs[1671] = (inputs[181]) ^ (inputs[158]);
    assign layer0_outputs[1672] = ~(inputs[215]) | (inputs[245]);
    assign layer0_outputs[1673] = ~((inputs[23]) ^ (inputs[144]));
    assign layer0_outputs[1674] = (inputs[135]) & ~(inputs[65]);
    assign layer0_outputs[1675] = ~(inputs[107]);
    assign layer0_outputs[1676] = ~(inputs[212]) | (inputs[14]);
    assign layer0_outputs[1677] = 1'b1;
    assign layer0_outputs[1678] = ~((inputs[85]) | (inputs[142]));
    assign layer0_outputs[1679] = ~(inputs[126]);
    assign layer0_outputs[1680] = ~(inputs[73]) | (inputs[243]);
    assign layer0_outputs[1681] = ~((inputs[69]) & (inputs[87]));
    assign layer0_outputs[1682] = ~((inputs[181]) | (inputs[53]));
    assign layer0_outputs[1683] = ~(inputs[234]) | (inputs[74]);
    assign layer0_outputs[1684] = ~(inputs[135]) | (inputs[38]);
    assign layer0_outputs[1685] = (inputs[59]) ^ (inputs[103]);
    assign layer0_outputs[1686] = (inputs[122]) & (inputs[73]);
    assign layer0_outputs[1687] = ~(inputs[68]);
    assign layer0_outputs[1688] = ~((inputs[123]) | (inputs[153]));
    assign layer0_outputs[1689] = inputs[142];
    assign layer0_outputs[1690] = (inputs[229]) ^ (inputs[25]);
    assign layer0_outputs[1691] = (inputs[217]) & ~(inputs[80]);
    assign layer0_outputs[1692] = (inputs[107]) & ~(inputs[0]);
    assign layer0_outputs[1693] = ~((inputs[173]) | (inputs[239]));
    assign layer0_outputs[1694] = 1'b0;
    assign layer0_outputs[1695] = (inputs[183]) ^ (inputs[16]);
    assign layer0_outputs[1696] = (inputs[125]) & ~(inputs[242]);
    assign layer0_outputs[1697] = (inputs[239]) | (inputs[209]);
    assign layer0_outputs[1698] = ~((inputs[127]) ^ (inputs[221]));
    assign layer0_outputs[1699] = ~(inputs[134]);
    assign layer0_outputs[1700] = ~((inputs[56]) ^ (inputs[63]));
    assign layer0_outputs[1701] = 1'b1;
    assign layer0_outputs[1702] = ~(inputs[91]);
    assign layer0_outputs[1703] = ~((inputs[139]) | (inputs[50]));
    assign layer0_outputs[1704] = (inputs[157]) & ~(inputs[129]);
    assign layer0_outputs[1705] = 1'b0;
    assign layer0_outputs[1706] = ~((inputs[26]) | (inputs[214]));
    assign layer0_outputs[1707] = (inputs[43]) & ~(inputs[62]);
    assign layer0_outputs[1708] = (inputs[200]) | (inputs[230]);
    assign layer0_outputs[1709] = ~((inputs[25]) | (inputs[107]));
    assign layer0_outputs[1710] = ~(inputs[179]);
    assign layer0_outputs[1711] = (inputs[234]) & ~(inputs[94]);
    assign layer0_outputs[1712] = ~(inputs[37]);
    assign layer0_outputs[1713] = ~(inputs[255]) | (inputs[255]);
    assign layer0_outputs[1714] = inputs[76];
    assign layer0_outputs[1715] = ~((inputs[244]) ^ (inputs[238]));
    assign layer0_outputs[1716] = ~((inputs[182]) | (inputs[21]));
    assign layer0_outputs[1717] = inputs[133];
    assign layer0_outputs[1718] = ~(inputs[205]) | (inputs[18]);
    assign layer0_outputs[1719] = 1'b0;
    assign layer0_outputs[1720] = ~(inputs[39]);
    assign layer0_outputs[1721] = inputs[167];
    assign layer0_outputs[1722] = ~((inputs[41]) | (inputs[140]));
    assign layer0_outputs[1723] = (inputs[218]) | (inputs[235]);
    assign layer0_outputs[1724] = 1'b1;
    assign layer0_outputs[1725] = inputs[94];
    assign layer0_outputs[1726] = ~(inputs[103]) | (inputs[2]);
    assign layer0_outputs[1727] = (inputs[138]) ^ (inputs[246]);
    assign layer0_outputs[1728] = inputs[191];
    assign layer0_outputs[1729] = ~((inputs[111]) | (inputs[179]));
    assign layer0_outputs[1730] = ~((inputs[6]) ^ (inputs[124]));
    assign layer0_outputs[1731] = ~((inputs[255]) | (inputs[97]));
    assign layer0_outputs[1732] = ~(inputs[213]);
    assign layer0_outputs[1733] = inputs[42];
    assign layer0_outputs[1734] = ~(inputs[102]) | (inputs[192]);
    assign layer0_outputs[1735] = (inputs[120]) & ~(inputs[239]);
    assign layer0_outputs[1736] = (inputs[242]) | (inputs[78]);
    assign layer0_outputs[1737] = 1'b0;
    assign layer0_outputs[1738] = (inputs[180]) & ~(inputs[248]);
    assign layer0_outputs[1739] = ~(inputs[173]);
    assign layer0_outputs[1740] = (inputs[100]) & ~(inputs[27]);
    assign layer0_outputs[1741] = (inputs[62]) & ~(inputs[65]);
    assign layer0_outputs[1742] = (inputs[121]) & ~(inputs[190]);
    assign layer0_outputs[1743] = (inputs[46]) & ~(inputs[89]);
    assign layer0_outputs[1744] = ~(inputs[85]) | (inputs[32]);
    assign layer0_outputs[1745] = ~(inputs[69]) | (inputs[43]);
    assign layer0_outputs[1746] = ~(inputs[179]) | (inputs[142]);
    assign layer0_outputs[1747] = ~(inputs[249]) | (inputs[47]);
    assign layer0_outputs[1748] = inputs[203];
    assign layer0_outputs[1749] = (inputs[47]) & (inputs[244]);
    assign layer0_outputs[1750] = (inputs[110]) & ~(inputs[96]);
    assign layer0_outputs[1751] = ~((inputs[74]) | (inputs[13]));
    assign layer0_outputs[1752] = ~((inputs[203]) | (inputs[23]));
    assign layer0_outputs[1753] = ~(inputs[61]) | (inputs[174]);
    assign layer0_outputs[1754] = (inputs[83]) ^ (inputs[32]);
    assign layer0_outputs[1755] = inputs[154];
    assign layer0_outputs[1756] = (inputs[49]) | (inputs[191]);
    assign layer0_outputs[1757] = ~(inputs[118]) | (inputs[190]);
    assign layer0_outputs[1758] = inputs[85];
    assign layer0_outputs[1759] = ~((inputs[104]) ^ (inputs[253]));
    assign layer0_outputs[1760] = (inputs[150]) & ~(inputs[93]);
    assign layer0_outputs[1761] = (inputs[39]) | (inputs[54]);
    assign layer0_outputs[1762] = (inputs[228]) | (inputs[105]);
    assign layer0_outputs[1763] = inputs[137];
    assign layer0_outputs[1764] = (inputs[188]) & ~(inputs[129]);
    assign layer0_outputs[1765] = ~(inputs[27]) | (inputs[208]);
    assign layer0_outputs[1766] = (inputs[34]) | (inputs[190]);
    assign layer0_outputs[1767] = ~((inputs[252]) ^ (inputs[222]));
    assign layer0_outputs[1768] = ~(inputs[254]) | (inputs[51]);
    assign layer0_outputs[1769] = ~((inputs[10]) ^ (inputs[22]));
    assign layer0_outputs[1770] = ~((inputs[121]) | (inputs[85]));
    assign layer0_outputs[1771] = (inputs[23]) & ~(inputs[227]);
    assign layer0_outputs[1772] = (inputs[175]) & (inputs[70]);
    assign layer0_outputs[1773] = (inputs[201]) & ~(inputs[131]);
    assign layer0_outputs[1774] = ~(inputs[157]) | (inputs[128]);
    assign layer0_outputs[1775] = (inputs[68]) | (inputs[54]);
    assign layer0_outputs[1776] = ~((inputs[6]) ^ (inputs[208]));
    assign layer0_outputs[1777] = (inputs[127]) | (inputs[23]);
    assign layer0_outputs[1778] = 1'b0;
    assign layer0_outputs[1779] = ~(inputs[163]);
    assign layer0_outputs[1780] = inputs[9];
    assign layer0_outputs[1781] = ~(inputs[181]) | (inputs[208]);
    assign layer0_outputs[1782] = ~(inputs[23]);
    assign layer0_outputs[1783] = (inputs[61]) & (inputs[15]);
    assign layer0_outputs[1784] = ~((inputs[80]) ^ (inputs[155]));
    assign layer0_outputs[1785] = ~(inputs[182]);
    assign layer0_outputs[1786] = inputs[151];
    assign layer0_outputs[1787] = inputs[135];
    assign layer0_outputs[1788] = ~((inputs[87]) ^ (inputs[5]));
    assign layer0_outputs[1789] = ~((inputs[62]) | (inputs[220]));
    assign layer0_outputs[1790] = ~(inputs[212]);
    assign layer0_outputs[1791] = ~((inputs[236]) | (inputs[30]));
    assign layer0_outputs[1792] = ~((inputs[42]) | (inputs[172]));
    assign layer0_outputs[1793] = inputs[206];
    assign layer0_outputs[1794] = ~(inputs[220]) | (inputs[161]);
    assign layer0_outputs[1795] = (inputs[6]) & ~(inputs[184]);
    assign layer0_outputs[1796] = ~(inputs[106]);
    assign layer0_outputs[1797] = (inputs[18]) ^ (inputs[32]);
    assign layer0_outputs[1798] = (inputs[121]) & ~(inputs[53]);
    assign layer0_outputs[1799] = ~(inputs[239]);
    assign layer0_outputs[1800] = inputs[157];
    assign layer0_outputs[1801] = ~(inputs[138]) | (inputs[19]);
    assign layer0_outputs[1802] = (inputs[13]) & ~(inputs[62]);
    assign layer0_outputs[1803] = ~((inputs[16]) ^ (inputs[68]));
    assign layer0_outputs[1804] = (inputs[233]) ^ (inputs[19]);
    assign layer0_outputs[1805] = ~((inputs[132]) ^ (inputs[12]));
    assign layer0_outputs[1806] = (inputs[54]) | (inputs[170]);
    assign layer0_outputs[1807] = ~(inputs[101]) | (inputs[226]);
    assign layer0_outputs[1808] = (inputs[87]) & ~(inputs[156]);
    assign layer0_outputs[1809] = (inputs[30]) & ~(inputs[187]);
    assign layer0_outputs[1810] = ~((inputs[184]) | (inputs[232]));
    assign layer0_outputs[1811] = (inputs[202]) ^ (inputs[218]);
    assign layer0_outputs[1812] = ~(inputs[91]);
    assign layer0_outputs[1813] = ~((inputs[255]) & (inputs[46]));
    assign layer0_outputs[1814] = ~(inputs[85]);
    assign layer0_outputs[1815] = (inputs[58]) & ~(inputs[252]);
    assign layer0_outputs[1816] = ~(inputs[157]);
    assign layer0_outputs[1817] = (inputs[137]) & ~(inputs[204]);
    assign layer0_outputs[1818] = (inputs[169]) & ~(inputs[47]);
    assign layer0_outputs[1819] = ~((inputs[152]) | (inputs[126]));
    assign layer0_outputs[1820] = (inputs[196]) & ~(inputs[232]);
    assign layer0_outputs[1821] = inputs[39];
    assign layer0_outputs[1822] = ~(inputs[210]) | (inputs[35]);
    assign layer0_outputs[1823] = inputs[3];
    assign layer0_outputs[1824] = (inputs[219]) | (inputs[163]);
    assign layer0_outputs[1825] = ~(inputs[171]) | (inputs[208]);
    assign layer0_outputs[1826] = (inputs[83]) | (inputs[98]);
    assign layer0_outputs[1827] = (inputs[170]) & ~(inputs[159]);
    assign layer0_outputs[1828] = inputs[255];
    assign layer0_outputs[1829] = inputs[64];
    assign layer0_outputs[1830] = inputs[194];
    assign layer0_outputs[1831] = (inputs[175]) ^ (inputs[163]);
    assign layer0_outputs[1832] = 1'b1;
    assign layer0_outputs[1833] = ~(inputs[168]);
    assign layer0_outputs[1834] = (inputs[28]) | (inputs[1]);
    assign layer0_outputs[1835] = (inputs[78]) | (inputs[209]);
    assign layer0_outputs[1836] = ~(inputs[251]);
    assign layer0_outputs[1837] = ~(inputs[185]) | (inputs[145]);
    assign layer0_outputs[1838] = ~(inputs[219]);
    assign layer0_outputs[1839] = ~((inputs[113]) | (inputs[97]));
    assign layer0_outputs[1840] = ~((inputs[244]) ^ (inputs[109]));
    assign layer0_outputs[1841] = (inputs[218]) | (inputs[55]);
    assign layer0_outputs[1842] = ~(inputs[221]) | (inputs[9]);
    assign layer0_outputs[1843] = ~(inputs[187]) | (inputs[125]);
    assign layer0_outputs[1844] = ~((inputs[170]) ^ (inputs[204]));
    assign layer0_outputs[1845] = inputs[172];
    assign layer0_outputs[1846] = (inputs[155]) & ~(inputs[249]);
    assign layer0_outputs[1847] = ~((inputs[212]) ^ (inputs[56]));
    assign layer0_outputs[1848] = (inputs[63]) & ~(inputs[91]);
    assign layer0_outputs[1849] = ~(inputs[54]) | (inputs[115]);
    assign layer0_outputs[1850] = ~((inputs[90]) | (inputs[206]));
    assign layer0_outputs[1851] = 1'b1;
    assign layer0_outputs[1852] = ~(inputs[102]) | (inputs[207]);
    assign layer0_outputs[1853] = ~(inputs[254]) | (inputs[45]);
    assign layer0_outputs[1854] = ~((inputs[250]) & (inputs[84]));
    assign layer0_outputs[1855] = ~(inputs[88]) | (inputs[126]);
    assign layer0_outputs[1856] = (inputs[76]) | (inputs[200]);
    assign layer0_outputs[1857] = ~((inputs[161]) | (inputs[67]));
    assign layer0_outputs[1858] = ~((inputs[114]) ^ (inputs[145]));
    assign layer0_outputs[1859] = (inputs[156]) ^ (inputs[78]);
    assign layer0_outputs[1860] = ~(inputs[230]);
    assign layer0_outputs[1861] = ~((inputs[151]) | (inputs[216]));
    assign layer0_outputs[1862] = ~(inputs[82]);
    assign layer0_outputs[1863] = (inputs[26]) & (inputs[129]);
    assign layer0_outputs[1864] = 1'b0;
    assign layer0_outputs[1865] = (inputs[87]) & ~(inputs[178]);
    assign layer0_outputs[1866] = inputs[72];
    assign layer0_outputs[1867] = ~(inputs[60]);
    assign layer0_outputs[1868] = ~(inputs[67]);
    assign layer0_outputs[1869] = (inputs[65]) | (inputs[234]);
    assign layer0_outputs[1870] = inputs[42];
    assign layer0_outputs[1871] = ~(inputs[184]) | (inputs[73]);
    assign layer0_outputs[1872] = ~((inputs[134]) ^ (inputs[162]));
    assign layer0_outputs[1873] = (inputs[184]) ^ (inputs[45]);
    assign layer0_outputs[1874] = (inputs[129]) | (inputs[165]);
    assign layer0_outputs[1875] = ~(inputs[2]);
    assign layer0_outputs[1876] = 1'b1;
    assign layer0_outputs[1877] = (inputs[119]) | (inputs[234]);
    assign layer0_outputs[1878] = ~(inputs[163]);
    assign layer0_outputs[1879] = ~(inputs[92]);
    assign layer0_outputs[1880] = ~((inputs[4]) ^ (inputs[105]));
    assign layer0_outputs[1881] = ~(inputs[89]);
    assign layer0_outputs[1882] = ~((inputs[180]) | (inputs[36]));
    assign layer0_outputs[1883] = ~(inputs[60]);
    assign layer0_outputs[1884] = (inputs[86]) | (inputs[229]);
    assign layer0_outputs[1885] = (inputs[40]) & ~(inputs[93]);
    assign layer0_outputs[1886] = ~((inputs[159]) & (inputs[191]));
    assign layer0_outputs[1887] = (inputs[220]) | (inputs[132]);
    assign layer0_outputs[1888] = (inputs[130]) | (inputs[223]);
    assign layer0_outputs[1889] = ~(inputs[182]) | (inputs[205]);
    assign layer0_outputs[1890] = ~(inputs[23]);
    assign layer0_outputs[1891] = ~((inputs[32]) ^ (inputs[19]));
    assign layer0_outputs[1892] = ~((inputs[180]) | (inputs[239]));
    assign layer0_outputs[1893] = ~(inputs[138]);
    assign layer0_outputs[1894] = ~(inputs[231]);
    assign layer0_outputs[1895] = (inputs[210]) & ~(inputs[237]);
    assign layer0_outputs[1896] = inputs[144];
    assign layer0_outputs[1897] = (inputs[10]) ^ (inputs[98]);
    assign layer0_outputs[1898] = ~(inputs[140]);
    assign layer0_outputs[1899] = ~(inputs[45]) | (inputs[174]);
    assign layer0_outputs[1900] = ~((inputs[185]) | (inputs[134]));
    assign layer0_outputs[1901] = ~(inputs[149]);
    assign layer0_outputs[1902] = inputs[180];
    assign layer0_outputs[1903] = (inputs[80]) ^ (inputs[186]);
    assign layer0_outputs[1904] = ~(inputs[32]);
    assign layer0_outputs[1905] = ~((inputs[22]) | (inputs[29]));
    assign layer0_outputs[1906] = 1'b0;
    assign layer0_outputs[1907] = ~((inputs[94]) ^ (inputs[18]));
    assign layer0_outputs[1908] = (inputs[74]) & ~(inputs[236]);
    assign layer0_outputs[1909] = (inputs[128]) & ~(inputs[241]);
    assign layer0_outputs[1910] = (inputs[39]) & ~(inputs[27]);
    assign layer0_outputs[1911] = ~(inputs[52]);
    assign layer0_outputs[1912] = (inputs[117]) & ~(inputs[97]);
    assign layer0_outputs[1913] = ~((inputs[37]) ^ (inputs[154]));
    assign layer0_outputs[1914] = ~(inputs[99]);
    assign layer0_outputs[1915] = inputs[108];
    assign layer0_outputs[1916] = ~((inputs[60]) | (inputs[59]));
    assign layer0_outputs[1917] = ~(inputs[175]);
    assign layer0_outputs[1918] = ~(inputs[88]) | (inputs[170]);
    assign layer0_outputs[1919] = ~((inputs[241]) ^ (inputs[167]));
    assign layer0_outputs[1920] = (inputs[66]) | (inputs[227]);
    assign layer0_outputs[1921] = (inputs[78]) & ~(inputs[97]);
    assign layer0_outputs[1922] = inputs[106];
    assign layer0_outputs[1923] = (inputs[203]) & ~(inputs[97]);
    assign layer0_outputs[1924] = (inputs[151]) & ~(inputs[175]);
    assign layer0_outputs[1925] = (inputs[84]) ^ (inputs[188]);
    assign layer0_outputs[1926] = ~((inputs[220]) | (inputs[247]));
    assign layer0_outputs[1927] = ~((inputs[178]) | (inputs[69]));
    assign layer0_outputs[1928] = inputs[92];
    assign layer0_outputs[1929] = ~(inputs[86]);
    assign layer0_outputs[1930] = ~(inputs[87]) | (inputs[162]);
    assign layer0_outputs[1931] = ~(inputs[209]) | (inputs[17]);
    assign layer0_outputs[1932] = ~((inputs[172]) | (inputs[9]));
    assign layer0_outputs[1933] = ~(inputs[53]) | (inputs[129]);
    assign layer0_outputs[1934] = ~((inputs[134]) | (inputs[156]));
    assign layer0_outputs[1935] = ~((inputs[34]) ^ (inputs[179]));
    assign layer0_outputs[1936] = inputs[120];
    assign layer0_outputs[1937] = ~((inputs[76]) | (inputs[160]));
    assign layer0_outputs[1938] = (inputs[15]) & ~(inputs[28]);
    assign layer0_outputs[1939] = inputs[210];
    assign layer0_outputs[1940] = inputs[55];
    assign layer0_outputs[1941] = ~((inputs[239]) ^ (inputs[5]));
    assign layer0_outputs[1942] = ~((inputs[101]) ^ (inputs[237]));
    assign layer0_outputs[1943] = ~(inputs[181]);
    assign layer0_outputs[1944] = (inputs[5]) ^ (inputs[208]);
    assign layer0_outputs[1945] = ~(inputs[6]) | (inputs[227]);
    assign layer0_outputs[1946] = ~((inputs[155]) | (inputs[179]));
    assign layer0_outputs[1947] = ~((inputs[199]) ^ (inputs[191]));
    assign layer0_outputs[1948] = (inputs[46]) ^ (inputs[67]);
    assign layer0_outputs[1949] = ~((inputs[210]) & (inputs[21]));
    assign layer0_outputs[1950] = ~(inputs[171]);
    assign layer0_outputs[1951] = (inputs[222]) | (inputs[252]);
    assign layer0_outputs[1952] = ~(inputs[232]) | (inputs[202]);
    assign layer0_outputs[1953] = (inputs[167]) & ~(inputs[18]);
    assign layer0_outputs[1954] = ~(inputs[133]) | (inputs[228]);
    assign layer0_outputs[1955] = inputs[189];
    assign layer0_outputs[1956] = ~(inputs[95]) | (inputs[194]);
    assign layer0_outputs[1957] = ~((inputs[15]) & (inputs[199]));
    assign layer0_outputs[1958] = ~(inputs[214]);
    assign layer0_outputs[1959] = inputs[201];
    assign layer0_outputs[1960] = (inputs[153]) ^ (inputs[5]);
    assign layer0_outputs[1961] = (inputs[123]) & ~(inputs[36]);
    assign layer0_outputs[1962] = 1'b1;
    assign layer0_outputs[1963] = ~((inputs[147]) | (inputs[122]));
    assign layer0_outputs[1964] = ~((inputs[4]) & (inputs[31]));
    assign layer0_outputs[1965] = ~((inputs[228]) | (inputs[70]));
    assign layer0_outputs[1966] = ~(inputs[25]);
    assign layer0_outputs[1967] = 1'b1;
    assign layer0_outputs[1968] = ~(inputs[148]) | (inputs[193]);
    assign layer0_outputs[1969] = ~((inputs[245]) & (inputs[79]));
    assign layer0_outputs[1970] = (inputs[218]) & ~(inputs[174]);
    assign layer0_outputs[1971] = ~((inputs[87]) ^ (inputs[145]));
    assign layer0_outputs[1972] = (inputs[33]) ^ (inputs[106]);
    assign layer0_outputs[1973] = inputs[183];
    assign layer0_outputs[1974] = (inputs[25]) & ~(inputs[93]);
    assign layer0_outputs[1975] = ~(inputs[186]) | (inputs[99]);
    assign layer0_outputs[1976] = ~((inputs[77]) | (inputs[94]));
    assign layer0_outputs[1977] = ~((inputs[16]) | (inputs[144]));
    assign layer0_outputs[1978] = (inputs[63]) | (inputs[231]);
    assign layer0_outputs[1979] = (inputs[11]) | (inputs[81]);
    assign layer0_outputs[1980] = ~((inputs[125]) | (inputs[47]));
    assign layer0_outputs[1981] = inputs[140];
    assign layer0_outputs[1982] = ~((inputs[194]) | (inputs[157]));
    assign layer0_outputs[1983] = inputs[77];
    assign layer0_outputs[1984] = ~((inputs[125]) ^ (inputs[139]));
    assign layer0_outputs[1985] = ~(inputs[193]);
    assign layer0_outputs[1986] = (inputs[22]) & (inputs[35]);
    assign layer0_outputs[1987] = (inputs[153]) & ~(inputs[18]);
    assign layer0_outputs[1988] = ~(inputs[111]);
    assign layer0_outputs[1989] = (inputs[49]) & (inputs[44]);
    assign layer0_outputs[1990] = ~(inputs[95]);
    assign layer0_outputs[1991] = ~(inputs[255]);
    assign layer0_outputs[1992] = ~(inputs[136]);
    assign layer0_outputs[1993] = ~(inputs[239]);
    assign layer0_outputs[1994] = ~((inputs[252]) ^ (inputs[148]));
    assign layer0_outputs[1995] = (inputs[252]) | (inputs[89]);
    assign layer0_outputs[1996] = ~(inputs[87]) | (inputs[43]);
    assign layer0_outputs[1997] = (inputs[42]) ^ (inputs[229]);
    assign layer0_outputs[1998] = ~((inputs[65]) | (inputs[148]));
    assign layer0_outputs[1999] = (inputs[82]) ^ (inputs[255]);
    assign layer0_outputs[2000] = (inputs[182]) ^ (inputs[41]);
    assign layer0_outputs[2001] = (inputs[216]) & ~(inputs[49]);
    assign layer0_outputs[2002] = inputs[166];
    assign layer0_outputs[2003] = ~(inputs[81]) | (inputs[24]);
    assign layer0_outputs[2004] = ~(inputs[104]) | (inputs[67]);
    assign layer0_outputs[2005] = ~(inputs[167]);
    assign layer0_outputs[2006] = (inputs[196]) & ~(inputs[253]);
    assign layer0_outputs[2007] = ~(inputs[253]);
    assign layer0_outputs[2008] = ~(inputs[239]) | (inputs[216]);
    assign layer0_outputs[2009] = (inputs[38]) | (inputs[239]);
    assign layer0_outputs[2010] = inputs[100];
    assign layer0_outputs[2011] = (inputs[227]) & ~(inputs[161]);
    assign layer0_outputs[2012] = inputs[153];
    assign layer0_outputs[2013] = inputs[152];
    assign layer0_outputs[2014] = ~(inputs[216]) | (inputs[111]);
    assign layer0_outputs[2015] = inputs[203];
    assign layer0_outputs[2016] = ~(inputs[186]);
    assign layer0_outputs[2017] = ~((inputs[163]) | (inputs[187]));
    assign layer0_outputs[2018] = ~((inputs[153]) | (inputs[25]));
    assign layer0_outputs[2019] = ~(inputs[38]) | (inputs[13]);
    assign layer0_outputs[2020] = (inputs[91]) | (inputs[238]);
    assign layer0_outputs[2021] = ~(inputs[188]);
    assign layer0_outputs[2022] = inputs[6];
    assign layer0_outputs[2023] = inputs[217];
    assign layer0_outputs[2024] = ~(inputs[189]) | (inputs[45]);
    assign layer0_outputs[2025] = (inputs[71]) | (inputs[204]);
    assign layer0_outputs[2026] = inputs[154];
    assign layer0_outputs[2027] = ~((inputs[140]) | (inputs[115]));
    assign layer0_outputs[2028] = inputs[100];
    assign layer0_outputs[2029] = 1'b0;
    assign layer0_outputs[2030] = ~(inputs[231]) | (inputs[13]);
    assign layer0_outputs[2031] = ~(inputs[132]);
    assign layer0_outputs[2032] = ~((inputs[245]) | (inputs[83]));
    assign layer0_outputs[2033] = ~(inputs[141]);
    assign layer0_outputs[2034] = (inputs[238]) ^ (inputs[212]);
    assign layer0_outputs[2035] = 1'b1;
    assign layer0_outputs[2036] = ~((inputs[160]) & (inputs[82]));
    assign layer0_outputs[2037] = ~(inputs[22]);
    assign layer0_outputs[2038] = (inputs[253]) & ~(inputs[207]);
    assign layer0_outputs[2039] = ~((inputs[194]) | (inputs[5]));
    assign layer0_outputs[2040] = ~(inputs[8]) | (inputs[220]);
    assign layer0_outputs[2041] = (inputs[165]) & ~(inputs[228]);
    assign layer0_outputs[2042] = (inputs[53]) | (inputs[65]);
    assign layer0_outputs[2043] = (inputs[142]) & (inputs[146]);
    assign layer0_outputs[2044] = inputs[203];
    assign layer0_outputs[2045] = ~((inputs[236]) | (inputs[61]));
    assign layer0_outputs[2046] = ~((inputs[57]) ^ (inputs[208]));
    assign layer0_outputs[2047] = (inputs[223]) ^ (inputs[105]);
    assign layer0_outputs[2048] = 1'b1;
    assign layer0_outputs[2049] = ~((inputs[143]) | (inputs[215]));
    assign layer0_outputs[2050] = (inputs[199]) | (inputs[127]);
    assign layer0_outputs[2051] = (inputs[105]) & ~(inputs[0]);
    assign layer0_outputs[2052] = ~((inputs[217]) | (inputs[104]));
    assign layer0_outputs[2053] = (inputs[106]) & ~(inputs[254]);
    assign layer0_outputs[2054] = ~((inputs[92]) | (inputs[93]));
    assign layer0_outputs[2055] = ~(inputs[34]);
    assign layer0_outputs[2056] = 1'b0;
    assign layer0_outputs[2057] = ~(inputs[107]);
    assign layer0_outputs[2058] = (inputs[86]) & ~(inputs[32]);
    assign layer0_outputs[2059] = ~(inputs[42]) | (inputs[94]);
    assign layer0_outputs[2060] = (inputs[131]) | (inputs[59]);
    assign layer0_outputs[2061] = ~(inputs[252]) | (inputs[49]);
    assign layer0_outputs[2062] = inputs[234];
    assign layer0_outputs[2063] = (inputs[146]) | (inputs[169]);
    assign layer0_outputs[2064] = (inputs[43]) & ~(inputs[254]);
    assign layer0_outputs[2065] = (inputs[189]) | (inputs[252]);
    assign layer0_outputs[2066] = (inputs[175]) & ~(inputs[245]);
    assign layer0_outputs[2067] = (inputs[158]) | (inputs[180]);
    assign layer0_outputs[2068] = (inputs[190]) | (inputs[250]);
    assign layer0_outputs[2069] = ~(inputs[96]) | (inputs[23]);
    assign layer0_outputs[2070] = ~((inputs[18]) | (inputs[103]));
    assign layer0_outputs[2071] = (inputs[170]) | (inputs[38]);
    assign layer0_outputs[2072] = ~(inputs[65]);
    assign layer0_outputs[2073] = ~((inputs[138]) | (inputs[81]));
    assign layer0_outputs[2074] = ~(inputs[123]);
    assign layer0_outputs[2075] = inputs[150];
    assign layer0_outputs[2076] = inputs[124];
    assign layer0_outputs[2077] = (inputs[86]) & ~(inputs[62]);
    assign layer0_outputs[2078] = (inputs[18]) | (inputs[182]);
    assign layer0_outputs[2079] = 1'b0;
    assign layer0_outputs[2080] = ~(inputs[247]) | (inputs[207]);
    assign layer0_outputs[2081] = 1'b1;
    assign layer0_outputs[2082] = inputs[68];
    assign layer0_outputs[2083] = ~(inputs[26]) | (inputs[62]);
    assign layer0_outputs[2084] = inputs[156];
    assign layer0_outputs[2085] = (inputs[198]) & ~(inputs[206]);
    assign layer0_outputs[2086] = (inputs[198]) | (inputs[80]);
    assign layer0_outputs[2087] = ~((inputs[34]) | (inputs[231]));
    assign layer0_outputs[2088] = ~((inputs[21]) | (inputs[14]));
    assign layer0_outputs[2089] = (inputs[84]) ^ (inputs[41]);
    assign layer0_outputs[2090] = ~((inputs[157]) | (inputs[132]));
    assign layer0_outputs[2091] = inputs[231];
    assign layer0_outputs[2092] = (inputs[219]) & ~(inputs[206]);
    assign layer0_outputs[2093] = (inputs[153]) & ~(inputs[182]);
    assign layer0_outputs[2094] = (inputs[128]) | (inputs[86]);
    assign layer0_outputs[2095] = (inputs[9]) | (inputs[194]);
    assign layer0_outputs[2096] = (inputs[18]) | (inputs[130]);
    assign layer0_outputs[2097] = (inputs[117]) & ~(inputs[80]);
    assign layer0_outputs[2098] = ~((inputs[54]) ^ (inputs[144]));
    assign layer0_outputs[2099] = ~((inputs[239]) ^ (inputs[228]));
    assign layer0_outputs[2100] = inputs[57];
    assign layer0_outputs[2101] = inputs[84];
    assign layer0_outputs[2102] = ~((inputs[211]) | (inputs[188]));
    assign layer0_outputs[2103] = (inputs[145]) ^ (inputs[166]);
    assign layer0_outputs[2104] = ~(inputs[179]);
    assign layer0_outputs[2105] = inputs[57];
    assign layer0_outputs[2106] = ~(inputs[242]);
    assign layer0_outputs[2107] = ~(inputs[100]) | (inputs[13]);
    assign layer0_outputs[2108] = ~((inputs[87]) ^ (inputs[70]));
    assign layer0_outputs[2109] = ~((inputs[35]) ^ (inputs[196]));
    assign layer0_outputs[2110] = inputs[41];
    assign layer0_outputs[2111] = ~(inputs[92]);
    assign layer0_outputs[2112] = (inputs[118]) & ~(inputs[38]);
    assign layer0_outputs[2113] = (inputs[25]) ^ (inputs[76]);
    assign layer0_outputs[2114] = 1'b0;
    assign layer0_outputs[2115] = ~((inputs[106]) | (inputs[150]));
    assign layer0_outputs[2116] = inputs[254];
    assign layer0_outputs[2117] = ~((inputs[206]) | (inputs[68]));
    assign layer0_outputs[2118] = (inputs[57]) | (inputs[37]);
    assign layer0_outputs[2119] = ~(inputs[47]);
    assign layer0_outputs[2120] = ~(inputs[182]);
    assign layer0_outputs[2121] = (inputs[107]) & ~(inputs[22]);
    assign layer0_outputs[2122] = ~((inputs[228]) & (inputs[7]));
    assign layer0_outputs[2123] = (inputs[71]) & ~(inputs[204]);
    assign layer0_outputs[2124] = 1'b0;
    assign layer0_outputs[2125] = inputs[182];
    assign layer0_outputs[2126] = inputs[207];
    assign layer0_outputs[2127] = inputs[214];
    assign layer0_outputs[2128] = inputs[40];
    assign layer0_outputs[2129] = (inputs[180]) | (inputs[251]);
    assign layer0_outputs[2130] = ~((inputs[91]) | (inputs[122]));
    assign layer0_outputs[2131] = ~(inputs[193]);
    assign layer0_outputs[2132] = 1'b1;
    assign layer0_outputs[2133] = ~(inputs[201]) | (inputs[32]);
    assign layer0_outputs[2134] = inputs[214];
    assign layer0_outputs[2135] = ~(inputs[52]) | (inputs[144]);
    assign layer0_outputs[2136] = (inputs[192]) & ~(inputs[2]);
    assign layer0_outputs[2137] = (inputs[179]) & ~(inputs[6]);
    assign layer0_outputs[2138] = 1'b0;
    assign layer0_outputs[2139] = (inputs[255]) & ~(inputs[143]);
    assign layer0_outputs[2140] = inputs[59];
    assign layer0_outputs[2141] = ~((inputs[76]) ^ (inputs[75]));
    assign layer0_outputs[2142] = inputs[82];
    assign layer0_outputs[2143] = ~(inputs[229]);
    assign layer0_outputs[2144] = inputs[118];
    assign layer0_outputs[2145] = 1'b1;
    assign layer0_outputs[2146] = (inputs[40]) & ~(inputs[90]);
    assign layer0_outputs[2147] = 1'b0;
    assign layer0_outputs[2148] = (inputs[203]) & ~(inputs[7]);
    assign layer0_outputs[2149] = ~(inputs[114]);
    assign layer0_outputs[2150] = ~((inputs[216]) ^ (inputs[240]));
    assign layer0_outputs[2151] = ~((inputs[158]) & (inputs[243]));
    assign layer0_outputs[2152] = ~((inputs[172]) | (inputs[187]));
    assign layer0_outputs[2153] = ~(inputs[217]);
    assign layer0_outputs[2154] = (inputs[106]) ^ (inputs[210]);
    assign layer0_outputs[2155] = ~(inputs[202]);
    assign layer0_outputs[2156] = ~((inputs[148]) ^ (inputs[4]));
    assign layer0_outputs[2157] = ~(inputs[151]) | (inputs[127]);
    assign layer0_outputs[2158] = ~((inputs[150]) | (inputs[220]));
    assign layer0_outputs[2159] = 1'b1;
    assign layer0_outputs[2160] = ~(inputs[132]);
    assign layer0_outputs[2161] = ~((inputs[108]) ^ (inputs[233]));
    assign layer0_outputs[2162] = ~((inputs[15]) ^ (inputs[150]));
    assign layer0_outputs[2163] = inputs[255];
    assign layer0_outputs[2164] = (inputs[116]) & ~(inputs[84]);
    assign layer0_outputs[2165] = (inputs[200]) & ~(inputs[31]);
    assign layer0_outputs[2166] = (inputs[12]) & (inputs[12]);
    assign layer0_outputs[2167] = ~(inputs[179]) | (inputs[64]);
    assign layer0_outputs[2168] = ~((inputs[84]) | (inputs[42]));
    assign layer0_outputs[2169] = (inputs[178]) & ~(inputs[15]);
    assign layer0_outputs[2170] = ~(inputs[188]) | (inputs[253]);
    assign layer0_outputs[2171] = (inputs[230]) | (inputs[106]);
    assign layer0_outputs[2172] = (inputs[198]) & ~(inputs[110]);
    assign layer0_outputs[2173] = ~((inputs[96]) | (inputs[221]));
    assign layer0_outputs[2174] = (inputs[167]) & ~(inputs[251]);
    assign layer0_outputs[2175] = ~((inputs[64]) | (inputs[234]));
    assign layer0_outputs[2176] = ~(inputs[186]) | (inputs[65]);
    assign layer0_outputs[2177] = ~((inputs[10]) | (inputs[110]));
    assign layer0_outputs[2178] = ~((inputs[96]) | (inputs[101]));
    assign layer0_outputs[2179] = inputs[119];
    assign layer0_outputs[2180] = 1'b0;
    assign layer0_outputs[2181] = ~(inputs[124]);
    assign layer0_outputs[2182] = (inputs[176]) & ~(inputs[245]);
    assign layer0_outputs[2183] = (inputs[23]) & ~(inputs[91]);
    assign layer0_outputs[2184] = 1'b0;
    assign layer0_outputs[2185] = (inputs[65]) | (inputs[177]);
    assign layer0_outputs[2186] = ~(inputs[158]) | (inputs[236]);
    assign layer0_outputs[2187] = (inputs[133]) & ~(inputs[38]);
    assign layer0_outputs[2188] = (inputs[193]) & ~(inputs[34]);
    assign layer0_outputs[2189] = ~(inputs[84]) | (inputs[194]);
    assign layer0_outputs[2190] = ~((inputs[173]) ^ (inputs[4]));
    assign layer0_outputs[2191] = ~(inputs[120]) | (inputs[62]);
    assign layer0_outputs[2192] = ~(inputs[164]) | (inputs[45]);
    assign layer0_outputs[2193] = ~(inputs[80]);
    assign layer0_outputs[2194] = ~(inputs[30]) | (inputs[240]);
    assign layer0_outputs[2195] = ~(inputs[44]);
    assign layer0_outputs[2196] = (inputs[250]) & ~(inputs[141]);
    assign layer0_outputs[2197] = ~((inputs[162]) ^ (inputs[190]));
    assign layer0_outputs[2198] = (inputs[186]) & ~(inputs[206]);
    assign layer0_outputs[2199] = 1'b1;
    assign layer0_outputs[2200] = (inputs[102]) & ~(inputs[251]);
    assign layer0_outputs[2201] = (inputs[239]) & (inputs[239]);
    assign layer0_outputs[2202] = (inputs[25]) ^ (inputs[114]);
    assign layer0_outputs[2203] = ~((inputs[184]) | (inputs[222]));
    assign layer0_outputs[2204] = (inputs[50]) & (inputs[110]);
    assign layer0_outputs[2205] = ~((inputs[214]) | (inputs[98]));
    assign layer0_outputs[2206] = (inputs[84]) | (inputs[250]);
    assign layer0_outputs[2207] = (inputs[254]) ^ (inputs[121]);
    assign layer0_outputs[2208] = ~((inputs[91]) ^ (inputs[12]));
    assign layer0_outputs[2209] = ~(inputs[123]);
    assign layer0_outputs[2210] = ~((inputs[110]) | (inputs[133]));
    assign layer0_outputs[2211] = ~((inputs[8]) ^ (inputs[169]));
    assign layer0_outputs[2212] = ~(inputs[183]);
    assign layer0_outputs[2213] = inputs[87];
    assign layer0_outputs[2214] = (inputs[170]) | (inputs[96]);
    assign layer0_outputs[2215] = ~(inputs[122]);
    assign layer0_outputs[2216] = inputs[182];
    assign layer0_outputs[2217] = ~(inputs[54]) | (inputs[117]);
    assign layer0_outputs[2218] = ~(inputs[177]) | (inputs[254]);
    assign layer0_outputs[2219] = (inputs[12]) | (inputs[183]);
    assign layer0_outputs[2220] = ~(inputs[74]);
    assign layer0_outputs[2221] = ~(inputs[40]) | (inputs[88]);
    assign layer0_outputs[2222] = 1'b0;
    assign layer0_outputs[2223] = ~(inputs[112]) | (inputs[21]);
    assign layer0_outputs[2224] = (inputs[3]) ^ (inputs[241]);
    assign layer0_outputs[2225] = (inputs[9]) & (inputs[144]);
    assign layer0_outputs[2226] = ~(inputs[51]) | (inputs[96]);
    assign layer0_outputs[2227] = (inputs[219]) | (inputs[178]);
    assign layer0_outputs[2228] = inputs[167];
    assign layer0_outputs[2229] = ~(inputs[71]);
    assign layer0_outputs[2230] = (inputs[143]) | (inputs[125]);
    assign layer0_outputs[2231] = (inputs[47]) & ~(inputs[31]);
    assign layer0_outputs[2232] = (inputs[251]) ^ (inputs[158]);
    assign layer0_outputs[2233] = 1'b0;
    assign layer0_outputs[2234] = (inputs[171]) & ~(inputs[175]);
    assign layer0_outputs[2235] = inputs[235];
    assign layer0_outputs[2236] = ~((inputs[87]) | (inputs[247]));
    assign layer0_outputs[2237] = (inputs[167]) & ~(inputs[196]);
    assign layer0_outputs[2238] = (inputs[7]) | (inputs[39]);
    assign layer0_outputs[2239] = ~(inputs[181]);
    assign layer0_outputs[2240] = ~(inputs[214]);
    assign layer0_outputs[2241] = (inputs[116]) & ~(inputs[44]);
    assign layer0_outputs[2242] = (inputs[138]) ^ (inputs[57]);
    assign layer0_outputs[2243] = (inputs[138]) & ~(inputs[210]);
    assign layer0_outputs[2244] = ~((inputs[22]) ^ (inputs[41]));
    assign layer0_outputs[2245] = (inputs[8]) | (inputs[31]);
    assign layer0_outputs[2246] = (inputs[251]) ^ (inputs[232]);
    assign layer0_outputs[2247] = (inputs[133]) & ~(inputs[14]);
    assign layer0_outputs[2248] = (inputs[244]) | (inputs[48]);
    assign layer0_outputs[2249] = ~(inputs[152]);
    assign layer0_outputs[2250] = inputs[166];
    assign layer0_outputs[2251] = ~(inputs[199]);
    assign layer0_outputs[2252] = (inputs[161]) & ~(inputs[111]);
    assign layer0_outputs[2253] = (inputs[16]) ^ (inputs[100]);
    assign layer0_outputs[2254] = ~((inputs[47]) & (inputs[81]));
    assign layer0_outputs[2255] = ~((inputs[181]) | (inputs[29]));
    assign layer0_outputs[2256] = (inputs[96]) | (inputs[42]);
    assign layer0_outputs[2257] = ~(inputs[207]);
    assign layer0_outputs[2258] = ~(inputs[89]);
    assign layer0_outputs[2259] = ~((inputs[38]) & (inputs[85]));
    assign layer0_outputs[2260] = inputs[104];
    assign layer0_outputs[2261] = inputs[131];
    assign layer0_outputs[2262] = (inputs[235]) | (inputs[137]);
    assign layer0_outputs[2263] = (inputs[122]) | (inputs[54]);
    assign layer0_outputs[2264] = ~((inputs[173]) | (inputs[219]));
    assign layer0_outputs[2265] = ~((inputs[197]) | (inputs[100]));
    assign layer0_outputs[2266] = ~((inputs[44]) | (inputs[180]));
    assign layer0_outputs[2267] = inputs[213];
    assign layer0_outputs[2268] = (inputs[54]) | (inputs[162]);
    assign layer0_outputs[2269] = (inputs[181]) | (inputs[149]);
    assign layer0_outputs[2270] = (inputs[70]) & ~(inputs[123]);
    assign layer0_outputs[2271] = ~((inputs[239]) | (inputs[176]));
    assign layer0_outputs[2272] = ~(inputs[195]);
    assign layer0_outputs[2273] = inputs[86];
    assign layer0_outputs[2274] = (inputs[153]) | (inputs[149]);
    assign layer0_outputs[2275] = (inputs[18]) ^ (inputs[187]);
    assign layer0_outputs[2276] = ~((inputs[125]) | (inputs[117]));
    assign layer0_outputs[2277] = ~((inputs[21]) | (inputs[95]));
    assign layer0_outputs[2278] = ~(inputs[215]) | (inputs[182]);
    assign layer0_outputs[2279] = ~((inputs[226]) ^ (inputs[52]));
    assign layer0_outputs[2280] = ~(inputs[73]);
    assign layer0_outputs[2281] = ~(inputs[246]);
    assign layer0_outputs[2282] = (inputs[34]) ^ (inputs[128]);
    assign layer0_outputs[2283] = ~(inputs[188]);
    assign layer0_outputs[2284] = ~((inputs[57]) ^ (inputs[247]));
    assign layer0_outputs[2285] = ~((inputs[43]) ^ (inputs[17]));
    assign layer0_outputs[2286] = ~(inputs[136]) | (inputs[108]);
    assign layer0_outputs[2287] = (inputs[169]) & ~(inputs[46]);
    assign layer0_outputs[2288] = ~((inputs[198]) | (inputs[53]));
    assign layer0_outputs[2289] = (inputs[87]) & ~(inputs[145]);
    assign layer0_outputs[2290] = (inputs[146]) & ~(inputs[112]);
    assign layer0_outputs[2291] = ~(inputs[131]) | (inputs[35]);
    assign layer0_outputs[2292] = ~((inputs[139]) ^ (inputs[71]));
    assign layer0_outputs[2293] = inputs[203];
    assign layer0_outputs[2294] = (inputs[131]) | (inputs[229]);
    assign layer0_outputs[2295] = ~((inputs[9]) | (inputs[100]));
    assign layer0_outputs[2296] = inputs[68];
    assign layer0_outputs[2297] = inputs[153];
    assign layer0_outputs[2298] = inputs[117];
    assign layer0_outputs[2299] = ~(inputs[158]);
    assign layer0_outputs[2300] = (inputs[54]) & ~(inputs[227]);
    assign layer0_outputs[2301] = (inputs[233]) | (inputs[9]);
    assign layer0_outputs[2302] = ~(inputs[167]);
    assign layer0_outputs[2303] = (inputs[242]) | (inputs[116]);
    assign layer0_outputs[2304] = (inputs[222]) | (inputs[184]);
    assign layer0_outputs[2305] = (inputs[217]) ^ (inputs[208]);
    assign layer0_outputs[2306] = ~(inputs[226]);
    assign layer0_outputs[2307] = ~(inputs[45]);
    assign layer0_outputs[2308] = ~((inputs[244]) | (inputs[123]));
    assign layer0_outputs[2309] = (inputs[151]) & ~(inputs[83]);
    assign layer0_outputs[2310] = ~(inputs[117]);
    assign layer0_outputs[2311] = (inputs[211]) & ~(inputs[44]);
    assign layer0_outputs[2312] = ~((inputs[53]) & (inputs[5]));
    assign layer0_outputs[2313] = (inputs[28]) ^ (inputs[217]);
    assign layer0_outputs[2314] = ~(inputs[79]) | (inputs[167]);
    assign layer0_outputs[2315] = ~(inputs[190]) | (inputs[9]);
    assign layer0_outputs[2316] = ~((inputs[208]) | (inputs[125]));
    assign layer0_outputs[2317] = ~((inputs[155]) | (inputs[140]));
    assign layer0_outputs[2318] = (inputs[20]) & (inputs[99]);
    assign layer0_outputs[2319] = ~((inputs[108]) | (inputs[56]));
    assign layer0_outputs[2320] = ~(inputs[199]);
    assign layer0_outputs[2321] = ~((inputs[1]) & (inputs[160]));
    assign layer0_outputs[2322] = ~(inputs[24]) | (inputs[17]);
    assign layer0_outputs[2323] = (inputs[142]) | (inputs[210]);
    assign layer0_outputs[2324] = ~(inputs[148]);
    assign layer0_outputs[2325] = ~(inputs[135]) | (inputs[233]);
    assign layer0_outputs[2326] = inputs[252];
    assign layer0_outputs[2327] = ~(inputs[229]) | (inputs[48]);
    assign layer0_outputs[2328] = (inputs[21]) & ~(inputs[41]);
    assign layer0_outputs[2329] = (inputs[118]) ^ (inputs[247]);
    assign layer0_outputs[2330] = (inputs[102]) & ~(inputs[198]);
    assign layer0_outputs[2331] = (inputs[4]) ^ (inputs[234]);
    assign layer0_outputs[2332] = ~(inputs[134]) | (inputs[41]);
    assign layer0_outputs[2333] = inputs[189];
    assign layer0_outputs[2334] = (inputs[98]) | (inputs[108]);
    assign layer0_outputs[2335] = inputs[194];
    assign layer0_outputs[2336] = ~(inputs[215]) | (inputs[16]);
    assign layer0_outputs[2337] = ~(inputs[86]);
    assign layer0_outputs[2338] = ~(inputs[96]);
    assign layer0_outputs[2339] = (inputs[189]) | (inputs[191]);
    assign layer0_outputs[2340] = ~((inputs[245]) ^ (inputs[85]));
    assign layer0_outputs[2341] = ~((inputs[57]) ^ (inputs[252]));
    assign layer0_outputs[2342] = inputs[58];
    assign layer0_outputs[2343] = ~((inputs[146]) ^ (inputs[134]));
    assign layer0_outputs[2344] = (inputs[78]) & ~(inputs[54]);
    assign layer0_outputs[2345] = (inputs[152]) | (inputs[151]);
    assign layer0_outputs[2346] = ~(inputs[69]);
    assign layer0_outputs[2347] = (inputs[127]) & ~(inputs[80]);
    assign layer0_outputs[2348] = ~(inputs[101]);
    assign layer0_outputs[2349] = (inputs[45]) & (inputs[12]);
    assign layer0_outputs[2350] = ~((inputs[34]) ^ (inputs[85]));
    assign layer0_outputs[2351] = ~(inputs[38]) | (inputs[227]);
    assign layer0_outputs[2352] = ~((inputs[144]) | (inputs[221]));
    assign layer0_outputs[2353] = (inputs[78]) ^ (inputs[99]);
    assign layer0_outputs[2354] = inputs[181];
    assign layer0_outputs[2355] = ~((inputs[44]) | (inputs[191]));
    assign layer0_outputs[2356] = (inputs[189]) | (inputs[187]);
    assign layer0_outputs[2357] = ~(inputs[150]);
    assign layer0_outputs[2358] = (inputs[206]) ^ (inputs[189]);
    assign layer0_outputs[2359] = inputs[98];
    assign layer0_outputs[2360] = inputs[234];
    assign layer0_outputs[2361] = (inputs[215]) | (inputs[61]);
    assign layer0_outputs[2362] = inputs[216];
    assign layer0_outputs[2363] = (inputs[78]) & ~(inputs[248]);
    assign layer0_outputs[2364] = inputs[164];
    assign layer0_outputs[2365] = ~(inputs[161]) | (inputs[158]);
    assign layer0_outputs[2366] = (inputs[95]) ^ (inputs[146]);
    assign layer0_outputs[2367] = ~(inputs[125]);
    assign layer0_outputs[2368] = inputs[165];
    assign layer0_outputs[2369] = ~((inputs[137]) | (inputs[99]));
    assign layer0_outputs[2370] = ~((inputs[8]) ^ (inputs[242]));
    assign layer0_outputs[2371] = (inputs[199]) & ~(inputs[224]);
    assign layer0_outputs[2372] = inputs[30];
    assign layer0_outputs[2373] = (inputs[1]) ^ (inputs[122]);
    assign layer0_outputs[2374] = ~(inputs[161]) | (inputs[12]);
    assign layer0_outputs[2375] = ~(inputs[142]) | (inputs[46]);
    assign layer0_outputs[2376] = ~((inputs[193]) | (inputs[201]));
    assign layer0_outputs[2377] = 1'b1;
    assign layer0_outputs[2378] = 1'b1;
    assign layer0_outputs[2379] = ~((inputs[253]) | (inputs[75]));
    assign layer0_outputs[2380] = ~(inputs[144]);
    assign layer0_outputs[2381] = ~(inputs[115]) | (inputs[192]);
    assign layer0_outputs[2382] = (inputs[139]) | (inputs[211]);
    assign layer0_outputs[2383] = inputs[206];
    assign layer0_outputs[2384] = ~((inputs[173]) & (inputs[227]));
    assign layer0_outputs[2385] = (inputs[165]) | (inputs[203]);
    assign layer0_outputs[2386] = inputs[66];
    assign layer0_outputs[2387] = (inputs[86]) & ~(inputs[197]);
    assign layer0_outputs[2388] = ~(inputs[90]) | (inputs[114]);
    assign layer0_outputs[2389] = ~((inputs[83]) ^ (inputs[40]));
    assign layer0_outputs[2390] = ~((inputs[106]) ^ (inputs[60]));
    assign layer0_outputs[2391] = (inputs[162]) & ~(inputs[158]);
    assign layer0_outputs[2392] = (inputs[70]) & ~(inputs[7]);
    assign layer0_outputs[2393] = ~(inputs[38]);
    assign layer0_outputs[2394] = ~((inputs[32]) ^ (inputs[130]));
    assign layer0_outputs[2395] = ~((inputs[238]) | (inputs[92]));
    assign layer0_outputs[2396] = ~((inputs[187]) | (inputs[160]));
    assign layer0_outputs[2397] = (inputs[249]) | (inputs[212]);
    assign layer0_outputs[2398] = inputs[180];
    assign layer0_outputs[2399] = (inputs[17]) & ~(inputs[127]);
    assign layer0_outputs[2400] = (inputs[203]) & ~(inputs[231]);
    assign layer0_outputs[2401] = ~((inputs[208]) ^ (inputs[206]));
    assign layer0_outputs[2402] = inputs[137];
    assign layer0_outputs[2403] = ~((inputs[251]) ^ (inputs[58]));
    assign layer0_outputs[2404] = ~(inputs[65]);
    assign layer0_outputs[2405] = inputs[253];
    assign layer0_outputs[2406] = inputs[99];
    assign layer0_outputs[2407] = (inputs[108]) | (inputs[221]);
    assign layer0_outputs[2408] = (inputs[205]) ^ (inputs[1]);
    assign layer0_outputs[2409] = ~(inputs[171]) | (inputs[147]);
    assign layer0_outputs[2410] = inputs[13];
    assign layer0_outputs[2411] = (inputs[45]) ^ (inputs[55]);
    assign layer0_outputs[2412] = (inputs[136]) & ~(inputs[142]);
    assign layer0_outputs[2413] = (inputs[126]) ^ (inputs[147]);
    assign layer0_outputs[2414] = (inputs[99]) & ~(inputs[236]);
    assign layer0_outputs[2415] = (inputs[53]) ^ (inputs[200]);
    assign layer0_outputs[2416] = (inputs[109]) & ~(inputs[21]);
    assign layer0_outputs[2417] = (inputs[110]) & (inputs[28]);
    assign layer0_outputs[2418] = inputs[219];
    assign layer0_outputs[2419] = 1'b0;
    assign layer0_outputs[2420] = (inputs[234]) ^ (inputs[18]);
    assign layer0_outputs[2421] = inputs[216];
    assign layer0_outputs[2422] = ~(inputs[102]);
    assign layer0_outputs[2423] = ~(inputs[9]) | (inputs[157]);
    assign layer0_outputs[2424] = (inputs[204]) | (inputs[71]);
    assign layer0_outputs[2425] = inputs[88];
    assign layer0_outputs[2426] = ~(inputs[170]);
    assign layer0_outputs[2427] = inputs[38];
    assign layer0_outputs[2428] = (inputs[110]) & ~(inputs[109]);
    assign layer0_outputs[2429] = ~((inputs[134]) ^ (inputs[32]));
    assign layer0_outputs[2430] = inputs[34];
    assign layer0_outputs[2431] = 1'b1;
    assign layer0_outputs[2432] = ~(inputs[154]) | (inputs[209]);
    assign layer0_outputs[2433] = ~(inputs[207]) | (inputs[175]);
    assign layer0_outputs[2434] = inputs[140];
    assign layer0_outputs[2435] = (inputs[182]) | (inputs[165]);
    assign layer0_outputs[2436] = ~((inputs[43]) & (inputs[81]));
    assign layer0_outputs[2437] = ~((inputs[56]) ^ (inputs[251]));
    assign layer0_outputs[2438] = (inputs[138]) & ~(inputs[42]);
    assign layer0_outputs[2439] = (inputs[50]) | (inputs[138]);
    assign layer0_outputs[2440] = ~((inputs[110]) & (inputs[41]));
    assign layer0_outputs[2441] = ~(inputs[217]) | (inputs[19]);
    assign layer0_outputs[2442] = ~((inputs[172]) | (inputs[171]));
    assign layer0_outputs[2443] = ~((inputs[63]) | (inputs[200]));
    assign layer0_outputs[2444] = inputs[137];
    assign layer0_outputs[2445] = ~(inputs[120]);
    assign layer0_outputs[2446] = ~(inputs[212]) | (inputs[62]);
    assign layer0_outputs[2447] = (inputs[155]) ^ (inputs[225]);
    assign layer0_outputs[2448] = (inputs[95]) & ~(inputs[1]);
    assign layer0_outputs[2449] = (inputs[23]) & ~(inputs[83]);
    assign layer0_outputs[2450] = ~((inputs[253]) | (inputs[91]));
    assign layer0_outputs[2451] = (inputs[63]) & (inputs[14]);
    assign layer0_outputs[2452] = (inputs[52]) & ~(inputs[246]);
    assign layer0_outputs[2453] = ~((inputs[201]) & (inputs[72]));
    assign layer0_outputs[2454] = (inputs[37]) ^ (inputs[169]);
    assign layer0_outputs[2455] = (inputs[220]) ^ (inputs[188]);
    assign layer0_outputs[2456] = ~((inputs[212]) ^ (inputs[75]));
    assign layer0_outputs[2457] = ~((inputs[45]) | (inputs[223]));
    assign layer0_outputs[2458] = (inputs[72]) & ~(inputs[220]);
    assign layer0_outputs[2459] = ~(inputs[233]);
    assign layer0_outputs[2460] = (inputs[86]) & ~(inputs[230]);
    assign layer0_outputs[2461] = (inputs[155]) & ~(inputs[46]);
    assign layer0_outputs[2462] = (inputs[181]) ^ (inputs[161]);
    assign layer0_outputs[2463] = ~(inputs[128]);
    assign layer0_outputs[2464] = ~((inputs[116]) | (inputs[24]));
    assign layer0_outputs[2465] = inputs[198];
    assign layer0_outputs[2466] = (inputs[48]) & ~(inputs[133]);
    assign layer0_outputs[2467] = (inputs[33]) & (inputs[3]);
    assign layer0_outputs[2468] = (inputs[88]) & ~(inputs[150]);
    assign layer0_outputs[2469] = inputs[164];
    assign layer0_outputs[2470] = 1'b1;
    assign layer0_outputs[2471] = ~(inputs[208]) | (inputs[205]);
    assign layer0_outputs[2472] = (inputs[184]) & ~(inputs[130]);
    assign layer0_outputs[2473] = (inputs[149]) | (inputs[167]);
    assign layer0_outputs[2474] = (inputs[26]) | (inputs[110]);
    assign layer0_outputs[2475] = (inputs[196]) ^ (inputs[34]);
    assign layer0_outputs[2476] = (inputs[45]) & (inputs[223]);
    assign layer0_outputs[2477] = ~(inputs[40]) | (inputs[231]);
    assign layer0_outputs[2478] = inputs[66];
    assign layer0_outputs[2479] = ~(inputs[217]) | (inputs[250]);
    assign layer0_outputs[2480] = (inputs[193]) & ~(inputs[142]);
    assign layer0_outputs[2481] = inputs[186];
    assign layer0_outputs[2482] = (inputs[146]) | (inputs[118]);
    assign layer0_outputs[2483] = ~((inputs[108]) ^ (inputs[68]));
    assign layer0_outputs[2484] = ~(inputs[71]) | (inputs[14]);
    assign layer0_outputs[2485] = (inputs[135]) | (inputs[143]);
    assign layer0_outputs[2486] = ~((inputs[208]) ^ (inputs[25]));
    assign layer0_outputs[2487] = (inputs[194]) | (inputs[166]);
    assign layer0_outputs[2488] = ~(inputs[155]) | (inputs[174]);
    assign layer0_outputs[2489] = ~(inputs[145]) | (inputs[7]);
    assign layer0_outputs[2490] = ~(inputs[42]) | (inputs[225]);
    assign layer0_outputs[2491] = inputs[41];
    assign layer0_outputs[2492] = (inputs[206]) ^ (inputs[6]);
    assign layer0_outputs[2493] = (inputs[167]) & ~(inputs[39]);
    assign layer0_outputs[2494] = inputs[40];
    assign layer0_outputs[2495] = ~((inputs[172]) | (inputs[23]));
    assign layer0_outputs[2496] = (inputs[243]) & (inputs[128]);
    assign layer0_outputs[2497] = ~(inputs[35]) | (inputs[81]);
    assign layer0_outputs[2498] = (inputs[116]) & ~(inputs[10]);
    assign layer0_outputs[2499] = ~((inputs[61]) | (inputs[133]));
    assign layer0_outputs[2500] = inputs[212];
    assign layer0_outputs[2501] = ~((inputs[99]) ^ (inputs[148]));
    assign layer0_outputs[2502] = ~(inputs[230]) | (inputs[145]);
    assign layer0_outputs[2503] = ~(inputs[123]);
    assign layer0_outputs[2504] = ~(inputs[76]) | (inputs[35]);
    assign layer0_outputs[2505] = ~((inputs[122]) ^ (inputs[249]));
    assign layer0_outputs[2506] = ~((inputs[204]) ^ (inputs[147]));
    assign layer0_outputs[2507] = (inputs[164]) & ~(inputs[177]);
    assign layer0_outputs[2508] = (inputs[192]) ^ (inputs[86]);
    assign layer0_outputs[2509] = inputs[128];
    assign layer0_outputs[2510] = 1'b0;
    assign layer0_outputs[2511] = inputs[1];
    assign layer0_outputs[2512] = (inputs[212]) & ~(inputs[79]);
    assign layer0_outputs[2513] = (inputs[228]) | (inputs[197]);
    assign layer0_outputs[2514] = inputs[173];
    assign layer0_outputs[2515] = ~((inputs[233]) | (inputs[209]));
    assign layer0_outputs[2516] = ~(inputs[200]) | (inputs[44]);
    assign layer0_outputs[2517] = ~((inputs[28]) | (inputs[138]));
    assign layer0_outputs[2518] = 1'b1;
    assign layer0_outputs[2519] = ~((inputs[235]) ^ (inputs[35]));
    assign layer0_outputs[2520] = ~(inputs[143]);
    assign layer0_outputs[2521] = ~(inputs[165]) | (inputs[6]);
    assign layer0_outputs[2522] = ~(inputs[122]) | (inputs[156]);
    assign layer0_outputs[2523] = ~((inputs[45]) & (inputs[244]));
    assign layer0_outputs[2524] = (inputs[131]) & ~(inputs[1]);
    assign layer0_outputs[2525] = inputs[147];
    assign layer0_outputs[2526] = (inputs[247]) & (inputs[235]);
    assign layer0_outputs[2527] = ~(inputs[227]);
    assign layer0_outputs[2528] = ~((inputs[34]) ^ (inputs[167]));
    assign layer0_outputs[2529] = (inputs[108]) | (inputs[172]);
    assign layer0_outputs[2530] = ~(inputs[116]);
    assign layer0_outputs[2531] = ~(inputs[50]) | (inputs[11]);
    assign layer0_outputs[2532] = inputs[214];
    assign layer0_outputs[2533] = ~(inputs[60]) | (inputs[15]);
    assign layer0_outputs[2534] = ~(inputs[33]) | (inputs[157]);
    assign layer0_outputs[2535] = (inputs[40]) | (inputs[253]);
    assign layer0_outputs[2536] = ~((inputs[123]) | (inputs[194]));
    assign layer0_outputs[2537] = (inputs[178]) | (inputs[224]);
    assign layer0_outputs[2538] = ~(inputs[174]);
    assign layer0_outputs[2539] = 1'b0;
    assign layer0_outputs[2540] = (inputs[114]) & ~(inputs[5]);
    assign layer0_outputs[2541] = (inputs[130]) ^ (inputs[47]);
    assign layer0_outputs[2542] = inputs[183];
    assign layer0_outputs[2543] = (inputs[222]) ^ (inputs[255]);
    assign layer0_outputs[2544] = ~((inputs[86]) | (inputs[28]));
    assign layer0_outputs[2545] = inputs[164];
    assign layer0_outputs[2546] = ~((inputs[174]) ^ (inputs[245]));
    assign layer0_outputs[2547] = ~(inputs[88]);
    assign layer0_outputs[2548] = (inputs[109]) | (inputs[4]);
    assign layer0_outputs[2549] = inputs[93];
    assign layer0_outputs[2550] = ~((inputs[0]) ^ (inputs[196]));
    assign layer0_outputs[2551] = (inputs[192]) & (inputs[156]);
    assign layer0_outputs[2552] = ~((inputs[191]) ^ (inputs[148]));
    assign layer0_outputs[2553] = ~((inputs[216]) | (inputs[211]));
    assign layer0_outputs[2554] = inputs[105];
    assign layer0_outputs[2555] = ~(inputs[71]) | (inputs[51]);
    assign layer0_outputs[2556] = 1'b1;
    assign layer0_outputs[2557] = (inputs[5]) ^ (inputs[68]);
    assign layer0_outputs[2558] = (inputs[123]) & ~(inputs[25]);
    assign layer0_outputs[2559] = (inputs[244]) & ~(inputs[65]);
    assign layer0_outputs[2560] = ~((inputs[217]) | (inputs[11]));
    assign layer0_outputs[2561] = (inputs[245]) | (inputs[58]);
    assign layer0_outputs[2562] = inputs[24];
    assign layer0_outputs[2563] = (inputs[169]) & ~(inputs[130]);
    assign layer0_outputs[2564] = (inputs[38]) & ~(inputs[20]);
    assign layer0_outputs[2565] = (inputs[230]) & ~(inputs[61]);
    assign layer0_outputs[2566] = inputs[109];
    assign layer0_outputs[2567] = inputs[35];
    assign layer0_outputs[2568] = (inputs[157]) & ~(inputs[19]);
    assign layer0_outputs[2569] = ~(inputs[250]);
    assign layer0_outputs[2570] = (inputs[107]) & ~(inputs[172]);
    assign layer0_outputs[2571] = ~(inputs[136]);
    assign layer0_outputs[2572] = ~(inputs[173]);
    assign layer0_outputs[2573] = (inputs[56]) & ~(inputs[125]);
    assign layer0_outputs[2574] = ~(inputs[139]) | (inputs[96]);
    assign layer0_outputs[2575] = (inputs[117]) & ~(inputs[89]);
    assign layer0_outputs[2576] = 1'b1;
    assign layer0_outputs[2577] = (inputs[90]) & ~(inputs[62]);
    assign layer0_outputs[2578] = ~((inputs[143]) ^ (inputs[46]));
    assign layer0_outputs[2579] = (inputs[114]) & ~(inputs[30]);
    assign layer0_outputs[2580] = ~((inputs[191]) ^ (inputs[211]));
    assign layer0_outputs[2581] = ~((inputs[115]) ^ (inputs[52]));
    assign layer0_outputs[2582] = ~((inputs[17]) & (inputs[0]));
    assign layer0_outputs[2583] = (inputs[49]) & (inputs[144]);
    assign layer0_outputs[2584] = (inputs[203]) & ~(inputs[200]);
    assign layer0_outputs[2585] = inputs[138];
    assign layer0_outputs[2586] = (inputs[34]) ^ (inputs[150]);
    assign layer0_outputs[2587] = (inputs[205]) | (inputs[22]);
    assign layer0_outputs[2588] = (inputs[71]) & ~(inputs[223]);
    assign layer0_outputs[2589] = ~((inputs[181]) | (inputs[190]));
    assign layer0_outputs[2590] = (inputs[83]) ^ (inputs[35]);
    assign layer0_outputs[2591] = (inputs[61]) & ~(inputs[75]);
    assign layer0_outputs[2592] = (inputs[91]) ^ (inputs[192]);
    assign layer0_outputs[2593] = (inputs[226]) & ~(inputs[203]);
    assign layer0_outputs[2594] = ~(inputs[246]) | (inputs[13]);
    assign layer0_outputs[2595] = ~((inputs[212]) & (inputs[158]));
    assign layer0_outputs[2596] = (inputs[130]) | (inputs[93]);
    assign layer0_outputs[2597] = inputs[55];
    assign layer0_outputs[2598] = ~((inputs[156]) | (inputs[94]));
    assign layer0_outputs[2599] = (inputs[151]) | (inputs[165]);
    assign layer0_outputs[2600] = (inputs[235]) & (inputs[235]);
    assign layer0_outputs[2601] = 1'b0;
    assign layer0_outputs[2602] = ~(inputs[248]);
    assign layer0_outputs[2603] = ~((inputs[240]) | (inputs[98]));
    assign layer0_outputs[2604] = ~((inputs[158]) ^ (inputs[40]));
    assign layer0_outputs[2605] = (inputs[139]) & ~(inputs[13]);
    assign layer0_outputs[2606] = ~(inputs[93]) | (inputs[28]);
    assign layer0_outputs[2607] = ~((inputs[78]) & (inputs[252]));
    assign layer0_outputs[2608] = (inputs[165]) & ~(inputs[116]);
    assign layer0_outputs[2609] = ~(inputs[207]);
    assign layer0_outputs[2610] = (inputs[167]) & ~(inputs[94]);
    assign layer0_outputs[2611] = ~(inputs[66]);
    assign layer0_outputs[2612] = ~((inputs[154]) | (inputs[129]));
    assign layer0_outputs[2613] = (inputs[118]) & ~(inputs[179]);
    assign layer0_outputs[2614] = inputs[195];
    assign layer0_outputs[2615] = (inputs[76]) ^ (inputs[178]);
    assign layer0_outputs[2616] = ~((inputs[116]) | (inputs[21]));
    assign layer0_outputs[2617] = (inputs[174]) ^ (inputs[241]);
    assign layer0_outputs[2618] = ~(inputs[248]);
    assign layer0_outputs[2619] = ~(inputs[189]);
    assign layer0_outputs[2620] = ~(inputs[108]) | (inputs[95]);
    assign layer0_outputs[2621] = ~(inputs[69]);
    assign layer0_outputs[2622] = (inputs[219]) ^ (inputs[229]);
    assign layer0_outputs[2623] = ~((inputs[244]) ^ (inputs[149]));
    assign layer0_outputs[2624] = 1'b0;
    assign layer0_outputs[2625] = ~(inputs[143]);
    assign layer0_outputs[2626] = inputs[30];
    assign layer0_outputs[2627] = (inputs[214]) | (inputs[103]);
    assign layer0_outputs[2628] = ~((inputs[182]) ^ (inputs[104]));
    assign layer0_outputs[2629] = ~((inputs[55]) | (inputs[214]));
    assign layer0_outputs[2630] = 1'b1;
    assign layer0_outputs[2631] = ~((inputs[157]) ^ (inputs[9]));
    assign layer0_outputs[2632] = (inputs[139]) & (inputs[177]);
    assign layer0_outputs[2633] = inputs[148];
    assign layer0_outputs[2634] = ~((inputs[238]) | (inputs[106]));
    assign layer0_outputs[2635] = 1'b1;
    assign layer0_outputs[2636] = inputs[251];
    assign layer0_outputs[2637] = (inputs[204]) & ~(inputs[146]);
    assign layer0_outputs[2638] = (inputs[103]) ^ (inputs[64]);
    assign layer0_outputs[2639] = (inputs[182]) | (inputs[234]);
    assign layer0_outputs[2640] = 1'b0;
    assign layer0_outputs[2641] = (inputs[87]) ^ (inputs[85]);
    assign layer0_outputs[2642] = ~((inputs[88]) | (inputs[78]));
    assign layer0_outputs[2643] = ~(inputs[151]);
    assign layer0_outputs[2644] = (inputs[1]) | (inputs[109]);
    assign layer0_outputs[2645] = (inputs[58]) ^ (inputs[192]);
    assign layer0_outputs[2646] = ~(inputs[93]);
    assign layer0_outputs[2647] = (inputs[106]) | (inputs[206]);
    assign layer0_outputs[2648] = (inputs[66]) ^ (inputs[181]);
    assign layer0_outputs[2649] = (inputs[47]) & ~(inputs[134]);
    assign layer0_outputs[2650] = inputs[148];
    assign layer0_outputs[2651] = (inputs[98]) & ~(inputs[82]);
    assign layer0_outputs[2652] = inputs[150];
    assign layer0_outputs[2653] = inputs[73];
    assign layer0_outputs[2654] = ~(inputs[93]);
    assign layer0_outputs[2655] = (inputs[72]) | (inputs[196]);
    assign layer0_outputs[2656] = (inputs[53]) & ~(inputs[11]);
    assign layer0_outputs[2657] = ~((inputs[84]) ^ (inputs[133]));
    assign layer0_outputs[2658] = ~(inputs[113]);
    assign layer0_outputs[2659] = (inputs[188]) | (inputs[75]);
    assign layer0_outputs[2660] = (inputs[162]) | (inputs[38]);
    assign layer0_outputs[2661] = (inputs[123]) | (inputs[82]);
    assign layer0_outputs[2662] = inputs[115];
    assign layer0_outputs[2663] = 1'b1;
    assign layer0_outputs[2664] = ~(inputs[218]);
    assign layer0_outputs[2665] = (inputs[152]) & (inputs[249]);
    assign layer0_outputs[2666] = ~((inputs[248]) | (inputs[10]));
    assign layer0_outputs[2667] = (inputs[64]) | (inputs[97]);
    assign layer0_outputs[2668] = ~((inputs[120]) ^ (inputs[43]));
    assign layer0_outputs[2669] = ~(inputs[152]);
    assign layer0_outputs[2670] = ~(inputs[33]) | (inputs[72]);
    assign layer0_outputs[2671] = ~((inputs[41]) | (inputs[244]));
    assign layer0_outputs[2672] = (inputs[74]) ^ (inputs[170]);
    assign layer0_outputs[2673] = (inputs[169]) & ~(inputs[253]);
    assign layer0_outputs[2674] = ~(inputs[95]);
    assign layer0_outputs[2675] = (inputs[9]) | (inputs[168]);
    assign layer0_outputs[2676] = 1'b0;
    assign layer0_outputs[2677] = ~(inputs[176]);
    assign layer0_outputs[2678] = 1'b0;
    assign layer0_outputs[2679] = (inputs[145]) ^ (inputs[170]);
    assign layer0_outputs[2680] = ~(inputs[37]) | (inputs[124]);
    assign layer0_outputs[2681] = ~(inputs[36]);
    assign layer0_outputs[2682] = ~(inputs[241]) | (inputs[19]);
    assign layer0_outputs[2683] = ~((inputs[74]) | (inputs[51]));
    assign layer0_outputs[2684] = ~((inputs[50]) ^ (inputs[99]));
    assign layer0_outputs[2685] = inputs[101];
    assign layer0_outputs[2686] = ~(inputs[61]);
    assign layer0_outputs[2687] = (inputs[29]) | (inputs[57]);
    assign layer0_outputs[2688] = (inputs[7]) | (inputs[197]);
    assign layer0_outputs[2689] = 1'b0;
    assign layer0_outputs[2690] = ~((inputs[224]) ^ (inputs[244]));
    assign layer0_outputs[2691] = ~(inputs[155]) | (inputs[219]);
    assign layer0_outputs[2692] = ~(inputs[133]) | (inputs[127]);
    assign layer0_outputs[2693] = inputs[120];
    assign layer0_outputs[2694] = (inputs[113]) | (inputs[54]);
    assign layer0_outputs[2695] = (inputs[202]) & ~(inputs[103]);
    assign layer0_outputs[2696] = inputs[86];
    assign layer0_outputs[2697] = 1'b0;
    assign layer0_outputs[2698] = (inputs[70]) & ~(inputs[216]);
    assign layer0_outputs[2699] = ~((inputs[70]) | (inputs[35]));
    assign layer0_outputs[2700] = ~((inputs[75]) ^ (inputs[45]));
    assign layer0_outputs[2701] = ~(inputs[141]) | (inputs[48]);
    assign layer0_outputs[2702] = (inputs[254]) & ~(inputs[228]);
    assign layer0_outputs[2703] = 1'b0;
    assign layer0_outputs[2704] = inputs[196];
    assign layer0_outputs[2705] = ~(inputs[225]);
    assign layer0_outputs[2706] = inputs[173];
    assign layer0_outputs[2707] = (inputs[13]) & ~(inputs[148]);
    assign layer0_outputs[2708] = ~((inputs[118]) ^ (inputs[70]));
    assign layer0_outputs[2709] = ~((inputs[220]) | (inputs[250]));
    assign layer0_outputs[2710] = ~(inputs[246]) | (inputs[144]);
    assign layer0_outputs[2711] = inputs[91];
    assign layer0_outputs[2712] = ~((inputs[232]) | (inputs[53]));
    assign layer0_outputs[2713] = ~((inputs[210]) | (inputs[147]));
    assign layer0_outputs[2714] = (inputs[146]) & ~(inputs[205]);
    assign layer0_outputs[2715] = (inputs[50]) | (inputs[223]);
    assign layer0_outputs[2716] = (inputs[54]) & ~(inputs[115]);
    assign layer0_outputs[2717] = ~(inputs[12]);
    assign layer0_outputs[2718] = ~((inputs[105]) | (inputs[243]));
    assign layer0_outputs[2719] = ~((inputs[164]) | (inputs[213]));
    assign layer0_outputs[2720] = ~((inputs[123]) & (inputs[124]));
    assign layer0_outputs[2721] = (inputs[250]) ^ (inputs[187]);
    assign layer0_outputs[2722] = ~((inputs[143]) ^ (inputs[59]));
    assign layer0_outputs[2723] = inputs[69];
    assign layer0_outputs[2724] = ~((inputs[188]) ^ (inputs[195]));
    assign layer0_outputs[2725] = ~(inputs[54]);
    assign layer0_outputs[2726] = ~((inputs[13]) | (inputs[171]));
    assign layer0_outputs[2727] = ~((inputs[28]) ^ (inputs[132]));
    assign layer0_outputs[2728] = ~(inputs[217]);
    assign layer0_outputs[2729] = (inputs[148]) | (inputs[247]);
    assign layer0_outputs[2730] = ~(inputs[12]);
    assign layer0_outputs[2731] = ~(inputs[166]);
    assign layer0_outputs[2732] = inputs[53];
    assign layer0_outputs[2733] = 1'b0;
    assign layer0_outputs[2734] = ~((inputs[149]) & (inputs[29]));
    assign layer0_outputs[2735] = (inputs[0]) ^ (inputs[245]);
    assign layer0_outputs[2736] = inputs[102];
    assign layer0_outputs[2737] = (inputs[70]) ^ (inputs[242]);
    assign layer0_outputs[2738] = (inputs[38]) | (inputs[156]);
    assign layer0_outputs[2739] = ~((inputs[240]) ^ (inputs[92]));
    assign layer0_outputs[2740] = ~((inputs[5]) ^ (inputs[131]));
    assign layer0_outputs[2741] = (inputs[132]) ^ (inputs[52]);
    assign layer0_outputs[2742] = inputs[246];
    assign layer0_outputs[2743] = ~((inputs[87]) | (inputs[132]));
    assign layer0_outputs[2744] = (inputs[35]) ^ (inputs[180]);
    assign layer0_outputs[2745] = ~((inputs[203]) & (inputs[38]));
    assign layer0_outputs[2746] = (inputs[115]) & ~(inputs[207]);
    assign layer0_outputs[2747] = inputs[206];
    assign layer0_outputs[2748] = ~(inputs[154]);
    assign layer0_outputs[2749] = inputs[121];
    assign layer0_outputs[2750] = ~((inputs[14]) & (inputs[60]));
    assign layer0_outputs[2751] = ~(inputs[207]);
    assign layer0_outputs[2752] = inputs[100];
    assign layer0_outputs[2753] = ~(inputs[184]) | (inputs[195]);
    assign layer0_outputs[2754] = ~(inputs[63]) | (inputs[65]);
    assign layer0_outputs[2755] = ~(inputs[184]);
    assign layer0_outputs[2756] = (inputs[8]) | (inputs[150]);
    assign layer0_outputs[2757] = (inputs[92]) | (inputs[225]);
    assign layer0_outputs[2758] = inputs[56];
    assign layer0_outputs[2759] = (inputs[86]) & ~(inputs[128]);
    assign layer0_outputs[2760] = inputs[173];
    assign layer0_outputs[2761] = 1'b0;
    assign layer0_outputs[2762] = ~((inputs[156]) | (inputs[170]));
    assign layer0_outputs[2763] = 1'b0;
    assign layer0_outputs[2764] = ~((inputs[137]) | (inputs[251]));
    assign layer0_outputs[2765] = ~(inputs[168]);
    assign layer0_outputs[2766] = (inputs[85]) | (inputs[137]);
    assign layer0_outputs[2767] = ~((inputs[200]) | (inputs[82]));
    assign layer0_outputs[2768] = (inputs[201]) & ~(inputs[190]);
    assign layer0_outputs[2769] = ~(inputs[103]) | (inputs[149]);
    assign layer0_outputs[2770] = ~((inputs[161]) | (inputs[216]));
    assign layer0_outputs[2771] = ~(inputs[121]) | (inputs[190]);
    assign layer0_outputs[2772] = 1'b0;
    assign layer0_outputs[2773] = inputs[161];
    assign layer0_outputs[2774] = inputs[168];
    assign layer0_outputs[2775] = ~(inputs[115]) | (inputs[200]);
    assign layer0_outputs[2776] = inputs[230];
    assign layer0_outputs[2777] = ~(inputs[37]);
    assign layer0_outputs[2778] = ~((inputs[163]) | (inputs[53]));
    assign layer0_outputs[2779] = (inputs[83]) ^ (inputs[79]);
    assign layer0_outputs[2780] = (inputs[179]) | (inputs[222]);
    assign layer0_outputs[2781] = ~(inputs[137]);
    assign layer0_outputs[2782] = (inputs[6]) & ~(inputs[25]);
    assign layer0_outputs[2783] = (inputs[67]) & (inputs[159]);
    assign layer0_outputs[2784] = ~(inputs[148]);
    assign layer0_outputs[2785] = ~((inputs[149]) ^ (inputs[254]));
    assign layer0_outputs[2786] = (inputs[27]) & ~(inputs[242]);
    assign layer0_outputs[2787] = ~(inputs[11]) | (inputs[15]);
    assign layer0_outputs[2788] = ~(inputs[164]) | (inputs[159]);
    assign layer0_outputs[2789] = (inputs[95]) | (inputs[148]);
    assign layer0_outputs[2790] = ~(inputs[164]);
    assign layer0_outputs[2791] = inputs[98];
    assign layer0_outputs[2792] = inputs[168];
    assign layer0_outputs[2793] = (inputs[253]) | (inputs[103]);
    assign layer0_outputs[2794] = ~((inputs[2]) & (inputs[75]));
    assign layer0_outputs[2795] = ~(inputs[134]) | (inputs[41]);
    assign layer0_outputs[2796] = (inputs[150]) ^ (inputs[159]);
    assign layer0_outputs[2797] = 1'b1;
    assign layer0_outputs[2798] = (inputs[136]) & ~(inputs[62]);
    assign layer0_outputs[2799] = inputs[109];
    assign layer0_outputs[2800] = (inputs[139]) ^ (inputs[109]);
    assign layer0_outputs[2801] = (inputs[92]) & ~(inputs[160]);
    assign layer0_outputs[2802] = (inputs[156]) ^ (inputs[6]);
    assign layer0_outputs[2803] = inputs[44];
    assign layer0_outputs[2804] = (inputs[223]) | (inputs[242]);
    assign layer0_outputs[2805] = ~((inputs[76]) | (inputs[75]));
    assign layer0_outputs[2806] = inputs[58];
    assign layer0_outputs[2807] = ~((inputs[116]) | (inputs[52]));
    assign layer0_outputs[2808] = ~(inputs[110]) | (inputs[175]);
    assign layer0_outputs[2809] = 1'b1;
    assign layer0_outputs[2810] = inputs[66];
    assign layer0_outputs[2811] = ~(inputs[203]) | (inputs[236]);
    assign layer0_outputs[2812] = (inputs[64]) & ~(inputs[7]);
    assign layer0_outputs[2813] = (inputs[78]) & ~(inputs[159]);
    assign layer0_outputs[2814] = (inputs[215]) & ~(inputs[242]);
    assign layer0_outputs[2815] = ~((inputs[40]) | (inputs[55]));
    assign layer0_outputs[2816] = inputs[133];
    assign layer0_outputs[2817] = ~((inputs[83]) | (inputs[249]));
    assign layer0_outputs[2818] = inputs[212];
    assign layer0_outputs[2819] = ~(inputs[60]);
    assign layer0_outputs[2820] = ~(inputs[6]) | (inputs[188]);
    assign layer0_outputs[2821] = (inputs[116]) & ~(inputs[9]);
    assign layer0_outputs[2822] = ~((inputs[177]) ^ (inputs[82]));
    assign layer0_outputs[2823] = inputs[119];
    assign layer0_outputs[2824] = ~(inputs[152]) | (inputs[84]);
    assign layer0_outputs[2825] = ~((inputs[245]) ^ (inputs[34]));
    assign layer0_outputs[2826] = inputs[167];
    assign layer0_outputs[2827] = (inputs[81]) & ~(inputs[35]);
    assign layer0_outputs[2828] = (inputs[216]) | (inputs[99]);
    assign layer0_outputs[2829] = ~((inputs[179]) ^ (inputs[244]));
    assign layer0_outputs[2830] = inputs[118];
    assign layer0_outputs[2831] = (inputs[88]) & ~(inputs[6]);
    assign layer0_outputs[2832] = inputs[250];
    assign layer0_outputs[2833] = (inputs[163]) | (inputs[78]);
    assign layer0_outputs[2834] = ~((inputs[233]) | (inputs[118]));
    assign layer0_outputs[2835] = inputs[224];
    assign layer0_outputs[2836] = ~(inputs[159]);
    assign layer0_outputs[2837] = (inputs[83]) & ~(inputs[64]);
    assign layer0_outputs[2838] = (inputs[146]) & ~(inputs[121]);
    assign layer0_outputs[2839] = ~(inputs[38]);
    assign layer0_outputs[2840] = inputs[100];
    assign layer0_outputs[2841] = (inputs[134]) & ~(inputs[30]);
    assign layer0_outputs[2842] = ~(inputs[95]) | (inputs[80]);
    assign layer0_outputs[2843] = (inputs[195]) | (inputs[177]);
    assign layer0_outputs[2844] = inputs[168];
    assign layer0_outputs[2845] = ~((inputs[31]) ^ (inputs[93]));
    assign layer0_outputs[2846] = ~(inputs[199]) | (inputs[37]);
    assign layer0_outputs[2847] = ~((inputs[159]) | (inputs[154]));
    assign layer0_outputs[2848] = (inputs[23]) | (inputs[116]);
    assign layer0_outputs[2849] = (inputs[180]) & ~(inputs[190]);
    assign layer0_outputs[2850] = 1'b1;
    assign layer0_outputs[2851] = (inputs[93]) & ~(inputs[241]);
    assign layer0_outputs[2852] = ~((inputs[161]) | (inputs[170]));
    assign layer0_outputs[2853] = inputs[55];
    assign layer0_outputs[2854] = ~((inputs[141]) | (inputs[105]));
    assign layer0_outputs[2855] = ~((inputs[223]) | (inputs[211]));
    assign layer0_outputs[2856] = ~(inputs[221]) | (inputs[31]);
    assign layer0_outputs[2857] = ~(inputs[70]);
    assign layer0_outputs[2858] = (inputs[70]) & ~(inputs[227]);
    assign layer0_outputs[2859] = (inputs[45]) | (inputs[118]);
    assign layer0_outputs[2860] = ~(inputs[108]);
    assign layer0_outputs[2861] = ~(inputs[205]);
    assign layer0_outputs[2862] = ~(inputs[56]) | (inputs[131]);
    assign layer0_outputs[2863] = ~((inputs[98]) ^ (inputs[64]));
    assign layer0_outputs[2864] = ~((inputs[81]) | (inputs[62]));
    assign layer0_outputs[2865] = ~((inputs[254]) | (inputs[15]));
    assign layer0_outputs[2866] = ~(inputs[112]);
    assign layer0_outputs[2867] = inputs[42];
    assign layer0_outputs[2868] = ~(inputs[71]) | (inputs[27]);
    assign layer0_outputs[2869] = inputs[219];
    assign layer0_outputs[2870] = ~(inputs[166]) | (inputs[98]);
    assign layer0_outputs[2871] = ~(inputs[134]) | (inputs[191]);
    assign layer0_outputs[2872] = ~(inputs[129]);
    assign layer0_outputs[2873] = ~((inputs[92]) | (inputs[202]));
    assign layer0_outputs[2874] = (inputs[101]) & (inputs[152]);
    assign layer0_outputs[2875] = (inputs[124]) | (inputs[34]);
    assign layer0_outputs[2876] = inputs[59];
    assign layer0_outputs[2877] = inputs[191];
    assign layer0_outputs[2878] = ~(inputs[226]);
    assign layer0_outputs[2879] = (inputs[165]) ^ (inputs[182]);
    assign layer0_outputs[2880] = ~(inputs[241]) | (inputs[24]);
    assign layer0_outputs[2881] = ~((inputs[115]) ^ (inputs[38]));
    assign layer0_outputs[2882] = (inputs[122]) & ~(inputs[169]);
    assign layer0_outputs[2883] = (inputs[203]) ^ (inputs[19]);
    assign layer0_outputs[2884] = ~((inputs[13]) | (inputs[164]));
    assign layer0_outputs[2885] = ~((inputs[67]) | (inputs[137]));
    assign layer0_outputs[2886] = ~((inputs[202]) & (inputs[252]));
    assign layer0_outputs[2887] = (inputs[207]) | (inputs[85]);
    assign layer0_outputs[2888] = (inputs[59]) | (inputs[161]);
    assign layer0_outputs[2889] = ~((inputs[206]) & (inputs[62]));
    assign layer0_outputs[2890] = ~((inputs[227]) & (inputs[193]));
    assign layer0_outputs[2891] = inputs[96];
    assign layer0_outputs[2892] = (inputs[140]) | (inputs[189]);
    assign layer0_outputs[2893] = ~(inputs[107]) | (inputs[244]);
    assign layer0_outputs[2894] = (inputs[76]) | (inputs[15]);
    assign layer0_outputs[2895] = ~((inputs[79]) & (inputs[221]));
    assign layer0_outputs[2896] = ~((inputs[248]) & (inputs[141]));
    assign layer0_outputs[2897] = ~(inputs[156]);
    assign layer0_outputs[2898] = 1'b1;
    assign layer0_outputs[2899] = (inputs[32]) ^ (inputs[42]);
    assign layer0_outputs[2900] = ~((inputs[127]) ^ (inputs[47]));
    assign layer0_outputs[2901] = ~(inputs[140]);
    assign layer0_outputs[2902] = (inputs[133]) | (inputs[62]);
    assign layer0_outputs[2903] = ~(inputs[230]) | (inputs[159]);
    assign layer0_outputs[2904] = (inputs[231]) & ~(inputs[219]);
    assign layer0_outputs[2905] = inputs[84];
    assign layer0_outputs[2906] = ~(inputs[65]) | (inputs[55]);
    assign layer0_outputs[2907] = ~((inputs[140]) | (inputs[170]));
    assign layer0_outputs[2908] = inputs[251];
    assign layer0_outputs[2909] = inputs[214];
    assign layer0_outputs[2910] = (inputs[154]) & ~(inputs[3]);
    assign layer0_outputs[2911] = ~((inputs[47]) & (inputs[130]));
    assign layer0_outputs[2912] = ~(inputs[119]);
    assign layer0_outputs[2913] = ~((inputs[210]) ^ (inputs[74]));
    assign layer0_outputs[2914] = ~((inputs[88]) | (inputs[227]));
    assign layer0_outputs[2915] = ~(inputs[97]);
    assign layer0_outputs[2916] = inputs[101];
    assign layer0_outputs[2917] = (inputs[211]) & ~(inputs[56]);
    assign layer0_outputs[2918] = ~(inputs[88]);
    assign layer0_outputs[2919] = ~(inputs[107]) | (inputs[8]);
    assign layer0_outputs[2920] = (inputs[182]) & ~(inputs[83]);
    assign layer0_outputs[2921] = (inputs[140]) | (inputs[25]);
    assign layer0_outputs[2922] = (inputs[42]) & ~(inputs[213]);
    assign layer0_outputs[2923] = inputs[177];
    assign layer0_outputs[2924] = ~((inputs[243]) ^ (inputs[108]));
    assign layer0_outputs[2925] = ~(inputs[196]);
    assign layer0_outputs[2926] = ~(inputs[43]) | (inputs[243]);
    assign layer0_outputs[2927] = (inputs[190]) | (inputs[253]);
    assign layer0_outputs[2928] = ~((inputs[39]) | (inputs[91]));
    assign layer0_outputs[2929] = ~((inputs[171]) | (inputs[123]));
    assign layer0_outputs[2930] = 1'b0;
    assign layer0_outputs[2931] = ~((inputs[184]) | (inputs[235]));
    assign layer0_outputs[2932] = (inputs[126]) ^ (inputs[159]);
    assign layer0_outputs[2933] = ~(inputs[148]);
    assign layer0_outputs[2934] = ~(inputs[42]);
    assign layer0_outputs[2935] = ~((inputs[155]) ^ (inputs[112]));
    assign layer0_outputs[2936] = ~((inputs[30]) | (inputs[117]));
    assign layer0_outputs[2937] = ~(inputs[70]);
    assign layer0_outputs[2938] = (inputs[8]) & (inputs[98]);
    assign layer0_outputs[2939] = ~(inputs[204]);
    assign layer0_outputs[2940] = ~(inputs[9]) | (inputs[18]);
    assign layer0_outputs[2941] = ~((inputs[177]) ^ (inputs[129]));
    assign layer0_outputs[2942] = ~((inputs[218]) ^ (inputs[212]));
    assign layer0_outputs[2943] = ~(inputs[105]) | (inputs[155]);
    assign layer0_outputs[2944] = ~((inputs[104]) ^ (inputs[254]));
    assign layer0_outputs[2945] = (inputs[149]) & ~(inputs[67]);
    assign layer0_outputs[2946] = (inputs[160]) & ~(inputs[174]);
    assign layer0_outputs[2947] = (inputs[195]) | (inputs[124]);
    assign layer0_outputs[2948] = ~(inputs[157]) | (inputs[229]);
    assign layer0_outputs[2949] = ~(inputs[14]);
    assign layer0_outputs[2950] = (inputs[154]) ^ (inputs[53]);
    assign layer0_outputs[2951] = ~((inputs[140]) & (inputs[189]));
    assign layer0_outputs[2952] = ~(inputs[118]) | (inputs[100]);
    assign layer0_outputs[2953] = (inputs[142]) ^ (inputs[60]);
    assign layer0_outputs[2954] = ~((inputs[126]) | (inputs[75]));
    assign layer0_outputs[2955] = (inputs[225]) ^ (inputs[210]);
    assign layer0_outputs[2956] = ~(inputs[97]);
    assign layer0_outputs[2957] = ~((inputs[66]) | (inputs[40]));
    assign layer0_outputs[2958] = ~(inputs[238]);
    assign layer0_outputs[2959] = (inputs[89]) | (inputs[36]);
    assign layer0_outputs[2960] = (inputs[66]) | (inputs[205]);
    assign layer0_outputs[2961] = inputs[136];
    assign layer0_outputs[2962] = inputs[64];
    assign layer0_outputs[2963] = inputs[184];
    assign layer0_outputs[2964] = ~(inputs[230]);
    assign layer0_outputs[2965] = (inputs[36]) & ~(inputs[131]);
    assign layer0_outputs[2966] = ~(inputs[86]);
    assign layer0_outputs[2967] = (inputs[238]) | (inputs[20]);
    assign layer0_outputs[2968] = (inputs[248]) & ~(inputs[208]);
    assign layer0_outputs[2969] = (inputs[245]) & (inputs[70]);
    assign layer0_outputs[2970] = (inputs[218]) | (inputs[100]);
    assign layer0_outputs[2971] = (inputs[170]) ^ (inputs[239]);
    assign layer0_outputs[2972] = (inputs[229]) | (inputs[74]);
    assign layer0_outputs[2973] = ~(inputs[184]) | (inputs[229]);
    assign layer0_outputs[2974] = (inputs[182]) ^ (inputs[164]);
    assign layer0_outputs[2975] = ~((inputs[173]) | (inputs[24]));
    assign layer0_outputs[2976] = ~(inputs[52]);
    assign layer0_outputs[2977] = ~((inputs[180]) & (inputs[91]));
    assign layer0_outputs[2978] = 1'b0;
    assign layer0_outputs[2979] = (inputs[135]) | (inputs[150]);
    assign layer0_outputs[2980] = (inputs[79]) | (inputs[145]);
    assign layer0_outputs[2981] = 1'b0;
    assign layer0_outputs[2982] = (inputs[95]) & ~(inputs[248]);
    assign layer0_outputs[2983] = inputs[213];
    assign layer0_outputs[2984] = 1'b0;
    assign layer0_outputs[2985] = 1'b1;
    assign layer0_outputs[2986] = (inputs[132]) & ~(inputs[191]);
    assign layer0_outputs[2987] = ~(inputs[201]) | (inputs[36]);
    assign layer0_outputs[2988] = ~((inputs[73]) ^ (inputs[128]));
    assign layer0_outputs[2989] = ~(inputs[195]);
    assign layer0_outputs[2990] = (inputs[184]) ^ (inputs[90]);
    assign layer0_outputs[2991] = ~((inputs[227]) ^ (inputs[9]));
    assign layer0_outputs[2992] = (inputs[103]) | (inputs[62]);
    assign layer0_outputs[2993] = 1'b0;
    assign layer0_outputs[2994] = ~((inputs[37]) ^ (inputs[4]));
    assign layer0_outputs[2995] = (inputs[185]) | (inputs[11]);
    assign layer0_outputs[2996] = (inputs[187]) ^ (inputs[24]);
    assign layer0_outputs[2997] = (inputs[163]) | (inputs[77]);
    assign layer0_outputs[2998] = (inputs[226]) ^ (inputs[86]);
    assign layer0_outputs[2999] = (inputs[152]) | (inputs[8]);
    assign layer0_outputs[3000] = ~(inputs[86]);
    assign layer0_outputs[3001] = ~((inputs[155]) | (inputs[65]));
    assign layer0_outputs[3002] = ~((inputs[243]) & (inputs[193]));
    assign layer0_outputs[3003] = (inputs[142]) ^ (inputs[41]);
    assign layer0_outputs[3004] = (inputs[229]) & ~(inputs[25]);
    assign layer0_outputs[3005] = ~(inputs[120]);
    assign layer0_outputs[3006] = inputs[173];
    assign layer0_outputs[3007] = (inputs[156]) & ~(inputs[149]);
    assign layer0_outputs[3008] = ~(inputs[217]) | (inputs[33]);
    assign layer0_outputs[3009] = ~(inputs[233]) | (inputs[191]);
    assign layer0_outputs[3010] = ~(inputs[125]) | (inputs[239]);
    assign layer0_outputs[3011] = (inputs[29]) | (inputs[123]);
    assign layer0_outputs[3012] = ~((inputs[31]) ^ (inputs[218]));
    assign layer0_outputs[3013] = ~(inputs[198]);
    assign layer0_outputs[3014] = (inputs[231]) ^ (inputs[33]);
    assign layer0_outputs[3015] = (inputs[36]) | (inputs[132]);
    assign layer0_outputs[3016] = inputs[203];
    assign layer0_outputs[3017] = ~((inputs[181]) | (inputs[23]));
    assign layer0_outputs[3018] = 1'b0;
    assign layer0_outputs[3019] = 1'b1;
    assign layer0_outputs[3020] = (inputs[200]) & ~(inputs[85]);
    assign layer0_outputs[3021] = ~(inputs[253]) | (inputs[129]);
    assign layer0_outputs[3022] = ~(inputs[200]);
    assign layer0_outputs[3023] = inputs[107];
    assign layer0_outputs[3024] = ~((inputs[198]) | (inputs[213]));
    assign layer0_outputs[3025] = ~(inputs[180]) | (inputs[226]);
    assign layer0_outputs[3026] = (inputs[50]) ^ (inputs[64]);
    assign layer0_outputs[3027] = (inputs[184]) ^ (inputs[50]);
    assign layer0_outputs[3028] = (inputs[228]) | (inputs[226]);
    assign layer0_outputs[3029] = (inputs[199]) | (inputs[21]);
    assign layer0_outputs[3030] = inputs[124];
    assign layer0_outputs[3031] = (inputs[208]) ^ (inputs[4]);
    assign layer0_outputs[3032] = 1'b0;
    assign layer0_outputs[3033] = (inputs[132]) & ~(inputs[126]);
    assign layer0_outputs[3034] = ~((inputs[146]) | (inputs[106]));
    assign layer0_outputs[3035] = 1'b1;
    assign layer0_outputs[3036] = ~((inputs[7]) ^ (inputs[73]));
    assign layer0_outputs[3037] = ~(inputs[69]) | (inputs[241]);
    assign layer0_outputs[3038] = ~((inputs[213]) | (inputs[49]));
    assign layer0_outputs[3039] = (inputs[112]) | (inputs[151]);
    assign layer0_outputs[3040] = ~(inputs[105]);
    assign layer0_outputs[3041] = ~((inputs[8]) ^ (inputs[119]));
    assign layer0_outputs[3042] = ~((inputs[46]) ^ (inputs[70]));
    assign layer0_outputs[3043] = (inputs[9]) ^ (inputs[182]);
    assign layer0_outputs[3044] = ~(inputs[90]);
    assign layer0_outputs[3045] = ~((inputs[106]) | (inputs[94]));
    assign layer0_outputs[3046] = inputs[167];
    assign layer0_outputs[3047] = (inputs[130]) | (inputs[147]);
    assign layer0_outputs[3048] = inputs[210];
    assign layer0_outputs[3049] = 1'b0;
    assign layer0_outputs[3050] = (inputs[72]) ^ (inputs[255]);
    assign layer0_outputs[3051] = ~(inputs[137]) | (inputs[62]);
    assign layer0_outputs[3052] = ~((inputs[179]) ^ (inputs[34]));
    assign layer0_outputs[3053] = ~((inputs[131]) | (inputs[228]));
    assign layer0_outputs[3054] = ~(inputs[236]);
    assign layer0_outputs[3055] = (inputs[106]) ^ (inputs[226]);
    assign layer0_outputs[3056] = (inputs[233]) & ~(inputs[211]);
    assign layer0_outputs[3057] = ~((inputs[160]) | (inputs[110]));
    assign layer0_outputs[3058] = ~((inputs[225]) ^ (inputs[37]));
    assign layer0_outputs[3059] = ~((inputs[181]) | (inputs[220]));
    assign layer0_outputs[3060] = ~(inputs[164]);
    assign layer0_outputs[3061] = ~((inputs[224]) | (inputs[18]));
    assign layer0_outputs[3062] = (inputs[41]) | (inputs[197]);
    assign layer0_outputs[3063] = ~((inputs[173]) | (inputs[68]));
    assign layer0_outputs[3064] = (inputs[15]) ^ (inputs[1]);
    assign layer0_outputs[3065] = ~(inputs[86]);
    assign layer0_outputs[3066] = ~((inputs[65]) | (inputs[99]));
    assign layer0_outputs[3067] = (inputs[174]) ^ (inputs[191]);
    assign layer0_outputs[3068] = ~(inputs[166]);
    assign layer0_outputs[3069] = (inputs[66]) | (inputs[55]);
    assign layer0_outputs[3070] = ~(inputs[230]);
    assign layer0_outputs[3071] = ~(inputs[119]);
    assign layer0_outputs[3072] = ~(inputs[217]) | (inputs[192]);
    assign layer0_outputs[3073] = ~(inputs[136]);
    assign layer0_outputs[3074] = ~((inputs[226]) & (inputs[99]));
    assign layer0_outputs[3075] = ~(inputs[185]) | (inputs[25]);
    assign layer0_outputs[3076] = 1'b1;
    assign layer0_outputs[3077] = inputs[4];
    assign layer0_outputs[3078] = inputs[151];
    assign layer0_outputs[3079] = (inputs[90]) & ~(inputs[177]);
    assign layer0_outputs[3080] = ~((inputs[230]) | (inputs[172]));
    assign layer0_outputs[3081] = ~(inputs[38]);
    assign layer0_outputs[3082] = (inputs[204]) & (inputs[164]);
    assign layer0_outputs[3083] = ~((inputs[221]) & (inputs[109]));
    assign layer0_outputs[3084] = ~(inputs[90]) | (inputs[254]);
    assign layer0_outputs[3085] = inputs[181];
    assign layer0_outputs[3086] = ~(inputs[21]) | (inputs[8]);
    assign layer0_outputs[3087] = ~(inputs[52]) | (inputs[19]);
    assign layer0_outputs[3088] = (inputs[5]) | (inputs[233]);
    assign layer0_outputs[3089] = (inputs[61]) | (inputs[232]);
    assign layer0_outputs[3090] = ~(inputs[125]);
    assign layer0_outputs[3091] = (inputs[195]) | (inputs[156]);
    assign layer0_outputs[3092] = 1'b1;
    assign layer0_outputs[3093] = ~(inputs[93]) | (inputs[219]);
    assign layer0_outputs[3094] = (inputs[57]) | (inputs[178]);
    assign layer0_outputs[3095] = inputs[120];
    assign layer0_outputs[3096] = ~(inputs[25]) | (inputs[49]);
    assign layer0_outputs[3097] = ~(inputs[150]) | (inputs[174]);
    assign layer0_outputs[3098] = inputs[139];
    assign layer0_outputs[3099] = ~(inputs[79]);
    assign layer0_outputs[3100] = ~((inputs[123]) | (inputs[183]));
    assign layer0_outputs[3101] = inputs[201];
    assign layer0_outputs[3102] = (inputs[3]) | (inputs[41]);
    assign layer0_outputs[3103] = (inputs[150]) & ~(inputs[214]);
    assign layer0_outputs[3104] = ~((inputs[1]) | (inputs[198]));
    assign layer0_outputs[3105] = inputs[117];
    assign layer0_outputs[3106] = 1'b0;
    assign layer0_outputs[3107] = 1'b1;
    assign layer0_outputs[3108] = (inputs[249]) ^ (inputs[68]);
    assign layer0_outputs[3109] = inputs[255];
    assign layer0_outputs[3110] = (inputs[194]) ^ (inputs[207]);
    assign layer0_outputs[3111] = ~((inputs[206]) & (inputs[67]));
    assign layer0_outputs[3112] = ~((inputs[177]) | (inputs[228]));
    assign layer0_outputs[3113] = (inputs[62]) ^ (inputs[82]);
    assign layer0_outputs[3114] = (inputs[212]) ^ (inputs[250]);
    assign layer0_outputs[3115] = ~((inputs[174]) | (inputs[6]));
    assign layer0_outputs[3116] = ~(inputs[250]);
    assign layer0_outputs[3117] = ~(inputs[171]) | (inputs[255]);
    assign layer0_outputs[3118] = inputs[197];
    assign layer0_outputs[3119] = (inputs[211]) ^ (inputs[156]);
    assign layer0_outputs[3120] = (inputs[232]) & ~(inputs[209]);
    assign layer0_outputs[3121] = 1'b1;
    assign layer0_outputs[3122] = (inputs[52]) ^ (inputs[81]);
    assign layer0_outputs[3123] = (inputs[118]) ^ (inputs[38]);
    assign layer0_outputs[3124] = (inputs[168]) ^ (inputs[105]);
    assign layer0_outputs[3125] = ~(inputs[212]);
    assign layer0_outputs[3126] = (inputs[196]) ^ (inputs[54]);
    assign layer0_outputs[3127] = (inputs[68]) & ~(inputs[37]);
    assign layer0_outputs[3128] = (inputs[104]) & ~(inputs[77]);
    assign layer0_outputs[3129] = (inputs[86]) & ~(inputs[20]);
    assign layer0_outputs[3130] = ~((inputs[169]) | (inputs[26]));
    assign layer0_outputs[3131] = (inputs[19]) | (inputs[190]);
    assign layer0_outputs[3132] = ~(inputs[152]);
    assign layer0_outputs[3133] = ~(inputs[134]) | (inputs[28]);
    assign layer0_outputs[3134] = ~((inputs[248]) | (inputs[174]));
    assign layer0_outputs[3135] = ~(inputs[5]);
    assign layer0_outputs[3136] = (inputs[162]) & ~(inputs[28]);
    assign layer0_outputs[3137] = ~(inputs[78]) | (inputs[36]);
    assign layer0_outputs[3138] = ~((inputs[83]) & (inputs[184]));
    assign layer0_outputs[3139] = (inputs[76]) | (inputs[190]);
    assign layer0_outputs[3140] = (inputs[199]) | (inputs[113]);
    assign layer0_outputs[3141] = ~(inputs[104]) | (inputs[29]);
    assign layer0_outputs[3142] = (inputs[242]) ^ (inputs[41]);
    assign layer0_outputs[3143] = ~(inputs[186]) | (inputs[27]);
    assign layer0_outputs[3144] = (inputs[118]) & (inputs[135]);
    assign layer0_outputs[3145] = (inputs[125]) & ~(inputs[253]);
    assign layer0_outputs[3146] = inputs[210];
    assign layer0_outputs[3147] = ~((inputs[144]) ^ (inputs[121]));
    assign layer0_outputs[3148] = (inputs[215]) & ~(inputs[45]);
    assign layer0_outputs[3149] = ~((inputs[110]) | (inputs[97]));
    assign layer0_outputs[3150] = ~(inputs[51]);
    assign layer0_outputs[3151] = ~((inputs[14]) & (inputs[179]));
    assign layer0_outputs[3152] = ~(inputs[214]) | (inputs[69]);
    assign layer0_outputs[3153] = (inputs[172]) | (inputs[17]);
    assign layer0_outputs[3154] = 1'b0;
    assign layer0_outputs[3155] = ~(inputs[208]) | (inputs[85]);
    assign layer0_outputs[3156] = ~(inputs[31]);
    assign layer0_outputs[3157] = inputs[151];
    assign layer0_outputs[3158] = (inputs[33]) & ~(inputs[94]);
    assign layer0_outputs[3159] = (inputs[223]) | (inputs[23]);
    assign layer0_outputs[3160] = (inputs[96]) ^ (inputs[180]);
    assign layer0_outputs[3161] = ~(inputs[27]);
    assign layer0_outputs[3162] = ~(inputs[193]);
    assign layer0_outputs[3163] = inputs[197];
    assign layer0_outputs[3164] = ~(inputs[114]) | (inputs[27]);
    assign layer0_outputs[3165] = inputs[149];
    assign layer0_outputs[3166] = ~(inputs[18]) | (inputs[127]);
    assign layer0_outputs[3167] = 1'b0;
    assign layer0_outputs[3168] = (inputs[24]) & ~(inputs[95]);
    assign layer0_outputs[3169] = inputs[102];
    assign layer0_outputs[3170] = inputs[245];
    assign layer0_outputs[3171] = (inputs[13]) & ~(inputs[146]);
    assign layer0_outputs[3172] = ~(inputs[226]) | (inputs[16]);
    assign layer0_outputs[3173] = ~(inputs[19]);
    assign layer0_outputs[3174] = (inputs[252]) ^ (inputs[229]);
    assign layer0_outputs[3175] = ~((inputs[133]) ^ (inputs[96]));
    assign layer0_outputs[3176] = ~(inputs[178]);
    assign layer0_outputs[3177] = inputs[78];
    assign layer0_outputs[3178] = (inputs[174]) | (inputs[140]);
    assign layer0_outputs[3179] = inputs[36];
    assign layer0_outputs[3180] = (inputs[185]) & ~(inputs[238]);
    assign layer0_outputs[3181] = ~((inputs[199]) | (inputs[187]));
    assign layer0_outputs[3182] = inputs[216];
    assign layer0_outputs[3183] = ~((inputs[58]) ^ (inputs[55]));
    assign layer0_outputs[3184] = (inputs[77]) & ~(inputs[247]);
    assign layer0_outputs[3185] = inputs[149];
    assign layer0_outputs[3186] = 1'b0;
    assign layer0_outputs[3187] = (inputs[71]) ^ (inputs[173]);
    assign layer0_outputs[3188] = ~((inputs[223]) & (inputs[0]));
    assign layer0_outputs[3189] = ~((inputs[141]) | (inputs[147]));
    assign layer0_outputs[3190] = 1'b1;
    assign layer0_outputs[3191] = (inputs[224]) & ~(inputs[63]);
    assign layer0_outputs[3192] = (inputs[183]) & ~(inputs[211]);
    assign layer0_outputs[3193] = ~(inputs[202]);
    assign layer0_outputs[3194] = ~(inputs[178]);
    assign layer0_outputs[3195] = 1'b1;
    assign layer0_outputs[3196] = (inputs[202]) ^ (inputs[185]);
    assign layer0_outputs[3197] = ~(inputs[36]) | (inputs[24]);
    assign layer0_outputs[3198] = (inputs[76]) & ~(inputs[244]);
    assign layer0_outputs[3199] = ~(inputs[57]);
    assign layer0_outputs[3200] = ~(inputs[165]);
    assign layer0_outputs[3201] = ~(inputs[217]);
    assign layer0_outputs[3202] = ~(inputs[66]) | (inputs[204]);
    assign layer0_outputs[3203] = ~((inputs[3]) ^ (inputs[76]));
    assign layer0_outputs[3204] = (inputs[105]) | (inputs[142]);
    assign layer0_outputs[3205] = ~(inputs[242]) | (inputs[254]);
    assign layer0_outputs[3206] = (inputs[178]) | (inputs[159]);
    assign layer0_outputs[3207] = (inputs[255]) & ~(inputs[226]);
    assign layer0_outputs[3208] = (inputs[163]) & ~(inputs[67]);
    assign layer0_outputs[3209] = (inputs[207]) & ~(inputs[2]);
    assign layer0_outputs[3210] = inputs[212];
    assign layer0_outputs[3211] = inputs[151];
    assign layer0_outputs[3212] = (inputs[185]) | (inputs[190]);
    assign layer0_outputs[3213] = (inputs[21]) & ~(inputs[40]);
    assign layer0_outputs[3214] = inputs[142];
    assign layer0_outputs[3215] = 1'b0;
    assign layer0_outputs[3216] = (inputs[86]) | (inputs[247]);
    assign layer0_outputs[3217] = (inputs[154]) ^ (inputs[69]);
    assign layer0_outputs[3218] = ~((inputs[93]) | (inputs[189]));
    assign layer0_outputs[3219] = (inputs[200]) & ~(inputs[36]);
    assign layer0_outputs[3220] = (inputs[59]) ^ (inputs[71]);
    assign layer0_outputs[3221] = 1'b0;
    assign layer0_outputs[3222] = (inputs[213]) & ~(inputs[188]);
    assign layer0_outputs[3223] = ~((inputs[117]) | (inputs[17]));
    assign layer0_outputs[3224] = ~((inputs[140]) | (inputs[184]));
    assign layer0_outputs[3225] = ~(inputs[136]);
    assign layer0_outputs[3226] = ~(inputs[143]);
    assign layer0_outputs[3227] = inputs[197];
    assign layer0_outputs[3228] = inputs[47];
    assign layer0_outputs[3229] = inputs[43];
    assign layer0_outputs[3230] = ~((inputs[128]) | (inputs[125]));
    assign layer0_outputs[3231] = 1'b0;
    assign layer0_outputs[3232] = ~((inputs[160]) | (inputs[23]));
    assign layer0_outputs[3233] = inputs[74];
    assign layer0_outputs[3234] = ~((inputs[43]) & (inputs[254]));
    assign layer0_outputs[3235] = ~(inputs[196]);
    assign layer0_outputs[3236] = (inputs[187]) & ~(inputs[229]);
    assign layer0_outputs[3237] = (inputs[214]) & ~(inputs[51]);
    assign layer0_outputs[3238] = (inputs[30]) | (inputs[231]);
    assign layer0_outputs[3239] = ~((inputs[85]) ^ (inputs[249]));
    assign layer0_outputs[3240] = (inputs[92]) & ~(inputs[1]);
    assign layer0_outputs[3241] = ~(inputs[139]) | (inputs[97]);
    assign layer0_outputs[3242] = (inputs[195]) | (inputs[209]);
    assign layer0_outputs[3243] = ~((inputs[233]) | (inputs[221]));
    assign layer0_outputs[3244] = inputs[191];
    assign layer0_outputs[3245] = ~((inputs[8]) ^ (inputs[128]));
    assign layer0_outputs[3246] = ~((inputs[128]) ^ (inputs[123]));
    assign layer0_outputs[3247] = ~((inputs[222]) ^ (inputs[51]));
    assign layer0_outputs[3248] = ~(inputs[93]);
    assign layer0_outputs[3249] = ~(inputs[155]);
    assign layer0_outputs[3250] = ~((inputs[107]) ^ (inputs[105]));
    assign layer0_outputs[3251] = ~((inputs[199]) ^ (inputs[50]));
    assign layer0_outputs[3252] = ~((inputs[10]) | (inputs[28]));
    assign layer0_outputs[3253] = ~(inputs[177]);
    assign layer0_outputs[3254] = inputs[144];
    assign layer0_outputs[3255] = ~(inputs[183]);
    assign layer0_outputs[3256] = inputs[149];
    assign layer0_outputs[3257] = ~((inputs[187]) ^ (inputs[71]));
    assign layer0_outputs[3258] = ~(inputs[199]) | (inputs[161]);
    assign layer0_outputs[3259] = (inputs[142]) & (inputs[49]);
    assign layer0_outputs[3260] = (inputs[255]) | (inputs[202]);
    assign layer0_outputs[3261] = (inputs[125]) | (inputs[108]);
    assign layer0_outputs[3262] = (inputs[82]) & ~(inputs[209]);
    assign layer0_outputs[3263] = ~(inputs[25]);
    assign layer0_outputs[3264] = ~((inputs[150]) | (inputs[21]));
    assign layer0_outputs[3265] = (inputs[37]) | (inputs[57]);
    assign layer0_outputs[3266] = inputs[22];
    assign layer0_outputs[3267] = (inputs[168]) & ~(inputs[48]);
    assign layer0_outputs[3268] = ~(inputs[86]) | (inputs[173]);
    assign layer0_outputs[3269] = inputs[105];
    assign layer0_outputs[3270] = (inputs[216]) & ~(inputs[9]);
    assign layer0_outputs[3271] = ~((inputs[13]) & (inputs[240]));
    assign layer0_outputs[3272] = ~(inputs[38]) | (inputs[241]);
    assign layer0_outputs[3273] = (inputs[14]) & ~(inputs[26]);
    assign layer0_outputs[3274] = inputs[87];
    assign layer0_outputs[3275] = inputs[208];
    assign layer0_outputs[3276] = (inputs[129]) | (inputs[186]);
    assign layer0_outputs[3277] = (inputs[20]) | (inputs[88]);
    assign layer0_outputs[3278] = (inputs[235]) | (inputs[115]);
    assign layer0_outputs[3279] = (inputs[138]) ^ (inputs[108]);
    assign layer0_outputs[3280] = (inputs[37]) ^ (inputs[234]);
    assign layer0_outputs[3281] = (inputs[215]) & ~(inputs[20]);
    assign layer0_outputs[3282] = ~(inputs[63]);
    assign layer0_outputs[3283] = (inputs[140]) ^ (inputs[10]);
    assign layer0_outputs[3284] = 1'b1;
    assign layer0_outputs[3285] = ~((inputs[28]) ^ (inputs[239]));
    assign layer0_outputs[3286] = ~(inputs[103]);
    assign layer0_outputs[3287] = ~(inputs[134]);
    assign layer0_outputs[3288] = ~((inputs[178]) | (inputs[174]));
    assign layer0_outputs[3289] = inputs[108];
    assign layer0_outputs[3290] = inputs[29];
    assign layer0_outputs[3291] = (inputs[156]) | (inputs[97]);
    assign layer0_outputs[3292] = (inputs[196]) | (inputs[197]);
    assign layer0_outputs[3293] = inputs[164];
    assign layer0_outputs[3294] = ~(inputs[160]);
    assign layer0_outputs[3295] = ~(inputs[44]) | (inputs[176]);
    assign layer0_outputs[3296] = ~((inputs[110]) ^ (inputs[11]));
    assign layer0_outputs[3297] = ~((inputs[242]) ^ (inputs[72]));
    assign layer0_outputs[3298] = ~((inputs[152]) & (inputs[141]));
    assign layer0_outputs[3299] = ~((inputs[100]) ^ (inputs[70]));
    assign layer0_outputs[3300] = ~((inputs[33]) ^ (inputs[30]));
    assign layer0_outputs[3301] = ~(inputs[59]) | (inputs[29]);
    assign layer0_outputs[3302] = ~((inputs[147]) ^ (inputs[24]));
    assign layer0_outputs[3303] = ~(inputs[12]);
    assign layer0_outputs[3304] = (inputs[86]) & ~(inputs[57]);
    assign layer0_outputs[3305] = 1'b1;
    assign layer0_outputs[3306] = inputs[102];
    assign layer0_outputs[3307] = inputs[20];
    assign layer0_outputs[3308] = (inputs[86]) ^ (inputs[117]);
    assign layer0_outputs[3309] = ~(inputs[27]);
    assign layer0_outputs[3310] = ~(inputs[137]);
    assign layer0_outputs[3311] = inputs[73];
    assign layer0_outputs[3312] = ~(inputs[85]);
    assign layer0_outputs[3313] = 1'b1;
    assign layer0_outputs[3314] = (inputs[191]) & ~(inputs[33]);
    assign layer0_outputs[3315] = ~((inputs[130]) & (inputs[162]));
    assign layer0_outputs[3316] = inputs[53];
    assign layer0_outputs[3317] = (inputs[98]) & (inputs[226]);
    assign layer0_outputs[3318] = (inputs[40]) ^ (inputs[30]);
    assign layer0_outputs[3319] = (inputs[95]) | (inputs[83]);
    assign layer0_outputs[3320] = (inputs[65]) & ~(inputs[78]);
    assign layer0_outputs[3321] = (inputs[45]) ^ (inputs[36]);
    assign layer0_outputs[3322] = (inputs[49]) ^ (inputs[61]);
    assign layer0_outputs[3323] = (inputs[177]) & ~(inputs[239]);
    assign layer0_outputs[3324] = ~(inputs[118]) | (inputs[2]);
    assign layer0_outputs[3325] = (inputs[17]) & (inputs[31]);
    assign layer0_outputs[3326] = inputs[158];
    assign layer0_outputs[3327] = ~((inputs[250]) | (inputs[25]));
    assign layer0_outputs[3328] = inputs[186];
    assign layer0_outputs[3329] = (inputs[83]) | (inputs[192]);
    assign layer0_outputs[3330] = ~((inputs[118]) | (inputs[110]));
    assign layer0_outputs[3331] = ~((inputs[139]) | (inputs[10]));
    assign layer0_outputs[3332] = inputs[41];
    assign layer0_outputs[3333] = (inputs[143]) & (inputs[20]);
    assign layer0_outputs[3334] = ~((inputs[52]) ^ (inputs[65]));
    assign layer0_outputs[3335] = (inputs[253]) | (inputs[85]);
    assign layer0_outputs[3336] = (inputs[117]) & ~(inputs[247]);
    assign layer0_outputs[3337] = ~(inputs[169]);
    assign layer0_outputs[3338] = (inputs[108]) & ~(inputs[64]);
    assign layer0_outputs[3339] = ~((inputs[209]) ^ (inputs[151]));
    assign layer0_outputs[3340] = ~(inputs[210]) | (inputs[68]);
    assign layer0_outputs[3341] = ~(inputs[74]);
    assign layer0_outputs[3342] = inputs[125];
    assign layer0_outputs[3343] = ~((inputs[159]) ^ (inputs[142]));
    assign layer0_outputs[3344] = (inputs[101]) ^ (inputs[223]);
    assign layer0_outputs[3345] = (inputs[175]) ^ (inputs[116]);
    assign layer0_outputs[3346] = ~(inputs[77]);
    assign layer0_outputs[3347] = ~((inputs[171]) ^ (inputs[71]));
    assign layer0_outputs[3348] = ~(inputs[236]) | (inputs[33]);
    assign layer0_outputs[3349] = (inputs[209]) ^ (inputs[238]);
    assign layer0_outputs[3350] = (inputs[217]) ^ (inputs[78]);
    assign layer0_outputs[3351] = 1'b1;
    assign layer0_outputs[3352] = (inputs[14]) ^ (inputs[235]);
    assign layer0_outputs[3353] = (inputs[230]) | (inputs[113]);
    assign layer0_outputs[3354] = (inputs[1]) & (inputs[28]);
    assign layer0_outputs[3355] = ~(inputs[239]) | (inputs[39]);
    assign layer0_outputs[3356] = inputs[63];
    assign layer0_outputs[3357] = ~(inputs[230]);
    assign layer0_outputs[3358] = (inputs[67]) | (inputs[149]);
    assign layer0_outputs[3359] = ~((inputs[122]) | (inputs[35]));
    assign layer0_outputs[3360] = ~(inputs[228]);
    assign layer0_outputs[3361] = (inputs[156]) | (inputs[141]);
    assign layer0_outputs[3362] = (inputs[145]) | (inputs[250]);
    assign layer0_outputs[3363] = ~((inputs[191]) & (inputs[108]));
    assign layer0_outputs[3364] = (inputs[188]) ^ (inputs[79]);
    assign layer0_outputs[3365] = ~((inputs[194]) | (inputs[119]));
    assign layer0_outputs[3366] = ~((inputs[111]) | (inputs[50]));
    assign layer0_outputs[3367] = (inputs[65]) | (inputs[158]);
    assign layer0_outputs[3368] = ~((inputs[226]) ^ (inputs[87]));
    assign layer0_outputs[3369] = inputs[58];
    assign layer0_outputs[3370] = (inputs[229]) ^ (inputs[139]);
    assign layer0_outputs[3371] = inputs[166];
    assign layer0_outputs[3372] = ~((inputs[78]) ^ (inputs[3]));
    assign layer0_outputs[3373] = 1'b1;
    assign layer0_outputs[3374] = ~(inputs[192]) | (inputs[240]);
    assign layer0_outputs[3375] = (inputs[55]) & ~(inputs[235]);
    assign layer0_outputs[3376] = ~((inputs[215]) | (inputs[246]));
    assign layer0_outputs[3377] = inputs[250];
    assign layer0_outputs[3378] = ~(inputs[135]);
    assign layer0_outputs[3379] = ~(inputs[110]);
    assign layer0_outputs[3380] = ~(inputs[187]) | (inputs[215]);
    assign layer0_outputs[3381] = ~((inputs[93]) | (inputs[248]));
    assign layer0_outputs[3382] = ~(inputs[194]);
    assign layer0_outputs[3383] = ~((inputs[162]) | (inputs[51]));
    assign layer0_outputs[3384] = inputs[148];
    assign layer0_outputs[3385] = inputs[16];
    assign layer0_outputs[3386] = (inputs[176]) & (inputs[52]);
    assign layer0_outputs[3387] = ~(inputs[248]);
    assign layer0_outputs[3388] = ~((inputs[215]) | (inputs[99]));
    assign layer0_outputs[3389] = ~((inputs[101]) | (inputs[60]));
    assign layer0_outputs[3390] = ~((inputs[169]) | (inputs[51]));
    assign layer0_outputs[3391] = ~(inputs[24]) | (inputs[189]);
    assign layer0_outputs[3392] = (inputs[107]) & ~(inputs[243]);
    assign layer0_outputs[3393] = inputs[3];
    assign layer0_outputs[3394] = (inputs[223]) ^ (inputs[102]);
    assign layer0_outputs[3395] = ~(inputs[58]) | (inputs[24]);
    assign layer0_outputs[3396] = (inputs[117]) | (inputs[224]);
    assign layer0_outputs[3397] = 1'b1;
    assign layer0_outputs[3398] = ~(inputs[89]);
    assign layer0_outputs[3399] = inputs[231];
    assign layer0_outputs[3400] = ~(inputs[182]) | (inputs[108]);
    assign layer0_outputs[3401] = 1'b1;
    assign layer0_outputs[3402] = ~((inputs[121]) ^ (inputs[225]));
    assign layer0_outputs[3403] = ~((inputs[45]) | (inputs[46]));
    assign layer0_outputs[3404] = ~((inputs[128]) | (inputs[173]));
    assign layer0_outputs[3405] = 1'b1;
    assign layer0_outputs[3406] = ~(inputs[99]) | (inputs[127]);
    assign layer0_outputs[3407] = (inputs[59]) | (inputs[88]);
    assign layer0_outputs[3408] = 1'b1;
    assign layer0_outputs[3409] = ~((inputs[12]) | (inputs[123]));
    assign layer0_outputs[3410] = ~((inputs[210]) ^ (inputs[75]));
    assign layer0_outputs[3411] = inputs[107];
    assign layer0_outputs[3412] = ~((inputs[186]) ^ (inputs[46]));
    assign layer0_outputs[3413] = (inputs[98]) | (inputs[184]);
    assign layer0_outputs[3414] = 1'b0;
    assign layer0_outputs[3415] = inputs[218];
    assign layer0_outputs[3416] = ~(inputs[172]) | (inputs[238]);
    assign layer0_outputs[3417] = 1'b1;
    assign layer0_outputs[3418] = 1'b0;
    assign layer0_outputs[3419] = (inputs[49]) | (inputs[192]);
    assign layer0_outputs[3420] = (inputs[68]) ^ (inputs[123]);
    assign layer0_outputs[3421] = (inputs[97]) | (inputs[75]);
    assign layer0_outputs[3422] = (inputs[89]) & (inputs[139]);
    assign layer0_outputs[3423] = ~((inputs[115]) | (inputs[83]));
    assign layer0_outputs[3424] = inputs[38];
    assign layer0_outputs[3425] = (inputs[185]) | (inputs[12]);
    assign layer0_outputs[3426] = inputs[95];
    assign layer0_outputs[3427] = ~((inputs[99]) ^ (inputs[16]));
    assign layer0_outputs[3428] = (inputs[177]) & (inputs[138]);
    assign layer0_outputs[3429] = ~(inputs[185]);
    assign layer0_outputs[3430] = (inputs[50]) ^ (inputs[230]);
    assign layer0_outputs[3431] = inputs[137];
    assign layer0_outputs[3432] = (inputs[138]) ^ (inputs[32]);
    assign layer0_outputs[3433] = inputs[85];
    assign layer0_outputs[3434] = (inputs[165]) ^ (inputs[85]);
    assign layer0_outputs[3435] = ~(inputs[201]);
    assign layer0_outputs[3436] = (inputs[7]) & ~(inputs[209]);
    assign layer0_outputs[3437] = ~(inputs[213]);
    assign layer0_outputs[3438] = ~(inputs[61]) | (inputs[82]);
    assign layer0_outputs[3439] = 1'b0;
    assign layer0_outputs[3440] = inputs[54];
    assign layer0_outputs[3441] = ~((inputs[168]) ^ (inputs[206]));
    assign layer0_outputs[3442] = ~(inputs[105]);
    assign layer0_outputs[3443] = 1'b1;
    assign layer0_outputs[3444] = ~(inputs[158]);
    assign layer0_outputs[3445] = 1'b0;
    assign layer0_outputs[3446] = ~(inputs[81]);
    assign layer0_outputs[3447] = (inputs[97]) & ~(inputs[7]);
    assign layer0_outputs[3448] = ~((inputs[170]) ^ (inputs[91]));
    assign layer0_outputs[3449] = inputs[86];
    assign layer0_outputs[3450] = (inputs[29]) & ~(inputs[218]);
    assign layer0_outputs[3451] = (inputs[37]) | (inputs[23]);
    assign layer0_outputs[3452] = (inputs[84]) & ~(inputs[174]);
    assign layer0_outputs[3453] = ~(inputs[226]);
    assign layer0_outputs[3454] = ~(inputs[94]) | (inputs[173]);
    assign layer0_outputs[3455] = ~(inputs[132]);
    assign layer0_outputs[3456] = ~(inputs[123]);
    assign layer0_outputs[3457] = inputs[106];
    assign layer0_outputs[3458] = ~((inputs[97]) & (inputs[11]));
    assign layer0_outputs[3459] = (inputs[183]) & ~(inputs[213]);
    assign layer0_outputs[3460] = (inputs[180]) & ~(inputs[222]);
    assign layer0_outputs[3461] = ~(inputs[162]);
    assign layer0_outputs[3462] = (inputs[140]) | (inputs[222]);
    assign layer0_outputs[3463] = ~(inputs[106]) | (inputs[141]);
    assign layer0_outputs[3464] = (inputs[198]) | (inputs[172]);
    assign layer0_outputs[3465] = (inputs[27]) & ~(inputs[240]);
    assign layer0_outputs[3466] = ~(inputs[121]);
    assign layer0_outputs[3467] = ~((inputs[2]) & (inputs[14]));
    assign layer0_outputs[3468] = (inputs[29]) & ~(inputs[111]);
    assign layer0_outputs[3469] = inputs[120];
    assign layer0_outputs[3470] = ~((inputs[82]) | (inputs[167]));
    assign layer0_outputs[3471] = inputs[60];
    assign layer0_outputs[3472] = ~(inputs[213]) | (inputs[37]);
    assign layer0_outputs[3473] = ~(inputs[172]);
    assign layer0_outputs[3474] = inputs[163];
    assign layer0_outputs[3475] = (inputs[204]) ^ (inputs[192]);
    assign layer0_outputs[3476] = ~(inputs[27]);
    assign layer0_outputs[3477] = inputs[124];
    assign layer0_outputs[3478] = ~((inputs[98]) ^ (inputs[26]));
    assign layer0_outputs[3479] = ~((inputs[227]) | (inputs[72]));
    assign layer0_outputs[3480] = 1'b0;
    assign layer0_outputs[3481] = inputs[131];
    assign layer0_outputs[3482] = (inputs[152]) | (inputs[135]);
    assign layer0_outputs[3483] = inputs[137];
    assign layer0_outputs[3484] = 1'b1;
    assign layer0_outputs[3485] = (inputs[197]) & ~(inputs[113]);
    assign layer0_outputs[3486] = inputs[110];
    assign layer0_outputs[3487] = ~(inputs[191]);
    assign layer0_outputs[3488] = (inputs[172]) | (inputs[109]);
    assign layer0_outputs[3489] = inputs[3];
    assign layer0_outputs[3490] = ~(inputs[63]) | (inputs[191]);
    assign layer0_outputs[3491] = 1'b1;
    assign layer0_outputs[3492] = ~(inputs[218]) | (inputs[95]);
    assign layer0_outputs[3493] = (inputs[32]) & ~(inputs[206]);
    assign layer0_outputs[3494] = (inputs[103]) & ~(inputs[193]);
    assign layer0_outputs[3495] = (inputs[95]) & ~(inputs[64]);
    assign layer0_outputs[3496] = 1'b0;
    assign layer0_outputs[3497] = ~((inputs[233]) ^ (inputs[177]));
    assign layer0_outputs[3498] = ~((inputs[203]) | (inputs[174]));
    assign layer0_outputs[3499] = (inputs[22]) & ~(inputs[2]);
    assign layer0_outputs[3500] = ~(inputs[141]) | (inputs[94]);
    assign layer0_outputs[3501] = ~(inputs[136]);
    assign layer0_outputs[3502] = ~((inputs[114]) & (inputs[127]));
    assign layer0_outputs[3503] = ~((inputs[148]) | (inputs[51]));
    assign layer0_outputs[3504] = ~(inputs[38]) | (inputs[29]);
    assign layer0_outputs[3505] = (inputs[208]) & ~(inputs[244]);
    assign layer0_outputs[3506] = ~((inputs[212]) | (inputs[231]));
    assign layer0_outputs[3507] = (inputs[74]) & ~(inputs[96]);
    assign layer0_outputs[3508] = ~(inputs[186]);
    assign layer0_outputs[3509] = (inputs[67]) & ~(inputs[246]);
    assign layer0_outputs[3510] = ~(inputs[152]) | (inputs[212]);
    assign layer0_outputs[3511] = ~((inputs[27]) ^ (inputs[178]));
    assign layer0_outputs[3512] = (inputs[69]) & ~(inputs[7]);
    assign layer0_outputs[3513] = (inputs[154]) ^ (inputs[245]);
    assign layer0_outputs[3514] = ~(inputs[225]);
    assign layer0_outputs[3515] = (inputs[152]) & ~(inputs[162]);
    assign layer0_outputs[3516] = (inputs[180]) & ~(inputs[98]);
    assign layer0_outputs[3517] = inputs[117];
    assign layer0_outputs[3518] = inputs[253];
    assign layer0_outputs[3519] = (inputs[6]) ^ (inputs[201]);
    assign layer0_outputs[3520] = ~((inputs[221]) ^ (inputs[224]));
    assign layer0_outputs[3521] = ~((inputs[139]) | (inputs[124]));
    assign layer0_outputs[3522] = (inputs[72]) | (inputs[48]);
    assign layer0_outputs[3523] = ~(inputs[12]) | (inputs[168]);
    assign layer0_outputs[3524] = ~(inputs[143]) | (inputs[2]);
    assign layer0_outputs[3525] = ~(inputs[101]);
    assign layer0_outputs[3526] = ~(inputs[200]);
    assign layer0_outputs[3527] = inputs[61];
    assign layer0_outputs[3528] = (inputs[20]) & ~(inputs[2]);
    assign layer0_outputs[3529] = inputs[200];
    assign layer0_outputs[3530] = (inputs[30]) ^ (inputs[23]);
    assign layer0_outputs[3531] = inputs[42];
    assign layer0_outputs[3532] = (inputs[159]) & (inputs[255]);
    assign layer0_outputs[3533] = (inputs[62]) & ~(inputs[6]);
    assign layer0_outputs[3534] = ~(inputs[91]);
    assign layer0_outputs[3535] = (inputs[92]) | (inputs[74]);
    assign layer0_outputs[3536] = ~((inputs[166]) ^ (inputs[243]));
    assign layer0_outputs[3537] = (inputs[26]) & ~(inputs[159]);
    assign layer0_outputs[3538] = (inputs[193]) | (inputs[232]);
    assign layer0_outputs[3539] = (inputs[92]) & ~(inputs[47]);
    assign layer0_outputs[3540] = (inputs[154]) | (inputs[202]);
    assign layer0_outputs[3541] = ~((inputs[141]) ^ (inputs[112]));
    assign layer0_outputs[3542] = (inputs[97]) ^ (inputs[147]);
    assign layer0_outputs[3543] = (inputs[125]) | (inputs[227]);
    assign layer0_outputs[3544] = (inputs[237]) ^ (inputs[56]);
    assign layer0_outputs[3545] = ~((inputs[227]) | (inputs[85]));
    assign layer0_outputs[3546] = ~((inputs[180]) & (inputs[42]));
    assign layer0_outputs[3547] = (inputs[118]) | (inputs[157]);
    assign layer0_outputs[3548] = (inputs[182]) & ~(inputs[30]);
    assign layer0_outputs[3549] = (inputs[228]) | (inputs[20]);
    assign layer0_outputs[3550] = (inputs[74]) | (inputs[219]);
    assign layer0_outputs[3551] = ~(inputs[233]) | (inputs[1]);
    assign layer0_outputs[3552] = ~((inputs[225]) ^ (inputs[71]));
    assign layer0_outputs[3553] = (inputs[152]) | (inputs[28]);
    assign layer0_outputs[3554] = ~((inputs[130]) ^ (inputs[249]));
    assign layer0_outputs[3555] = ~((inputs[117]) ^ (inputs[130]));
    assign layer0_outputs[3556] = (inputs[145]) | (inputs[38]);
    assign layer0_outputs[3557] = ~(inputs[90]) | (inputs[195]);
    assign layer0_outputs[3558] = ~(inputs[202]) | (inputs[115]);
    assign layer0_outputs[3559] = (inputs[188]) ^ (inputs[238]);
    assign layer0_outputs[3560] = ~(inputs[108]);
    assign layer0_outputs[3561] = ~((inputs[50]) ^ (inputs[48]));
    assign layer0_outputs[3562] = ~((inputs[95]) | (inputs[75]));
    assign layer0_outputs[3563] = 1'b1;
    assign layer0_outputs[3564] = (inputs[114]) & (inputs[190]);
    assign layer0_outputs[3565] = inputs[66];
    assign layer0_outputs[3566] = ~(inputs[132]) | (inputs[24]);
    assign layer0_outputs[3567] = inputs[215];
    assign layer0_outputs[3568] = (inputs[223]) & (inputs[43]);
    assign layer0_outputs[3569] = ~((inputs[148]) | (inputs[83]));
    assign layer0_outputs[3570] = ~(inputs[53]) | (inputs[115]);
    assign layer0_outputs[3571] = 1'b1;
    assign layer0_outputs[3572] = (inputs[217]) ^ (inputs[28]);
    assign layer0_outputs[3573] = (inputs[156]) | (inputs[102]);
    assign layer0_outputs[3574] = ~(inputs[223]);
    assign layer0_outputs[3575] = ~((inputs[82]) | (inputs[80]));
    assign layer0_outputs[3576] = inputs[75];
    assign layer0_outputs[3577] = ~(inputs[239]);
    assign layer0_outputs[3578] = ~((inputs[85]) | (inputs[212]));
    assign layer0_outputs[3579] = ~(inputs[138]) | (inputs[220]);
    assign layer0_outputs[3580] = ~(inputs[119]);
    assign layer0_outputs[3581] = ~(inputs[102]) | (inputs[248]);
    assign layer0_outputs[3582] = ~((inputs[199]) & (inputs[185]));
    assign layer0_outputs[3583] = inputs[82];
    assign layer0_outputs[3584] = (inputs[138]) & ~(inputs[175]);
    assign layer0_outputs[3585] = ~(inputs[50]) | (inputs[19]);
    assign layer0_outputs[3586] = (inputs[27]) ^ (inputs[175]);
    assign layer0_outputs[3587] = ~((inputs[103]) | (inputs[222]));
    assign layer0_outputs[3588] = inputs[111];
    assign layer0_outputs[3589] = (inputs[52]) ^ (inputs[140]);
    assign layer0_outputs[3590] = ~(inputs[162]) | (inputs[64]);
    assign layer0_outputs[3591] = (inputs[20]) & ~(inputs[128]);
    assign layer0_outputs[3592] = ~(inputs[55]) | (inputs[132]);
    assign layer0_outputs[3593] = (inputs[153]) & ~(inputs[6]);
    assign layer0_outputs[3594] = ~((inputs[104]) | (inputs[130]));
    assign layer0_outputs[3595] = (inputs[221]) | (inputs[249]);
    assign layer0_outputs[3596] = 1'b0;
    assign layer0_outputs[3597] = (inputs[58]) ^ (inputs[238]);
    assign layer0_outputs[3598] = ~(inputs[72]) | (inputs[183]);
    assign layer0_outputs[3599] = inputs[54];
    assign layer0_outputs[3600] = ~((inputs[98]) ^ (inputs[35]));
    assign layer0_outputs[3601] = (inputs[197]) & ~(inputs[160]);
    assign layer0_outputs[3602] = ~(inputs[170]) | (inputs[211]);
    assign layer0_outputs[3603] = (inputs[87]) | (inputs[7]);
    assign layer0_outputs[3604] = inputs[142];
    assign layer0_outputs[3605] = (inputs[181]) | (inputs[83]);
    assign layer0_outputs[3606] = (inputs[65]) & (inputs[3]);
    assign layer0_outputs[3607] = (inputs[176]) & (inputs[21]);
    assign layer0_outputs[3608] = inputs[74];
    assign layer0_outputs[3609] = ~((inputs[14]) | (inputs[37]));
    assign layer0_outputs[3610] = ~(inputs[166]);
    assign layer0_outputs[3611] = inputs[88];
    assign layer0_outputs[3612] = ~((inputs[141]) | (inputs[77]));
    assign layer0_outputs[3613] = inputs[120];
    assign layer0_outputs[3614] = (inputs[177]) ^ (inputs[171]);
    assign layer0_outputs[3615] = (inputs[43]) | (inputs[4]);
    assign layer0_outputs[3616] = (inputs[152]) | (inputs[23]);
    assign layer0_outputs[3617] = (inputs[206]) ^ (inputs[176]);
    assign layer0_outputs[3618] = ~((inputs[60]) | (inputs[188]));
    assign layer0_outputs[3619] = (inputs[12]) ^ (inputs[36]);
    assign layer0_outputs[3620] = ~(inputs[203]);
    assign layer0_outputs[3621] = (inputs[107]) ^ (inputs[49]);
    assign layer0_outputs[3622] = ~(inputs[203]) | (inputs[161]);
    assign layer0_outputs[3623] = 1'b0;
    assign layer0_outputs[3624] = ~(inputs[249]) | (inputs[20]);
    assign layer0_outputs[3625] = ~((inputs[208]) ^ (inputs[86]));
    assign layer0_outputs[3626] = (inputs[62]) & ~(inputs[33]);
    assign layer0_outputs[3627] = (inputs[175]) & ~(inputs[12]);
    assign layer0_outputs[3628] = (inputs[241]) ^ (inputs[60]);
    assign layer0_outputs[3629] = (inputs[160]) & ~(inputs[22]);
    assign layer0_outputs[3630] = ~(inputs[52]);
    assign layer0_outputs[3631] = ~((inputs[169]) & (inputs[232]));
    assign layer0_outputs[3632] = (inputs[122]) & ~(inputs[49]);
    assign layer0_outputs[3633] = inputs[120];
    assign layer0_outputs[3634] = ~(inputs[205]);
    assign layer0_outputs[3635] = inputs[126];
    assign layer0_outputs[3636] = inputs[241];
    assign layer0_outputs[3637] = (inputs[50]) & ~(inputs[219]);
    assign layer0_outputs[3638] = (inputs[228]) | (inputs[251]);
    assign layer0_outputs[3639] = ~(inputs[136]);
    assign layer0_outputs[3640] = (inputs[20]) & (inputs[173]);
    assign layer0_outputs[3641] = ~((inputs[74]) ^ (inputs[114]));
    assign layer0_outputs[3642] = ~(inputs[233]);
    assign layer0_outputs[3643] = ~((inputs[222]) ^ (inputs[236]));
    assign layer0_outputs[3644] = ~(inputs[229]);
    assign layer0_outputs[3645] = inputs[214];
    assign layer0_outputs[3646] = ~((inputs[26]) | (inputs[185]));
    assign layer0_outputs[3647] = (inputs[58]) | (inputs[33]);
    assign layer0_outputs[3648] = (inputs[58]) & ~(inputs[154]);
    assign layer0_outputs[3649] = ~((inputs[125]) ^ (inputs[97]));
    assign layer0_outputs[3650] = (inputs[175]) ^ (inputs[175]);
    assign layer0_outputs[3651] = (inputs[226]) ^ (inputs[31]);
    assign layer0_outputs[3652] = (inputs[209]) ^ (inputs[107]);
    assign layer0_outputs[3653] = ~((inputs[201]) | (inputs[253]));
    assign layer0_outputs[3654] = (inputs[186]) | (inputs[91]);
    assign layer0_outputs[3655] = inputs[120];
    assign layer0_outputs[3656] = (inputs[10]) | (inputs[84]);
    assign layer0_outputs[3657] = inputs[9];
    assign layer0_outputs[3658] = inputs[139];
    assign layer0_outputs[3659] = inputs[137];
    assign layer0_outputs[3660] = (inputs[120]) & (inputs[105]);
    assign layer0_outputs[3661] = 1'b1;
    assign layer0_outputs[3662] = (inputs[106]) & ~(inputs[73]);
    assign layer0_outputs[3663] = inputs[84];
    assign layer0_outputs[3664] = (inputs[219]) & ~(inputs[51]);
    assign layer0_outputs[3665] = ~((inputs[149]) | (inputs[205]));
    assign layer0_outputs[3666] = (inputs[255]) | (inputs[205]);
    assign layer0_outputs[3667] = (inputs[207]) | (inputs[198]);
    assign layer0_outputs[3668] = ~((inputs[208]) | (inputs[73]));
    assign layer0_outputs[3669] = (inputs[133]) & ~(inputs[191]);
    assign layer0_outputs[3670] = (inputs[198]) & ~(inputs[15]);
    assign layer0_outputs[3671] = inputs[237];
    assign layer0_outputs[3672] = ~((inputs[19]) ^ (inputs[205]));
    assign layer0_outputs[3673] = ~((inputs[16]) | (inputs[235]));
    assign layer0_outputs[3674] = (inputs[246]) | (inputs[233]);
    assign layer0_outputs[3675] = ~((inputs[204]) | (inputs[181]));
    assign layer0_outputs[3676] = ~((inputs[223]) & (inputs[65]));
    assign layer0_outputs[3677] = ~(inputs[71]) | (inputs[68]);
    assign layer0_outputs[3678] = ~((inputs[2]) | (inputs[83]));
    assign layer0_outputs[3679] = (inputs[131]) & ~(inputs[6]);
    assign layer0_outputs[3680] = ~(inputs[102]);
    assign layer0_outputs[3681] = inputs[161];
    assign layer0_outputs[3682] = (inputs[187]) & ~(inputs[157]);
    assign layer0_outputs[3683] = (inputs[133]) & ~(inputs[240]);
    assign layer0_outputs[3684] = (inputs[121]) & ~(inputs[119]);
    assign layer0_outputs[3685] = (inputs[172]) | (inputs[22]);
    assign layer0_outputs[3686] = ~(inputs[203]);
    assign layer0_outputs[3687] = 1'b1;
    assign layer0_outputs[3688] = ~(inputs[100]) | (inputs[156]);
    assign layer0_outputs[3689] = ~((inputs[211]) | (inputs[26]));
    assign layer0_outputs[3690] = (inputs[51]) | (inputs[168]);
    assign layer0_outputs[3691] = (inputs[37]) | (inputs[70]);
    assign layer0_outputs[3692] = (inputs[11]) & (inputs[144]);
    assign layer0_outputs[3693] = ~(inputs[116]) | (inputs[246]);
    assign layer0_outputs[3694] = ~((inputs[161]) | (inputs[195]));
    assign layer0_outputs[3695] = (inputs[45]) | (inputs[133]);
    assign layer0_outputs[3696] = ~(inputs[204]) | (inputs[66]);
    assign layer0_outputs[3697] = ~(inputs[254]);
    assign layer0_outputs[3698] = inputs[56];
    assign layer0_outputs[3699] = (inputs[169]) | (inputs[205]);
    assign layer0_outputs[3700] = ~(inputs[167]) | (inputs[81]);
    assign layer0_outputs[3701] = (inputs[151]) & ~(inputs[173]);
    assign layer0_outputs[3702] = (inputs[82]) | (inputs[114]);
    assign layer0_outputs[3703] = inputs[183];
    assign layer0_outputs[3704] = (inputs[242]) | (inputs[56]);
    assign layer0_outputs[3705] = inputs[187];
    assign layer0_outputs[3706] = (inputs[137]) ^ (inputs[33]);
    assign layer0_outputs[3707] = (inputs[59]) & ~(inputs[2]);
    assign layer0_outputs[3708] = 1'b1;
    assign layer0_outputs[3709] = ~((inputs[221]) | (inputs[133]));
    assign layer0_outputs[3710] = ~(inputs[134]);
    assign layer0_outputs[3711] = inputs[21];
    assign layer0_outputs[3712] = (inputs[209]) ^ (inputs[201]);
    assign layer0_outputs[3713] = ~((inputs[15]) & (inputs[242]));
    assign layer0_outputs[3714] = ~(inputs[156]) | (inputs[13]);
    assign layer0_outputs[3715] = inputs[72];
    assign layer0_outputs[3716] = ~((inputs[4]) & (inputs[95]));
    assign layer0_outputs[3717] = (inputs[55]) & (inputs[119]);
    assign layer0_outputs[3718] = 1'b1;
    assign layer0_outputs[3719] = ~(inputs[68]) | (inputs[149]);
    assign layer0_outputs[3720] = (inputs[200]) & (inputs[76]);
    assign layer0_outputs[3721] = (inputs[79]) | (inputs[252]);
    assign layer0_outputs[3722] = ~(inputs[32]);
    assign layer0_outputs[3723] = ~((inputs[203]) | (inputs[36]));
    assign layer0_outputs[3724] = ~((inputs[80]) | (inputs[26]));
    assign layer0_outputs[3725] = ~((inputs[204]) & (inputs[11]));
    assign layer0_outputs[3726] = ~((inputs[28]) ^ (inputs[82]));
    assign layer0_outputs[3727] = (inputs[236]) ^ (inputs[232]);
    assign layer0_outputs[3728] = (inputs[220]) | (inputs[175]);
    assign layer0_outputs[3729] = ~((inputs[212]) | (inputs[196]));
    assign layer0_outputs[3730] = inputs[150];
    assign layer0_outputs[3731] = 1'b0;
    assign layer0_outputs[3732] = (inputs[77]) | (inputs[197]);
    assign layer0_outputs[3733] = (inputs[214]) ^ (inputs[77]);
    assign layer0_outputs[3734] = (inputs[0]) & ~(inputs[107]);
    assign layer0_outputs[3735] = (inputs[249]) & ~(inputs[207]);
    assign layer0_outputs[3736] = inputs[104];
    assign layer0_outputs[3737] = (inputs[219]) | (inputs[75]);
    assign layer0_outputs[3738] = (inputs[167]) & ~(inputs[163]);
    assign layer0_outputs[3739] = (inputs[16]) ^ (inputs[230]);
    assign layer0_outputs[3740] = ~(inputs[164]) | (inputs[211]);
    assign layer0_outputs[3741] = ~(inputs[125]);
    assign layer0_outputs[3742] = (inputs[217]) & ~(inputs[113]);
    assign layer0_outputs[3743] = ~(inputs[231]);
    assign layer0_outputs[3744] = (inputs[205]) & ~(inputs[1]);
    assign layer0_outputs[3745] = (inputs[233]) ^ (inputs[111]);
    assign layer0_outputs[3746] = (inputs[27]) ^ (inputs[1]);
    assign layer0_outputs[3747] = (inputs[165]) ^ (inputs[15]);
    assign layer0_outputs[3748] = (inputs[84]) ^ (inputs[214]);
    assign layer0_outputs[3749] = inputs[28];
    assign layer0_outputs[3750] = (inputs[62]) & ~(inputs[64]);
    assign layer0_outputs[3751] = ~(inputs[180]);
    assign layer0_outputs[3752] = ~(inputs[99]);
    assign layer0_outputs[3753] = inputs[233];
    assign layer0_outputs[3754] = (inputs[199]) & (inputs[196]);
    assign layer0_outputs[3755] = (inputs[159]) | (inputs[127]);
    assign layer0_outputs[3756] = (inputs[61]) & ~(inputs[24]);
    assign layer0_outputs[3757] = (inputs[126]) & ~(inputs[137]);
    assign layer0_outputs[3758] = ~(inputs[57]) | (inputs[18]);
    assign layer0_outputs[3759] = ~((inputs[92]) ^ (inputs[14]));
    assign layer0_outputs[3760] = ~((inputs[0]) | (inputs[7]));
    assign layer0_outputs[3761] = inputs[109];
    assign layer0_outputs[3762] = (inputs[212]) | (inputs[79]);
    assign layer0_outputs[3763] = ~((inputs[4]) ^ (inputs[77]));
    assign layer0_outputs[3764] = ~((inputs[142]) ^ (inputs[188]));
    assign layer0_outputs[3765] = ~((inputs[130]) & (inputs[49]));
    assign layer0_outputs[3766] = ~(inputs[172]);
    assign layer0_outputs[3767] = ~((inputs[99]) & (inputs[95]));
    assign layer0_outputs[3768] = inputs[248];
    assign layer0_outputs[3769] = ~((inputs[153]) | (inputs[154]));
    assign layer0_outputs[3770] = ~(inputs[116]) | (inputs[21]);
    assign layer0_outputs[3771] = ~((inputs[25]) | (inputs[52]));
    assign layer0_outputs[3772] = ~((inputs[17]) | (inputs[238]));
    assign layer0_outputs[3773] = (inputs[27]) | (inputs[87]);
    assign layer0_outputs[3774] = ~(inputs[71]) | (inputs[223]);
    assign layer0_outputs[3775] = inputs[120];
    assign layer0_outputs[3776] = (inputs[246]) & ~(inputs[12]);
    assign layer0_outputs[3777] = (inputs[149]) | (inputs[123]);
    assign layer0_outputs[3778] = (inputs[97]) | (inputs[73]);
    assign layer0_outputs[3779] = (inputs[184]) & (inputs[154]);
    assign layer0_outputs[3780] = ~(inputs[156]);
    assign layer0_outputs[3781] = (inputs[248]) ^ (inputs[27]);
    assign layer0_outputs[3782] = inputs[81];
    assign layer0_outputs[3783] = ~((inputs[138]) | (inputs[66]));
    assign layer0_outputs[3784] = inputs[168];
    assign layer0_outputs[3785] = inputs[130];
    assign layer0_outputs[3786] = ~((inputs[189]) ^ (inputs[149]));
    assign layer0_outputs[3787] = ~(inputs[79]);
    assign layer0_outputs[3788] = 1'b1;
    assign layer0_outputs[3789] = inputs[2];
    assign layer0_outputs[3790] = ~((inputs[84]) ^ (inputs[43]));
    assign layer0_outputs[3791] = (inputs[25]) | (inputs[114]);
    assign layer0_outputs[3792] = ~((inputs[157]) | (inputs[166]));
    assign layer0_outputs[3793] = ~(inputs[60]);
    assign layer0_outputs[3794] = 1'b0;
    assign layer0_outputs[3795] = (inputs[166]) | (inputs[129]);
    assign layer0_outputs[3796] = (inputs[138]) & ~(inputs[132]);
    assign layer0_outputs[3797] = ~(inputs[124]);
    assign layer0_outputs[3798] = (inputs[73]) | (inputs[48]);
    assign layer0_outputs[3799] = (inputs[47]) ^ (inputs[227]);
    assign layer0_outputs[3800] = (inputs[126]) | (inputs[156]);
    assign layer0_outputs[3801] = (inputs[26]) & ~(inputs[145]);
    assign layer0_outputs[3802] = (inputs[202]) & ~(inputs[46]);
    assign layer0_outputs[3803] = (inputs[91]) & ~(inputs[156]);
    assign layer0_outputs[3804] = ~(inputs[162]) | (inputs[184]);
    assign layer0_outputs[3805] = ~((inputs[196]) ^ (inputs[92]));
    assign layer0_outputs[3806] = ~(inputs[201]) | (inputs[68]);
    assign layer0_outputs[3807] = ~(inputs[173]) | (inputs[250]);
    assign layer0_outputs[3808] = ~((inputs[192]) ^ (inputs[105]));
    assign layer0_outputs[3809] = (inputs[12]) & ~(inputs[79]);
    assign layer0_outputs[3810] = ~((inputs[37]) ^ (inputs[20]));
    assign layer0_outputs[3811] = ~((inputs[132]) | (inputs[205]));
    assign layer0_outputs[3812] = ~(inputs[88]);
    assign layer0_outputs[3813] = ~(inputs[202]) | (inputs[24]);
    assign layer0_outputs[3814] = (inputs[240]) & (inputs[252]);
    assign layer0_outputs[3815] = ~(inputs[202]) | (inputs[88]);
    assign layer0_outputs[3816] = (inputs[97]) ^ (inputs[29]);
    assign layer0_outputs[3817] = inputs[186];
    assign layer0_outputs[3818] = (inputs[157]) | (inputs[153]);
    assign layer0_outputs[3819] = 1'b0;
    assign layer0_outputs[3820] = ~(inputs[39]) | (inputs[63]);
    assign layer0_outputs[3821] = inputs[45];
    assign layer0_outputs[3822] = (inputs[218]) & (inputs[135]);
    assign layer0_outputs[3823] = ~((inputs[95]) ^ (inputs[166]));
    assign layer0_outputs[3824] = (inputs[116]) & ~(inputs[230]);
    assign layer0_outputs[3825] = inputs[195];
    assign layer0_outputs[3826] = inputs[185];
    assign layer0_outputs[3827] = ~((inputs[241]) & (inputs[146]));
    assign layer0_outputs[3828] = ~(inputs[204]);
    assign layer0_outputs[3829] = 1'b0;
    assign layer0_outputs[3830] = inputs[56];
    assign layer0_outputs[3831] = ~((inputs[192]) | (inputs[147]));
    assign layer0_outputs[3832] = inputs[119];
    assign layer0_outputs[3833] = ~((inputs[186]) | (inputs[35]));
    assign layer0_outputs[3834] = ~(inputs[213]) | (inputs[81]);
    assign layer0_outputs[3835] = (inputs[122]) & ~(inputs[151]);
    assign layer0_outputs[3836] = ~((inputs[92]) | (inputs[77]));
    assign layer0_outputs[3837] = ~(inputs[210]) | (inputs[208]);
    assign layer0_outputs[3838] = (inputs[66]) | (inputs[90]);
    assign layer0_outputs[3839] = inputs[133];
    assign layer0_outputs[3840] = ~((inputs[134]) | (inputs[202]));
    assign layer0_outputs[3841] = (inputs[55]) ^ (inputs[63]);
    assign layer0_outputs[3842] = ~((inputs[176]) ^ (inputs[167]));
    assign layer0_outputs[3843] = (inputs[216]) | (inputs[28]);
    assign layer0_outputs[3844] = inputs[66];
    assign layer0_outputs[3845] = ~(inputs[100]) | (inputs[240]);
    assign layer0_outputs[3846] = ~(inputs[109]) | (inputs[205]);
    assign layer0_outputs[3847] = inputs[94];
    assign layer0_outputs[3848] = ~(inputs[61]) | (inputs[113]);
    assign layer0_outputs[3849] = (inputs[157]) & ~(inputs[46]);
    assign layer0_outputs[3850] = ~((inputs[246]) ^ (inputs[88]));
    assign layer0_outputs[3851] = 1'b1;
    assign layer0_outputs[3852] = (inputs[186]) & ~(inputs[99]);
    assign layer0_outputs[3853] = inputs[58];
    assign layer0_outputs[3854] = (inputs[218]) & (inputs[206]);
    assign layer0_outputs[3855] = (inputs[93]) ^ (inputs[192]);
    assign layer0_outputs[3856] = 1'b1;
    assign layer0_outputs[3857] = ~((inputs[174]) | (inputs[152]));
    assign layer0_outputs[3858] = ~(inputs[55]);
    assign layer0_outputs[3859] = ~((inputs[233]) | (inputs[178]));
    assign layer0_outputs[3860] = ~(inputs[83]) | (inputs[245]);
    assign layer0_outputs[3861] = ~(inputs[155]) | (inputs[251]);
    assign layer0_outputs[3862] = (inputs[179]) | (inputs[254]);
    assign layer0_outputs[3863] = ~(inputs[225]);
    assign layer0_outputs[3864] = (inputs[28]) ^ (inputs[81]);
    assign layer0_outputs[3865] = ~((inputs[6]) | (inputs[251]));
    assign layer0_outputs[3866] = ~((inputs[104]) | (inputs[235]));
    assign layer0_outputs[3867] = (inputs[78]) | (inputs[77]);
    assign layer0_outputs[3868] = ~(inputs[135]);
    assign layer0_outputs[3869] = ~(inputs[133]);
    assign layer0_outputs[3870] = (inputs[49]) ^ (inputs[105]);
    assign layer0_outputs[3871] = inputs[166];
    assign layer0_outputs[3872] = (inputs[243]) & ~(inputs[250]);
    assign layer0_outputs[3873] = ~((inputs[147]) | (inputs[37]));
    assign layer0_outputs[3874] = ~((inputs[147]) ^ (inputs[36]));
    assign layer0_outputs[3875] = inputs[198];
    assign layer0_outputs[3876] = (inputs[95]) & (inputs[210]);
    assign layer0_outputs[3877] = (inputs[130]) | (inputs[138]);
    assign layer0_outputs[3878] = ~((inputs[81]) | (inputs[124]));
    assign layer0_outputs[3879] = 1'b1;
    assign layer0_outputs[3880] = ~((inputs[112]) | (inputs[184]));
    assign layer0_outputs[3881] = (inputs[70]) & ~(inputs[235]);
    assign layer0_outputs[3882] = ~(inputs[197]) | (inputs[158]);
    assign layer0_outputs[3883] = ~((inputs[197]) ^ (inputs[228]));
    assign layer0_outputs[3884] = ~((inputs[22]) ^ (inputs[108]));
    assign layer0_outputs[3885] = inputs[78];
    assign layer0_outputs[3886] = ~((inputs[246]) & (inputs[20]));
    assign layer0_outputs[3887] = ~(inputs[47]);
    assign layer0_outputs[3888] = (inputs[126]) | (inputs[55]);
    assign layer0_outputs[3889] = ~(inputs[104]);
    assign layer0_outputs[3890] = 1'b0;
    assign layer0_outputs[3891] = inputs[120];
    assign layer0_outputs[3892] = ~(inputs[125]);
    assign layer0_outputs[3893] = ~(inputs[116]);
    assign layer0_outputs[3894] = ~((inputs[21]) ^ (inputs[64]));
    assign layer0_outputs[3895] = inputs[85];
    assign layer0_outputs[3896] = ~(inputs[12]) | (inputs[176]);
    assign layer0_outputs[3897] = (inputs[87]) & ~(inputs[82]);
    assign layer0_outputs[3898] = (inputs[109]) ^ (inputs[215]);
    assign layer0_outputs[3899] = ~((inputs[203]) ^ (inputs[222]));
    assign layer0_outputs[3900] = ~((inputs[116]) | (inputs[236]));
    assign layer0_outputs[3901] = (inputs[240]) | (inputs[184]);
    assign layer0_outputs[3902] = (inputs[80]) ^ (inputs[172]);
    assign layer0_outputs[3903] = inputs[253];
    assign layer0_outputs[3904] = (inputs[206]) | (inputs[194]);
    assign layer0_outputs[3905] = (inputs[250]) & ~(inputs[243]);
    assign layer0_outputs[3906] = (inputs[83]) | (inputs[114]);
    assign layer0_outputs[3907] = (inputs[76]) | (inputs[180]);
    assign layer0_outputs[3908] = ~(inputs[140]);
    assign layer0_outputs[3909] = ~((inputs[233]) ^ (inputs[232]));
    assign layer0_outputs[3910] = inputs[5];
    assign layer0_outputs[3911] = (inputs[67]) | (inputs[182]);
    assign layer0_outputs[3912] = ~((inputs[129]) ^ (inputs[145]));
    assign layer0_outputs[3913] = (inputs[17]) ^ (inputs[201]);
    assign layer0_outputs[3914] = ~((inputs[37]) | (inputs[171]));
    assign layer0_outputs[3915] = inputs[122];
    assign layer0_outputs[3916] = (inputs[48]) | (inputs[188]);
    assign layer0_outputs[3917] = (inputs[183]) & ~(inputs[211]);
    assign layer0_outputs[3918] = ~((inputs[110]) | (inputs[255]));
    assign layer0_outputs[3919] = ~((inputs[15]) | (inputs[144]));
    assign layer0_outputs[3920] = ~((inputs[62]) ^ (inputs[47]));
    assign layer0_outputs[3921] = ~(inputs[24]) | (inputs[128]);
    assign layer0_outputs[3922] = inputs[219];
    assign layer0_outputs[3923] = ~(inputs[138]);
    assign layer0_outputs[3924] = inputs[234];
    assign layer0_outputs[3925] = ~((inputs[125]) ^ (inputs[235]));
    assign layer0_outputs[3926] = (inputs[125]) & ~(inputs[33]);
    assign layer0_outputs[3927] = (inputs[72]) | (inputs[38]);
    assign layer0_outputs[3928] = ~(inputs[144]) | (inputs[19]);
    assign layer0_outputs[3929] = (inputs[94]) ^ (inputs[59]);
    assign layer0_outputs[3930] = 1'b0;
    assign layer0_outputs[3931] = (inputs[190]) & ~(inputs[2]);
    assign layer0_outputs[3932] = ~(inputs[159]);
    assign layer0_outputs[3933] = ~((inputs[129]) ^ (inputs[2]));
    assign layer0_outputs[3934] = ~((inputs[143]) & (inputs[111]));
    assign layer0_outputs[3935] = ~(inputs[219]);
    assign layer0_outputs[3936] = (inputs[243]) & ~(inputs[224]);
    assign layer0_outputs[3937] = ~(inputs[17]);
    assign layer0_outputs[3938] = ~((inputs[213]) & (inputs[249]));
    assign layer0_outputs[3939] = (inputs[255]) ^ (inputs[160]);
    assign layer0_outputs[3940] = ~((inputs[41]) | (inputs[228]));
    assign layer0_outputs[3941] = inputs[211];
    assign layer0_outputs[3942] = (inputs[71]) ^ (inputs[64]);
    assign layer0_outputs[3943] = ~(inputs[93]);
    assign layer0_outputs[3944] = (inputs[179]) | (inputs[195]);
    assign layer0_outputs[3945] = inputs[133];
    assign layer0_outputs[3946] = ~(inputs[116]) | (inputs[33]);
    assign layer0_outputs[3947] = ~(inputs[203]);
    assign layer0_outputs[3948] = (inputs[121]) & ~(inputs[93]);
    assign layer0_outputs[3949] = (inputs[169]) & ~(inputs[247]);
    assign layer0_outputs[3950] = inputs[132];
    assign layer0_outputs[3951] = ~((inputs[43]) | (inputs[61]));
    assign layer0_outputs[3952] = ~((inputs[131]) ^ (inputs[8]));
    assign layer0_outputs[3953] = ~(inputs[165]);
    assign layer0_outputs[3954] = ~(inputs[71]) | (inputs[246]);
    assign layer0_outputs[3955] = ~((inputs[195]) & (inputs[114]));
    assign layer0_outputs[3956] = ~(inputs[116]) | (inputs[226]);
    assign layer0_outputs[3957] = ~(inputs[135]) | (inputs[24]);
    assign layer0_outputs[3958] = ~(inputs[149]) | (inputs[234]);
    assign layer0_outputs[3959] = (inputs[195]) | (inputs[44]);
    assign layer0_outputs[3960] = (inputs[6]) | (inputs[199]);
    assign layer0_outputs[3961] = ~(inputs[5]);
    assign layer0_outputs[3962] = 1'b0;
    assign layer0_outputs[3963] = ~(inputs[163]);
    assign layer0_outputs[3964] = ~(inputs[167]) | (inputs[5]);
    assign layer0_outputs[3965] = ~(inputs[71]) | (inputs[8]);
    assign layer0_outputs[3966] = inputs[165];
    assign layer0_outputs[3967] = ~(inputs[141]) | (inputs[14]);
    assign layer0_outputs[3968] = ~((inputs[9]) & (inputs[242]));
    assign layer0_outputs[3969] = ~(inputs[73]);
    assign layer0_outputs[3970] = inputs[30];
    assign layer0_outputs[3971] = (inputs[175]) ^ (inputs[25]);
    assign layer0_outputs[3972] = (inputs[69]) | (inputs[85]);
    assign layer0_outputs[3973] = ~(inputs[23]);
    assign layer0_outputs[3974] = ~(inputs[66]);
    assign layer0_outputs[3975] = inputs[101];
    assign layer0_outputs[3976] = ~(inputs[58]) | (inputs[175]);
    assign layer0_outputs[3977] = ~(inputs[90]);
    assign layer0_outputs[3978] = ~(inputs[74]);
    assign layer0_outputs[3979] = (inputs[84]) & ~(inputs[94]);
    assign layer0_outputs[3980] = (inputs[37]) | (inputs[51]);
    assign layer0_outputs[3981] = ~(inputs[138]);
    assign layer0_outputs[3982] = ~((inputs[111]) | (inputs[181]));
    assign layer0_outputs[3983] = ~(inputs[166]);
    assign layer0_outputs[3984] = ~(inputs[144]);
    assign layer0_outputs[3985] = ~(inputs[116]) | (inputs[96]);
    assign layer0_outputs[3986] = ~((inputs[36]) & (inputs[145]));
    assign layer0_outputs[3987] = (inputs[38]) | (inputs[19]);
    assign layer0_outputs[3988] = (inputs[179]) | (inputs[60]);
    assign layer0_outputs[3989] = ~((inputs[76]) | (inputs[155]));
    assign layer0_outputs[3990] = ~(inputs[76]) | (inputs[224]);
    assign layer0_outputs[3991] = (inputs[212]) ^ (inputs[19]);
    assign layer0_outputs[3992] = (inputs[176]) & (inputs[193]);
    assign layer0_outputs[3993] = 1'b0;
    assign layer0_outputs[3994] = ~(inputs[81]) | (inputs[105]);
    assign layer0_outputs[3995] = ~((inputs[249]) & (inputs[130]));
    assign layer0_outputs[3996] = (inputs[229]) & ~(inputs[223]);
    assign layer0_outputs[3997] = inputs[227];
    assign layer0_outputs[3998] = ~(inputs[21]) | (inputs[79]);
    assign layer0_outputs[3999] = ~((inputs[126]) & (inputs[50]));
    assign layer0_outputs[4000] = inputs[100];
    assign layer0_outputs[4001] = (inputs[80]) & ~(inputs[12]);
    assign layer0_outputs[4002] = ~((inputs[43]) | (inputs[173]));
    assign layer0_outputs[4003] = ~((inputs[83]) | (inputs[248]));
    assign layer0_outputs[4004] = ~(inputs[106]) | (inputs[240]);
    assign layer0_outputs[4005] = (inputs[13]) & (inputs[113]);
    assign layer0_outputs[4006] = ~(inputs[48]);
    assign layer0_outputs[4007] = ~((inputs[233]) ^ (inputs[61]));
    assign layer0_outputs[4008] = (inputs[247]) | (inputs[183]);
    assign layer0_outputs[4009] = ~((inputs[192]) | (inputs[33]));
    assign layer0_outputs[4010] = (inputs[37]) | (inputs[63]);
    assign layer0_outputs[4011] = ~(inputs[22]);
    assign layer0_outputs[4012] = ~(inputs[80]);
    assign layer0_outputs[4013] = ~(inputs[72]);
    assign layer0_outputs[4014] = (inputs[111]) ^ (inputs[240]);
    assign layer0_outputs[4015] = inputs[195];
    assign layer0_outputs[4016] = (inputs[55]) ^ (inputs[230]);
    assign layer0_outputs[4017] = (inputs[36]) ^ (inputs[89]);
    assign layer0_outputs[4018] = ~((inputs[78]) | (inputs[106]));
    assign layer0_outputs[4019] = 1'b0;
    assign layer0_outputs[4020] = ~(inputs[65]);
    assign layer0_outputs[4021] = (inputs[155]) & ~(inputs[36]);
    assign layer0_outputs[4022] = inputs[101];
    assign layer0_outputs[4023] = (inputs[111]) & ~(inputs[227]);
    assign layer0_outputs[4024] = ~((inputs[101]) | (inputs[77]));
    assign layer0_outputs[4025] = ~((inputs[40]) | (inputs[26]));
    assign layer0_outputs[4026] = inputs[86];
    assign layer0_outputs[4027] = ~(inputs[88]);
    assign layer0_outputs[4028] = (inputs[176]) & ~(inputs[35]);
    assign layer0_outputs[4029] = (inputs[120]) & ~(inputs[16]);
    assign layer0_outputs[4030] = (inputs[216]) & ~(inputs[248]);
    assign layer0_outputs[4031] = inputs[3];
    assign layer0_outputs[4032] = ~(inputs[114]);
    assign layer0_outputs[4033] = (inputs[134]) & ~(inputs[108]);
    assign layer0_outputs[4034] = ~(inputs[213]);
    assign layer0_outputs[4035] = ~(inputs[137]);
    assign layer0_outputs[4036] = (inputs[73]) | (inputs[97]);
    assign layer0_outputs[4037] = ~(inputs[18]) | (inputs[161]);
    assign layer0_outputs[4038] = inputs[190];
    assign layer0_outputs[4039] = (inputs[104]) & ~(inputs[167]);
    assign layer0_outputs[4040] = (inputs[32]) & (inputs[60]);
    assign layer0_outputs[4041] = (inputs[58]) & ~(inputs[38]);
    assign layer0_outputs[4042] = 1'b0;
    assign layer0_outputs[4043] = inputs[139];
    assign layer0_outputs[4044] = (inputs[69]) | (inputs[196]);
    assign layer0_outputs[4045] = ~((inputs[34]) | (inputs[164]));
    assign layer0_outputs[4046] = (inputs[124]) | (inputs[87]);
    assign layer0_outputs[4047] = ~(inputs[75]) | (inputs[162]);
    assign layer0_outputs[4048] = ~(inputs[105]);
    assign layer0_outputs[4049] = inputs[140];
    assign layer0_outputs[4050] = ~(inputs[230]);
    assign layer0_outputs[4051] = ~(inputs[196]);
    assign layer0_outputs[4052] = (inputs[199]) & ~(inputs[249]);
    assign layer0_outputs[4053] = (inputs[252]) ^ (inputs[148]);
    assign layer0_outputs[4054] = (inputs[172]) | (inputs[176]);
    assign layer0_outputs[4055] = ~((inputs[8]) & (inputs[10]));
    assign layer0_outputs[4056] = ~(inputs[245]) | (inputs[191]);
    assign layer0_outputs[4057] = ~(inputs[11]) | (inputs[18]);
    assign layer0_outputs[4058] = ~(inputs[85]) | (inputs[163]);
    assign layer0_outputs[4059] = ~(inputs[100]) | (inputs[5]);
    assign layer0_outputs[4060] = ~(inputs[71]) | (inputs[111]);
    assign layer0_outputs[4061] = ~((inputs[114]) & (inputs[228]));
    assign layer0_outputs[4062] = (inputs[242]) & ~(inputs[176]);
    assign layer0_outputs[4063] = ~(inputs[75]) | (inputs[66]);
    assign layer0_outputs[4064] = (inputs[107]) | (inputs[176]);
    assign layer0_outputs[4065] = ~((inputs[135]) | (inputs[120]));
    assign layer0_outputs[4066] = ~(inputs[221]);
    assign layer0_outputs[4067] = 1'b1;
    assign layer0_outputs[4068] = ~(inputs[193]);
    assign layer0_outputs[4069] = inputs[170];
    assign layer0_outputs[4070] = inputs[249];
    assign layer0_outputs[4071] = (inputs[224]) & ~(inputs[140]);
    assign layer0_outputs[4072] = ~((inputs[95]) | (inputs[155]));
    assign layer0_outputs[4073] = ~(inputs[152]);
    assign layer0_outputs[4074] = ~(inputs[196]);
    assign layer0_outputs[4075] = ~((inputs[26]) ^ (inputs[225]));
    assign layer0_outputs[4076] = (inputs[204]) | (inputs[177]);
    assign layer0_outputs[4077] = ~((inputs[230]) ^ (inputs[67]));
    assign layer0_outputs[4078] = ~((inputs[48]) ^ (inputs[153]));
    assign layer0_outputs[4079] = ~((inputs[199]) | (inputs[156]));
    assign layer0_outputs[4080] = inputs[88];
    assign layer0_outputs[4081] = 1'b1;
    assign layer0_outputs[4082] = ~(inputs[46]);
    assign layer0_outputs[4083] = (inputs[1]) & ~(inputs[250]);
    assign layer0_outputs[4084] = (inputs[193]) ^ (inputs[57]);
    assign layer0_outputs[4085] = (inputs[79]) ^ (inputs[135]);
    assign layer0_outputs[4086] = (inputs[84]) ^ (inputs[133]);
    assign layer0_outputs[4087] = ~(inputs[198]) | (inputs[35]);
    assign layer0_outputs[4088] = ~(inputs[159]) | (inputs[33]);
    assign layer0_outputs[4089] = ~(inputs[162]);
    assign layer0_outputs[4090] = ~(inputs[221]);
    assign layer0_outputs[4091] = (inputs[13]) & (inputs[204]);
    assign layer0_outputs[4092] = ~(inputs[198]) | (inputs[105]);
    assign layer0_outputs[4093] = ~((inputs[68]) | (inputs[181]));
    assign layer0_outputs[4094] = (inputs[137]) & ~(inputs[204]);
    assign layer0_outputs[4095] = (inputs[209]) & ~(inputs[63]);
    assign layer0_outputs[4096] = ~((inputs[123]) | (inputs[109]));
    assign layer0_outputs[4097] = ~(inputs[43]) | (inputs[92]);
    assign layer0_outputs[4098] = ~((inputs[35]) & (inputs[241]));
    assign layer0_outputs[4099] = (inputs[231]) & ~(inputs[155]);
    assign layer0_outputs[4100] = inputs[60];
    assign layer0_outputs[4101] = (inputs[98]) | (inputs[253]);
    assign layer0_outputs[4102] = inputs[204];
    assign layer0_outputs[4103] = ~((inputs[134]) | (inputs[10]));
    assign layer0_outputs[4104] = (inputs[36]) ^ (inputs[36]);
    assign layer0_outputs[4105] = ~(inputs[235]);
    assign layer0_outputs[4106] = ~((inputs[134]) | (inputs[116]));
    assign layer0_outputs[4107] = ~(inputs[117]) | (inputs[109]);
    assign layer0_outputs[4108] = ~(inputs[129]) | (inputs[99]);
    assign layer0_outputs[4109] = ~((inputs[56]) | (inputs[114]));
    assign layer0_outputs[4110] = 1'b0;
    assign layer0_outputs[4111] = ~((inputs[180]) | (inputs[204]));
    assign layer0_outputs[4112] = (inputs[81]) ^ (inputs[240]);
    assign layer0_outputs[4113] = inputs[59];
    assign layer0_outputs[4114] = (inputs[112]) ^ (inputs[254]);
    assign layer0_outputs[4115] = ~(inputs[119]) | (inputs[148]);
    assign layer0_outputs[4116] = ~((inputs[149]) | (inputs[164]));
    assign layer0_outputs[4117] = ~((inputs[119]) | (inputs[63]));
    assign layer0_outputs[4118] = ~(inputs[84]) | (inputs[227]);
    assign layer0_outputs[4119] = ~(inputs[5]) | (inputs[207]);
    assign layer0_outputs[4120] = ~(inputs[163]) | (inputs[109]);
    assign layer0_outputs[4121] = ~((inputs[43]) ^ (inputs[218]));
    assign layer0_outputs[4122] = ~(inputs[106]);
    assign layer0_outputs[4123] = inputs[196];
    assign layer0_outputs[4124] = inputs[187];
    assign layer0_outputs[4125] = ~((inputs[113]) ^ (inputs[132]));
    assign layer0_outputs[4126] = (inputs[192]) & (inputs[127]);
    assign layer0_outputs[4127] = ~((inputs[217]) | (inputs[177]));
    assign layer0_outputs[4128] = inputs[83];
    assign layer0_outputs[4129] = ~((inputs[226]) & (inputs[211]));
    assign layer0_outputs[4130] = ~(inputs[62]);
    assign layer0_outputs[4131] = ~((inputs[173]) | (inputs[43]));
    assign layer0_outputs[4132] = ~(inputs[180]);
    assign layer0_outputs[4133] = ~(inputs[81]);
    assign layer0_outputs[4134] = ~(inputs[83]);
    assign layer0_outputs[4135] = (inputs[171]) & ~(inputs[82]);
    assign layer0_outputs[4136] = inputs[183];
    assign layer0_outputs[4137] = (inputs[174]) ^ (inputs[14]);
    assign layer0_outputs[4138] = inputs[145];
    assign layer0_outputs[4139] = (inputs[168]) & ~(inputs[19]);
    assign layer0_outputs[4140] = ~(inputs[187]) | (inputs[51]);
    assign layer0_outputs[4141] = ~((inputs[200]) | (inputs[207]));
    assign layer0_outputs[4142] = ~(inputs[69]) | (inputs[122]);
    assign layer0_outputs[4143] = ~(inputs[122]) | (inputs[57]);
    assign layer0_outputs[4144] = inputs[52];
    assign layer0_outputs[4145] = ~((inputs[87]) ^ (inputs[125]));
    assign layer0_outputs[4146] = ~((inputs[2]) | (inputs[151]));
    assign layer0_outputs[4147] = ~((inputs[26]) & (inputs[130]));
    assign layer0_outputs[4148] = ~(inputs[141]);
    assign layer0_outputs[4149] = ~((inputs[23]) | (inputs[75]));
    assign layer0_outputs[4150] = ~((inputs[170]) | (inputs[231]));
    assign layer0_outputs[4151] = (inputs[161]) ^ (inputs[81]);
    assign layer0_outputs[4152] = ~(inputs[181]);
    assign layer0_outputs[4153] = ~((inputs[87]) | (inputs[192]));
    assign layer0_outputs[4154] = ~((inputs[225]) & (inputs[81]));
    assign layer0_outputs[4155] = ~((inputs[242]) ^ (inputs[246]));
    assign layer0_outputs[4156] = ~(inputs[133]) | (inputs[39]);
    assign layer0_outputs[4157] = inputs[209];
    assign layer0_outputs[4158] = (inputs[172]) ^ (inputs[6]);
    assign layer0_outputs[4159] = ~(inputs[48]);
    assign layer0_outputs[4160] = ~((inputs[174]) & (inputs[26]));
    assign layer0_outputs[4161] = ~((inputs[123]) ^ (inputs[115]));
    assign layer0_outputs[4162] = ~(inputs[46]) | (inputs[66]);
    assign layer0_outputs[4163] = ~((inputs[4]) | (inputs[107]));
    assign layer0_outputs[4164] = ~(inputs[136]) | (inputs[106]);
    assign layer0_outputs[4165] = ~(inputs[40]);
    assign layer0_outputs[4166] = ~((inputs[211]) | (inputs[15]));
    assign layer0_outputs[4167] = ~((inputs[47]) | (inputs[89]));
    assign layer0_outputs[4168] = (inputs[117]) & ~(inputs[129]);
    assign layer0_outputs[4169] = (inputs[1]) & ~(inputs[27]);
    assign layer0_outputs[4170] = (inputs[89]) ^ (inputs[33]);
    assign layer0_outputs[4171] = (inputs[48]) | (inputs[102]);
    assign layer0_outputs[4172] = ~((inputs[177]) | (inputs[202]));
    assign layer0_outputs[4173] = (inputs[56]) & ~(inputs[202]);
    assign layer0_outputs[4174] = ~(inputs[90]) | (inputs[7]);
    assign layer0_outputs[4175] = (inputs[196]) & ~(inputs[115]);
    assign layer0_outputs[4176] = ~((inputs[149]) | (inputs[92]));
    assign layer0_outputs[4177] = ~(inputs[116]) | (inputs[5]);
    assign layer0_outputs[4178] = (inputs[134]) ^ (inputs[44]);
    assign layer0_outputs[4179] = ~((inputs[90]) ^ (inputs[145]));
    assign layer0_outputs[4180] = ~(inputs[88]) | (inputs[63]);
    assign layer0_outputs[4181] = ~(inputs[121]) | (inputs[113]);
    assign layer0_outputs[4182] = (inputs[29]) & ~(inputs[226]);
    assign layer0_outputs[4183] = ~((inputs[58]) ^ (inputs[243]));
    assign layer0_outputs[4184] = ~(inputs[133]);
    assign layer0_outputs[4185] = (inputs[21]) | (inputs[223]);
    assign layer0_outputs[4186] = ~(inputs[135]);
    assign layer0_outputs[4187] = ~(inputs[168]) | (inputs[108]);
    assign layer0_outputs[4188] = (inputs[75]) | (inputs[190]);
    assign layer0_outputs[4189] = (inputs[121]) & ~(inputs[53]);
    assign layer0_outputs[4190] = ~(inputs[137]) | (inputs[109]);
    assign layer0_outputs[4191] = (inputs[21]) & (inputs[248]);
    assign layer0_outputs[4192] = (inputs[234]) ^ (inputs[146]);
    assign layer0_outputs[4193] = (inputs[206]) | (inputs[196]);
    assign layer0_outputs[4194] = 1'b0;
    assign layer0_outputs[4195] = ~(inputs[198]);
    assign layer0_outputs[4196] = (inputs[133]) | (inputs[101]);
    assign layer0_outputs[4197] = (inputs[162]) & ~(inputs[65]);
    assign layer0_outputs[4198] = inputs[198];
    assign layer0_outputs[4199] = (inputs[34]) & (inputs[47]);
    assign layer0_outputs[4200] = ~((inputs[232]) ^ (inputs[40]));
    assign layer0_outputs[4201] = (inputs[244]) & ~(inputs[26]);
    assign layer0_outputs[4202] = (inputs[188]) & ~(inputs[48]);
    assign layer0_outputs[4203] = ~(inputs[201]);
    assign layer0_outputs[4204] = ~(inputs[123]) | (inputs[94]);
    assign layer0_outputs[4205] = 1'b0;
    assign layer0_outputs[4206] = ~((inputs[108]) ^ (inputs[106]));
    assign layer0_outputs[4207] = (inputs[32]) & (inputs[226]);
    assign layer0_outputs[4208] = ~(inputs[93]);
    assign layer0_outputs[4209] = (inputs[117]) ^ (inputs[65]);
    assign layer0_outputs[4210] = (inputs[209]) ^ (inputs[40]);
    assign layer0_outputs[4211] = ~((inputs[213]) | (inputs[70]));
    assign layer0_outputs[4212] = ~(inputs[49]);
    assign layer0_outputs[4213] = (inputs[141]) | (inputs[41]);
    assign layer0_outputs[4214] = ~(inputs[72]);
    assign layer0_outputs[4215] = ~(inputs[88]) | (inputs[10]);
    assign layer0_outputs[4216] = ~((inputs[135]) ^ (inputs[141]));
    assign layer0_outputs[4217] = ~((inputs[243]) | (inputs[126]));
    assign layer0_outputs[4218] = ~(inputs[56]) | (inputs[255]);
    assign layer0_outputs[4219] = inputs[232];
    assign layer0_outputs[4220] = ~(inputs[92]);
    assign layer0_outputs[4221] = (inputs[67]) & ~(inputs[126]);
    assign layer0_outputs[4222] = ~(inputs[117]);
    assign layer0_outputs[4223] = (inputs[183]) | (inputs[205]);
    assign layer0_outputs[4224] = (inputs[199]) | (inputs[111]);
    assign layer0_outputs[4225] = inputs[120];
    assign layer0_outputs[4226] = ~(inputs[220]) | (inputs[97]);
    assign layer0_outputs[4227] = inputs[164];
    assign layer0_outputs[4228] = (inputs[116]) & ~(inputs[231]);
    assign layer0_outputs[4229] = ~((inputs[149]) | (inputs[117]));
    assign layer0_outputs[4230] = (inputs[19]) | (inputs[142]);
    assign layer0_outputs[4231] = (inputs[71]) | (inputs[204]);
    assign layer0_outputs[4232] = ~(inputs[39]) | (inputs[113]);
    assign layer0_outputs[4233] = 1'b0;
    assign layer0_outputs[4234] = ~(inputs[86]);
    assign layer0_outputs[4235] = ~(inputs[133]);
    assign layer0_outputs[4236] = inputs[182];
    assign layer0_outputs[4237] = ~(inputs[89]);
    assign layer0_outputs[4238] = (inputs[89]) | (inputs[253]);
    assign layer0_outputs[4239] = ~((inputs[12]) & (inputs[180]));
    assign layer0_outputs[4240] = (inputs[231]) ^ (inputs[46]);
    assign layer0_outputs[4241] = (inputs[176]) ^ (inputs[131]);
    assign layer0_outputs[4242] = ~((inputs[52]) | (inputs[134]));
    assign layer0_outputs[4243] = inputs[25];
    assign layer0_outputs[4244] = (inputs[185]) & ~(inputs[94]);
    assign layer0_outputs[4245] = (inputs[99]) & ~(inputs[60]);
    assign layer0_outputs[4246] = (inputs[37]) | (inputs[242]);
    assign layer0_outputs[4247] = ~((inputs[76]) | (inputs[216]));
    assign layer0_outputs[4248] = (inputs[253]) & ~(inputs[34]);
    assign layer0_outputs[4249] = (inputs[48]) ^ (inputs[151]);
    assign layer0_outputs[4250] = (inputs[213]) & ~(inputs[52]);
    assign layer0_outputs[4251] = ~((inputs[77]) | (inputs[1]));
    assign layer0_outputs[4252] = ~((inputs[73]) ^ (inputs[121]));
    assign layer0_outputs[4253] = inputs[135];
    assign layer0_outputs[4254] = (inputs[25]) | (inputs[186]);
    assign layer0_outputs[4255] = (inputs[150]) & ~(inputs[31]);
    assign layer0_outputs[4256] = ~(inputs[214]) | (inputs[249]);
    assign layer0_outputs[4257] = (inputs[1]) & ~(inputs[35]);
    assign layer0_outputs[4258] = ~((inputs[162]) | (inputs[215]));
    assign layer0_outputs[4259] = inputs[239];
    assign layer0_outputs[4260] = inputs[91];
    assign layer0_outputs[4261] = 1'b1;
    assign layer0_outputs[4262] = (inputs[225]) ^ (inputs[157]);
    assign layer0_outputs[4263] = inputs[200];
    assign layer0_outputs[4264] = (inputs[250]) | (inputs[189]);
    assign layer0_outputs[4265] = ~(inputs[24]);
    assign layer0_outputs[4266] = (inputs[150]) & ~(inputs[213]);
    assign layer0_outputs[4267] = (inputs[157]) | (inputs[47]);
    assign layer0_outputs[4268] = ~(inputs[69]) | (inputs[209]);
    assign layer0_outputs[4269] = (inputs[0]) | (inputs[150]);
    assign layer0_outputs[4270] = (inputs[58]) ^ (inputs[179]);
    assign layer0_outputs[4271] = ~(inputs[135]) | (inputs[27]);
    assign layer0_outputs[4272] = ~((inputs[232]) ^ (inputs[45]));
    assign layer0_outputs[4273] = ~(inputs[61]) | (inputs[175]);
    assign layer0_outputs[4274] = ~((inputs[215]) ^ (inputs[80]));
    assign layer0_outputs[4275] = ~(inputs[58]) | (inputs[39]);
    assign layer0_outputs[4276] = ~(inputs[39]);
    assign layer0_outputs[4277] = (inputs[157]) ^ (inputs[184]);
    assign layer0_outputs[4278] = (inputs[171]) | (inputs[154]);
    assign layer0_outputs[4279] = (inputs[122]) & ~(inputs[45]);
    assign layer0_outputs[4280] = (inputs[19]) | (inputs[87]);
    assign layer0_outputs[4281] = ~((inputs[104]) ^ (inputs[20]));
    assign layer0_outputs[4282] = ~(inputs[219]) | (inputs[35]);
    assign layer0_outputs[4283] = ~(inputs[213]) | (inputs[252]);
    assign layer0_outputs[4284] = ~(inputs[38]);
    assign layer0_outputs[4285] = ~((inputs[168]) ^ (inputs[112]));
    assign layer0_outputs[4286] = ~(inputs[107]);
    assign layer0_outputs[4287] = ~(inputs[4]) | (inputs[63]);
    assign layer0_outputs[4288] = (inputs[37]) | (inputs[193]);
    assign layer0_outputs[4289] = 1'b1;
    assign layer0_outputs[4290] = ~(inputs[56]) | (inputs[235]);
    assign layer0_outputs[4291] = inputs[218];
    assign layer0_outputs[4292] = (inputs[196]) & ~(inputs[225]);
    assign layer0_outputs[4293] = ~(inputs[153]) | (inputs[255]);
    assign layer0_outputs[4294] = ~((inputs[51]) | (inputs[192]));
    assign layer0_outputs[4295] = (inputs[51]) | (inputs[149]);
    assign layer0_outputs[4296] = (inputs[151]) | (inputs[230]);
    assign layer0_outputs[4297] = (inputs[243]) | (inputs[215]);
    assign layer0_outputs[4298] = (inputs[72]) & ~(inputs[161]);
    assign layer0_outputs[4299] = 1'b0;
    assign layer0_outputs[4300] = (inputs[79]) | (inputs[230]);
    assign layer0_outputs[4301] = ~(inputs[49]);
    assign layer0_outputs[4302] = 1'b0;
    assign layer0_outputs[4303] = ~((inputs[14]) ^ (inputs[169]));
    assign layer0_outputs[4304] = (inputs[113]) ^ (inputs[67]);
    assign layer0_outputs[4305] = ~(inputs[12]);
    assign layer0_outputs[4306] = (inputs[121]) ^ (inputs[254]);
    assign layer0_outputs[4307] = (inputs[71]) & ~(inputs[187]);
    assign layer0_outputs[4308] = (inputs[78]) | (inputs[107]);
    assign layer0_outputs[4309] = ~(inputs[10]) | (inputs[33]);
    assign layer0_outputs[4310] = (inputs[233]) | (inputs[10]);
    assign layer0_outputs[4311] = (inputs[187]) & ~(inputs[160]);
    assign layer0_outputs[4312] = (inputs[117]) | (inputs[86]);
    assign layer0_outputs[4313] = inputs[92];
    assign layer0_outputs[4314] = ~((inputs[192]) | (inputs[182]));
    assign layer0_outputs[4315] = ~((inputs[104]) ^ (inputs[201]));
    assign layer0_outputs[4316] = inputs[160];
    assign layer0_outputs[4317] = ~(inputs[23]);
    assign layer0_outputs[4318] = ~(inputs[50]);
    assign layer0_outputs[4319] = (inputs[173]) ^ (inputs[152]);
    assign layer0_outputs[4320] = ~((inputs[124]) ^ (inputs[62]));
    assign layer0_outputs[4321] = ~((inputs[157]) | (inputs[212]));
    assign layer0_outputs[4322] = (inputs[168]) & ~(inputs[195]);
    assign layer0_outputs[4323] = inputs[229];
    assign layer0_outputs[4324] = ~(inputs[153]);
    assign layer0_outputs[4325] = ~(inputs[160]);
    assign layer0_outputs[4326] = ~((inputs[59]) | (inputs[205]));
    assign layer0_outputs[4327] = (inputs[123]) & ~(inputs[2]);
    assign layer0_outputs[4328] = ~(inputs[229]) | (inputs[157]);
    assign layer0_outputs[4329] = ~(inputs[187]);
    assign layer0_outputs[4330] = inputs[101];
    assign layer0_outputs[4331] = (inputs[103]) & ~(inputs[130]);
    assign layer0_outputs[4332] = inputs[222];
    assign layer0_outputs[4333] = (inputs[99]) & ~(inputs[69]);
    assign layer0_outputs[4334] = (inputs[109]) & ~(inputs[51]);
    assign layer0_outputs[4335] = (inputs[53]) | (inputs[55]);
    assign layer0_outputs[4336] = inputs[102];
    assign layer0_outputs[4337] = ~((inputs[130]) | (inputs[18]));
    assign layer0_outputs[4338] = ~(inputs[8]);
    assign layer0_outputs[4339] = ~((inputs[151]) ^ (inputs[49]));
    assign layer0_outputs[4340] = 1'b1;
    assign layer0_outputs[4341] = (inputs[31]) ^ (inputs[112]);
    assign layer0_outputs[4342] = (inputs[74]) & (inputs[33]);
    assign layer0_outputs[4343] = ~(inputs[179]) | (inputs[38]);
    assign layer0_outputs[4344] = (inputs[20]) & ~(inputs[104]);
    assign layer0_outputs[4345] = ~((inputs[172]) ^ (inputs[255]));
    assign layer0_outputs[4346] = ~(inputs[122]) | (inputs[205]);
    assign layer0_outputs[4347] = (inputs[106]) & ~(inputs[115]);
    assign layer0_outputs[4348] = (inputs[79]) & (inputs[174]);
    assign layer0_outputs[4349] = (inputs[15]) & ~(inputs[17]);
    assign layer0_outputs[4350] = (inputs[254]) & ~(inputs[176]);
    assign layer0_outputs[4351] = ~(inputs[65]);
    assign layer0_outputs[4352] = inputs[67];
    assign layer0_outputs[4353] = (inputs[151]) & ~(inputs[45]);
    assign layer0_outputs[4354] = ~((inputs[169]) ^ (inputs[183]));
    assign layer0_outputs[4355] = (inputs[244]) ^ (inputs[122]);
    assign layer0_outputs[4356] = (inputs[90]) & ~(inputs[68]);
    assign layer0_outputs[4357] = ~((inputs[141]) | (inputs[200]));
    assign layer0_outputs[4358] = ~((inputs[142]) ^ (inputs[0]));
    assign layer0_outputs[4359] = (inputs[187]) | (inputs[80]);
    assign layer0_outputs[4360] = ~((inputs[121]) ^ (inputs[242]));
    assign layer0_outputs[4361] = ~(inputs[107]) | (inputs[149]);
    assign layer0_outputs[4362] = ~(inputs[56]) | (inputs[100]);
    assign layer0_outputs[4363] = ~(inputs[194]) | (inputs[25]);
    assign layer0_outputs[4364] = ~((inputs[10]) | (inputs[90]));
    assign layer0_outputs[4365] = ~((inputs[234]) ^ (inputs[252]));
    assign layer0_outputs[4366] = ~(inputs[42]);
    assign layer0_outputs[4367] = ~((inputs[55]) ^ (inputs[195]));
    assign layer0_outputs[4368] = (inputs[246]) | (inputs[103]);
    assign layer0_outputs[4369] = ~((inputs[153]) ^ (inputs[13]));
    assign layer0_outputs[4370] = ~(inputs[92]) | (inputs[22]);
    assign layer0_outputs[4371] = (inputs[95]) | (inputs[182]);
    assign layer0_outputs[4372] = inputs[178];
    assign layer0_outputs[4373] = ~(inputs[36]) | (inputs[109]);
    assign layer0_outputs[4374] = ~(inputs[57]);
    assign layer0_outputs[4375] = (inputs[145]) | (inputs[85]);
    assign layer0_outputs[4376] = (inputs[83]) | (inputs[91]);
    assign layer0_outputs[4377] = ~((inputs[125]) | (inputs[180]));
    assign layer0_outputs[4378] = (inputs[137]) & ~(inputs[225]);
    assign layer0_outputs[4379] = ~(inputs[120]);
    assign layer0_outputs[4380] = ~((inputs[91]) | (inputs[98]));
    assign layer0_outputs[4381] = ~((inputs[186]) | (inputs[181]));
    assign layer0_outputs[4382] = 1'b0;
    assign layer0_outputs[4383] = (inputs[117]) | (inputs[62]);
    assign layer0_outputs[4384] = ~(inputs[146]);
    assign layer0_outputs[4385] = (inputs[200]) ^ (inputs[169]);
    assign layer0_outputs[4386] = (inputs[17]) & ~(inputs[228]);
    assign layer0_outputs[4387] = (inputs[117]) | (inputs[13]);
    assign layer0_outputs[4388] = (inputs[59]) & ~(inputs[247]);
    assign layer0_outputs[4389] = ~((inputs[180]) ^ (inputs[34]));
    assign layer0_outputs[4390] = (inputs[37]) | (inputs[25]);
    assign layer0_outputs[4391] = (inputs[32]) & (inputs[35]);
    assign layer0_outputs[4392] = (inputs[67]) & ~(inputs[0]);
    assign layer0_outputs[4393] = (inputs[24]) & ~(inputs[44]);
    assign layer0_outputs[4394] = (inputs[186]) ^ (inputs[33]);
    assign layer0_outputs[4395] = ~(inputs[54]);
    assign layer0_outputs[4396] = ~(inputs[198]);
    assign layer0_outputs[4397] = ~(inputs[106]);
    assign layer0_outputs[4398] = ~(inputs[186]) | (inputs[183]);
    assign layer0_outputs[4399] = ~((inputs[51]) | (inputs[217]));
    assign layer0_outputs[4400] = ~(inputs[80]);
    assign layer0_outputs[4401] = ~(inputs[3]);
    assign layer0_outputs[4402] = ~(inputs[67]);
    assign layer0_outputs[4403] = ~((inputs[113]) & (inputs[224]));
    assign layer0_outputs[4404] = ~(inputs[163]) | (inputs[3]);
    assign layer0_outputs[4405] = inputs[45];
    assign layer0_outputs[4406] = ~((inputs[248]) & (inputs[57]));
    assign layer0_outputs[4407] = inputs[189];
    assign layer0_outputs[4408] = (inputs[118]) & ~(inputs[17]);
    assign layer0_outputs[4409] = ~(inputs[181]);
    assign layer0_outputs[4410] = ~((inputs[131]) ^ (inputs[244]));
    assign layer0_outputs[4411] = ~((inputs[167]) ^ (inputs[147]));
    assign layer0_outputs[4412] = ~((inputs[29]) | (inputs[60]));
    assign layer0_outputs[4413] = (inputs[121]) & ~(inputs[62]);
    assign layer0_outputs[4414] = ~(inputs[181]) | (inputs[103]);
    assign layer0_outputs[4415] = ~((inputs[149]) | (inputs[247]));
    assign layer0_outputs[4416] = ~((inputs[90]) ^ (inputs[213]));
    assign layer0_outputs[4417] = ~(inputs[84]) | (inputs[4]);
    assign layer0_outputs[4418] = (inputs[170]) & ~(inputs[42]);
    assign layer0_outputs[4419] = inputs[245];
    assign layer0_outputs[4420] = ~(inputs[162]) | (inputs[125]);
    assign layer0_outputs[4421] = ~((inputs[195]) | (inputs[158]));
    assign layer0_outputs[4422] = ~(inputs[113]);
    assign layer0_outputs[4423] = (inputs[239]) ^ (inputs[101]);
    assign layer0_outputs[4424] = inputs[55];
    assign layer0_outputs[4425] = inputs[35];
    assign layer0_outputs[4426] = ~((inputs[83]) | (inputs[36]));
    assign layer0_outputs[4427] = ~((inputs[106]) | (inputs[215]));
    assign layer0_outputs[4428] = ~(inputs[23]) | (inputs[222]);
    assign layer0_outputs[4429] = ~((inputs[163]) | (inputs[189]));
    assign layer0_outputs[4430] = inputs[56];
    assign layer0_outputs[4431] = inputs[131];
    assign layer0_outputs[4432] = ~(inputs[112]) | (inputs[142]);
    assign layer0_outputs[4433] = ~(inputs[90]);
    assign layer0_outputs[4434] = inputs[172];
    assign layer0_outputs[4435] = ~((inputs[102]) ^ (inputs[209]));
    assign layer0_outputs[4436] = ~(inputs[135]);
    assign layer0_outputs[4437] = ~(inputs[244]);
    assign layer0_outputs[4438] = inputs[73];
    assign layer0_outputs[4439] = ~((inputs[194]) ^ (inputs[32]));
    assign layer0_outputs[4440] = ~((inputs[210]) | (inputs[205]));
    assign layer0_outputs[4441] = ~(inputs[225]);
    assign layer0_outputs[4442] = ~(inputs[113]);
    assign layer0_outputs[4443] = inputs[165];
    assign layer0_outputs[4444] = ~(inputs[135]) | (inputs[52]);
    assign layer0_outputs[4445] = (inputs[32]) & (inputs[51]);
    assign layer0_outputs[4446] = inputs[245];
    assign layer0_outputs[4447] = ~(inputs[220]) | (inputs[21]);
    assign layer0_outputs[4448] = ~((inputs[61]) | (inputs[32]));
    assign layer0_outputs[4449] = ~(inputs[181]);
    assign layer0_outputs[4450] = (inputs[238]) | (inputs[134]);
    assign layer0_outputs[4451] = ~((inputs[94]) ^ (inputs[233]));
    assign layer0_outputs[4452] = ~(inputs[216]);
    assign layer0_outputs[4453] = ~((inputs[99]) ^ (inputs[1]));
    assign layer0_outputs[4454] = 1'b0;
    assign layer0_outputs[4455] = ~((inputs[158]) | (inputs[22]));
    assign layer0_outputs[4456] = inputs[166];
    assign layer0_outputs[4457] = (inputs[127]) | (inputs[251]);
    assign layer0_outputs[4458] = (inputs[238]) & (inputs[89]);
    assign layer0_outputs[4459] = inputs[119];
    assign layer0_outputs[4460] = (inputs[210]) ^ (inputs[231]);
    assign layer0_outputs[4461] = (inputs[93]) | (inputs[198]);
    assign layer0_outputs[4462] = ~(inputs[68]) | (inputs[235]);
    assign layer0_outputs[4463] = (inputs[21]) & (inputs[51]);
    assign layer0_outputs[4464] = inputs[105];
    assign layer0_outputs[4465] = ~(inputs[155]) | (inputs[109]);
    assign layer0_outputs[4466] = (inputs[15]) | (inputs[217]);
    assign layer0_outputs[4467] = (inputs[153]) & ~(inputs[177]);
    assign layer0_outputs[4468] = ~(inputs[160]);
    assign layer0_outputs[4469] = (inputs[94]) & ~(inputs[10]);
    assign layer0_outputs[4470] = ~((inputs[253]) ^ (inputs[3]));
    assign layer0_outputs[4471] = ~((inputs[78]) & (inputs[254]));
    assign layer0_outputs[4472] = inputs[190];
    assign layer0_outputs[4473] = ~((inputs[154]) & (inputs[27]));
    assign layer0_outputs[4474] = ~(inputs[81]);
    assign layer0_outputs[4475] = inputs[182];
    assign layer0_outputs[4476] = (inputs[36]) | (inputs[122]);
    assign layer0_outputs[4477] = ~((inputs[28]) | (inputs[170]));
    assign layer0_outputs[4478] = (inputs[3]) | (inputs[134]);
    assign layer0_outputs[4479] = inputs[57];
    assign layer0_outputs[4480] = ~(inputs[111]);
    assign layer0_outputs[4481] = (inputs[78]) ^ (inputs[195]);
    assign layer0_outputs[4482] = ~(inputs[59]);
    assign layer0_outputs[4483] = inputs[95];
    assign layer0_outputs[4484] = (inputs[58]) & ~(inputs[231]);
    assign layer0_outputs[4485] = ~(inputs[205]);
    assign layer0_outputs[4486] = (inputs[89]) ^ (inputs[159]);
    assign layer0_outputs[4487] = ~(inputs[19]);
    assign layer0_outputs[4488] = 1'b1;
    assign layer0_outputs[4489] = ~(inputs[93]) | (inputs[46]);
    assign layer0_outputs[4490] = (inputs[122]) ^ (inputs[49]);
    assign layer0_outputs[4491] = ~(inputs[121]);
    assign layer0_outputs[4492] = ~((inputs[102]) | (inputs[87]));
    assign layer0_outputs[4493] = ~(inputs[168]) | (inputs[220]);
    assign layer0_outputs[4494] = (inputs[166]) ^ (inputs[103]);
    assign layer0_outputs[4495] = (inputs[34]) ^ (inputs[217]);
    assign layer0_outputs[4496] = ~(inputs[213]) | (inputs[189]);
    assign layer0_outputs[4497] = ~(inputs[39]);
    assign layer0_outputs[4498] = (inputs[163]) | (inputs[52]);
    assign layer0_outputs[4499] = ~(inputs[255]) | (inputs[29]);
    assign layer0_outputs[4500] = ~(inputs[87]) | (inputs[147]);
    assign layer0_outputs[4501] = ~((inputs[237]) ^ (inputs[232]));
    assign layer0_outputs[4502] = (inputs[154]) | (inputs[211]);
    assign layer0_outputs[4503] = (inputs[67]) & ~(inputs[124]);
    assign layer0_outputs[4504] = ~((inputs[203]) ^ (inputs[34]));
    assign layer0_outputs[4505] = ~((inputs[41]) | (inputs[119]));
    assign layer0_outputs[4506] = inputs[114];
    assign layer0_outputs[4507] = inputs[198];
    assign layer0_outputs[4508] = ~(inputs[170]);
    assign layer0_outputs[4509] = ~((inputs[118]) ^ (inputs[222]));
    assign layer0_outputs[4510] = (inputs[226]) ^ (inputs[157]);
    assign layer0_outputs[4511] = ~(inputs[57]);
    assign layer0_outputs[4512] = inputs[239];
    assign layer0_outputs[4513] = ~(inputs[102]) | (inputs[213]);
    assign layer0_outputs[4514] = ~(inputs[133]);
    assign layer0_outputs[4515] = (inputs[214]) & ~(inputs[25]);
    assign layer0_outputs[4516] = ~((inputs[176]) ^ (inputs[23]));
    assign layer0_outputs[4517] = ~(inputs[122]) | (inputs[61]);
    assign layer0_outputs[4518] = 1'b1;
    assign layer0_outputs[4519] = 1'b0;
    assign layer0_outputs[4520] = (inputs[167]) ^ (inputs[0]);
    assign layer0_outputs[4521] = ~(inputs[183]) | (inputs[227]);
    assign layer0_outputs[4522] = ~((inputs[132]) & (inputs[73]));
    assign layer0_outputs[4523] = ~((inputs[39]) | (inputs[53]));
    assign layer0_outputs[4524] = ~((inputs[133]) & (inputs[139]));
    assign layer0_outputs[4525] = (inputs[222]) & (inputs[4]);
    assign layer0_outputs[4526] = ~((inputs[53]) | (inputs[39]));
    assign layer0_outputs[4527] = ~((inputs[193]) ^ (inputs[75]));
    assign layer0_outputs[4528] = (inputs[181]) & ~(inputs[145]);
    assign layer0_outputs[4529] = (inputs[190]) | (inputs[186]);
    assign layer0_outputs[4530] = ~(inputs[121]);
    assign layer0_outputs[4531] = ~((inputs[41]) | (inputs[210]));
    assign layer0_outputs[4532] = ~(inputs[122]);
    assign layer0_outputs[4533] = inputs[197];
    assign layer0_outputs[4534] = inputs[116];
    assign layer0_outputs[4535] = ~(inputs[207]);
    assign layer0_outputs[4536] = ~((inputs[30]) ^ (inputs[151]));
    assign layer0_outputs[4537] = 1'b0;
    assign layer0_outputs[4538] = (inputs[210]) | (inputs[76]);
    assign layer0_outputs[4539] = ~((inputs[64]) & (inputs[48]));
    assign layer0_outputs[4540] = ~(inputs[218]) | (inputs[238]);
    assign layer0_outputs[4541] = ~((inputs[63]) ^ (inputs[199]));
    assign layer0_outputs[4542] = inputs[165];
    assign layer0_outputs[4543] = ~(inputs[57]) | (inputs[192]);
    assign layer0_outputs[4544] = (inputs[70]) | (inputs[66]);
    assign layer0_outputs[4545] = (inputs[150]) & ~(inputs[50]);
    assign layer0_outputs[4546] = ~(inputs[151]) | (inputs[231]);
    assign layer0_outputs[4547] = (inputs[146]) & ~(inputs[61]);
    assign layer0_outputs[4548] = (inputs[216]) ^ (inputs[140]);
    assign layer0_outputs[4549] = (inputs[184]) & ~(inputs[133]);
    assign layer0_outputs[4550] = ~(inputs[54]);
    assign layer0_outputs[4551] = (inputs[58]) & ~(inputs[35]);
    assign layer0_outputs[4552] = inputs[207];
    assign layer0_outputs[4553] = ~((inputs[2]) | (inputs[206]));
    assign layer0_outputs[4554] = inputs[120];
    assign layer0_outputs[4555] = ~((inputs[177]) ^ (inputs[53]));
    assign layer0_outputs[4556] = (inputs[201]) ^ (inputs[237]);
    assign layer0_outputs[4557] = ~((inputs[187]) ^ (inputs[154]));
    assign layer0_outputs[4558] = (inputs[255]) | (inputs[60]);
    assign layer0_outputs[4559] = ~((inputs[20]) ^ (inputs[179]));
    assign layer0_outputs[4560] = ~(inputs[119]) | (inputs[232]);
    assign layer0_outputs[4561] = (inputs[57]) ^ (inputs[194]);
    assign layer0_outputs[4562] = 1'b0;
    assign layer0_outputs[4563] = inputs[148];
    assign layer0_outputs[4564] = ~((inputs[248]) ^ (inputs[242]));
    assign layer0_outputs[4565] = ~(inputs[59]);
    assign layer0_outputs[4566] = (inputs[142]) ^ (inputs[94]);
    assign layer0_outputs[4567] = ~(inputs[249]) | (inputs[250]);
    assign layer0_outputs[4568] = 1'b1;
    assign layer0_outputs[4569] = ~((inputs[84]) | (inputs[238]));
    assign layer0_outputs[4570] = (inputs[90]) & ~(inputs[178]);
    assign layer0_outputs[4571] = (inputs[108]) | (inputs[184]);
    assign layer0_outputs[4572] = ~((inputs[230]) ^ (inputs[206]));
    assign layer0_outputs[4573] = ~((inputs[60]) ^ (inputs[69]));
    assign layer0_outputs[4574] = ~(inputs[148]);
    assign layer0_outputs[4575] = ~((inputs[76]) ^ (inputs[247]));
    assign layer0_outputs[4576] = ~(inputs[16]) | (inputs[80]);
    assign layer0_outputs[4577] = ~(inputs[82]);
    assign layer0_outputs[4578] = (inputs[13]) & (inputs[251]);
    assign layer0_outputs[4579] = ~(inputs[162]) | (inputs[233]);
    assign layer0_outputs[4580] = (inputs[116]) | (inputs[214]);
    assign layer0_outputs[4581] = ~((inputs[47]) ^ (inputs[100]));
    assign layer0_outputs[4582] = (inputs[67]) | (inputs[237]);
    assign layer0_outputs[4583] = inputs[117];
    assign layer0_outputs[4584] = 1'b0;
    assign layer0_outputs[4585] = inputs[233];
    assign layer0_outputs[4586] = ~((inputs[45]) ^ (inputs[249]));
    assign layer0_outputs[4587] = ~((inputs[69]) & (inputs[136]));
    assign layer0_outputs[4588] = inputs[48];
    assign layer0_outputs[4589] = ~(inputs[138]);
    assign layer0_outputs[4590] = ~((inputs[146]) | (inputs[160]));
    assign layer0_outputs[4591] = ~(inputs[121]);
    assign layer0_outputs[4592] = inputs[197];
    assign layer0_outputs[4593] = ~((inputs[201]) & (inputs[215]));
    assign layer0_outputs[4594] = (inputs[219]) | (inputs[59]);
    assign layer0_outputs[4595] = (inputs[134]) | (inputs[230]);
    assign layer0_outputs[4596] = (inputs[232]) | (inputs[52]);
    assign layer0_outputs[4597] = (inputs[138]) ^ (inputs[145]);
    assign layer0_outputs[4598] = (inputs[89]) & ~(inputs[8]);
    assign layer0_outputs[4599] = (inputs[134]) & ~(inputs[3]);
    assign layer0_outputs[4600] = (inputs[77]) & ~(inputs[22]);
    assign layer0_outputs[4601] = ~((inputs[198]) ^ (inputs[77]));
    assign layer0_outputs[4602] = (inputs[112]) & ~(inputs[158]);
    assign layer0_outputs[4603] = inputs[147];
    assign layer0_outputs[4604] = ~(inputs[222]) | (inputs[194]);
    assign layer0_outputs[4605] = (inputs[232]) & ~(inputs[175]);
    assign layer0_outputs[4606] = inputs[216];
    assign layer0_outputs[4607] = ~((inputs[171]) ^ (inputs[18]));
    assign layer0_outputs[4608] = (inputs[219]) | (inputs[124]);
    assign layer0_outputs[4609] = (inputs[199]) & ~(inputs[9]);
    assign layer0_outputs[4610] = ~(inputs[54]);
    assign layer0_outputs[4611] = (inputs[241]) | (inputs[179]);
    assign layer0_outputs[4612] = ~((inputs[187]) | (inputs[189]));
    assign layer0_outputs[4613] = inputs[56];
    assign layer0_outputs[4614] = inputs[170];
    assign layer0_outputs[4615] = inputs[100];
    assign layer0_outputs[4616] = inputs[18];
    assign layer0_outputs[4617] = ~(inputs[207]) | (inputs[248]);
    assign layer0_outputs[4618] = (inputs[11]) & ~(inputs[2]);
    assign layer0_outputs[4619] = ~(inputs[165]);
    assign layer0_outputs[4620] = ~((inputs[69]) ^ (inputs[141]));
    assign layer0_outputs[4621] = (inputs[90]) & ~(inputs[204]);
    assign layer0_outputs[4622] = inputs[92];
    assign layer0_outputs[4623] = 1'b0;
    assign layer0_outputs[4624] = ~((inputs[11]) | (inputs[67]));
    assign layer0_outputs[4625] = ~(inputs[78]);
    assign layer0_outputs[4626] = inputs[212];
    assign layer0_outputs[4627] = ~(inputs[107]);
    assign layer0_outputs[4628] = ~((inputs[53]) | (inputs[67]));
    assign layer0_outputs[4629] = (inputs[159]) | (inputs[127]);
    assign layer0_outputs[4630] = (inputs[12]) ^ (inputs[15]);
    assign layer0_outputs[4631] = ~((inputs[41]) | (inputs[157]));
    assign layer0_outputs[4632] = (inputs[4]) & ~(inputs[193]);
    assign layer0_outputs[4633] = ~(inputs[213]);
    assign layer0_outputs[4634] = (inputs[132]) & ~(inputs[55]);
    assign layer0_outputs[4635] = (inputs[185]) | (inputs[23]);
    assign layer0_outputs[4636] = (inputs[52]) & ~(inputs[33]);
    assign layer0_outputs[4637] = inputs[133];
    assign layer0_outputs[4638] = (inputs[136]) | (inputs[79]);
    assign layer0_outputs[4639] = ~(inputs[80]) | (inputs[206]);
    assign layer0_outputs[4640] = ~(inputs[216]);
    assign layer0_outputs[4641] = (inputs[54]) & ~(inputs[254]);
    assign layer0_outputs[4642] = (inputs[49]) | (inputs[170]);
    assign layer0_outputs[4643] = ~(inputs[238]);
    assign layer0_outputs[4644] = inputs[116];
    assign layer0_outputs[4645] = inputs[116];
    assign layer0_outputs[4646] = ~(inputs[107]) | (inputs[175]);
    assign layer0_outputs[4647] = ~(inputs[51]);
    assign layer0_outputs[4648] = (inputs[194]) | (inputs[177]);
    assign layer0_outputs[4649] = ~(inputs[25]);
    assign layer0_outputs[4650] = (inputs[150]) & ~(inputs[188]);
    assign layer0_outputs[4651] = (inputs[91]) & ~(inputs[226]);
    assign layer0_outputs[4652] = ~((inputs[88]) | (inputs[162]));
    assign layer0_outputs[4653] = ~(inputs[164]) | (inputs[18]);
    assign layer0_outputs[4654] = inputs[57];
    assign layer0_outputs[4655] = inputs[4];
    assign layer0_outputs[4656] = (inputs[179]) & ~(inputs[93]);
    assign layer0_outputs[4657] = inputs[117];
    assign layer0_outputs[4658] = ~(inputs[125]);
    assign layer0_outputs[4659] = ~(inputs[77]) | (inputs[253]);
    assign layer0_outputs[4660] = (inputs[225]) & (inputs[83]);
    assign layer0_outputs[4661] = ~(inputs[245]);
    assign layer0_outputs[4662] = ~(inputs[244]) | (inputs[224]);
    assign layer0_outputs[4663] = inputs[39];
    assign layer0_outputs[4664] = (inputs[67]) ^ (inputs[243]);
    assign layer0_outputs[4665] = inputs[117];
    assign layer0_outputs[4666] = (inputs[107]) & ~(inputs[136]);
    assign layer0_outputs[4667] = (inputs[246]) & ~(inputs[246]);
    assign layer0_outputs[4668] = (inputs[109]) ^ (inputs[172]);
    assign layer0_outputs[4669] = ~(inputs[189]);
    assign layer0_outputs[4670] = ~(inputs[165]) | (inputs[25]);
    assign layer0_outputs[4671] = ~(inputs[162]) | (inputs[159]);
    assign layer0_outputs[4672] = ~(inputs[169]) | (inputs[215]);
    assign layer0_outputs[4673] = (inputs[243]) & ~(inputs[220]);
    assign layer0_outputs[4674] = inputs[207];
    assign layer0_outputs[4675] = (inputs[244]) & ~(inputs[176]);
    assign layer0_outputs[4676] = (inputs[31]) | (inputs[66]);
    assign layer0_outputs[4677] = ~(inputs[57]) | (inputs[88]);
    assign layer0_outputs[4678] = 1'b0;
    assign layer0_outputs[4679] = (inputs[66]) | (inputs[37]);
    assign layer0_outputs[4680] = (inputs[105]) & ~(inputs[162]);
    assign layer0_outputs[4681] = (inputs[187]) | (inputs[80]);
    assign layer0_outputs[4682] = ~((inputs[1]) | (inputs[226]));
    assign layer0_outputs[4683] = ~(inputs[146]);
    assign layer0_outputs[4684] = 1'b0;
    assign layer0_outputs[4685] = ~((inputs[225]) ^ (inputs[68]));
    assign layer0_outputs[4686] = (inputs[67]) & ~(inputs[19]);
    assign layer0_outputs[4687] = ~((inputs[203]) & (inputs[108]));
    assign layer0_outputs[4688] = ~((inputs[211]) | (inputs[228]));
    assign layer0_outputs[4689] = 1'b1;
    assign layer0_outputs[4690] = inputs[219];
    assign layer0_outputs[4691] = ~((inputs[65]) & (inputs[78]));
    assign layer0_outputs[4692] = ~(inputs[186]);
    assign layer0_outputs[4693] = (inputs[72]) ^ (inputs[40]);
    assign layer0_outputs[4694] = (inputs[118]) & ~(inputs[236]);
    assign layer0_outputs[4695] = (inputs[105]) | (inputs[177]);
    assign layer0_outputs[4696] = inputs[55];
    assign layer0_outputs[4697] = inputs[89];
    assign layer0_outputs[4698] = ~(inputs[121]);
    assign layer0_outputs[4699] = inputs[99];
    assign layer0_outputs[4700] = ~((inputs[136]) | (inputs[204]));
    assign layer0_outputs[4701] = (inputs[251]) | (inputs[156]);
    assign layer0_outputs[4702] = (inputs[70]) ^ (inputs[49]);
    assign layer0_outputs[4703] = ~((inputs[162]) | (inputs[217]));
    assign layer0_outputs[4704] = inputs[227];
    assign layer0_outputs[4705] = ~(inputs[36]) | (inputs[18]);
    assign layer0_outputs[4706] = inputs[211];
    assign layer0_outputs[4707] = (inputs[236]) & ~(inputs[107]);
    assign layer0_outputs[4708] = ~(inputs[63]) | (inputs[161]);
    assign layer0_outputs[4709] = ~(inputs[45]) | (inputs[225]);
    assign layer0_outputs[4710] = ~((inputs[98]) ^ (inputs[211]));
    assign layer0_outputs[4711] = ~(inputs[7]) | (inputs[17]);
    assign layer0_outputs[4712] = inputs[138];
    assign layer0_outputs[4713] = ~((inputs[54]) | (inputs[221]));
    assign layer0_outputs[4714] = ~((inputs[198]) | (inputs[206]));
    assign layer0_outputs[4715] = (inputs[168]) & ~(inputs[85]);
    assign layer0_outputs[4716] = inputs[231];
    assign layer0_outputs[4717] = ~(inputs[152]) | (inputs[156]);
    assign layer0_outputs[4718] = ~((inputs[86]) & (inputs[83]));
    assign layer0_outputs[4719] = (inputs[180]) | (inputs[11]);
    assign layer0_outputs[4720] = (inputs[213]) | (inputs[38]);
    assign layer0_outputs[4721] = (inputs[235]) & ~(inputs[66]);
    assign layer0_outputs[4722] = (inputs[107]) | (inputs[236]);
    assign layer0_outputs[4723] = inputs[147];
    assign layer0_outputs[4724] = inputs[220];
    assign layer0_outputs[4725] = (inputs[63]) & (inputs[29]);
    assign layer0_outputs[4726] = (inputs[197]) ^ (inputs[11]);
    assign layer0_outputs[4727] = inputs[102];
    assign layer0_outputs[4728] = (inputs[234]) & ~(inputs[30]);
    assign layer0_outputs[4729] = inputs[139];
    assign layer0_outputs[4730] = inputs[225];
    assign layer0_outputs[4731] = (inputs[48]) ^ (inputs[60]);
    assign layer0_outputs[4732] = (inputs[117]) & ~(inputs[40]);
    assign layer0_outputs[4733] = (inputs[89]) | (inputs[40]);
    assign layer0_outputs[4734] = ~((inputs[101]) | (inputs[5]));
    assign layer0_outputs[4735] = ~((inputs[165]) ^ (inputs[192]));
    assign layer0_outputs[4736] = ~(inputs[147]);
    assign layer0_outputs[4737] = ~(inputs[228]);
    assign layer0_outputs[4738] = ~(inputs[34]);
    assign layer0_outputs[4739] = (inputs[44]) | (inputs[41]);
    assign layer0_outputs[4740] = ~((inputs[115]) | (inputs[42]));
    assign layer0_outputs[4741] = (inputs[111]) & (inputs[51]);
    assign layer0_outputs[4742] = ~(inputs[186]) | (inputs[204]);
    assign layer0_outputs[4743] = inputs[122];
    assign layer0_outputs[4744] = ~((inputs[139]) ^ (inputs[140]));
    assign layer0_outputs[4745] = ~(inputs[134]);
    assign layer0_outputs[4746] = (inputs[215]) & ~(inputs[127]);
    assign layer0_outputs[4747] = ~(inputs[197]);
    assign layer0_outputs[4748] = ~((inputs[93]) ^ (inputs[90]));
    assign layer0_outputs[4749] = inputs[25];
    assign layer0_outputs[4750] = ~(inputs[148]) | (inputs[193]);
    assign layer0_outputs[4751] = inputs[104];
    assign layer0_outputs[4752] = ~((inputs[179]) | (inputs[174]));
    assign layer0_outputs[4753] = ~(inputs[107]) | (inputs[227]);
    assign layer0_outputs[4754] = ~((inputs[43]) | (inputs[228]));
    assign layer0_outputs[4755] = inputs[199];
    assign layer0_outputs[4756] = ~(inputs[166]) | (inputs[11]);
    assign layer0_outputs[4757] = ~((inputs[164]) ^ (inputs[191]));
    assign layer0_outputs[4758] = ~((inputs[18]) ^ (inputs[183]));
    assign layer0_outputs[4759] = (inputs[46]) & ~(inputs[209]);
    assign layer0_outputs[4760] = (inputs[173]) & ~(inputs[29]);
    assign layer0_outputs[4761] = ~(inputs[242]);
    assign layer0_outputs[4762] = ~(inputs[29]) | (inputs[91]);
    assign layer0_outputs[4763] = (inputs[44]) ^ (inputs[135]);
    assign layer0_outputs[4764] = (inputs[219]) & ~(inputs[238]);
    assign layer0_outputs[4765] = (inputs[138]) | (inputs[179]);
    assign layer0_outputs[4766] = (inputs[121]) ^ (inputs[24]);
    assign layer0_outputs[4767] = inputs[222];
    assign layer0_outputs[4768] = ~((inputs[68]) | (inputs[193]));
    assign layer0_outputs[4769] = (inputs[105]) | (inputs[45]);
    assign layer0_outputs[4770] = (inputs[133]) | (inputs[204]);
    assign layer0_outputs[4771] = inputs[217];
    assign layer0_outputs[4772] = inputs[242];
    assign layer0_outputs[4773] = ~(inputs[170]);
    assign layer0_outputs[4774] = ~(inputs[86]) | (inputs[50]);
    assign layer0_outputs[4775] = ~(inputs[217]) | (inputs[222]);
    assign layer0_outputs[4776] = ~(inputs[208]);
    assign layer0_outputs[4777] = ~((inputs[61]) | (inputs[160]));
    assign layer0_outputs[4778] = inputs[147];
    assign layer0_outputs[4779] = ~(inputs[185]) | (inputs[145]);
    assign layer0_outputs[4780] = 1'b1;
    assign layer0_outputs[4781] = (inputs[144]) ^ (inputs[211]);
    assign layer0_outputs[4782] = ~((inputs[21]) & (inputs[236]));
    assign layer0_outputs[4783] = ~((inputs[185]) & (inputs[252]));
    assign layer0_outputs[4784] = 1'b0;
    assign layer0_outputs[4785] = ~(inputs[40]);
    assign layer0_outputs[4786] = inputs[198];
    assign layer0_outputs[4787] = ~(inputs[226]) | (inputs[178]);
    assign layer0_outputs[4788] = ~((inputs[235]) | (inputs[36]));
    assign layer0_outputs[4789] = inputs[73];
    assign layer0_outputs[4790] = 1'b1;
    assign layer0_outputs[4791] = (inputs[225]) | (inputs[91]);
    assign layer0_outputs[4792] = inputs[213];
    assign layer0_outputs[4793] = ~(inputs[49]) | (inputs[254]);
    assign layer0_outputs[4794] = (inputs[27]) & ~(inputs[189]);
    assign layer0_outputs[4795] = inputs[37];
    assign layer0_outputs[4796] = ~(inputs[214]) | (inputs[174]);
    assign layer0_outputs[4797] = (inputs[41]) | (inputs[165]);
    assign layer0_outputs[4798] = inputs[69];
    assign layer0_outputs[4799] = (inputs[68]) & ~(inputs[12]);
    assign layer0_outputs[4800] = inputs[22];
    assign layer0_outputs[4801] = ~((inputs[137]) ^ (inputs[20]));
    assign layer0_outputs[4802] = ~((inputs[42]) | (inputs[62]));
    assign layer0_outputs[4803] = ~((inputs[183]) | (inputs[171]));
    assign layer0_outputs[4804] = inputs[196];
    assign layer0_outputs[4805] = (inputs[85]) & ~(inputs[12]);
    assign layer0_outputs[4806] = inputs[155];
    assign layer0_outputs[4807] = (inputs[5]) ^ (inputs[15]);
    assign layer0_outputs[4808] = (inputs[120]) & ~(inputs[97]);
    assign layer0_outputs[4809] = inputs[164];
    assign layer0_outputs[4810] = inputs[89];
    assign layer0_outputs[4811] = ~((inputs[30]) | (inputs[86]));
    assign layer0_outputs[4812] = ~(inputs[84]);
    assign layer0_outputs[4813] = ~(inputs[252]);
    assign layer0_outputs[4814] = inputs[41];
    assign layer0_outputs[4815] = ~(inputs[85]) | (inputs[223]);
    assign layer0_outputs[4816] = (inputs[176]) ^ (inputs[151]);
    assign layer0_outputs[4817] = inputs[200];
    assign layer0_outputs[4818] = (inputs[68]) ^ (inputs[140]);
    assign layer0_outputs[4819] = (inputs[108]) & ~(inputs[61]);
    assign layer0_outputs[4820] = (inputs[187]) ^ (inputs[91]);
    assign layer0_outputs[4821] = ~(inputs[16]) | (inputs[241]);
    assign layer0_outputs[4822] = (inputs[168]) & ~(inputs[81]);
    assign layer0_outputs[4823] = ~((inputs[31]) | (inputs[146]));
    assign layer0_outputs[4824] = (inputs[213]) | (inputs[215]);
    assign layer0_outputs[4825] = ~(inputs[119]);
    assign layer0_outputs[4826] = (inputs[224]) ^ (inputs[186]);
    assign layer0_outputs[4827] = (inputs[164]) ^ (inputs[71]);
    assign layer0_outputs[4828] = (inputs[167]) & ~(inputs[192]);
    assign layer0_outputs[4829] = (inputs[199]) & ~(inputs[250]);
    assign layer0_outputs[4830] = (inputs[96]) | (inputs[200]);
    assign layer0_outputs[4831] = (inputs[121]) & ~(inputs[220]);
    assign layer0_outputs[4832] = ~(inputs[109]) | (inputs[62]);
    assign layer0_outputs[4833] = (inputs[3]) | (inputs[103]);
    assign layer0_outputs[4834] = (inputs[64]) ^ (inputs[233]);
    assign layer0_outputs[4835] = (inputs[39]) | (inputs[95]);
    assign layer0_outputs[4836] = ~((inputs[46]) ^ (inputs[200]));
    assign layer0_outputs[4837] = (inputs[111]) ^ (inputs[86]);
    assign layer0_outputs[4838] = (inputs[254]) ^ (inputs[75]);
    assign layer0_outputs[4839] = ~((inputs[104]) | (inputs[246]));
    assign layer0_outputs[4840] = (inputs[155]) | (inputs[252]);
    assign layer0_outputs[4841] = ~((inputs[182]) | (inputs[188]));
    assign layer0_outputs[4842] = ~(inputs[55]) | (inputs[102]);
    assign layer0_outputs[4843] = ~((inputs[147]) ^ (inputs[249]));
    assign layer0_outputs[4844] = ~((inputs[6]) ^ (inputs[8]));
    assign layer0_outputs[4845] = (inputs[203]) & ~(inputs[234]);
    assign layer0_outputs[4846] = ~((inputs[54]) | (inputs[31]));
    assign layer0_outputs[4847] = ~((inputs[61]) ^ (inputs[28]));
    assign layer0_outputs[4848] = ~(inputs[255]);
    assign layer0_outputs[4849] = ~(inputs[59]) | (inputs[96]);
    assign layer0_outputs[4850] = ~((inputs[115]) | (inputs[221]));
    assign layer0_outputs[4851] = 1'b1;
    assign layer0_outputs[4852] = ~((inputs[65]) | (inputs[93]));
    assign layer0_outputs[4853] = (inputs[17]) ^ (inputs[18]);
    assign layer0_outputs[4854] = ~(inputs[77]) | (inputs[15]);
    assign layer0_outputs[4855] = ~((inputs[230]) ^ (inputs[173]));
    assign layer0_outputs[4856] = (inputs[185]) ^ (inputs[18]);
    assign layer0_outputs[4857] = inputs[24];
    assign layer0_outputs[4858] = (inputs[100]) | (inputs[4]);
    assign layer0_outputs[4859] = inputs[220];
    assign layer0_outputs[4860] = ~(inputs[237]) | (inputs[76]);
    assign layer0_outputs[4861] = (inputs[195]) & ~(inputs[223]);
    assign layer0_outputs[4862] = inputs[226];
    assign layer0_outputs[4863] = inputs[91];
    assign layer0_outputs[4864] = (inputs[137]) | (inputs[113]);
    assign layer0_outputs[4865] = ~((inputs[123]) ^ (inputs[95]));
    assign layer0_outputs[4866] = ~(inputs[188]);
    assign layer0_outputs[4867] = ~(inputs[166]) | (inputs[195]);
    assign layer0_outputs[4868] = 1'b0;
    assign layer0_outputs[4869] = ~(inputs[151]);
    assign layer0_outputs[4870] = (inputs[16]) & ~(inputs[18]);
    assign layer0_outputs[4871] = inputs[144];
    assign layer0_outputs[4872] = (inputs[136]) & ~(inputs[124]);
    assign layer0_outputs[4873] = (inputs[39]) & ~(inputs[252]);
    assign layer0_outputs[4874] = ~((inputs[2]) | (inputs[14]));
    assign layer0_outputs[4875] = 1'b1;
    assign layer0_outputs[4876] = (inputs[71]) & ~(inputs[235]);
    assign layer0_outputs[4877] = (inputs[108]) & ~(inputs[146]);
    assign layer0_outputs[4878] = ~((inputs[55]) | (inputs[172]));
    assign layer0_outputs[4879] = (inputs[166]) & ~(inputs[195]);
    assign layer0_outputs[4880] = (inputs[120]) & ~(inputs[70]);
    assign layer0_outputs[4881] = (inputs[159]) & ~(inputs[248]);
    assign layer0_outputs[4882] = (inputs[153]) | (inputs[207]);
    assign layer0_outputs[4883] = (inputs[138]) & ~(inputs[171]);
    assign layer0_outputs[4884] = (inputs[169]) | (inputs[145]);
    assign layer0_outputs[4885] = ~(inputs[174]);
    assign layer0_outputs[4886] = (inputs[252]) ^ (inputs[214]);
    assign layer0_outputs[4887] = ~(inputs[133]);
    assign layer0_outputs[4888] = (inputs[142]) & ~(inputs[237]);
    assign layer0_outputs[4889] = (inputs[45]) & ~(inputs[6]);
    assign layer0_outputs[4890] = (inputs[40]) | (inputs[150]);
    assign layer0_outputs[4891] = ~(inputs[115]);
    assign layer0_outputs[4892] = inputs[140];
    assign layer0_outputs[4893] = (inputs[1]) & (inputs[1]);
    assign layer0_outputs[4894] = (inputs[136]) | (inputs[145]);
    assign layer0_outputs[4895] = (inputs[93]) | (inputs[244]);
    assign layer0_outputs[4896] = ~(inputs[179]);
    assign layer0_outputs[4897] = ~((inputs[129]) & (inputs[210]));
    assign layer0_outputs[4898] = (inputs[204]) ^ (inputs[158]);
    assign layer0_outputs[4899] = (inputs[108]) | (inputs[83]);
    assign layer0_outputs[4900] = ~((inputs[73]) ^ (inputs[251]));
    assign layer0_outputs[4901] = inputs[35];
    assign layer0_outputs[4902] = ~(inputs[108]) | (inputs[112]);
    assign layer0_outputs[4903] = ~(inputs[88]) | (inputs[92]);
    assign layer0_outputs[4904] = ~((inputs[61]) | (inputs[120]));
    assign layer0_outputs[4905] = ~(inputs[157]);
    assign layer0_outputs[4906] = inputs[211];
    assign layer0_outputs[4907] = ~((inputs[130]) ^ (inputs[132]));
    assign layer0_outputs[4908] = inputs[83];
    assign layer0_outputs[4909] = (inputs[151]) & ~(inputs[45]);
    assign layer0_outputs[4910] = inputs[196];
    assign layer0_outputs[4911] = inputs[105];
    assign layer0_outputs[4912] = ~(inputs[239]);
    assign layer0_outputs[4913] = ~((inputs[104]) | (inputs[177]));
    assign layer0_outputs[4914] = 1'b0;
    assign layer0_outputs[4915] = ~(inputs[215]);
    assign layer0_outputs[4916] = ~((inputs[232]) | (inputs[131]));
    assign layer0_outputs[4917] = ~(inputs[134]) | (inputs[70]);
    assign layer0_outputs[4918] = ~(inputs[198]);
    assign layer0_outputs[4919] = (inputs[101]) | (inputs[176]);
    assign layer0_outputs[4920] = (inputs[191]) & (inputs[236]);
    assign layer0_outputs[4921] = (inputs[186]) & ~(inputs[46]);
    assign layer0_outputs[4922] = inputs[163];
    assign layer0_outputs[4923] = ~((inputs[201]) & (inputs[133]));
    assign layer0_outputs[4924] = (inputs[18]) & (inputs[49]);
    assign layer0_outputs[4925] = ~((inputs[204]) | (inputs[164]));
    assign layer0_outputs[4926] = ~(inputs[172]) | (inputs[189]);
    assign layer0_outputs[4927] = ~(inputs[121]) | (inputs[157]);
    assign layer0_outputs[4928] = ~((inputs[243]) & (inputs[37]));
    assign layer0_outputs[4929] = ~(inputs[219]);
    assign layer0_outputs[4930] = ~(inputs[125]) | (inputs[63]);
    assign layer0_outputs[4931] = ~((inputs[64]) | (inputs[240]));
    assign layer0_outputs[4932] = (inputs[70]) & ~(inputs[64]);
    assign layer0_outputs[4933] = ~(inputs[165]) | (inputs[146]);
    assign layer0_outputs[4934] = ~((inputs[237]) ^ (inputs[229]));
    assign layer0_outputs[4935] = inputs[185];
    assign layer0_outputs[4936] = 1'b0;
    assign layer0_outputs[4937] = (inputs[16]) & ~(inputs[241]);
    assign layer0_outputs[4938] = (inputs[210]) ^ (inputs[217]);
    assign layer0_outputs[4939] = (inputs[79]) | (inputs[153]);
    assign layer0_outputs[4940] = ~(inputs[216]);
    assign layer0_outputs[4941] = inputs[40];
    assign layer0_outputs[4942] = ~(inputs[98]);
    assign layer0_outputs[4943] = ~((inputs[109]) ^ (inputs[225]));
    assign layer0_outputs[4944] = (inputs[51]) | (inputs[96]);
    assign layer0_outputs[4945] = ~((inputs[143]) ^ (inputs[191]));
    assign layer0_outputs[4946] = ~(inputs[16]) | (inputs[190]);
    assign layer0_outputs[4947] = ~(inputs[53]);
    assign layer0_outputs[4948] = ~(inputs[171]) | (inputs[30]);
    assign layer0_outputs[4949] = ~(inputs[26]);
    assign layer0_outputs[4950] = ~(inputs[0]);
    assign layer0_outputs[4951] = 1'b0;
    assign layer0_outputs[4952] = ~(inputs[136]) | (inputs[230]);
    assign layer0_outputs[4953] = ~(inputs[42]);
    assign layer0_outputs[4954] = inputs[49];
    assign layer0_outputs[4955] = (inputs[158]) | (inputs[9]);
    assign layer0_outputs[4956] = ~((inputs[129]) & (inputs[185]));
    assign layer0_outputs[4957] = inputs[178];
    assign layer0_outputs[4958] = ~(inputs[40]) | (inputs[160]);
    assign layer0_outputs[4959] = ~((inputs[167]) | (inputs[58]));
    assign layer0_outputs[4960] = ~(inputs[186]);
    assign layer0_outputs[4961] = ~(inputs[118]) | (inputs[230]);
    assign layer0_outputs[4962] = (inputs[66]) & ~(inputs[14]);
    assign layer0_outputs[4963] = ~(inputs[41]);
    assign layer0_outputs[4964] = ~((inputs[23]) | (inputs[103]));
    assign layer0_outputs[4965] = inputs[164];
    assign layer0_outputs[4966] = ~(inputs[69]) | (inputs[24]);
    assign layer0_outputs[4967] = (inputs[69]) & ~(inputs[116]);
    assign layer0_outputs[4968] = ~((inputs[78]) ^ (inputs[46]));
    assign layer0_outputs[4969] = inputs[163];
    assign layer0_outputs[4970] = inputs[138];
    assign layer0_outputs[4971] = ~(inputs[54]);
    assign layer0_outputs[4972] = ~(inputs[242]);
    assign layer0_outputs[4973] = ~(inputs[84]) | (inputs[205]);
    assign layer0_outputs[4974] = ~((inputs[252]) | (inputs[8]));
    assign layer0_outputs[4975] = ~((inputs[112]) ^ (inputs[145]));
    assign layer0_outputs[4976] = (inputs[54]) & ~(inputs[6]);
    assign layer0_outputs[4977] = ~(inputs[133]) | (inputs[62]);
    assign layer0_outputs[4978] = ~(inputs[156]);
    assign layer0_outputs[4979] = ~(inputs[197]);
    assign layer0_outputs[4980] = ~(inputs[10]);
    assign layer0_outputs[4981] = (inputs[93]) ^ (inputs[221]);
    assign layer0_outputs[4982] = inputs[18];
    assign layer0_outputs[4983] = inputs[166];
    assign layer0_outputs[4984] = ~(inputs[184]);
    assign layer0_outputs[4985] = ~(inputs[141]) | (inputs[65]);
    assign layer0_outputs[4986] = (inputs[11]) | (inputs[231]);
    assign layer0_outputs[4987] = (inputs[35]) ^ (inputs[169]);
    assign layer0_outputs[4988] = 1'b0;
    assign layer0_outputs[4989] = ~((inputs[246]) ^ (inputs[131]));
    assign layer0_outputs[4990] = ~((inputs[26]) | (inputs[191]));
    assign layer0_outputs[4991] = ~((inputs[109]) | (inputs[61]));
    assign layer0_outputs[4992] = ~(inputs[105]);
    assign layer0_outputs[4993] = (inputs[182]) & ~(inputs[44]);
    assign layer0_outputs[4994] = (inputs[178]) ^ (inputs[248]);
    assign layer0_outputs[4995] = ~(inputs[207]);
    assign layer0_outputs[4996] = (inputs[140]) ^ (inputs[20]);
    assign layer0_outputs[4997] = ~((inputs[61]) ^ (inputs[80]));
    assign layer0_outputs[4998] = ~(inputs[60]) | (inputs[28]);
    assign layer0_outputs[4999] = (inputs[70]) & ~(inputs[22]);
    assign layer0_outputs[5000] = ~(inputs[125]);
    assign layer0_outputs[5001] = (inputs[22]) & ~(inputs[146]);
    assign layer0_outputs[5002] = inputs[202];
    assign layer0_outputs[5003] = (inputs[27]) | (inputs[185]);
    assign layer0_outputs[5004] = (inputs[170]) & ~(inputs[175]);
    assign layer0_outputs[5005] = ~(inputs[209]);
    assign layer0_outputs[5006] = (inputs[191]) & ~(inputs[144]);
    assign layer0_outputs[5007] = inputs[131];
    assign layer0_outputs[5008] = ~((inputs[135]) & (inputs[57]));
    assign layer0_outputs[5009] = (inputs[84]) & ~(inputs[54]);
    assign layer0_outputs[5010] = ~((inputs[28]) ^ (inputs[12]));
    assign layer0_outputs[5011] = inputs[69];
    assign layer0_outputs[5012] = (inputs[98]) | (inputs[183]);
    assign layer0_outputs[5013] = (inputs[220]) ^ (inputs[251]);
    assign layer0_outputs[5014] = (inputs[157]) | (inputs[255]);
    assign layer0_outputs[5015] = ~((inputs[78]) ^ (inputs[49]));
    assign layer0_outputs[5016] = (inputs[50]) & (inputs[241]);
    assign layer0_outputs[5017] = ~(inputs[173]) | (inputs[21]);
    assign layer0_outputs[5018] = ~((inputs[107]) ^ (inputs[115]));
    assign layer0_outputs[5019] = (inputs[225]) & ~(inputs[148]);
    assign layer0_outputs[5020] = ~(inputs[120]) | (inputs[17]);
    assign layer0_outputs[5021] = 1'b0;
    assign layer0_outputs[5022] = (inputs[127]) | (inputs[181]);
    assign layer0_outputs[5023] = ~((inputs[174]) | (inputs[20]));
    assign layer0_outputs[5024] = (inputs[77]) & ~(inputs[69]);
    assign layer0_outputs[5025] = 1'b1;
    assign layer0_outputs[5026] = 1'b0;
    assign layer0_outputs[5027] = (inputs[83]) ^ (inputs[179]);
    assign layer0_outputs[5028] = 1'b0;
    assign layer0_outputs[5029] = ~(inputs[114]) | (inputs[70]);
    assign layer0_outputs[5030] = ~(inputs[55]);
    assign layer0_outputs[5031] = ~(inputs[164]);
    assign layer0_outputs[5032] = (inputs[44]) | (inputs[196]);
    assign layer0_outputs[5033] = inputs[197];
    assign layer0_outputs[5034] = ~((inputs[245]) ^ (inputs[155]));
    assign layer0_outputs[5035] = 1'b0;
    assign layer0_outputs[5036] = (inputs[154]) | (inputs[15]);
    assign layer0_outputs[5037] = inputs[167];
    assign layer0_outputs[5038] = ~((inputs[124]) | (inputs[89]));
    assign layer0_outputs[5039] = (inputs[61]) ^ (inputs[150]);
    assign layer0_outputs[5040] = ~((inputs[169]) | (inputs[16]));
    assign layer0_outputs[5041] = ~(inputs[25]);
    assign layer0_outputs[5042] = ~(inputs[90]) | (inputs[141]);
    assign layer0_outputs[5043] = ~((inputs[0]) ^ (inputs[111]));
    assign layer0_outputs[5044] = ~(inputs[244]);
    assign layer0_outputs[5045] = ~(inputs[55]) | (inputs[64]);
    assign layer0_outputs[5046] = ~(inputs[166]);
    assign layer0_outputs[5047] = inputs[117];
    assign layer0_outputs[5048] = ~(inputs[89]);
    assign layer0_outputs[5049] = (inputs[93]) ^ (inputs[17]);
    assign layer0_outputs[5050] = (inputs[112]) | (inputs[60]);
    assign layer0_outputs[5051] = (inputs[56]) | (inputs[247]);
    assign layer0_outputs[5052] = 1'b1;
    assign layer0_outputs[5053] = ~(inputs[134]) | (inputs[220]);
    assign layer0_outputs[5054] = inputs[39];
    assign layer0_outputs[5055] = ~(inputs[10]) | (inputs[60]);
    assign layer0_outputs[5056] = ~(inputs[22]) | (inputs[80]);
    assign layer0_outputs[5057] = ~((inputs[208]) | (inputs[97]));
    assign layer0_outputs[5058] = (inputs[89]) & ~(inputs[171]);
    assign layer0_outputs[5059] = ~(inputs[227]) | (inputs[192]);
    assign layer0_outputs[5060] = inputs[156];
    assign layer0_outputs[5061] = (inputs[161]) & ~(inputs[223]);
    assign layer0_outputs[5062] = 1'b1;
    assign layer0_outputs[5063] = ~((inputs[10]) ^ (inputs[149]));
    assign layer0_outputs[5064] = ~(inputs[157]) | (inputs[2]);
    assign layer0_outputs[5065] = ~(inputs[231]) | (inputs[190]);
    assign layer0_outputs[5066] = ~((inputs[223]) ^ (inputs[41]));
    assign layer0_outputs[5067] = (inputs[97]) ^ (inputs[188]);
    assign layer0_outputs[5068] = 1'b0;
    assign layer0_outputs[5069] = ~(inputs[187]) | (inputs[82]);
    assign layer0_outputs[5070] = (inputs[136]) & (inputs[136]);
    assign layer0_outputs[5071] = inputs[43];
    assign layer0_outputs[5072] = (inputs[110]) & ~(inputs[243]);
    assign layer0_outputs[5073] = ~(inputs[176]);
    assign layer0_outputs[5074] = 1'b0;
    assign layer0_outputs[5075] = ~((inputs[172]) | (inputs[96]));
    assign layer0_outputs[5076] = (inputs[215]) | (inputs[40]);
    assign layer0_outputs[5077] = inputs[54];
    assign layer0_outputs[5078] = ~(inputs[22]);
    assign layer0_outputs[5079] = (inputs[1]) & ~(inputs[62]);
    assign layer0_outputs[5080] = ~((inputs[97]) | (inputs[187]));
    assign layer0_outputs[5081] = 1'b0;
    assign layer0_outputs[5082] = (inputs[137]) & ~(inputs[68]);
    assign layer0_outputs[5083] = (inputs[167]) & ~(inputs[224]);
    assign layer0_outputs[5084] = (inputs[224]) | (inputs[205]);
    assign layer0_outputs[5085] = ~((inputs[138]) | (inputs[146]));
    assign layer0_outputs[5086] = ~(inputs[23]);
    assign layer0_outputs[5087] = (inputs[112]) ^ (inputs[105]);
    assign layer0_outputs[5088] = (inputs[124]) & ~(inputs[234]);
    assign layer0_outputs[5089] = ~(inputs[170]);
    assign layer0_outputs[5090] = ~((inputs[90]) ^ (inputs[189]));
    assign layer0_outputs[5091] = (inputs[177]) | (inputs[211]);
    assign layer0_outputs[5092] = inputs[22];
    assign layer0_outputs[5093] = ~((inputs[195]) ^ (inputs[5]));
    assign layer0_outputs[5094] = ~(inputs[119]);
    assign layer0_outputs[5095] = (inputs[247]) ^ (inputs[224]);
    assign layer0_outputs[5096] = (inputs[2]) | (inputs[76]);
    assign layer0_outputs[5097] = ~((inputs[161]) ^ (inputs[57]));
    assign layer0_outputs[5098] = (inputs[40]) | (inputs[163]);
    assign layer0_outputs[5099] = inputs[165];
    assign layer0_outputs[5100] = inputs[181];
    assign layer0_outputs[5101] = ~(inputs[5]) | (inputs[147]);
    assign layer0_outputs[5102] = ~(inputs[193]) | (inputs[238]);
    assign layer0_outputs[5103] = (inputs[254]) | (inputs[90]);
    assign layer0_outputs[5104] = ~(inputs[200]) | (inputs[11]);
    assign layer0_outputs[5105] = ~((inputs[235]) | (inputs[237]));
    assign layer0_outputs[5106] = ~((inputs[156]) | (inputs[139]));
    assign layer0_outputs[5107] = ~(inputs[140]);
    assign layer0_outputs[5108] = inputs[55];
    assign layer0_outputs[5109] = ~((inputs[101]) ^ (inputs[114]));
    assign layer0_outputs[5110] = ~(inputs[32]);
    assign layer0_outputs[5111] = inputs[164];
    assign layer0_outputs[5112] = (inputs[122]) ^ (inputs[142]);
    assign layer0_outputs[5113] = ~(inputs[150]);
    assign layer0_outputs[5114] = (inputs[171]) & ~(inputs[114]);
    assign layer0_outputs[5115] = (inputs[131]) & ~(inputs[247]);
    assign layer0_outputs[5116] = (inputs[22]) ^ (inputs[143]);
    assign layer0_outputs[5117] = ~(inputs[174]);
    assign layer0_outputs[5118] = ~(inputs[139]) | (inputs[32]);
    assign layer0_outputs[5119] = (inputs[3]) & ~(inputs[144]);
    assign outputs[0] = (layer0_outputs[4090]) ^ (layer0_outputs[4751]);
    assign outputs[1] = (layer0_outputs[2188]) ^ (layer0_outputs[3085]);
    assign outputs[2] = ~(layer0_outputs[1224]);
    assign outputs[3] = (layer0_outputs[3792]) ^ (layer0_outputs[4442]);
    assign outputs[4] = (layer0_outputs[801]) ^ (layer0_outputs[1110]);
    assign outputs[5] = (layer0_outputs[2215]) & (layer0_outputs[5059]);
    assign outputs[6] = layer0_outputs[2519];
    assign outputs[7] = (layer0_outputs[2540]) ^ (layer0_outputs[4021]);
    assign outputs[8] = ~(layer0_outputs[4223]);
    assign outputs[9] = (layer0_outputs[1615]) ^ (layer0_outputs[3363]);
    assign outputs[10] = ~((layer0_outputs[3077]) | (layer0_outputs[1829]));
    assign outputs[11] = ~(layer0_outputs[2953]);
    assign outputs[12] = ~((layer0_outputs[4386]) ^ (layer0_outputs[2901]));
    assign outputs[13] = layer0_outputs[3311];
    assign outputs[14] = ~((layer0_outputs[4459]) | (layer0_outputs[3662]));
    assign outputs[15] = layer0_outputs[2241];
    assign outputs[16] = layer0_outputs[4526];
    assign outputs[17] = (layer0_outputs[4228]) & (layer0_outputs[3554]);
    assign outputs[18] = (layer0_outputs[3989]) ^ (layer0_outputs[4590]);
    assign outputs[19] = layer0_outputs[2187];
    assign outputs[20] = ~((layer0_outputs[3928]) & (layer0_outputs[4995]));
    assign outputs[21] = layer0_outputs[4146];
    assign outputs[22] = ~(layer0_outputs[4832]);
    assign outputs[23] = ~((layer0_outputs[5079]) ^ (layer0_outputs[5018]));
    assign outputs[24] = ~(layer0_outputs[206]) | (layer0_outputs[489]);
    assign outputs[25] = ~(layer0_outputs[1980]) | (layer0_outputs[712]);
    assign outputs[26] = ~(layer0_outputs[748]) | (layer0_outputs[526]);
    assign outputs[27] = (layer0_outputs[2853]) | (layer0_outputs[950]);
    assign outputs[28] = ~(layer0_outputs[1329]) | (layer0_outputs[927]);
    assign outputs[29] = ~((layer0_outputs[2739]) ^ (layer0_outputs[999]));
    assign outputs[30] = ~((layer0_outputs[1720]) ^ (layer0_outputs[2535]));
    assign outputs[31] = ~(layer0_outputs[3203]) | (layer0_outputs[886]);
    assign outputs[32] = ~((layer0_outputs[4155]) & (layer0_outputs[2271]));
    assign outputs[33] = (layer0_outputs[5019]) | (layer0_outputs[2744]);
    assign outputs[34] = (layer0_outputs[2404]) ^ (layer0_outputs[3532]);
    assign outputs[35] = ~(layer0_outputs[1162]);
    assign outputs[36] = ~((layer0_outputs[4648]) ^ (layer0_outputs[3109]));
    assign outputs[37] = (layer0_outputs[2218]) ^ (layer0_outputs[3727]);
    assign outputs[38] = ~(layer0_outputs[4322]);
    assign outputs[39] = ~(layer0_outputs[1197]);
    assign outputs[40] = (layer0_outputs[453]) ^ (layer0_outputs[3061]);
    assign outputs[41] = (layer0_outputs[1917]) & (layer0_outputs[4025]);
    assign outputs[42] = (layer0_outputs[4868]) | (layer0_outputs[4755]);
    assign outputs[43] = ~((layer0_outputs[1736]) | (layer0_outputs[3528]));
    assign outputs[44] = (layer0_outputs[1469]) ^ (layer0_outputs[3460]);
    assign outputs[45] = layer0_outputs[4997];
    assign outputs[46] = ~(layer0_outputs[1626]) | (layer0_outputs[364]);
    assign outputs[47] = layer0_outputs[67];
    assign outputs[48] = ~(layer0_outputs[3258]);
    assign outputs[49] = ~(layer0_outputs[1206]);
    assign outputs[50] = ~(layer0_outputs[4977]);
    assign outputs[51] = ~(layer0_outputs[5087]) | (layer0_outputs[407]);
    assign outputs[52] = ~((layer0_outputs[5093]) ^ (layer0_outputs[2858]));
    assign outputs[53] = ~(layer0_outputs[256]);
    assign outputs[54] = (layer0_outputs[1067]) & (layer0_outputs[4455]);
    assign outputs[55] = ~((layer0_outputs[3453]) & (layer0_outputs[4100]));
    assign outputs[56] = ~(layer0_outputs[1066]);
    assign outputs[57] = ~((layer0_outputs[3437]) ^ (layer0_outputs[103]));
    assign outputs[58] = layer0_outputs[531];
    assign outputs[59] = ~(layer0_outputs[1258]);
    assign outputs[60] = ~(layer0_outputs[3482]);
    assign outputs[61] = layer0_outputs[3610];
    assign outputs[62] = layer0_outputs[624];
    assign outputs[63] = ~(layer0_outputs[4522]);
    assign outputs[64] = ~((layer0_outputs[4670]) & (layer0_outputs[2348]));
    assign outputs[65] = layer0_outputs[176];
    assign outputs[66] = (layer0_outputs[3130]) ^ (layer0_outputs[2773]);
    assign outputs[67] = ~((layer0_outputs[2227]) ^ (layer0_outputs[3699]));
    assign outputs[68] = ~((layer0_outputs[3307]) | (layer0_outputs[2882]));
    assign outputs[69] = layer0_outputs[416];
    assign outputs[70] = (layer0_outputs[1712]) ^ (layer0_outputs[3924]);
    assign outputs[71] = layer0_outputs[1079];
    assign outputs[72] = ~(layer0_outputs[2940]) | (layer0_outputs[342]);
    assign outputs[73] = ~(layer0_outputs[2220]);
    assign outputs[74] = ~(layer0_outputs[798]);
    assign outputs[75] = layer0_outputs[3592];
    assign outputs[76] = (layer0_outputs[4818]) & ~(layer0_outputs[4636]);
    assign outputs[77] = layer0_outputs[3501];
    assign outputs[78] = ~(layer0_outputs[1896]) | (layer0_outputs[993]);
    assign outputs[79] = layer0_outputs[3830];
    assign outputs[80] = ~((layer0_outputs[3585]) ^ (layer0_outputs[1450]));
    assign outputs[81] = ~(layer0_outputs[820]);
    assign outputs[82] = (layer0_outputs[4135]) & ~(layer0_outputs[3430]);
    assign outputs[83] = 1'b1;
    assign outputs[84] = ~(layer0_outputs[386]);
    assign outputs[85] = layer0_outputs[4892];
    assign outputs[86] = ~(layer0_outputs[833]) | (layer0_outputs[726]);
    assign outputs[87] = layer0_outputs[4561];
    assign outputs[88] = ~((layer0_outputs[3123]) ^ (layer0_outputs[1187]));
    assign outputs[89] = ~((layer0_outputs[1805]) ^ (layer0_outputs[759]));
    assign outputs[90] = ~(layer0_outputs[2111]);
    assign outputs[91] = ~(layer0_outputs[3759]);
    assign outputs[92] = layer0_outputs[4563];
    assign outputs[93] = ~(layer0_outputs[5034]);
    assign outputs[94] = layer0_outputs[836];
    assign outputs[95] = (layer0_outputs[3310]) | (layer0_outputs[4042]);
    assign outputs[96] = ~(layer0_outputs[1303]) | (layer0_outputs[2084]);
    assign outputs[97] = ~(layer0_outputs[3249]);
    assign outputs[98] = ~((layer0_outputs[1161]) & (layer0_outputs[3910]));
    assign outputs[99] = ~((layer0_outputs[2367]) & (layer0_outputs[4736]));
    assign outputs[100] = ~(layer0_outputs[2889]) | (layer0_outputs[1253]);
    assign outputs[101] = ~((layer0_outputs[4092]) ^ (layer0_outputs[4472]));
    assign outputs[102] = layer0_outputs[1314];
    assign outputs[103] = ~(layer0_outputs[1138]);
    assign outputs[104] = ~((layer0_outputs[1610]) ^ (layer0_outputs[4232]));
    assign outputs[105] = ~(layer0_outputs[2547]) | (layer0_outputs[4018]);
    assign outputs[106] = ~(layer0_outputs[2719]);
    assign outputs[107] = ~(layer0_outputs[4793]) | (layer0_outputs[2144]);
    assign outputs[108] = ~(layer0_outputs[960]);
    assign outputs[109] = ~(layer0_outputs[1580]);
    assign outputs[110] = (layer0_outputs[957]) | (layer0_outputs[1834]);
    assign outputs[111] = ~(layer0_outputs[1538]) | (layer0_outputs[4172]);
    assign outputs[112] = ~((layer0_outputs[3920]) ^ (layer0_outputs[4713]));
    assign outputs[113] = ~((layer0_outputs[2825]) ^ (layer0_outputs[3126]));
    assign outputs[114] = ~((layer0_outputs[5109]) ^ (layer0_outputs[1536]));
    assign outputs[115] = ~(layer0_outputs[4898]);
    assign outputs[116] = ~(layer0_outputs[4392]);
    assign outputs[117] = layer0_outputs[3700];
    assign outputs[118] = 1'b1;
    assign outputs[119] = layer0_outputs[1137];
    assign outputs[120] = ~(layer0_outputs[3976]);
    assign outputs[121] = (layer0_outputs[3292]) ^ (layer0_outputs[4951]);
    assign outputs[122] = layer0_outputs[3667];
    assign outputs[123] = (layer0_outputs[2389]) & (layer0_outputs[4394]);
    assign outputs[124] = layer0_outputs[1961];
    assign outputs[125] = (layer0_outputs[2900]) | (layer0_outputs[3916]);
    assign outputs[126] = layer0_outputs[3178];
    assign outputs[127] = ~((layer0_outputs[312]) | (layer0_outputs[905]));
    assign outputs[128] = ~(layer0_outputs[4176]);
    assign outputs[129] = (layer0_outputs[766]) & ~(layer0_outputs[4799]);
    assign outputs[130] = ~((layer0_outputs[676]) ^ (layer0_outputs[511]));
    assign outputs[131] = ~(layer0_outputs[3483]) | (layer0_outputs[2640]);
    assign outputs[132] = layer0_outputs[4510];
    assign outputs[133] = layer0_outputs[2398];
    assign outputs[134] = ~(layer0_outputs[1642]) | (layer0_outputs[1526]);
    assign outputs[135] = ~((layer0_outputs[3367]) ^ (layer0_outputs[3016]));
    assign outputs[136] = layer0_outputs[400];
    assign outputs[137] = (layer0_outputs[4425]) ^ (layer0_outputs[3403]);
    assign outputs[138] = ~((layer0_outputs[3680]) ^ (layer0_outputs[2632]));
    assign outputs[139] = layer0_outputs[606];
    assign outputs[140] = layer0_outputs[2525];
    assign outputs[141] = (layer0_outputs[1239]) ^ (layer0_outputs[3533]);
    assign outputs[142] = (layer0_outputs[3335]) & (layer0_outputs[516]);
    assign outputs[143] = ~(layer0_outputs[453]);
    assign outputs[144] = layer0_outputs[685];
    assign outputs[145] = ~(layer0_outputs[977]);
    assign outputs[146] = ~((layer0_outputs[1654]) ^ (layer0_outputs[2447]));
    assign outputs[147] = layer0_outputs[4733];
    assign outputs[148] = (layer0_outputs[4838]) & ~(layer0_outputs[1]);
    assign outputs[149] = (layer0_outputs[3194]) & ~(layer0_outputs[2954]);
    assign outputs[150] = (layer0_outputs[2730]) & ~(layer0_outputs[2860]);
    assign outputs[151] = (layer0_outputs[2457]) ^ (layer0_outputs[3795]);
    assign outputs[152] = (layer0_outputs[2169]) ^ (layer0_outputs[1518]);
    assign outputs[153] = ~(layer0_outputs[2740]);
    assign outputs[154] = ~(layer0_outputs[1550]);
    assign outputs[155] = ~(layer0_outputs[1881]) | (layer0_outputs[1679]);
    assign outputs[156] = ~(layer0_outputs[5031]);
    assign outputs[157] = ~(layer0_outputs[120]);
    assign outputs[158] = (layer0_outputs[4936]) ^ (layer0_outputs[4052]);
    assign outputs[159] = ~((layer0_outputs[3259]) ^ (layer0_outputs[2694]));
    assign outputs[160] = ~(layer0_outputs[2403]);
    assign outputs[161] = ~(layer0_outputs[3590]) | (layer0_outputs[1161]);
    assign outputs[162] = layer0_outputs[702];
    assign outputs[163] = ~((layer0_outputs[673]) | (layer0_outputs[1291]));
    assign outputs[164] = (layer0_outputs[221]) & ~(layer0_outputs[2399]);
    assign outputs[165] = ~((layer0_outputs[3112]) ^ (layer0_outputs[3149]));
    assign outputs[166] = ~(layer0_outputs[4496]);
    assign outputs[167] = ~(layer0_outputs[3456]) | (layer0_outputs[1666]);
    assign outputs[168] = ~(layer0_outputs[4967]);
    assign outputs[169] = (layer0_outputs[2603]) | (layer0_outputs[1503]);
    assign outputs[170] = (layer0_outputs[3310]) & ~(layer0_outputs[4101]);
    assign outputs[171] = ~((layer0_outputs[4605]) ^ (layer0_outputs[3549]));
    assign outputs[172] = ~((layer0_outputs[4931]) & (layer0_outputs[2295]));
    assign outputs[173] = ~((layer0_outputs[687]) ^ (layer0_outputs[4777]));
    assign outputs[174] = (layer0_outputs[2860]) ^ (layer0_outputs[708]);
    assign outputs[175] = ~(layer0_outputs[747]);
    assign outputs[176] = ~((layer0_outputs[2218]) ^ (layer0_outputs[2856]));
    assign outputs[177] = layer0_outputs[2769];
    assign outputs[178] = layer0_outputs[652];
    assign outputs[179] = layer0_outputs[1638];
    assign outputs[180] = ~(layer0_outputs[1877]);
    assign outputs[181] = ~(layer0_outputs[4137]) | (layer0_outputs[3762]);
    assign outputs[182] = ~((layer0_outputs[645]) & (layer0_outputs[3521]));
    assign outputs[183] = (layer0_outputs[5105]) & (layer0_outputs[1132]);
    assign outputs[184] = ~((layer0_outputs[3617]) & (layer0_outputs[4233]));
    assign outputs[185] = ~(layer0_outputs[1987]);
    assign outputs[186] = ~((layer0_outputs[5017]) & (layer0_outputs[1715]));
    assign outputs[187] = ~(layer0_outputs[984]);
    assign outputs[188] = ~(layer0_outputs[4255]);
    assign outputs[189] = (layer0_outputs[569]) & ~(layer0_outputs[2335]);
    assign outputs[190] = (layer0_outputs[4627]) ^ (layer0_outputs[1078]);
    assign outputs[191] = ~((layer0_outputs[127]) & (layer0_outputs[1546]));
    assign outputs[192] = ~(layer0_outputs[966]) | (layer0_outputs[2974]);
    assign outputs[193] = ~(layer0_outputs[1731]) | (layer0_outputs[988]);
    assign outputs[194] = layer0_outputs[2429];
    assign outputs[195] = (layer0_outputs[2338]) & ~(layer0_outputs[3591]);
    assign outputs[196] = layer0_outputs[5088];
    assign outputs[197] = ~(layer0_outputs[4907]);
    assign outputs[198] = (layer0_outputs[1598]) & ~(layer0_outputs[2501]);
    assign outputs[199] = (layer0_outputs[498]) & ~(layer0_outputs[1923]);
    assign outputs[200] = ~((layer0_outputs[3273]) ^ (layer0_outputs[394]));
    assign outputs[201] = layer0_outputs[778];
    assign outputs[202] = (layer0_outputs[4950]) & ~(layer0_outputs[3211]);
    assign outputs[203] = ~(layer0_outputs[1002]);
    assign outputs[204] = layer0_outputs[639];
    assign outputs[205] = ~((layer0_outputs[4988]) ^ (layer0_outputs[2708]));
    assign outputs[206] = layer0_outputs[2752];
    assign outputs[207] = ~(layer0_outputs[1700]);
    assign outputs[208] = ~((layer0_outputs[4667]) ^ (layer0_outputs[1384]));
    assign outputs[209] = (layer0_outputs[3219]) | (layer0_outputs[5060]);
    assign outputs[210] = ~((layer0_outputs[1123]) & (layer0_outputs[3189]));
    assign outputs[211] = ~((layer0_outputs[4902]) ^ (layer0_outputs[81]));
    assign outputs[212] = ~(layer0_outputs[1612]);
    assign outputs[213] = (layer0_outputs[1400]) & (layer0_outputs[869]);
    assign outputs[214] = ~((layer0_outputs[4055]) ^ (layer0_outputs[3464]));
    assign outputs[215] = layer0_outputs[2507];
    assign outputs[216] = ~(layer0_outputs[5075]) | (layer0_outputs[4083]);
    assign outputs[217] = layer0_outputs[3748];
    assign outputs[218] = layer0_outputs[4048];
    assign outputs[219] = (layer0_outputs[2189]) ^ (layer0_outputs[3110]);
    assign outputs[220] = layer0_outputs[311];
    assign outputs[221] = layer0_outputs[516];
    assign outputs[222] = layer0_outputs[968];
    assign outputs[223] = ~(layer0_outputs[872]);
    assign outputs[224] = ~(layer0_outputs[1888]);
    assign outputs[225] = ~(layer0_outputs[1063]) | (layer0_outputs[75]);
    assign outputs[226] = layer0_outputs[808];
    assign outputs[227] = layer0_outputs[750];
    assign outputs[228] = ~(layer0_outputs[1085]) | (layer0_outputs[705]);
    assign outputs[229] = layer0_outputs[295];
    assign outputs[230] = (layer0_outputs[3966]) & ~(layer0_outputs[0]);
    assign outputs[231] = ~(layer0_outputs[4923]) | (layer0_outputs[3273]);
    assign outputs[232] = ~((layer0_outputs[3692]) ^ (layer0_outputs[3200]));
    assign outputs[233] = ~(layer0_outputs[189]);
    assign outputs[234] = layer0_outputs[3140];
    assign outputs[235] = (layer0_outputs[1801]) ^ (layer0_outputs[1535]);
    assign outputs[236] = ~((layer0_outputs[1073]) & (layer0_outputs[3892]));
    assign outputs[237] = ~((layer0_outputs[2268]) ^ (layer0_outputs[2341]));
    assign outputs[238] = ~((layer0_outputs[1546]) & (layer0_outputs[1847]));
    assign outputs[239] = layer0_outputs[4965];
    assign outputs[240] = (layer0_outputs[4604]) & (layer0_outputs[2752]);
    assign outputs[241] = 1'b1;
    assign outputs[242] = layer0_outputs[4532];
    assign outputs[243] = (layer0_outputs[779]) & ~(layer0_outputs[688]);
    assign outputs[244] = layer0_outputs[4969];
    assign outputs[245] = (layer0_outputs[492]) | (layer0_outputs[3514]);
    assign outputs[246] = (layer0_outputs[2365]) & (layer0_outputs[4090]);
    assign outputs[247] = layer0_outputs[4651];
    assign outputs[248] = ~(layer0_outputs[4907]);
    assign outputs[249] = ~((layer0_outputs[3730]) ^ (layer0_outputs[1635]));
    assign outputs[250] = ~((layer0_outputs[614]) ^ (layer0_outputs[2731]));
    assign outputs[251] = ~(layer0_outputs[1816]);
    assign outputs[252] = (layer0_outputs[1340]) ^ (layer0_outputs[295]);
    assign outputs[253] = ~((layer0_outputs[2724]) & (layer0_outputs[914]));
    assign outputs[254] = (layer0_outputs[665]) & ~(layer0_outputs[4392]);
    assign outputs[255] = (layer0_outputs[4196]) & (layer0_outputs[2162]);
    assign outputs[256] = ~(layer0_outputs[4129]) | (layer0_outputs[1634]);
    assign outputs[257] = layer0_outputs[1513];
    assign outputs[258] = (layer0_outputs[3390]) ^ (layer0_outputs[2179]);
    assign outputs[259] = ~((layer0_outputs[2931]) ^ (layer0_outputs[2682]));
    assign outputs[260] = (layer0_outputs[1458]) & (layer0_outputs[2279]);
    assign outputs[261] = (layer0_outputs[1608]) ^ (layer0_outputs[3984]);
    assign outputs[262] = layer0_outputs[2558];
    assign outputs[263] = ~((layer0_outputs[4128]) | (layer0_outputs[2388]));
    assign outputs[264] = (layer0_outputs[1186]) & ~(layer0_outputs[297]);
    assign outputs[265] = layer0_outputs[4080];
    assign outputs[266] = layer0_outputs[4628];
    assign outputs[267] = layer0_outputs[4295];
    assign outputs[268] = (layer0_outputs[4838]) & (layer0_outputs[240]);
    assign outputs[269] = ~(layer0_outputs[4374]);
    assign outputs[270] = ~(layer0_outputs[3811]);
    assign outputs[271] = (layer0_outputs[4201]) | (layer0_outputs[1472]);
    assign outputs[272] = ~(layer0_outputs[2893]);
    assign outputs[273] = (layer0_outputs[4789]) & (layer0_outputs[3160]);
    assign outputs[274] = ~(layer0_outputs[2988]);
    assign outputs[275] = 1'b1;
    assign outputs[276] = (layer0_outputs[735]) ^ (layer0_outputs[3173]);
    assign outputs[277] = layer0_outputs[2566];
    assign outputs[278] = (layer0_outputs[1156]) ^ (layer0_outputs[3698]);
    assign outputs[279] = layer0_outputs[401];
    assign outputs[280] = ~(layer0_outputs[737]);
    assign outputs[281] = ~((layer0_outputs[64]) ^ (layer0_outputs[3329]));
    assign outputs[282] = ~(layer0_outputs[1380]);
    assign outputs[283] = layer0_outputs[4847];
    assign outputs[284] = ~(layer0_outputs[1720]) | (layer0_outputs[746]);
    assign outputs[285] = layer0_outputs[311];
    assign outputs[286] = ~((layer0_outputs[1296]) ^ (layer0_outputs[4277]));
    assign outputs[287] = ~((layer0_outputs[1884]) ^ (layer0_outputs[3845]));
    assign outputs[288] = (layer0_outputs[2222]) | (layer0_outputs[3185]);
    assign outputs[289] = (layer0_outputs[4551]) & ~(layer0_outputs[3755]);
    assign outputs[290] = ~((layer0_outputs[2516]) | (layer0_outputs[3786]));
    assign outputs[291] = ~(layer0_outputs[2716]);
    assign outputs[292] = (layer0_outputs[3888]) & ~(layer0_outputs[4288]);
    assign outputs[293] = (layer0_outputs[505]) & ~(layer0_outputs[4585]);
    assign outputs[294] = (layer0_outputs[4474]) & ~(layer0_outputs[3775]);
    assign outputs[295] = ~(layer0_outputs[118]);
    assign outputs[296] = ~((layer0_outputs[774]) | (layer0_outputs[636]));
    assign outputs[297] = ~((layer0_outputs[3742]) & (layer0_outputs[4470]));
    assign outputs[298] = ~(layer0_outputs[3834]) | (layer0_outputs[4054]);
    assign outputs[299] = layer0_outputs[838];
    assign outputs[300] = (layer0_outputs[122]) ^ (layer0_outputs[1025]);
    assign outputs[301] = layer0_outputs[3923];
    assign outputs[302] = ~((layer0_outputs[5097]) & (layer0_outputs[1779]));
    assign outputs[303] = (layer0_outputs[3380]) & ~(layer0_outputs[1642]);
    assign outputs[304] = ~(layer0_outputs[2260]);
    assign outputs[305] = (layer0_outputs[3045]) | (layer0_outputs[3256]);
    assign outputs[306] = layer0_outputs[3384];
    assign outputs[307] = ~(layer0_outputs[59]);
    assign outputs[308] = ~(layer0_outputs[3967]);
    assign outputs[309] = layer0_outputs[4904];
    assign outputs[310] = layer0_outputs[3783];
    assign outputs[311] = (layer0_outputs[196]) ^ (layer0_outputs[1288]);
    assign outputs[312] = layer0_outputs[1311];
    assign outputs[313] = ~(layer0_outputs[704]);
    assign outputs[314] = layer0_outputs[1106];
    assign outputs[315] = ~(layer0_outputs[4859]);
    assign outputs[316] = ~((layer0_outputs[4206]) | (layer0_outputs[62]));
    assign outputs[317] = (layer0_outputs[2362]) | (layer0_outputs[1264]);
    assign outputs[318] = ~(layer0_outputs[4766]);
    assign outputs[319] = layer0_outputs[4356];
    assign outputs[320] = ~((layer0_outputs[3075]) & (layer0_outputs[833]));
    assign outputs[321] = ~(layer0_outputs[2692]) | (layer0_outputs[3007]);
    assign outputs[322] = ~(layer0_outputs[5070]);
    assign outputs[323] = ~(layer0_outputs[2301]);
    assign outputs[324] = ~(layer0_outputs[2181]);
    assign outputs[325] = ~(layer0_outputs[4983]);
    assign outputs[326] = ~((layer0_outputs[4360]) ^ (layer0_outputs[1966]));
    assign outputs[327] = (layer0_outputs[702]) | (layer0_outputs[2138]);
    assign outputs[328] = ~((layer0_outputs[692]) | (layer0_outputs[1479]));
    assign outputs[329] = layer0_outputs[4696];
    assign outputs[330] = ~((layer0_outputs[1428]) ^ (layer0_outputs[2227]));
    assign outputs[331] = ~(layer0_outputs[1273]);
    assign outputs[332] = layer0_outputs[3147];
    assign outputs[333] = (layer0_outputs[4388]) ^ (layer0_outputs[2201]);
    assign outputs[334] = (layer0_outputs[2662]) | (layer0_outputs[2959]);
    assign outputs[335] = (layer0_outputs[1232]) ^ (layer0_outputs[876]);
    assign outputs[336] = layer0_outputs[3481];
    assign outputs[337] = (layer0_outputs[3277]) | (layer0_outputs[18]);
    assign outputs[338] = layer0_outputs[4651];
    assign outputs[339] = ~(layer0_outputs[678]) | (layer0_outputs[1532]);
    assign outputs[340] = layer0_outputs[5111];
    assign outputs[341] = ~((layer0_outputs[1469]) ^ (layer0_outputs[4060]));
    assign outputs[342] = ~(layer0_outputs[1391]) | (layer0_outputs[4327]);
    assign outputs[343] = ~(layer0_outputs[2161]);
    assign outputs[344] = ~(layer0_outputs[2877]);
    assign outputs[345] = (layer0_outputs[3507]) & ~(layer0_outputs[803]);
    assign outputs[346] = ~(layer0_outputs[1710]) | (layer0_outputs[1186]);
    assign outputs[347] = ~((layer0_outputs[4834]) | (layer0_outputs[4900]));
    assign outputs[348] = (layer0_outputs[2283]) & (layer0_outputs[1569]);
    assign outputs[349] = (layer0_outputs[2757]) & (layer0_outputs[2645]);
    assign outputs[350] = (layer0_outputs[1749]) | (layer0_outputs[2261]);
    assign outputs[351] = ~((layer0_outputs[2657]) & (layer0_outputs[3248]));
    assign outputs[352] = ~((layer0_outputs[4161]) | (layer0_outputs[820]));
    assign outputs[353] = ~(layer0_outputs[180]) | (layer0_outputs[3707]);
    assign outputs[354] = ~((layer0_outputs[2046]) | (layer0_outputs[765]));
    assign outputs[355] = ~(layer0_outputs[811]) | (layer0_outputs[959]);
    assign outputs[356] = ~((layer0_outputs[3690]) | (layer0_outputs[733]));
    assign outputs[357] = ~((layer0_outputs[4001]) ^ (layer0_outputs[1594]));
    assign outputs[358] = (layer0_outputs[4369]) & (layer0_outputs[711]);
    assign outputs[359] = ~((layer0_outputs[2276]) | (layer0_outputs[1920]));
    assign outputs[360] = ~((layer0_outputs[3128]) | (layer0_outputs[2472]));
    assign outputs[361] = ~((layer0_outputs[1860]) ^ (layer0_outputs[1014]));
    assign outputs[362] = (layer0_outputs[1701]) & (layer0_outputs[4608]);
    assign outputs[363] = (layer0_outputs[2585]) ^ (layer0_outputs[652]);
    assign outputs[364] = ~((layer0_outputs[3637]) | (layer0_outputs[1476]));
    assign outputs[365] = layer0_outputs[4726];
    assign outputs[366] = ~(layer0_outputs[4290]);
    assign outputs[367] = layer0_outputs[3094];
    assign outputs[368] = layer0_outputs[4387];
    assign outputs[369] = ~(layer0_outputs[4541]);
    assign outputs[370] = layer0_outputs[4913];
    assign outputs[371] = layer0_outputs[2230];
    assign outputs[372] = (layer0_outputs[2260]) ^ (layer0_outputs[1301]);
    assign outputs[373] = (layer0_outputs[1232]) ^ (layer0_outputs[2527]);
    assign outputs[374] = ~(layer0_outputs[178]);
    assign outputs[375] = layer0_outputs[2679];
    assign outputs[376] = (layer0_outputs[2786]) ^ (layer0_outputs[4318]);
    assign outputs[377] = ~(layer0_outputs[1028]);
    assign outputs[378] = ~(layer0_outputs[795]);
    assign outputs[379] = ~(layer0_outputs[3473]) | (layer0_outputs[4817]);
    assign outputs[380] = layer0_outputs[4914];
    assign outputs[381] = (layer0_outputs[2355]) ^ (layer0_outputs[3321]);
    assign outputs[382] = ~(layer0_outputs[210]);
    assign outputs[383] = (layer0_outputs[3535]) & (layer0_outputs[3732]);
    assign outputs[384] = ~(layer0_outputs[4735]) | (layer0_outputs[823]);
    assign outputs[385] = ~(layer0_outputs[187]);
    assign outputs[386] = layer0_outputs[1565];
    assign outputs[387] = ~((layer0_outputs[1158]) & (layer0_outputs[1558]));
    assign outputs[388] = ~(layer0_outputs[4520]);
    assign outputs[389] = ~((layer0_outputs[37]) & (layer0_outputs[1818]));
    assign outputs[390] = layer0_outputs[4797];
    assign outputs[391] = ~(layer0_outputs[456]) | (layer0_outputs[2475]);
    assign outputs[392] = ~((layer0_outputs[496]) & (layer0_outputs[3500]));
    assign outputs[393] = layer0_outputs[4443];
    assign outputs[394] = layer0_outputs[3808];
    assign outputs[395] = layer0_outputs[2121];
    assign outputs[396] = layer0_outputs[3935];
    assign outputs[397] = ~((layer0_outputs[445]) & (layer0_outputs[1501]));
    assign outputs[398] = ~(layer0_outputs[2552]) | (layer0_outputs[548]);
    assign outputs[399] = ~(layer0_outputs[264]) | (layer0_outputs[3418]);
    assign outputs[400] = (layer0_outputs[7]) ^ (layer0_outputs[2173]);
    assign outputs[401] = ~(layer0_outputs[806]);
    assign outputs[402] = layer0_outputs[4501];
    assign outputs[403] = ~((layer0_outputs[3527]) | (layer0_outputs[1480]));
    assign outputs[404] = (layer0_outputs[4507]) & (layer0_outputs[2177]);
    assign outputs[405] = (layer0_outputs[2059]) & ~(layer0_outputs[4185]);
    assign outputs[406] = (layer0_outputs[371]) & ~(layer0_outputs[3882]);
    assign outputs[407] = ~(layer0_outputs[1637]);
    assign outputs[408] = layer0_outputs[2019];
    assign outputs[409] = ~(layer0_outputs[5000]);
    assign outputs[410] = (layer0_outputs[4661]) & ~(layer0_outputs[307]);
    assign outputs[411] = ~(layer0_outputs[3075]);
    assign outputs[412] = layer0_outputs[344];
    assign outputs[413] = ~(layer0_outputs[1774]) | (layer0_outputs[4394]);
    assign outputs[414] = ~(layer0_outputs[3192]);
    assign outputs[415] = layer0_outputs[4354];
    assign outputs[416] = ~(layer0_outputs[2049]);
    assign outputs[417] = ~((layer0_outputs[4923]) & (layer0_outputs[3976]));
    assign outputs[418] = ~(layer0_outputs[610]);
    assign outputs[419] = layer0_outputs[296];
    assign outputs[420] = (layer0_outputs[2105]) ^ (layer0_outputs[953]);
    assign outputs[421] = ~(layer0_outputs[4248]) | (layer0_outputs[2480]);
    assign outputs[422] = layer0_outputs[4560];
    assign outputs[423] = ~((layer0_outputs[206]) | (layer0_outputs[2406]));
    assign outputs[424] = layer0_outputs[1420];
    assign outputs[425] = ~(layer0_outputs[2132]) | (layer0_outputs[4491]);
    assign outputs[426] = (layer0_outputs[3290]) ^ (layer0_outputs[4046]);
    assign outputs[427] = (layer0_outputs[3222]) & ~(layer0_outputs[228]);
    assign outputs[428] = (layer0_outputs[4425]) | (layer0_outputs[1005]);
    assign outputs[429] = (layer0_outputs[2920]) & ~(layer0_outputs[4179]);
    assign outputs[430] = ~((layer0_outputs[3846]) & (layer0_outputs[2987]));
    assign outputs[431] = ~((layer0_outputs[3509]) | (layer0_outputs[4757]));
    assign outputs[432] = layer0_outputs[4166];
    assign outputs[433] = layer0_outputs[2213];
    assign outputs[434] = ~(layer0_outputs[3395]) | (layer0_outputs[4205]);
    assign outputs[435] = layer0_outputs[42];
    assign outputs[436] = (layer0_outputs[4050]) & ~(layer0_outputs[3152]);
    assign outputs[437] = layer0_outputs[906];
    assign outputs[438] = layer0_outputs[4424];
    assign outputs[439] = layer0_outputs[1304];
    assign outputs[440] = (layer0_outputs[2997]) & (layer0_outputs[591]);
    assign outputs[441] = layer0_outputs[353];
    assign outputs[442] = ~(layer0_outputs[1140]);
    assign outputs[443] = ~(layer0_outputs[44]);
    assign outputs[444] = ~((layer0_outputs[3846]) & (layer0_outputs[4496]));
    assign outputs[445] = ~(layer0_outputs[3908]);
    assign outputs[446] = ~(layer0_outputs[764]) | (layer0_outputs[4754]);
    assign outputs[447] = ~(layer0_outputs[4943]) | (layer0_outputs[3289]);
    assign outputs[448] = ~(layer0_outputs[2300]);
    assign outputs[449] = 1'b0;
    assign outputs[450] = ~((layer0_outputs[2865]) & (layer0_outputs[1279]));
    assign outputs[451] = (layer0_outputs[684]) | (layer0_outputs[588]);
    assign outputs[452] = (layer0_outputs[4017]) ^ (layer0_outputs[3003]);
    assign outputs[453] = ~((layer0_outputs[2886]) ^ (layer0_outputs[3253]));
    assign outputs[454] = ~((layer0_outputs[4553]) ^ (layer0_outputs[4723]));
    assign outputs[455] = (layer0_outputs[763]) ^ (layer0_outputs[5005]);
    assign outputs[456] = ~(layer0_outputs[2228]);
    assign outputs[457] = ~(layer0_outputs[3591]) | (layer0_outputs[723]);
    assign outputs[458] = (layer0_outputs[3676]) ^ (layer0_outputs[3917]);
    assign outputs[459] = (layer0_outputs[2688]) | (layer0_outputs[5040]);
    assign outputs[460] = layer0_outputs[858];
    assign outputs[461] = (layer0_outputs[3442]) ^ (layer0_outputs[1086]);
    assign outputs[462] = ~(layer0_outputs[4882]);
    assign outputs[463] = layer0_outputs[4628];
    assign outputs[464] = layer0_outputs[4103];
    assign outputs[465] = ~(layer0_outputs[2600]);
    assign outputs[466] = layer0_outputs[5100];
    assign outputs[467] = ~((layer0_outputs[1837]) & (layer0_outputs[2898]));
    assign outputs[468] = layer0_outputs[2802];
    assign outputs[469] = layer0_outputs[3091];
    assign outputs[470] = ~(layer0_outputs[3850]);
    assign outputs[471] = (layer0_outputs[4306]) ^ (layer0_outputs[4709]);
    assign outputs[472] = layer0_outputs[3225];
    assign outputs[473] = ~((layer0_outputs[14]) | (layer0_outputs[4970]));
    assign outputs[474] = ~(layer0_outputs[661]) | (layer0_outputs[3172]);
    assign outputs[475] = ~(layer0_outputs[2693]);
    assign outputs[476] = ~(layer0_outputs[683]) | (layer0_outputs[4227]);
    assign outputs[477] = ~((layer0_outputs[4460]) ^ (layer0_outputs[3468]));
    assign outputs[478] = ~(layer0_outputs[1786]);
    assign outputs[479] = ~(layer0_outputs[3467]) | (layer0_outputs[2717]);
    assign outputs[480] = layer0_outputs[2789];
    assign outputs[481] = ~(layer0_outputs[2805]);
    assign outputs[482] = ~((layer0_outputs[2328]) ^ (layer0_outputs[4800]));
    assign outputs[483] = ~(layer0_outputs[3483]);
    assign outputs[484] = ~((layer0_outputs[2193]) & (layer0_outputs[1614]));
    assign outputs[485] = ~(layer0_outputs[1332]);
    assign outputs[486] = (layer0_outputs[2577]) | (layer0_outputs[1471]);
    assign outputs[487] = layer0_outputs[3492];
    assign outputs[488] = layer0_outputs[477];
    assign outputs[489] = layer0_outputs[4121];
    assign outputs[490] = layer0_outputs[4922];
    assign outputs[491] = ~((layer0_outputs[1422]) ^ (layer0_outputs[3072]));
    assign outputs[492] = (layer0_outputs[4855]) & (layer0_outputs[1414]);
    assign outputs[493] = (layer0_outputs[4665]) & ~(layer0_outputs[3224]);
    assign outputs[494] = ~(layer0_outputs[519]);
    assign outputs[495] = ~(layer0_outputs[815]) | (layer0_outputs[1390]);
    assign outputs[496] = ~(layer0_outputs[1760]);
    assign outputs[497] = layer0_outputs[804];
    assign outputs[498] = ~(layer0_outputs[3325]);
    assign outputs[499] = (layer0_outputs[418]) | (layer0_outputs[2460]);
    assign outputs[500] = (layer0_outputs[4019]) | (layer0_outputs[3354]);
    assign outputs[501] = ~((layer0_outputs[2487]) | (layer0_outputs[4692]));
    assign outputs[502] = ~(layer0_outputs[1955]);
    assign outputs[503] = (layer0_outputs[32]) & ~(layer0_outputs[3452]);
    assign outputs[504] = layer0_outputs[319];
    assign outputs[505] = ~(layer0_outputs[2552]);
    assign outputs[506] = ~((layer0_outputs[3331]) ^ (layer0_outputs[3671]));
    assign outputs[507] = layer0_outputs[230];
    assign outputs[508] = ~(layer0_outputs[1520]);
    assign outputs[509] = ~(layer0_outputs[3152]);
    assign outputs[510] = ~(layer0_outputs[4541]);
    assign outputs[511] = ~((layer0_outputs[2340]) & (layer0_outputs[2452]));
    assign outputs[512] = layer0_outputs[2060];
    assign outputs[513] = (layer0_outputs[4677]) & (layer0_outputs[253]);
    assign outputs[514] = layer0_outputs[1998];
    assign outputs[515] = layer0_outputs[2764];
    assign outputs[516] = (layer0_outputs[850]) ^ (layer0_outputs[368]);
    assign outputs[517] = (layer0_outputs[961]) ^ (layer0_outputs[1566]);
    assign outputs[518] = (layer0_outputs[2108]) & ~(layer0_outputs[2892]);
    assign outputs[519] = ~((layer0_outputs[3400]) | (layer0_outputs[363]));
    assign outputs[520] = (layer0_outputs[3245]) & (layer0_outputs[3287]);
    assign outputs[521] = (layer0_outputs[3884]) & (layer0_outputs[2470]);
    assign outputs[522] = ~(layer0_outputs[4383]);
    assign outputs[523] = (layer0_outputs[241]) & (layer0_outputs[4211]);
    assign outputs[524] = (layer0_outputs[3287]) & ~(layer0_outputs[908]);
    assign outputs[525] = ~(layer0_outputs[127]);
    assign outputs[526] = ~((layer0_outputs[4827]) | (layer0_outputs[2044]));
    assign outputs[527] = ~(layer0_outputs[1421]);
    assign outputs[528] = (layer0_outputs[4190]) & (layer0_outputs[3766]);
    assign outputs[529] = (layer0_outputs[4555]) & ~(layer0_outputs[3706]);
    assign outputs[530] = (layer0_outputs[3381]) & (layer0_outputs[1019]);
    assign outputs[531] = (layer0_outputs[3740]) & (layer0_outputs[405]);
    assign outputs[532] = (layer0_outputs[3086]) ^ (layer0_outputs[4312]);
    assign outputs[533] = ~((layer0_outputs[3099]) | (layer0_outputs[4447]));
    assign outputs[534] = ~((layer0_outputs[475]) ^ (layer0_outputs[393]));
    assign outputs[535] = (layer0_outputs[3498]) & ~(layer0_outputs[4359]);
    assign outputs[536] = ~(layer0_outputs[4467]) | (layer0_outputs[4001]);
    assign outputs[537] = 1'b0;
    assign outputs[538] = (layer0_outputs[2264]) & ~(layer0_outputs[1455]);
    assign outputs[539] = layer0_outputs[1189];
    assign outputs[540] = (layer0_outputs[397]) & ~(layer0_outputs[3184]);
    assign outputs[541] = (layer0_outputs[4072]) & ~(layer0_outputs[4884]);
    assign outputs[542] = (layer0_outputs[4235]) & ~(layer0_outputs[2166]);
    assign outputs[543] = ~((layer0_outputs[4036]) ^ (layer0_outputs[1552]));
    assign outputs[544] = layer0_outputs[981];
    assign outputs[545] = 1'b0;
    assign outputs[546] = (layer0_outputs[4935]) ^ (layer0_outputs[1379]);
    assign outputs[547] = ~((layer0_outputs[3289]) | (layer0_outputs[1087]));
    assign outputs[548] = ~((layer0_outputs[898]) ^ (layer0_outputs[163]));
    assign outputs[549] = (layer0_outputs[425]) & (layer0_outputs[2450]);
    assign outputs[550] = (layer0_outputs[1786]) & (layer0_outputs[1592]);
    assign outputs[551] = (layer0_outputs[2920]) & (layer0_outputs[1014]);
    assign outputs[552] = (layer0_outputs[309]) & (layer0_outputs[367]);
    assign outputs[553] = (layer0_outputs[2140]) ^ (layer0_outputs[1770]);
    assign outputs[554] = ~(layer0_outputs[3304]) | (layer0_outputs[2962]);
    assign outputs[555] = (layer0_outputs[112]) & ~(layer0_outputs[3430]);
    assign outputs[556] = ~((layer0_outputs[2993]) ^ (layer0_outputs[2737]));
    assign outputs[557] = ~(layer0_outputs[459]);
    assign outputs[558] = ~(layer0_outputs[2787]);
    assign outputs[559] = ~((layer0_outputs[2702]) | (layer0_outputs[2753]));
    assign outputs[560] = (layer0_outputs[1814]) ^ (layer0_outputs[3629]);
    assign outputs[561] = ~(layer0_outputs[2672]);
    assign outputs[562] = 1'b0;
    assign outputs[563] = ~((layer0_outputs[135]) ^ (layer0_outputs[1182]));
    assign outputs[564] = ~(layer0_outputs[4044]);
    assign outputs[565] = layer0_outputs[4815];
    assign outputs[566] = (layer0_outputs[1058]) ^ (layer0_outputs[2424]);
    assign outputs[567] = ~((layer0_outputs[2520]) | (layer0_outputs[3292]));
    assign outputs[568] = ~((layer0_outputs[3614]) & (layer0_outputs[3351]));
    assign outputs[569] = ~((layer0_outputs[1831]) | (layer0_outputs[269]));
    assign outputs[570] = layer0_outputs[5071];
    assign outputs[571] = (layer0_outputs[243]) & (layer0_outputs[1381]);
    assign outputs[572] = (layer0_outputs[3020]) & ~(layer0_outputs[4731]);
    assign outputs[573] = layer0_outputs[3910];
    assign outputs[574] = ~((layer0_outputs[3750]) | (layer0_outputs[508]));
    assign outputs[575] = (layer0_outputs[1963]) & ~(layer0_outputs[1300]);
    assign outputs[576] = (layer0_outputs[3079]) ^ (layer0_outputs[4133]);
    assign outputs[577] = (layer0_outputs[2417]) & ~(layer0_outputs[1473]);
    assign outputs[578] = layer0_outputs[1784];
    assign outputs[579] = (layer0_outputs[1710]) & ~(layer0_outputs[4636]);
    assign outputs[580] = (layer0_outputs[5078]) & ~(layer0_outputs[1474]);
    assign outputs[581] = (layer0_outputs[2143]) & (layer0_outputs[577]);
    assign outputs[582] = (layer0_outputs[821]) & (layer0_outputs[818]);
    assign outputs[583] = (layer0_outputs[4772]) & ~(layer0_outputs[2982]);
    assign outputs[584] = (layer0_outputs[131]) & (layer0_outputs[601]);
    assign outputs[585] = (layer0_outputs[1579]) & ~(layer0_outputs[882]);
    assign outputs[586] = (layer0_outputs[354]) & ~(layer0_outputs[4921]);
    assign outputs[587] = (layer0_outputs[3423]) & ~(layer0_outputs[700]);
    assign outputs[588] = (layer0_outputs[3709]) & ~(layer0_outputs[2263]);
    assign outputs[589] = ~((layer0_outputs[4556]) | (layer0_outputs[2247]));
    assign outputs[590] = layer0_outputs[1056];
    assign outputs[591] = (layer0_outputs[4444]) ^ (layer0_outputs[2797]);
    assign outputs[592] = ~((layer0_outputs[128]) | (layer0_outputs[1432]));
    assign outputs[593] = ~(layer0_outputs[4877]);
    assign outputs[594] = ~(layer0_outputs[2444]);
    assign outputs[595] = layer0_outputs[4429];
    assign outputs[596] = (layer0_outputs[1489]) & ~(layer0_outputs[3419]);
    assign outputs[597] = (layer0_outputs[4736]) & ~(layer0_outputs[3474]);
    assign outputs[598] = layer0_outputs[2829];
    assign outputs[599] = ~(layer0_outputs[1492]);
    assign outputs[600] = (layer0_outputs[1977]) & ~(layer0_outputs[2298]);
    assign outputs[601] = (layer0_outputs[2864]) & ~(layer0_outputs[5047]);
    assign outputs[602] = (layer0_outputs[4462]) & ~(layer0_outputs[906]);
    assign outputs[603] = (layer0_outputs[4380]) & ~(layer0_outputs[3659]);
    assign outputs[604] = ~(layer0_outputs[3141]);
    assign outputs[605] = (layer0_outputs[1261]) ^ (layer0_outputs[3408]);
    assign outputs[606] = layer0_outputs[4091];
    assign outputs[607] = ~((layer0_outputs[694]) | (layer0_outputs[548]));
    assign outputs[608] = 1'b0;
    assign outputs[609] = ~(layer0_outputs[750]);
    assign outputs[610] = ~((layer0_outputs[2353]) | (layer0_outputs[2378]));
    assign outputs[611] = ~((layer0_outputs[4972]) & (layer0_outputs[1467]));
    assign outputs[612] = ~((layer0_outputs[5089]) ^ (layer0_outputs[291]));
    assign outputs[613] = ~((layer0_outputs[3196]) | (layer0_outputs[4436]));
    assign outputs[614] = ~(layer0_outputs[4536]);
    assign outputs[615] = layer0_outputs[2621];
    assign outputs[616] = layer0_outputs[4324];
    assign outputs[617] = (layer0_outputs[2748]) & ~(layer0_outputs[4826]);
    assign outputs[618] = (layer0_outputs[4035]) & (layer0_outputs[302]);
    assign outputs[619] = layer0_outputs[2309];
    assign outputs[620] = (layer0_outputs[4673]) & ~(layer0_outputs[3661]);
    assign outputs[621] = (layer0_outputs[766]) & (layer0_outputs[3080]);
    assign outputs[622] = (layer0_outputs[970]) & ~(layer0_outputs[2571]);
    assign outputs[623] = (layer0_outputs[2806]) & (layer0_outputs[1198]);
    assign outputs[624] = (layer0_outputs[3128]) & ~(layer0_outputs[834]);
    assign outputs[625] = (layer0_outputs[2879]) ^ (layer0_outputs[2025]);
    assign outputs[626] = ~((layer0_outputs[2020]) | (layer0_outputs[4954]));
    assign outputs[627] = 1'b0;
    assign outputs[628] = layer0_outputs[4132];
    assign outputs[629] = layer0_outputs[4357];
    assign outputs[630] = ~((layer0_outputs[1125]) | (layer0_outputs[3038]));
    assign outputs[631] = (layer0_outputs[3708]) & ~(layer0_outputs[2828]);
    assign outputs[632] = ~((layer0_outputs[3107]) | (layer0_outputs[136]));
    assign outputs[633] = (layer0_outputs[4919]) ^ (layer0_outputs[2880]);
    assign outputs[634] = ~(layer0_outputs[3912]);
    assign outputs[635] = ~((layer0_outputs[1778]) | (layer0_outputs[1173]));
    assign outputs[636] = (layer0_outputs[4139]) & ~(layer0_outputs[463]);
    assign outputs[637] = ~(layer0_outputs[3639]);
    assign outputs[638] = ~((layer0_outputs[3685]) | (layer0_outputs[693]));
    assign outputs[639] = ~(layer0_outputs[3335]);
    assign outputs[640] = (layer0_outputs[4734]) & ~(layer0_outputs[4010]);
    assign outputs[641] = (layer0_outputs[1259]) & (layer0_outputs[3878]);
    assign outputs[642] = ~((layer0_outputs[3745]) | (layer0_outputs[2044]));
    assign outputs[643] = ~((layer0_outputs[1903]) | (layer0_outputs[279]));
    assign outputs[644] = (layer0_outputs[3025]) & ~(layer0_outputs[3398]);
    assign outputs[645] = (layer0_outputs[3553]) & (layer0_outputs[2611]);
    assign outputs[646] = ~((layer0_outputs[952]) ^ (layer0_outputs[888]));
    assign outputs[647] = ~(layer0_outputs[782]);
    assign outputs[648] = layer0_outputs[339];
    assign outputs[649] = layer0_outputs[3429];
    assign outputs[650] = layer0_outputs[1120];
    assign outputs[651] = layer0_outputs[1181];
    assign outputs[652] = ~((layer0_outputs[184]) | (layer0_outputs[3984]));
    assign outputs[653] = (layer0_outputs[2014]) & ~(layer0_outputs[3988]);
    assign outputs[654] = ~(layer0_outputs[4164]);
    assign outputs[655] = ~(layer0_outputs[1467]);
    assign outputs[656] = (layer0_outputs[3400]) ^ (layer0_outputs[2267]);
    assign outputs[657] = ~(layer0_outputs[3522]);
    assign outputs[658] = layer0_outputs[4248];
    assign outputs[659] = ~(layer0_outputs[4069]);
    assign outputs[660] = (layer0_outputs[93]) & ~(layer0_outputs[1599]);
    assign outputs[661] = ~(layer0_outputs[1887]);
    assign outputs[662] = (layer0_outputs[3518]) & (layer0_outputs[4807]);
    assign outputs[663] = ~(layer0_outputs[2508]);
    assign outputs[664] = (layer0_outputs[1976]) & ~(layer0_outputs[720]);
    assign outputs[665] = layer0_outputs[4751];
    assign outputs[666] = (layer0_outputs[4903]) ^ (layer0_outputs[4586]);
    assign outputs[667] = layer0_outputs[2785];
    assign outputs[668] = (layer0_outputs[1718]) & ~(layer0_outputs[2097]);
    assign outputs[669] = (layer0_outputs[3815]) & (layer0_outputs[1872]);
    assign outputs[670] = (layer0_outputs[2483]) & ~(layer0_outputs[4158]);
    assign outputs[671] = (layer0_outputs[3810]) & (layer0_outputs[2152]);
    assign outputs[672] = (layer0_outputs[354]) & ~(layer0_outputs[1285]);
    assign outputs[673] = (layer0_outputs[4795]) ^ (layer0_outputs[2937]);
    assign outputs[674] = (layer0_outputs[3758]) & ~(layer0_outputs[4618]);
    assign outputs[675] = ~(layer0_outputs[3894]);
    assign outputs[676] = ~((layer0_outputs[3415]) | (layer0_outputs[179]));
    assign outputs[677] = ~(layer0_outputs[2122]);
    assign outputs[678] = layer0_outputs[4537];
    assign outputs[679] = ~((layer0_outputs[4899]) | (layer0_outputs[4431]));
    assign outputs[680] = (layer0_outputs[2130]) & ~(layer0_outputs[175]);
    assign outputs[681] = ~((layer0_outputs[4818]) | (layer0_outputs[48]));
    assign outputs[682] = (layer0_outputs[2151]) & ~(layer0_outputs[869]);
    assign outputs[683] = (layer0_outputs[790]) & (layer0_outputs[313]);
    assign outputs[684] = ~(layer0_outputs[1651]) | (layer0_outputs[1135]);
    assign outputs[685] = (layer0_outputs[3032]) & ~(layer0_outputs[3526]);
    assign outputs[686] = layer0_outputs[1788];
    assign outputs[687] = layer0_outputs[4040];
    assign outputs[688] = 1'b0;
    assign outputs[689] = (layer0_outputs[1085]) | (layer0_outputs[3211]);
    assign outputs[690] = (layer0_outputs[938]) & (layer0_outputs[197]);
    assign outputs[691] = ~((layer0_outputs[2070]) ^ (layer0_outputs[5094]));
    assign outputs[692] = ~(layer0_outputs[2286]);
    assign outputs[693] = ~(layer0_outputs[1094]) | (layer0_outputs[2219]);
    assign outputs[694] = ~(layer0_outputs[4478]);
    assign outputs[695] = (layer0_outputs[2464]) & ~(layer0_outputs[846]);
    assign outputs[696] = (layer0_outputs[2863]) & ~(layer0_outputs[2570]);
    assign outputs[697] = layer0_outputs[2211];
    assign outputs[698] = ~(layer0_outputs[232]);
    assign outputs[699] = (layer0_outputs[1735]) & (layer0_outputs[1838]);
    assign outputs[700] = ~((layer0_outputs[2095]) | (layer0_outputs[4086]));
    assign outputs[701] = (layer0_outputs[4846]) & ~(layer0_outputs[2498]);
    assign outputs[702] = (layer0_outputs[1037]) & ~(layer0_outputs[4423]);
    assign outputs[703] = ~(layer0_outputs[4932]);
    assign outputs[704] = ~(layer0_outputs[2529]);
    assign outputs[705] = (layer0_outputs[3718]) & ~(layer0_outputs[4945]);
    assign outputs[706] = (layer0_outputs[1683]) & ~(layer0_outputs[4538]);
    assign outputs[707] = (layer0_outputs[3633]) ^ (layer0_outputs[2163]);
    assign outputs[708] = (layer0_outputs[3967]) & (layer0_outputs[1963]);
    assign outputs[709] = (layer0_outputs[1672]) & (layer0_outputs[1374]);
    assign outputs[710] = (layer0_outputs[2369]) & (layer0_outputs[156]);
    assign outputs[711] = ~(layer0_outputs[1325]);
    assign outputs[712] = (layer0_outputs[3859]) & ~(layer0_outputs[627]);
    assign outputs[713] = layer0_outputs[3740];
    assign outputs[714] = (layer0_outputs[1958]) & ~(layer0_outputs[316]);
    assign outputs[715] = ~((layer0_outputs[4771]) | (layer0_outputs[1119]));
    assign outputs[716] = (layer0_outputs[415]) & (layer0_outputs[2395]);
    assign outputs[717] = ~(layer0_outputs[635]);
    assign outputs[718] = (layer0_outputs[1730]) & (layer0_outputs[4808]);
    assign outputs[719] = (layer0_outputs[292]) & ~(layer0_outputs[2659]);
    assign outputs[720] = ~(layer0_outputs[1603]);
    assign outputs[721] = (layer0_outputs[4138]) & (layer0_outputs[433]);
    assign outputs[722] = ~(layer0_outputs[686]) | (layer0_outputs[4324]);
    assign outputs[723] = (layer0_outputs[137]) ^ (layer0_outputs[1676]);
    assign outputs[724] = ~(layer0_outputs[1195]);
    assign outputs[725] = (layer0_outputs[1932]) & ~(layer0_outputs[3056]);
    assign outputs[726] = (layer0_outputs[2178]) & (layer0_outputs[1907]);
    assign outputs[727] = ~(layer0_outputs[2741]);
    assign outputs[728] = ~(layer0_outputs[2824]);
    assign outputs[729] = (layer0_outputs[1029]) & ~(layer0_outputs[2009]);
    assign outputs[730] = (layer0_outputs[1313]) & ~(layer0_outputs[2906]);
    assign outputs[731] = (layer0_outputs[1631]) & (layer0_outputs[2379]);
    assign outputs[732] = layer0_outputs[774];
    assign outputs[733] = (layer0_outputs[2670]) ^ (layer0_outputs[1525]);
    assign outputs[734] = ~(layer0_outputs[2223]);
    assign outputs[735] = ~(layer0_outputs[4701]);
    assign outputs[736] = ~(layer0_outputs[2528]);
    assign outputs[737] = layer0_outputs[149];
    assign outputs[738] = layer0_outputs[4286];
    assign outputs[739] = (layer0_outputs[2619]) & (layer0_outputs[1695]);
    assign outputs[740] = (layer0_outputs[3921]) & (layer0_outputs[2782]);
    assign outputs[741] = (layer0_outputs[1719]) & ~(layer0_outputs[4291]);
    assign outputs[742] = ~(layer0_outputs[5108]);
    assign outputs[743] = ~(layer0_outputs[4586]);
    assign outputs[744] = ~((layer0_outputs[4642]) | (layer0_outputs[3543]));
    assign outputs[745] = ~(layer0_outputs[860]);
    assign outputs[746] = (layer0_outputs[3598]) & ~(layer0_outputs[3033]);
    assign outputs[747] = 1'b0;
    assign outputs[748] = (layer0_outputs[603]) & (layer0_outputs[2817]);
    assign outputs[749] = (layer0_outputs[3790]) ^ (layer0_outputs[1605]);
    assign outputs[750] = (layer0_outputs[2767]) ^ (layer0_outputs[4548]);
    assign outputs[751] = (layer0_outputs[5057]) ^ (layer0_outputs[4693]);
    assign outputs[752] = layer0_outputs[2174];
    assign outputs[753] = ~(layer0_outputs[5112]);
    assign outputs[754] = (layer0_outputs[1789]) & ~(layer0_outputs[3432]);
    assign outputs[755] = (layer0_outputs[1033]) & ~(layer0_outputs[1603]);
    assign outputs[756] = ~((layer0_outputs[493]) ^ (layer0_outputs[1733]));
    assign outputs[757] = (layer0_outputs[4163]) & ~(layer0_outputs[293]);
    assign outputs[758] = layer0_outputs[2790];
    assign outputs[759] = (layer0_outputs[1411]) & (layer0_outputs[4682]);
    assign outputs[760] = (layer0_outputs[3878]) & ~(layer0_outputs[1919]);
    assign outputs[761] = layer0_outputs[3114];
    assign outputs[762] = layer0_outputs[690];
    assign outputs[763] = (layer0_outputs[666]) & (layer0_outputs[1926]);
    assign outputs[764] = ~(layer0_outputs[2058]);
    assign outputs[765] = (layer0_outputs[3302]) & ~(layer0_outputs[3031]);
    assign outputs[766] = ~((layer0_outputs[356]) | (layer0_outputs[2883]));
    assign outputs[767] = (layer0_outputs[759]) & ~(layer0_outputs[198]);
    assign outputs[768] = (layer0_outputs[379]) & (layer0_outputs[3642]);
    assign outputs[769] = (layer0_outputs[2393]) & (layer0_outputs[2798]);
    assign outputs[770] = (layer0_outputs[5090]) & ~(layer0_outputs[1895]);
    assign outputs[771] = (layer0_outputs[1422]) & (layer0_outputs[1164]);
    assign outputs[772] = ~((layer0_outputs[1780]) | (layer0_outputs[2648]));
    assign outputs[773] = (layer0_outputs[3381]) & (layer0_outputs[1527]);
    assign outputs[774] = (layer0_outputs[2074]) & ~(layer0_outputs[4542]);
    assign outputs[775] = (layer0_outputs[3736]) ^ (layer0_outputs[2827]);
    assign outputs[776] = (layer0_outputs[435]) & (layer0_outputs[3406]);
    assign outputs[777] = layer0_outputs[1286];
    assign outputs[778] = layer0_outputs[1596];
    assign outputs[779] = ~((layer0_outputs[2069]) | (layer0_outputs[4198]));
    assign outputs[780] = 1'b0;
    assign outputs[781] = (layer0_outputs[4872]) & ~(layer0_outputs[1530]);
    assign outputs[782] = layer0_outputs[2831];
    assign outputs[783] = layer0_outputs[4660];
    assign outputs[784] = (layer0_outputs[1081]) & (layer0_outputs[398]);
    assign outputs[785] = ~((layer0_outputs[4837]) | (layer0_outputs[1221]));
    assign outputs[786] = (layer0_outputs[1554]) & ~(layer0_outputs[4255]);
    assign outputs[787] = (layer0_outputs[2468]) & (layer0_outputs[3845]);
    assign outputs[788] = ~((layer0_outputs[3968]) | (layer0_outputs[3904]));
    assign outputs[789] = (layer0_outputs[578]) & ~(layer0_outputs[3547]);
    assign outputs[790] = ~((layer0_outputs[3820]) & (layer0_outputs[4488]));
    assign outputs[791] = ~((layer0_outputs[521]) | (layer0_outputs[4264]));
    assign outputs[792] = (layer0_outputs[1055]) & ~(layer0_outputs[1775]);
    assign outputs[793] = (layer0_outputs[4364]) & ~(layer0_outputs[5072]);
    assign outputs[794] = (layer0_outputs[3039]) & ~(layer0_outputs[3488]);
    assign outputs[795] = layer0_outputs[1452];
    assign outputs[796] = (layer0_outputs[1039]) & ~(layer0_outputs[3800]);
    assign outputs[797] = ~((layer0_outputs[1032]) | (layer0_outputs[1479]));
    assign outputs[798] = layer0_outputs[1061];
    assign outputs[799] = layer0_outputs[5085];
    assign outputs[800] = layer0_outputs[1016];
    assign outputs[801] = layer0_outputs[2885];
    assign outputs[802] = ~(layer0_outputs[3877]);
    assign outputs[803] = (layer0_outputs[2536]) & ~(layer0_outputs[2718]);
    assign outputs[804] = ~((layer0_outputs[1270]) | (layer0_outputs[1316]));
    assign outputs[805] = (layer0_outputs[1436]) & ~(layer0_outputs[2113]);
    assign outputs[806] = layer0_outputs[1251];
    assign outputs[807] = ~(layer0_outputs[830]);
    assign outputs[808] = ~((layer0_outputs[1559]) | (layer0_outputs[653]));
    assign outputs[809] = (layer0_outputs[3162]) & ~(layer0_outputs[714]);
    assign outputs[810] = ~((layer0_outputs[3942]) ^ (layer0_outputs[4183]));
    assign outputs[811] = ~((layer0_outputs[4375]) | (layer0_outputs[2026]));
    assign outputs[812] = ~((layer0_outputs[1093]) | (layer0_outputs[1336]));
    assign outputs[813] = (layer0_outputs[29]) & ~(layer0_outputs[3997]);
    assign outputs[814] = (layer0_outputs[4773]) & ~(layer0_outputs[3361]);
    assign outputs[815] = (layer0_outputs[2019]) & ~(layer0_outputs[3294]);
    assign outputs[816] = ~((layer0_outputs[5022]) | (layer0_outputs[2685]));
    assign outputs[817] = (layer0_outputs[3300]) & (layer0_outputs[3052]);
    assign outputs[818] = ~((layer0_outputs[1736]) | (layer0_outputs[4595]));
    assign outputs[819] = (layer0_outputs[687]) & ~(layer0_outputs[1293]);
    assign outputs[820] = (layer0_outputs[1417]) & ~(layer0_outputs[499]);
    assign outputs[821] = ~((layer0_outputs[2655]) ^ (layer0_outputs[3013]));
    assign outputs[822] = ~((layer0_outputs[3139]) | (layer0_outputs[1306]));
    assign outputs[823] = (layer0_outputs[2985]) & (layer0_outputs[3359]);
    assign outputs[824] = (layer0_outputs[2872]) ^ (layer0_outputs[3652]);
    assign outputs[825] = (layer0_outputs[3701]) & ~(layer0_outputs[2633]);
    assign outputs[826] = ~(layer0_outputs[2738]);
    assign outputs[827] = ~((layer0_outputs[4988]) | (layer0_outputs[2947]));
    assign outputs[828] = (layer0_outputs[949]) & (layer0_outputs[2712]);
    assign outputs[829] = ~(layer0_outputs[4432]);
    assign outputs[830] = (layer0_outputs[3797]) & ~(layer0_outputs[2874]);
    assign outputs[831] = layer0_outputs[2923];
    assign outputs[832] = layer0_outputs[4242];
    assign outputs[833] = ~((layer0_outputs[4318]) ^ (layer0_outputs[3163]));
    assign outputs[834] = (layer0_outputs[4142]) & ~(layer0_outputs[4285]);
    assign outputs[835] = ~(layer0_outputs[245]);
    assign outputs[836] = ~((layer0_outputs[943]) | (layer0_outputs[4600]));
    assign outputs[837] = (layer0_outputs[3620]) & (layer0_outputs[185]);
    assign outputs[838] = (layer0_outputs[2700]) & (layer0_outputs[2143]);
    assign outputs[839] = ~(layer0_outputs[3392]);
    assign outputs[840] = ~((layer0_outputs[2284]) ^ (layer0_outputs[745]));
    assign outputs[841] = ~((layer0_outputs[4679]) | (layer0_outputs[1129]));
    assign outputs[842] = (layer0_outputs[1688]) & ~(layer0_outputs[5054]);
    assign outputs[843] = (layer0_outputs[854]) & (layer0_outputs[1482]);
    assign outputs[844] = (layer0_outputs[2624]) & ~(layer0_outputs[3801]);
    assign outputs[845] = (layer0_outputs[1628]) & ~(layer0_outputs[2706]);
    assign outputs[846] = ~(layer0_outputs[1496]);
    assign outputs[847] = (layer0_outputs[4106]) & (layer0_outputs[2847]);
    assign outputs[848] = (layer0_outputs[1294]) & ~(layer0_outputs[4725]);
    assign outputs[849] = layer0_outputs[2412];
    assign outputs[850] = ~((layer0_outputs[3216]) | (layer0_outputs[4834]));
    assign outputs[851] = (layer0_outputs[1986]) ^ (layer0_outputs[258]);
    assign outputs[852] = layer0_outputs[3861];
    assign outputs[853] = ~(layer0_outputs[4903]);
    assign outputs[854] = ~(layer0_outputs[154]) | (layer0_outputs[3436]);
    assign outputs[855] = ~(layer0_outputs[52]);
    assign outputs[856] = ~((layer0_outputs[3384]) | (layer0_outputs[2154]));
    assign outputs[857] = layer0_outputs[3062];
    assign outputs[858] = (layer0_outputs[655]) ^ (layer0_outputs[4216]);
    assign outputs[859] = layer0_outputs[2017];
    assign outputs[860] = (layer0_outputs[2991]) & ~(layer0_outputs[4529]);
    assign outputs[861] = ~((layer0_outputs[327]) | (layer0_outputs[3476]));
    assign outputs[862] = (layer0_outputs[194]) & (layer0_outputs[4889]);
    assign outputs[863] = ~(layer0_outputs[4490]);
    assign outputs[864] = (layer0_outputs[2764]) & ~(layer0_outputs[1269]);
    assign outputs[865] = (layer0_outputs[769]) & ~(layer0_outputs[2036]);
    assign outputs[866] = ~((layer0_outputs[2482]) | (layer0_outputs[2015]));
    assign outputs[867] = ~((layer0_outputs[2171]) | (layer0_outputs[1293]));
    assign outputs[868] = layer0_outputs[3655];
    assign outputs[869] = ~((layer0_outputs[3055]) ^ (layer0_outputs[1665]));
    assign outputs[870] = ~((layer0_outputs[4746]) | (layer0_outputs[950]));
    assign outputs[871] = ~((layer0_outputs[4595]) | (layer0_outputs[3108]));
    assign outputs[872] = (layer0_outputs[3077]) & ~(layer0_outputs[2569]);
    assign outputs[873] = (layer0_outputs[3314]) & ~(layer0_outputs[2648]);
    assign outputs[874] = (layer0_outputs[3473]) & ~(layer0_outputs[1776]);
    assign outputs[875] = (layer0_outputs[3791]) & ~(layer0_outputs[777]);
    assign outputs[876] = ~((layer0_outputs[1400]) | (layer0_outputs[2068]));
    assign outputs[877] = (layer0_outputs[5058]) & (layer0_outputs[987]);
    assign outputs[878] = layer0_outputs[2390];
    assign outputs[879] = ~(layer0_outputs[794]);
    assign outputs[880] = ~((layer0_outputs[1551]) | (layer0_outputs[2363]));
    assign outputs[881] = (layer0_outputs[3644]) & ~(layer0_outputs[1755]);
    assign outputs[882] = (layer0_outputs[213]) & (layer0_outputs[4960]);
    assign outputs[883] = ~((layer0_outputs[4635]) | (layer0_outputs[4372]));
    assign outputs[884] = (layer0_outputs[212]) & (layer0_outputs[1797]);
    assign outputs[885] = (layer0_outputs[2812]) & (layer0_outputs[1557]);
    assign outputs[886] = ~((layer0_outputs[2528]) | (layer0_outputs[319]));
    assign outputs[887] = (layer0_outputs[111]) & (layer0_outputs[4110]);
    assign outputs[888] = layer0_outputs[178];
    assign outputs[889] = (layer0_outputs[1590]) & ~(layer0_outputs[4681]);
    assign outputs[890] = (layer0_outputs[4343]) & ~(layer0_outputs[4198]);
    assign outputs[891] = ~((layer0_outputs[17]) | (layer0_outputs[3972]));
    assign outputs[892] = layer0_outputs[3769];
    assign outputs[893] = layer0_outputs[2442];
    assign outputs[894] = (layer0_outputs[4182]) & (layer0_outputs[1053]);
    assign outputs[895] = layer0_outputs[4191];
    assign outputs[896] = ~(layer0_outputs[2607]) | (layer0_outputs[3158]);
    assign outputs[897] = (layer0_outputs[4050]) & ~(layer0_outputs[2368]);
    assign outputs[898] = ~(layer0_outputs[4240]);
    assign outputs[899] = (layer0_outputs[792]) & (layer0_outputs[3993]);
    assign outputs[900] = ~((layer0_outputs[2191]) | (layer0_outputs[4185]));
    assign outputs[901] = layer0_outputs[3636];
    assign outputs[902] = (layer0_outputs[5006]) & ~(layer0_outputs[3816]);
    assign outputs[903] = layer0_outputs[3989];
    assign outputs[904] = (layer0_outputs[1965]) & ~(layer0_outputs[2274]);
    assign outputs[905] = ~((layer0_outputs[4957]) | (layer0_outputs[1841]));
    assign outputs[906] = (layer0_outputs[2088]) & ~(layer0_outputs[1042]);
    assign outputs[907] = (layer0_outputs[372]) & ~(layer0_outputs[1771]);
    assign outputs[908] = (layer0_outputs[1338]) & (layer0_outputs[3012]);
    assign outputs[909] = ~(layer0_outputs[2557]);
    assign outputs[910] = ~(layer0_outputs[805]);
    assign outputs[911] = ~(layer0_outputs[3767]);
    assign outputs[912] = ~((layer0_outputs[524]) | (layer0_outputs[2214]));
    assign outputs[913] = ~(layer0_outputs[4133]) | (layer0_outputs[5037]);
    assign outputs[914] = 1'b0;
    assign outputs[915] = (layer0_outputs[2284]) & ~(layer0_outputs[3071]);
    assign outputs[916] = ~((layer0_outputs[4355]) | (layer0_outputs[1105]));
    assign outputs[917] = ~((layer0_outputs[329]) ^ (layer0_outputs[1664]));
    assign outputs[918] = layer0_outputs[4416];
    assign outputs[919] = (layer0_outputs[2495]) & ~(layer0_outputs[2403]);
    assign outputs[920] = ~(layer0_outputs[762]);
    assign outputs[921] = (layer0_outputs[4774]) & ~(layer0_outputs[1925]);
    assign outputs[922] = ~(layer0_outputs[2757]);
    assign outputs[923] = ~((layer0_outputs[3539]) | (layer0_outputs[3842]));
    assign outputs[924] = layer0_outputs[1267];
    assign outputs[925] = (layer0_outputs[2518]) ^ (layer0_outputs[3834]);
    assign outputs[926] = ~((layer0_outputs[4091]) | (layer0_outputs[2148]));
    assign outputs[927] = ~(layer0_outputs[1213]);
    assign outputs[928] = layer0_outputs[2057];
    assign outputs[929] = (layer0_outputs[4381]) & (layer0_outputs[1752]);
    assign outputs[930] = layer0_outputs[2884];
    assign outputs[931] = (layer0_outputs[3207]) & (layer0_outputs[4908]);
    assign outputs[932] = (layer0_outputs[3448]) & (layer0_outputs[1765]);
    assign outputs[933] = (layer0_outputs[3034]) & ~(layer0_outputs[4944]);
    assign outputs[934] = ~((layer0_outputs[668]) ^ (layer0_outputs[570]));
    assign outputs[935] = (layer0_outputs[4500]) & ~(layer0_outputs[1648]);
    assign outputs[936] = ~((layer0_outputs[2026]) | (layer0_outputs[1948]));
    assign outputs[937] = ~(layer0_outputs[2171]) | (layer0_outputs[4126]);
    assign outputs[938] = layer0_outputs[1796];
    assign outputs[939] = layer0_outputs[2237];
    assign outputs[940] = layer0_outputs[2054];
    assign outputs[941] = layer0_outputs[983];
    assign outputs[942] = (layer0_outputs[2051]) & (layer0_outputs[743]);
    assign outputs[943] = (layer0_outputs[3243]) & ~(layer0_outputs[570]);
    assign outputs[944] = ~((layer0_outputs[4645]) | (layer0_outputs[956]));
    assign outputs[945] = layer0_outputs[4302];
    assign outputs[946] = (layer0_outputs[3241]) & (layer0_outputs[4268]);
    assign outputs[947] = ~((layer0_outputs[434]) ^ (layer0_outputs[390]));
    assign outputs[948] = (layer0_outputs[2239]) & ~(layer0_outputs[4760]);
    assign outputs[949] = ~(layer0_outputs[1079]);
    assign outputs[950] = (layer0_outputs[299]) & ~(layer0_outputs[2154]);
    assign outputs[951] = (layer0_outputs[4494]) & ~(layer0_outputs[1625]);
    assign outputs[952] = ~(layer0_outputs[4851]) | (layer0_outputs[1323]);
    assign outputs[953] = ~(layer0_outputs[2992]);
    assign outputs[954] = layer0_outputs[4229];
    assign outputs[955] = ~((layer0_outputs[1737]) ^ (layer0_outputs[1421]));
    assign outputs[956] = (layer0_outputs[2271]) & ~(layer0_outputs[2524]);
    assign outputs[957] = (layer0_outputs[2505]) & (layer0_outputs[4742]);
    assign outputs[958] = (layer0_outputs[2493]) ^ (layer0_outputs[2526]);
    assign outputs[959] = (layer0_outputs[2713]) & ~(layer0_outputs[5115]);
    assign outputs[960] = (layer0_outputs[2226]) & (layer0_outputs[4428]);
    assign outputs[961] = (layer0_outputs[985]) ^ (layer0_outputs[164]);
    assign outputs[962] = ~(layer0_outputs[145]);
    assign outputs[963] = (layer0_outputs[3701]) & ~(layer0_outputs[3238]);
    assign outputs[964] = (layer0_outputs[608]) & ~(layer0_outputs[1690]);
    assign outputs[965] = (layer0_outputs[2598]) & (layer0_outputs[965]);
    assign outputs[966] = ~((layer0_outputs[3240]) | (layer0_outputs[1308]));
    assign outputs[967] = ~(layer0_outputs[4746]);
    assign outputs[968] = ~((layer0_outputs[2996]) | (layer0_outputs[2588]));
    assign outputs[969] = (layer0_outputs[1211]) & ~(layer0_outputs[3345]);
    assign outputs[970] = ~(layer0_outputs[3174]);
    assign outputs[971] = (layer0_outputs[2856]) & (layer0_outputs[3977]);
    assign outputs[972] = (layer0_outputs[507]) & (layer0_outputs[3859]);
    assign outputs[973] = ~((layer0_outputs[2958]) ^ (layer0_outputs[907]));
    assign outputs[974] = layer0_outputs[2047];
    assign outputs[975] = ~(layer0_outputs[3654]);
    assign outputs[976] = layer0_outputs[1946];
    assign outputs[977] = ~((layer0_outputs[4594]) ^ (layer0_outputs[4703]));
    assign outputs[978] = ~(layer0_outputs[4498]);
    assign outputs[979] = (layer0_outputs[2426]) & ~(layer0_outputs[3632]);
    assign outputs[980] = (layer0_outputs[1950]) & ~(layer0_outputs[4292]);
    assign outputs[981] = ~(layer0_outputs[2375]);
    assign outputs[982] = (layer0_outputs[3810]) & (layer0_outputs[2027]);
    assign outputs[983] = ~((layer0_outputs[3295]) | (layer0_outputs[3715]));
    assign outputs[984] = ~((layer0_outputs[2090]) ^ (layer0_outputs[2080]));
    assign outputs[985] = (layer0_outputs[3002]) & (layer0_outputs[277]);
    assign outputs[986] = (layer0_outputs[698]) & ~(layer0_outputs[411]);
    assign outputs[987] = layer0_outputs[2372];
    assign outputs[988] = ~((layer0_outputs[2322]) | (layer0_outputs[35]));
    assign outputs[989] = (layer0_outputs[1585]) & ~(layer0_outputs[3333]);
    assign outputs[990] = ~(layer0_outputs[552]);
    assign outputs[991] = (layer0_outputs[1210]) & ~(layer0_outputs[4196]);
    assign outputs[992] = ~((layer0_outputs[664]) | (layer0_outputs[2053]));
    assign outputs[993] = (layer0_outputs[44]) & ~(layer0_outputs[4798]);
    assign outputs[994] = ~((layer0_outputs[266]) | (layer0_outputs[4662]));
    assign outputs[995] = ~(layer0_outputs[2134]);
    assign outputs[996] = ~(layer0_outputs[1806]);
    assign outputs[997] = (layer0_outputs[1215]) & ~(layer0_outputs[3852]);
    assign outputs[998] = ~(layer0_outputs[2481]);
    assign outputs[999] = (layer0_outputs[2436]) & (layer0_outputs[3359]);
    assign outputs[1000] = (layer0_outputs[1918]) ^ (layer0_outputs[1385]);
    assign outputs[1001] = (layer0_outputs[2314]) & (layer0_outputs[4880]);
    assign outputs[1002] = layer0_outputs[358];
    assign outputs[1003] = (layer0_outputs[1352]) & (layer0_outputs[862]);
    assign outputs[1004] = ~(layer0_outputs[151]);
    assign outputs[1005] = (layer0_outputs[406]) & ~(layer0_outputs[5011]);
    assign outputs[1006] = layer0_outputs[4176];
    assign outputs[1007] = (layer0_outputs[2616]) & ~(layer0_outputs[4308]);
    assign outputs[1008] = (layer0_outputs[1240]) & ~(layer0_outputs[1847]);
    assign outputs[1009] = (layer0_outputs[5040]) ^ (layer0_outputs[2201]);
    assign outputs[1010] = ~((layer0_outputs[4870]) ^ (layer0_outputs[1657]));
    assign outputs[1011] = ~(layer0_outputs[1031]);
    assign outputs[1012] = ~((layer0_outputs[2421]) | (layer0_outputs[585]));
    assign outputs[1013] = 1'b0;
    assign outputs[1014] = (layer0_outputs[4150]) & (layer0_outputs[4891]);
    assign outputs[1015] = (layer0_outputs[2161]) & ~(layer0_outputs[63]);
    assign outputs[1016] = layer0_outputs[4116];
    assign outputs[1017] = layer0_outputs[1272];
    assign outputs[1018] = (layer0_outputs[1202]) | (layer0_outputs[275]);
    assign outputs[1019] = (layer0_outputs[4619]) & (layer0_outputs[539]);
    assign outputs[1020] = ~(layer0_outputs[3960]);
    assign outputs[1021] = ~((layer0_outputs[1369]) | (layer0_outputs[190]));
    assign outputs[1022] = (layer0_outputs[3053]) & ~(layer0_outputs[1050]);
    assign outputs[1023] = ~(layer0_outputs[2247]);
    assign outputs[1024] = ~(layer0_outputs[2522]) | (layer0_outputs[1783]);
    assign outputs[1025] = ~((layer0_outputs[1853]) ^ (layer0_outputs[4259]));
    assign outputs[1026] = ~(layer0_outputs[258]);
    assign outputs[1027] = ~((layer0_outputs[2120]) | (layer0_outputs[3832]));
    assign outputs[1028] = layer0_outputs[1175];
    assign outputs[1029] = ~(layer0_outputs[4363]) | (layer0_outputs[3065]);
    assign outputs[1030] = ~(layer0_outputs[3433]);
    assign outputs[1031] = ~(layer0_outputs[324]);
    assign outputs[1032] = ~(layer0_outputs[510]);
    assign outputs[1033] = layer0_outputs[1118];
    assign outputs[1034] = layer0_outputs[4115];
    assign outputs[1035] = ~(layer0_outputs[1117]) | (layer0_outputs[4888]);
    assign outputs[1036] = ~(layer0_outputs[1171]) | (layer0_outputs[2654]);
    assign outputs[1037] = ~(layer0_outputs[4250]) | (layer0_outputs[1486]);
    assign outputs[1038] = ~(layer0_outputs[2203]) | (layer0_outputs[2245]);
    assign outputs[1039] = (layer0_outputs[3223]) | (layer0_outputs[345]);
    assign outputs[1040] = ~((layer0_outputs[2680]) & (layer0_outputs[878]));
    assign outputs[1041] = (layer0_outputs[2568]) ^ (layer0_outputs[2491]);
    assign outputs[1042] = (layer0_outputs[2740]) & ~(layer0_outputs[4959]);
    assign outputs[1043] = ~((layer0_outputs[54]) & (layer0_outputs[1030]));
    assign outputs[1044] = ~((layer0_outputs[1622]) ^ (layer0_outputs[2832]));
    assign outputs[1045] = ~(layer0_outputs[4637]);
    assign outputs[1046] = ~(layer0_outputs[3748]);
    assign outputs[1047] = layer0_outputs[3485];
    assign outputs[1048] = ~((layer0_outputs[3168]) ^ (layer0_outputs[989]));
    assign outputs[1049] = layer0_outputs[2356];
    assign outputs[1050] = (layer0_outputs[1571]) ^ (layer0_outputs[1179]);
    assign outputs[1051] = (layer0_outputs[3568]) ^ (layer0_outputs[4]);
    assign outputs[1052] = ~((layer0_outputs[2542]) ^ (layer0_outputs[2099]));
    assign outputs[1053] = ~(layer0_outputs[1000]);
    assign outputs[1054] = ~(layer0_outputs[3150]);
    assign outputs[1055] = ~((layer0_outputs[3177]) ^ (layer0_outputs[1627]));
    assign outputs[1056] = (layer0_outputs[777]) & ~(layer0_outputs[564]);
    assign outputs[1057] = layer0_outputs[2228];
    assign outputs[1058] = (layer0_outputs[3027]) | (layer0_outputs[823]);
    assign outputs[1059] = ~(layer0_outputs[1445]);
    assign outputs[1060] = (layer0_outputs[4314]) ^ (layer0_outputs[2690]);
    assign outputs[1061] = layer0_outputs[1373];
    assign outputs[1062] = layer0_outputs[4222];
    assign outputs[1063] = ~(layer0_outputs[2681]) | (layer0_outputs[3784]);
    assign outputs[1064] = layer0_outputs[2698];
    assign outputs[1065] = layer0_outputs[5099];
    assign outputs[1066] = (layer0_outputs[3949]) & ~(layer0_outputs[2541]);
    assign outputs[1067] = layer0_outputs[4451];
    assign outputs[1068] = (layer0_outputs[1824]) | (layer0_outputs[4514]);
    assign outputs[1069] = ~(layer0_outputs[2094]);
    assign outputs[1070] = (layer0_outputs[593]) ^ (layer0_outputs[2957]);
    assign outputs[1071] = ~((layer0_outputs[4632]) | (layer0_outputs[1178]));
    assign outputs[1072] = (layer0_outputs[2880]) & (layer0_outputs[3605]);
    assign outputs[1073] = ~(layer0_outputs[730]) | (layer0_outputs[2625]);
    assign outputs[1074] = ~(layer0_outputs[4408]);
    assign outputs[1075] = layer0_outputs[2758];
    assign outputs[1076] = ~(layer0_outputs[213]);
    assign outputs[1077] = ~(layer0_outputs[2211]);
    assign outputs[1078] = ~(layer0_outputs[3182]);
    assign outputs[1079] = ~(layer0_outputs[1843]);
    assign outputs[1080] = ~((layer0_outputs[1248]) ^ (layer0_outputs[4303]));
    assign outputs[1081] = (layer0_outputs[5059]) & ~(layer0_outputs[133]);
    assign outputs[1082] = ~(layer0_outputs[1978]) | (layer0_outputs[636]);
    assign outputs[1083] = layer0_outputs[187];
    assign outputs[1084] = (layer0_outputs[1661]) & ~(layer0_outputs[3729]);
    assign outputs[1085] = ~(layer0_outputs[30]);
    assign outputs[1086] = layer0_outputs[4993];
    assign outputs[1087] = ~(layer0_outputs[3843]);
    assign outputs[1088] = ~((layer0_outputs[2919]) ^ (layer0_outputs[4702]));
    assign outputs[1089] = ~(layer0_outputs[3609]);
    assign outputs[1090] = layer0_outputs[1924];
    assign outputs[1091] = ~(layer0_outputs[4653]) | (layer0_outputs[409]);
    assign outputs[1092] = layer0_outputs[3649];
    assign outputs[1093] = ~(layer0_outputs[3144]);
    assign outputs[1094] = (layer0_outputs[5109]) & ~(layer0_outputs[1003]);
    assign outputs[1095] = ~(layer0_outputs[3095]) | (layer0_outputs[117]);
    assign outputs[1096] = layer0_outputs[935];
    assign outputs[1097] = ~(layer0_outputs[4307]);
    assign outputs[1098] = (layer0_outputs[574]) ^ (layer0_outputs[505]);
    assign outputs[1099] = ~((layer0_outputs[359]) ^ (layer0_outputs[3978]));
    assign outputs[1100] = ~(layer0_outputs[4131]) | (layer0_outputs[4229]);
    assign outputs[1101] = ~(layer0_outputs[3344]);
    assign outputs[1102] = ~((layer0_outputs[1168]) | (layer0_outputs[2165]));
    assign outputs[1103] = (layer0_outputs[3993]) | (layer0_outputs[4539]);
    assign outputs[1104] = layer0_outputs[1148];
    assign outputs[1105] = ~((layer0_outputs[1937]) & (layer0_outputs[2938]));
    assign outputs[1106] = layer0_outputs[1348];
    assign outputs[1107] = layer0_outputs[1545];
    assign outputs[1108] = ~(layer0_outputs[4669]);
    assign outputs[1109] = (layer0_outputs[507]) ^ (layer0_outputs[4301]);
    assign outputs[1110] = ~(layer0_outputs[2861]) | (layer0_outputs[437]);
    assign outputs[1111] = ~(layer0_outputs[3197]) | (layer0_outputs[975]);
    assign outputs[1112] = layer0_outputs[3559];
    assign outputs[1113] = ~((layer0_outputs[2112]) & (layer0_outputs[2144]));
    assign outputs[1114] = (layer0_outputs[272]) & ~(layer0_outputs[1662]);
    assign outputs[1115] = ~(layer0_outputs[4971]);
    assign outputs[1116] = ~(layer0_outputs[4550]);
    assign outputs[1117] = ~(layer0_outputs[1641]);
    assign outputs[1118] = ~(layer0_outputs[654]);
    assign outputs[1119] = ~(layer0_outputs[4218]);
    assign outputs[1120] = (layer0_outputs[2574]) & ~(layer0_outputs[742]);
    assign outputs[1121] = ~(layer0_outputs[3350]);
    assign outputs[1122] = ~(layer0_outputs[840]);
    assign outputs[1123] = (layer0_outputs[2232]) | (layer0_outputs[5092]);
    assign outputs[1124] = ~(layer0_outputs[931]);
    assign outputs[1125] = ~((layer0_outputs[381]) | (layer0_outputs[2246]));
    assign outputs[1126] = ~(layer0_outputs[2985]) | (layer0_outputs[1761]);
    assign outputs[1127] = layer0_outputs[4592];
    assign outputs[1128] = ~(layer0_outputs[1835]) | (layer0_outputs[3110]);
    assign outputs[1129] = layer0_outputs[1636];
    assign outputs[1130] = (layer0_outputs[696]) | (layer0_outputs[3424]);
    assign outputs[1131] = ~(layer0_outputs[3679]);
    assign outputs[1132] = ~(layer0_outputs[2802]) | (layer0_outputs[4598]);
    assign outputs[1133] = (layer0_outputs[2544]) & ~(layer0_outputs[200]);
    assign outputs[1134] = ~((layer0_outputs[1168]) & (layer0_outputs[3562]));
    assign outputs[1135] = ~((layer0_outputs[4885]) ^ (layer0_outputs[1509]));
    assign outputs[1136] = layer0_outputs[5067];
    assign outputs[1137] = layer0_outputs[3802];
    assign outputs[1138] = (layer0_outputs[4569]) & ~(layer0_outputs[4925]);
    assign outputs[1139] = ~((layer0_outputs[4699]) ^ (layer0_outputs[1164]));
    assign outputs[1140] = layer0_outputs[4180];
    assign outputs[1141] = ~((layer0_outputs[1170]) ^ (layer0_outputs[1219]));
    assign outputs[1142] = ~(layer0_outputs[1781]) | (layer0_outputs[4236]);
    assign outputs[1143] = ~((layer0_outputs[1910]) ^ (layer0_outputs[3074]));
    assign outputs[1144] = ~(layer0_outputs[1098]);
    assign outputs[1145] = (layer0_outputs[3577]) & ~(layer0_outputs[2541]);
    assign outputs[1146] = ~(layer0_outputs[19]) | (layer0_outputs[4807]);
    assign outputs[1147] = (layer0_outputs[4734]) & (layer0_outputs[4581]);
    assign outputs[1148] = ~(layer0_outputs[2619]) | (layer0_outputs[1628]);
    assign outputs[1149] = ~(layer0_outputs[1892]);
    assign outputs[1150] = ~(layer0_outputs[1687]);
    assign outputs[1151] = ~(layer0_outputs[94]) | (layer0_outputs[275]);
    assign outputs[1152] = (layer0_outputs[3153]) | (layer0_outputs[2385]);
    assign outputs[1153] = layer0_outputs[1885];
    assign outputs[1154] = ~(layer0_outputs[1208]);
    assign outputs[1155] = layer0_outputs[2427];
    assign outputs[1156] = layer0_outputs[5037];
    assign outputs[1157] = layer0_outputs[4549];
    assign outputs[1158] = (layer0_outputs[1714]) ^ (layer0_outputs[1233]);
    assign outputs[1159] = (layer0_outputs[4999]) | (layer0_outputs[919]);
    assign outputs[1160] = ~((layer0_outputs[1484]) | (layer0_outputs[2840]));
    assign outputs[1161] = ~(layer0_outputs[4415]);
    assign outputs[1162] = (layer0_outputs[3204]) ^ (layer0_outputs[4597]);
    assign outputs[1163] = ~(layer0_outputs[204]) | (layer0_outputs[4246]);
    assign outputs[1164] = ~((layer0_outputs[4003]) & (layer0_outputs[1742]));
    assign outputs[1165] = layer0_outputs[2944];
    assign outputs[1166] = ~((layer0_outputs[842]) ^ (layer0_outputs[847]));
    assign outputs[1167] = ~(layer0_outputs[2989]);
    assign outputs[1168] = ~(layer0_outputs[984]) | (layer0_outputs[1452]);
    assign outputs[1169] = layer0_outputs[3046];
    assign outputs[1170] = ~(layer0_outputs[230]) | (layer0_outputs[4457]);
    assign outputs[1171] = ~(layer0_outputs[1284]);
    assign outputs[1172] = (layer0_outputs[4568]) & ~(layer0_outputs[3609]);
    assign outputs[1173] = ~(layer0_outputs[4219]);
    assign outputs[1174] = (layer0_outputs[788]) | (layer0_outputs[5077]);
    assign outputs[1175] = ~(layer0_outputs[5117]) | (layer0_outputs[1103]);
    assign outputs[1176] = (layer0_outputs[3671]) ^ (layer0_outputs[3103]);
    assign outputs[1177] = ~(layer0_outputs[2828]);
    assign outputs[1178] = ~(layer0_outputs[2186]);
    assign outputs[1179] = (layer0_outputs[1237]) & ~(layer0_outputs[2183]);
    assign outputs[1180] = (layer0_outputs[1783]) | (layer0_outputs[4991]);
    assign outputs[1181] = (layer0_outputs[2819]) ^ (layer0_outputs[3481]);
    assign outputs[1182] = (layer0_outputs[3680]) & (layer0_outputs[922]);
    assign outputs[1183] = (layer0_outputs[3421]) ^ (layer0_outputs[3720]);
    assign outputs[1184] = (layer0_outputs[4701]) ^ (layer0_outputs[3101]);
    assign outputs[1185] = (layer0_outputs[4641]) | (layer0_outputs[989]);
    assign outputs[1186] = layer0_outputs[4498];
    assign outputs[1187] = layer0_outputs[4679];
    assign outputs[1188] = ~(layer0_outputs[3958]) | (layer0_outputs[4359]);
    assign outputs[1189] = ~(layer0_outputs[3341]);
    assign outputs[1190] = ~(layer0_outputs[2627]);
    assign outputs[1191] = layer0_outputs[4873];
    assign outputs[1192] = (layer0_outputs[4238]) | (layer0_outputs[2525]);
    assign outputs[1193] = ~((layer0_outputs[3537]) | (layer0_outputs[3068]));
    assign outputs[1194] = layer0_outputs[1078];
    assign outputs[1195] = layer0_outputs[250];
    assign outputs[1196] = (layer0_outputs[4400]) & ~(layer0_outputs[4323]);
    assign outputs[1197] = ~(layer0_outputs[414]) | (layer0_outputs[4292]);
    assign outputs[1198] = layer0_outputs[958];
    assign outputs[1199] = ~(layer0_outputs[4420]);
    assign outputs[1200] = layer0_outputs[4715];
    assign outputs[1201] = ~(layer0_outputs[698]);
    assign outputs[1202] = ~((layer0_outputs[2842]) ^ (layer0_outputs[4946]));
    assign outputs[1203] = (layer0_outputs[2313]) ^ (layer0_outputs[2035]);
    assign outputs[1204] = ~(layer0_outputs[4276]);
    assign outputs[1205] = ~(layer0_outputs[3669]);
    assign outputs[1206] = ~((layer0_outputs[4574]) & (layer0_outputs[4093]));
    assign outputs[1207] = layer0_outputs[3286];
    assign outputs[1208] = layer0_outputs[571];
    assign outputs[1209] = ~((layer0_outputs[255]) & (layer0_outputs[1382]));
    assign outputs[1210] = ~(layer0_outputs[2762]) | (layer0_outputs[2169]);
    assign outputs[1211] = ~((layer0_outputs[978]) ^ (layer0_outputs[1936]));
    assign outputs[1212] = layer0_outputs[848];
    assign outputs[1213] = ~((layer0_outputs[4262]) ^ (layer0_outputs[1817]));
    assign outputs[1214] = (layer0_outputs[1768]) & (layer0_outputs[1308]);
    assign outputs[1215] = ~(layer0_outputs[1283]);
    assign outputs[1216] = ~(layer0_outputs[980]);
    assign outputs[1217] = (layer0_outputs[5102]) | (layer0_outputs[278]);
    assign outputs[1218] = ~(layer0_outputs[3571]) | (layer0_outputs[4158]);
    assign outputs[1219] = ~(layer0_outputs[3932]) | (layer0_outputs[2598]);
    assign outputs[1220] = (layer0_outputs[73]) ^ (layer0_outputs[515]);
    assign outputs[1221] = ~(layer0_outputs[3487]) | (layer0_outputs[5002]);
    assign outputs[1222] = layer0_outputs[2423];
    assign outputs[1223] = (layer0_outputs[2618]) & ~(layer0_outputs[2360]);
    assign outputs[1224] = ~(layer0_outputs[4704]);
    assign outputs[1225] = (layer0_outputs[280]) & (layer0_outputs[4032]);
    assign outputs[1226] = (layer0_outputs[1848]) | (layer0_outputs[1402]);
    assign outputs[1227] = ~(layer0_outputs[1755]) | (layer0_outputs[3691]);
    assign outputs[1228] = ~((layer0_outputs[878]) & (layer0_outputs[2319]));
    assign outputs[1229] = layer0_outputs[1430];
    assign outputs[1230] = ~(layer0_outputs[2207]);
    assign outputs[1231] = (layer0_outputs[902]) | (layer0_outputs[5110]);
    assign outputs[1232] = (layer0_outputs[2189]) & (layer0_outputs[2903]);
    assign outputs[1233] = ~(layer0_outputs[3734]) | (layer0_outputs[3596]);
    assign outputs[1234] = layer0_outputs[3236];
    assign outputs[1235] = layer0_outputs[4193];
    assign outputs[1236] = ~(layer0_outputs[3504]);
    assign outputs[1237] = (layer0_outputs[2455]) ^ (layer0_outputs[4302]);
    assign outputs[1238] = layer0_outputs[1345];
    assign outputs[1239] = ~(layer0_outputs[3974]) | (layer0_outputs[3293]);
    assign outputs[1240] = layer0_outputs[1065];
    assign outputs[1241] = ~(layer0_outputs[1507]);
    assign outputs[1242] = ~(layer0_outputs[1843]);
    assign outputs[1243] = ~(layer0_outputs[1170]) | (layer0_outputs[2149]);
    assign outputs[1244] = ~((layer0_outputs[3320]) ^ (layer0_outputs[1595]));
    assign outputs[1245] = (layer0_outputs[1672]) & ~(layer0_outputs[4868]);
    assign outputs[1246] = (layer0_outputs[1353]) ^ (layer0_outputs[502]);
    assign outputs[1247] = ~(layer0_outputs[4049]);
    assign outputs[1248] = (layer0_outputs[4456]) | (layer0_outputs[3482]);
    assign outputs[1249] = layer0_outputs[42];
    assign outputs[1250] = ~((layer0_outputs[3753]) | (layer0_outputs[995]));
    assign outputs[1251] = (layer0_outputs[1105]) | (layer0_outputs[3841]);
    assign outputs[1252] = layer0_outputs[3869];
    assign outputs[1253] = ~(layer0_outputs[3831]) | (layer0_outputs[602]);
    assign outputs[1254] = (layer0_outputs[3555]) & ~(layer0_outputs[404]);
    assign outputs[1255] = (layer0_outputs[912]) ^ (layer0_outputs[2756]);
    assign outputs[1256] = (layer0_outputs[1548]) ^ (layer0_outputs[4167]);
    assign outputs[1257] = (layer0_outputs[4277]) | (layer0_outputs[694]);
    assign outputs[1258] = layer0_outputs[2845];
    assign outputs[1259] = 1'b1;
    assign outputs[1260] = layer0_outputs[3316];
    assign outputs[1261] = ~(layer0_outputs[2200]);
    assign outputs[1262] = layer0_outputs[2679];
    assign outputs[1263] = layer0_outputs[2004];
    assign outputs[1264] = (layer0_outputs[2651]) ^ (layer0_outputs[2926]);
    assign outputs[1265] = ~((layer0_outputs[4979]) | (layer0_outputs[4300]));
    assign outputs[1266] = layer0_outputs[1294];
    assign outputs[1267] = ~(layer0_outputs[3098]);
    assign outputs[1268] = ~(layer0_outputs[2253]);
    assign outputs[1269] = layer0_outputs[3046];
    assign outputs[1270] = ~(layer0_outputs[1361]);
    assign outputs[1271] = layer0_outputs[2128];
    assign outputs[1272] = ~(layer0_outputs[736]) | (layer0_outputs[1858]);
    assign outputs[1273] = ~(layer0_outputs[2226]) | (layer0_outputs[1173]);
    assign outputs[1274] = (layer0_outputs[3251]) | (layer0_outputs[1062]);
    assign outputs[1275] = ~(layer0_outputs[488]);
    assign outputs[1276] = ~(layer0_outputs[3914]) | (layer0_outputs[5065]);
    assign outputs[1277] = ~(layer0_outputs[3342]);
    assign outputs[1278] = (layer0_outputs[3014]) ^ (layer0_outputs[4305]);
    assign outputs[1279] = ~((layer0_outputs[3665]) & (layer0_outputs[3382]));
    assign outputs[1280] = ~(layer0_outputs[3463]) | (layer0_outputs[1157]);
    assign outputs[1281] = (layer0_outputs[2608]) | (layer0_outputs[2514]);
    assign outputs[1282] = (layer0_outputs[3217]) | (layer0_outputs[3604]);
    assign outputs[1283] = ~(layer0_outputs[3821]) | (layer0_outputs[705]);
    assign outputs[1284] = (layer0_outputs[1036]) & (layer0_outputs[3525]);
    assign outputs[1285] = layer0_outputs[2564];
    assign outputs[1286] = layer0_outputs[696];
    assign outputs[1287] = ~((layer0_outputs[2001]) | (layer0_outputs[793]));
    assign outputs[1288] = layer0_outputs[1930];
    assign outputs[1289] = layer0_outputs[4084];
    assign outputs[1290] = layer0_outputs[2758];
    assign outputs[1291] = layer0_outputs[2327];
    assign outputs[1292] = ~(layer0_outputs[1622]) | (layer0_outputs[2064]);
    assign outputs[1293] = (layer0_outputs[4317]) ^ (layer0_outputs[4382]);
    assign outputs[1294] = ~(layer0_outputs[1241]) | (layer0_outputs[4856]);
    assign outputs[1295] = (layer0_outputs[1233]) & ~(layer0_outputs[4209]);
    assign outputs[1296] = ~((layer0_outputs[4358]) ^ (layer0_outputs[2901]));
    assign outputs[1297] = layer0_outputs[4443];
    assign outputs[1298] = ~(layer0_outputs[2005]);
    assign outputs[1299] = (layer0_outputs[2009]) | (layer0_outputs[3420]);
    assign outputs[1300] = layer0_outputs[1541];
    assign outputs[1301] = layer0_outputs[3371];
    assign outputs[1302] = (layer0_outputs[328]) ^ (layer0_outputs[637]);
    assign outputs[1303] = (layer0_outputs[1365]) | (layer0_outputs[2309]);
    assign outputs[1304] = ~(layer0_outputs[2490]);
    assign outputs[1305] = layer0_outputs[3580];
    assign outputs[1306] = (layer0_outputs[4104]) ^ (layer0_outputs[286]);
    assign outputs[1307] = (layer0_outputs[1379]) & (layer0_outputs[659]);
    assign outputs[1308] = (layer0_outputs[1281]) ^ (layer0_outputs[629]);
    assign outputs[1309] = (layer0_outputs[4682]) & ~(layer0_outputs[1305]);
    assign outputs[1310] = layer0_outputs[4296];
    assign outputs[1311] = (layer0_outputs[3206]) | (layer0_outputs[4969]);
    assign outputs[1312] = (layer0_outputs[675]) & (layer0_outputs[4910]);
    assign outputs[1313] = layer0_outputs[4865];
    assign outputs[1314] = ~(layer0_outputs[3237]);
    assign outputs[1315] = layer0_outputs[2073];
    assign outputs[1316] = layer0_outputs[1639];
    assign outputs[1317] = ~((layer0_outputs[2024]) & (layer0_outputs[2641]));
    assign outputs[1318] = (layer0_outputs[4106]) & ~(layer0_outputs[2508]);
    assign outputs[1319] = (layer0_outputs[4317]) ^ (layer0_outputs[2778]);
    assign outputs[1320] = layer0_outputs[1002];
    assign outputs[1321] = (layer0_outputs[3067]) ^ (layer0_outputs[751]);
    assign outputs[1322] = layer0_outputs[3455];
    assign outputs[1323] = ~(layer0_outputs[1483]);
    assign outputs[1324] = layer0_outputs[4398];
    assign outputs[1325] = layer0_outputs[4059];
    assign outputs[1326] = layer0_outputs[3102];
    assign outputs[1327] = (layer0_outputs[2614]) & ~(layer0_outputs[2363]);
    assign outputs[1328] = (layer0_outputs[4825]) & ~(layer0_outputs[1741]);
    assign outputs[1329] = layer0_outputs[3944];
    assign outputs[1330] = ~(layer0_outputs[1106]);
    assign outputs[1331] = ~(layer0_outputs[436]);
    assign outputs[1332] = ~(layer0_outputs[4823]) | (layer0_outputs[3424]);
    assign outputs[1333] = ~(layer0_outputs[3695]);
    assign outputs[1334] = ~(layer0_outputs[2785]);
    assign outputs[1335] = ~(layer0_outputs[1850]) | (layer0_outputs[596]);
    assign outputs[1336] = (layer0_outputs[3348]) & (layer0_outputs[2051]);
    assign outputs[1337] = (layer0_outputs[3157]) & ~(layer0_outputs[4986]);
    assign outputs[1338] = (layer0_outputs[4783]) & ~(layer0_outputs[1488]);
    assign outputs[1339] = layer0_outputs[4269];
    assign outputs[1340] = ~(layer0_outputs[4414]);
    assign outputs[1341] = ~(layer0_outputs[450]) | (layer0_outputs[2650]);
    assign outputs[1342] = (layer0_outputs[3348]) & ~(layer0_outputs[2986]);
    assign outputs[1343] = (layer0_outputs[3434]) & (layer0_outputs[3908]);
    assign outputs[1344] = ~(layer0_outputs[4268]);
    assign outputs[1345] = ~(layer0_outputs[3030]);
    assign outputs[1346] = layer0_outputs[173];
    assign outputs[1347] = (layer0_outputs[972]) ^ (layer0_outputs[4207]);
    assign outputs[1348] = ~(layer0_outputs[4329]);
    assign outputs[1349] = ~(layer0_outputs[205]);
    assign outputs[1350] = ~((layer0_outputs[3024]) ^ (layer0_outputs[4426]));
    assign outputs[1351] = ~(layer0_outputs[2192]);
    assign outputs[1352] = ~(layer0_outputs[1474]);
    assign outputs[1353] = layer0_outputs[157];
    assign outputs[1354] = ~((layer0_outputs[2185]) | (layer0_outputs[3120]));
    assign outputs[1355] = (layer0_outputs[4475]) & ~(layer0_outputs[1299]);
    assign outputs[1356] = ~(layer0_outputs[1309]) | (layer0_outputs[4456]);
    assign outputs[1357] = ~((layer0_outputs[757]) ^ (layer0_outputs[36]));
    assign outputs[1358] = ~((layer0_outputs[4043]) | (layer0_outputs[417]));
    assign outputs[1359] = ~(layer0_outputs[284]) | (layer0_outputs[5053]);
    assign outputs[1360] = layer0_outputs[300];
    assign outputs[1361] = layer0_outputs[4890];
    assign outputs[1362] = layer0_outputs[2070];
    assign outputs[1363] = ~(layer0_outputs[2115]);
    assign outputs[1364] = ~(layer0_outputs[2778]);
    assign outputs[1365] = layer0_outputs[326];
    assign outputs[1366] = ~(layer0_outputs[2866]) | (layer0_outputs[3744]);
    assign outputs[1367] = ~(layer0_outputs[2939]);
    assign outputs[1368] = ~(layer0_outputs[1177]) | (layer0_outputs[1897]);
    assign outputs[1369] = ~((layer0_outputs[4775]) ^ (layer0_outputs[3125]));
    assign outputs[1370] = ~((layer0_outputs[3484]) & (layer0_outputs[4714]));
    assign outputs[1371] = (layer0_outputs[4693]) & ~(layer0_outputs[1112]);
    assign outputs[1372] = ~(layer0_outputs[4179]);
    assign outputs[1373] = ~(layer0_outputs[2613]);
    assign outputs[1374] = ~(layer0_outputs[1049]) | (layer0_outputs[2454]);
    assign outputs[1375] = ~((layer0_outputs[346]) ^ (layer0_outputs[2749]));
    assign outputs[1376] = ~((layer0_outputs[4336]) & (layer0_outputs[5025]));
    assign outputs[1377] = ~(layer0_outputs[4880]);
    assign outputs[1378] = ~(layer0_outputs[2916]);
    assign outputs[1379] = ~(layer0_outputs[5097]);
    assign outputs[1380] = ~(layer0_outputs[4030]);
    assign outputs[1381] = layer0_outputs[2610];
    assign outputs[1382] = ~(layer0_outputs[3926]);
    assign outputs[1383] = (layer0_outputs[1629]) & (layer0_outputs[853]);
    assign outputs[1384] = (layer0_outputs[4489]) & ~(layer0_outputs[2800]);
    assign outputs[1385] = (layer0_outputs[3008]) & ~(layer0_outputs[3733]);
    assign outputs[1386] = layer0_outputs[2846];
    assign outputs[1387] = layer0_outputs[2944];
    assign outputs[1388] = ~(layer0_outputs[2190]);
    assign outputs[1389] = ~(layer0_outputs[472]);
    assign outputs[1390] = layer0_outputs[2462];
    assign outputs[1391] = (layer0_outputs[3460]) | (layer0_outputs[2065]);
    assign outputs[1392] = ~(layer0_outputs[3675]);
    assign outputs[1393] = ~(layer0_outputs[175]);
    assign outputs[1394] = ~(layer0_outputs[819]);
    assign outputs[1395] = layer0_outputs[1442];
    assign outputs[1396] = ~(layer0_outputs[632]);
    assign outputs[1397] = ~(layer0_outputs[753]);
    assign outputs[1398] = ~(layer0_outputs[1162]) | (layer0_outputs[5006]);
    assign outputs[1399] = layer0_outputs[4760];
    assign outputs[1400] = layer0_outputs[3065];
    assign outputs[1401] = 1'b1;
    assign outputs[1402] = (layer0_outputs[369]) ^ (layer0_outputs[1495]);
    assign outputs[1403] = ~(layer0_outputs[1310]);
    assign outputs[1404] = ~((layer0_outputs[2830]) | (layer0_outputs[4316]));
    assign outputs[1405] = ~(layer0_outputs[4508]);
    assign outputs[1406] = ~(layer0_outputs[1152]);
    assign outputs[1407] = (layer0_outputs[222]) ^ (layer0_outputs[1481]);
    assign outputs[1408] = (layer0_outputs[1103]) & ~(layer0_outputs[2414]);
    assign outputs[1409] = ~((layer0_outputs[3063]) & (layer0_outputs[4497]));
    assign outputs[1410] = ~((layer0_outputs[212]) & (layer0_outputs[1718]));
    assign outputs[1411] = layer0_outputs[3078];
    assign outputs[1412] = (layer0_outputs[11]) & ~(layer0_outputs[2212]);
    assign outputs[1413] = layer0_outputs[5118];
    assign outputs[1414] = layer0_outputs[1365];
    assign outputs[1415] = (layer0_outputs[3924]) ^ (layer0_outputs[4946]);
    assign outputs[1416] = ~(layer0_outputs[3111]) | (layer0_outputs[3451]);
    assign outputs[1417] = (layer0_outputs[3485]) & ~(layer0_outputs[3450]);
    assign outputs[1418] = (layer0_outputs[798]) & ~(layer0_outputs[2360]);
    assign outputs[1419] = layer0_outputs[107];
    assign outputs[1420] = ~(layer0_outputs[3169]);
    assign outputs[1421] = layer0_outputs[2129];
    assign outputs[1422] = ~((layer0_outputs[3266]) ^ (layer0_outputs[1341]));
    assign outputs[1423] = ~(layer0_outputs[4824]);
    assign outputs[1424] = ~(layer0_outputs[2973]) | (layer0_outputs[4870]);
    assign outputs[1425] = ~((layer0_outputs[4698]) ^ (layer0_outputs[760]));
    assign outputs[1426] = ~(layer0_outputs[2059]) | (layer0_outputs[441]);
    assign outputs[1427] = ~(layer0_outputs[758]);
    assign outputs[1428] = layer0_outputs[4295];
    assign outputs[1429] = ~((layer0_outputs[2312]) & (layer0_outputs[1882]));
    assign outputs[1430] = (layer0_outputs[1402]) | (layer0_outputs[2473]);
    assign outputs[1431] = (layer0_outputs[3599]) & (layer0_outputs[1967]);
    assign outputs[1432] = layer0_outputs[4127];
    assign outputs[1433] = (layer0_outputs[3286]) | (layer0_outputs[3916]);
    assign outputs[1434] = ~(layer0_outputs[2313]);
    assign outputs[1435] = layer0_outputs[3927];
    assign outputs[1436] = ~(layer0_outputs[567]);
    assign outputs[1437] = (layer0_outputs[2055]) & ~(layer0_outputs[728]);
    assign outputs[1438] = (layer0_outputs[3995]) & ~(layer0_outputs[341]);
    assign outputs[1439] = (layer0_outputs[643]) & ~(layer0_outputs[1311]);
    assign outputs[1440] = layer0_outputs[2364];
    assign outputs[1441] = ~(layer0_outputs[1912]);
    assign outputs[1442] = (layer0_outputs[3066]) & ~(layer0_outputs[793]);
    assign outputs[1443] = layer0_outputs[2514];
    assign outputs[1444] = ~((layer0_outputs[130]) | (layer0_outputs[3983]));
    assign outputs[1445] = ~(layer0_outputs[2943]) | (layer0_outputs[2066]);
    assign outputs[1446] = ~(layer0_outputs[617]) | (layer0_outputs[4814]);
    assign outputs[1447] = ~(layer0_outputs[4120]);
    assign outputs[1448] = (layer0_outputs[4758]) ^ (layer0_outputs[3714]);
    assign outputs[1449] = ~(layer0_outputs[1904]) | (layer0_outputs[3806]);
    assign outputs[1450] = (layer0_outputs[1821]) | (layer0_outputs[2270]);
    assign outputs[1451] = ~(layer0_outputs[2921]);
    assign outputs[1452] = layer0_outputs[2599];
    assign outputs[1453] = ~(layer0_outputs[3416]) | (layer0_outputs[5020]);
    assign outputs[1454] = layer0_outputs[914];
    assign outputs[1455] = ~(layer0_outputs[1490]) | (layer0_outputs[157]);
    assign outputs[1456] = ~(layer0_outputs[2299]) | (layer0_outputs[2278]);
    assign outputs[1457] = (layer0_outputs[4659]) ^ (layer0_outputs[1505]);
    assign outputs[1458] = ~(layer0_outputs[1663]);
    assign outputs[1459] = ~(layer0_outputs[2483]) | (layer0_outputs[3598]);
    assign outputs[1460] = layer0_outputs[1625];
    assign outputs[1461] = 1'b1;
    assign outputs[1462] = ~(layer0_outputs[3955]) | (layer0_outputs[2770]);
    assign outputs[1463] = ~(layer0_outputs[1470]);
    assign outputs[1464] = layer0_outputs[1673];
    assign outputs[1465] = ~((layer0_outputs[2685]) ^ (layer0_outputs[3114]));
    assign outputs[1466] = ~(layer0_outputs[4841]) | (layer0_outputs[4054]);
    assign outputs[1467] = layer0_outputs[125];
    assign outputs[1468] = layer0_outputs[5107];
    assign outputs[1469] = (layer0_outputs[760]) & (layer0_outputs[3752]);
    assign outputs[1470] = ~((layer0_outputs[4304]) ^ (layer0_outputs[4422]));
    assign outputs[1471] = layer0_outputs[1435];
    assign outputs[1472] = layer0_outputs[1200];
    assign outputs[1473] = layer0_outputs[2769];
    assign outputs[1474] = (layer0_outputs[4305]) ^ (layer0_outputs[4749]);
    assign outputs[1475] = (layer0_outputs[2485]) & ~(layer0_outputs[3756]);
    assign outputs[1476] = ~((layer0_outputs[23]) & (layer0_outputs[1839]));
    assign outputs[1477] = ~(layer0_outputs[3573]);
    assign outputs[1478] = ~((layer0_outputs[4615]) | (layer0_outputs[2765]));
    assign outputs[1479] = (layer0_outputs[214]) & ~(layer0_outputs[976]);
    assign outputs[1480] = (layer0_outputs[589]) | (layer0_outputs[3136]);
    assign outputs[1481] = (layer0_outputs[2405]) | (layer0_outputs[4264]);
    assign outputs[1482] = ~((layer0_outputs[2630]) & (layer0_outputs[3068]));
    assign outputs[1483] = ~((layer0_outputs[2351]) & (layer0_outputs[4757]));
    assign outputs[1484] = ~(layer0_outputs[1133]);
    assign outputs[1485] = ~(layer0_outputs[3084]);
    assign outputs[1486] = ~((layer0_outputs[3858]) | (layer0_outputs[4580]));
    assign outputs[1487] = layer0_outputs[4710];
    assign outputs[1488] = ~(layer0_outputs[3350]);
    assign outputs[1489] = ~((layer0_outputs[1959]) & (layer0_outputs[489]));
    assign outputs[1490] = layer0_outputs[814];
    assign outputs[1491] = layer0_outputs[4252];
    assign outputs[1492] = (layer0_outputs[4280]) ^ (layer0_outputs[1891]);
    assign outputs[1493] = ~(layer0_outputs[1587]);
    assign outputs[1494] = ~(layer0_outputs[3773]);
    assign outputs[1495] = (layer0_outputs[3636]) ^ (layer0_outputs[152]);
    assign outputs[1496] = ~(layer0_outputs[305]) | (layer0_outputs[1650]);
    assign outputs[1497] = ~(layer0_outputs[2434]);
    assign outputs[1498] = (layer0_outputs[1121]) ^ (layer0_outputs[3607]);
    assign outputs[1499] = ~(layer0_outputs[3572]);
    assign outputs[1500] = ~(layer0_outputs[2873]) | (layer0_outputs[4839]);
    assign outputs[1501] = (layer0_outputs[2834]) & (layer0_outputs[3889]);
    assign outputs[1502] = ~(layer0_outputs[2176]);
    assign outputs[1503] = layer0_outputs[4492];
    assign outputs[1504] = ~(layer0_outputs[1832]) | (layer0_outputs[827]);
    assign outputs[1505] = ~((layer0_outputs[3611]) | (layer0_outputs[1466]));
    assign outputs[1506] = ~(layer0_outputs[1263]);
    assign outputs[1507] = ~(layer0_outputs[21]) | (layer0_outputs[1113]);
    assign outputs[1508] = ~(layer0_outputs[395]);
    assign outputs[1509] = (layer0_outputs[4968]) ^ (layer0_outputs[1287]);
    assign outputs[1510] = ~(layer0_outputs[1604]);
    assign outputs[1511] = ~(layer0_outputs[3081]);
    assign outputs[1512] = ~((layer0_outputs[2823]) ^ (layer0_outputs[2372]));
    assign outputs[1513] = ~((layer0_outputs[2001]) | (layer0_outputs[2840]));
    assign outputs[1514] = ~((layer0_outputs[4956]) & (layer0_outputs[378]));
    assign outputs[1515] = ~(layer0_outputs[873]) | (layer0_outputs[5021]);
    assign outputs[1516] = ~(layer0_outputs[3344]) | (layer0_outputs[4781]);
    assign outputs[1517] = (layer0_outputs[3227]) | (layer0_outputs[3179]);
    assign outputs[1518] = ~((layer0_outputs[767]) | (layer0_outputs[4449]));
    assign outputs[1519] = (layer0_outputs[3697]) ^ (layer0_outputs[2804]);
    assign outputs[1520] = layer0_outputs[170];
    assign outputs[1521] = (layer0_outputs[2321]) & ~(layer0_outputs[85]);
    assign outputs[1522] = layer0_outputs[1759];
    assign outputs[1523] = (layer0_outputs[69]) ^ (layer0_outputs[2214]);
    assign outputs[1524] = (layer0_outputs[2263]) & (layer0_outputs[2337]);
    assign outputs[1525] = (layer0_outputs[4234]) & ~(layer0_outputs[3407]);
    assign outputs[1526] = ~((layer0_outputs[3964]) | (layer0_outputs[4099]));
    assign outputs[1527] = layer0_outputs[3647];
    assign outputs[1528] = ~(layer0_outputs[3394]);
    assign outputs[1529] = layer0_outputs[565];
    assign outputs[1530] = layer0_outputs[4208];
    assign outputs[1531] = (layer0_outputs[3644]) & ~(layer0_outputs[898]);
    assign outputs[1532] = layer0_outputs[554];
    assign outputs[1533] = layer0_outputs[2912];
    assign outputs[1534] = ~(layer0_outputs[1522]);
    assign outputs[1535] = (layer0_outputs[720]) & ~(layer0_outputs[2800]);
    assign outputs[1536] = ~(layer0_outputs[3435]);
    assign outputs[1537] = ~(layer0_outputs[4232]);
    assign outputs[1538] = layer0_outputs[2731];
    assign outputs[1539] = ~(layer0_outputs[3784]);
    assign outputs[1540] = (layer0_outputs[2755]) ^ (layer0_outputs[969]);
    assign outputs[1541] = (layer0_outputs[3672]) | (layer0_outputs[4192]);
    assign outputs[1542] = (layer0_outputs[867]) & ~(layer0_outputs[285]);
    assign outputs[1543] = ~(layer0_outputs[429]) | (layer0_outputs[1939]);
    assign outputs[1544] = ~(layer0_outputs[2748]);
    assign outputs[1545] = layer0_outputs[3893];
    assign outputs[1546] = layer0_outputs[3704];
    assign outputs[1547] = layer0_outputs[4378];
    assign outputs[1548] = ~(layer0_outputs[2855]) | (layer0_outputs[4503]);
    assign outputs[1549] = (layer0_outputs[3583]) ^ (layer0_outputs[317]);
    assign outputs[1550] = (layer0_outputs[4584]) | (layer0_outputs[3633]);
    assign outputs[1551] = (layer0_outputs[3897]) ^ (layer0_outputs[4066]);
    assign outputs[1552] = ~(layer0_outputs[3561]) | (layer0_outputs[1771]);
    assign outputs[1553] = ~(layer0_outputs[1319]);
    assign outputs[1554] = ~(layer0_outputs[543]) | (layer0_outputs[4874]);
    assign outputs[1555] = (layer0_outputs[74]) ^ (layer0_outputs[2254]);
    assign outputs[1556] = ~(layer0_outputs[4398]);
    assign outputs[1557] = (layer0_outputs[39]) & ~(layer0_outputs[3666]);
    assign outputs[1558] = (layer0_outputs[249]) & ~(layer0_outputs[2869]);
    assign outputs[1559] = ~(layer0_outputs[524]);
    assign outputs[1560] = layer0_outputs[3100];
    assign outputs[1561] = (layer0_outputs[4854]) & ~(layer0_outputs[4038]);
    assign outputs[1562] = ~(layer0_outputs[1167]);
    assign outputs[1563] = ~(layer0_outputs[2834]);
    assign outputs[1564] = (layer0_outputs[4502]) & ~(layer0_outputs[463]);
    assign outputs[1565] = ~(layer0_outputs[3365]);
    assign outputs[1566] = ~(layer0_outputs[1751]);
    assign outputs[1567] = layer0_outputs[4039];
    assign outputs[1568] = (layer0_outputs[3628]) ^ (layer0_outputs[1331]);
    assign outputs[1569] = ~(layer0_outputs[4689]) | (layer0_outputs[525]);
    assign outputs[1570] = ~(layer0_outputs[4666]);
    assign outputs[1571] = layer0_outputs[2721];
    assign outputs[1572] = (layer0_outputs[889]) ^ (layer0_outputs[2282]);
    assign outputs[1573] = ~(layer0_outputs[2028]);
    assign outputs[1574] = ~(layer0_outputs[2575]);
    assign outputs[1575] = (layer0_outputs[2919]) & (layer0_outputs[4670]);
    assign outputs[1576] = ~(layer0_outputs[4506]);
    assign outputs[1577] = (layer0_outputs[2195]) & (layer0_outputs[2198]);
    assign outputs[1578] = ~(layer0_outputs[3458]) | (layer0_outputs[2623]);
    assign outputs[1579] = (layer0_outputs[5048]) ^ (layer0_outputs[3643]);
    assign outputs[1580] = ~(layer0_outputs[80]);
    assign outputs[1581] = (layer0_outputs[1926]) ^ (layer0_outputs[336]);
    assign outputs[1582] = ~((layer0_outputs[392]) | (layer0_outputs[2318]));
    assign outputs[1583] = layer0_outputs[4740];
    assign outputs[1584] = (layer0_outputs[81]) ^ (layer0_outputs[390]);
    assign outputs[1585] = ~(layer0_outputs[2445]);
    assign outputs[1586] = ~((layer0_outputs[3871]) | (layer0_outputs[412]));
    assign outputs[1587] = ~(layer0_outputs[3906]) | (layer0_outputs[751]);
    assign outputs[1588] = ~(layer0_outputs[405]);
    assign outputs[1589] = (layer0_outputs[885]) & ~(layer0_outputs[4822]);
    assign outputs[1590] = layer0_outputs[3951];
    assign outputs[1591] = (layer0_outputs[3094]) & ~(layer0_outputs[2852]);
    assign outputs[1592] = layer0_outputs[1038];
    assign outputs[1593] = (layer0_outputs[3514]) & ~(layer0_outputs[4637]);
    assign outputs[1594] = ~(layer0_outputs[2437]);
    assign outputs[1595] = ~(layer0_outputs[2446]);
    assign outputs[1596] = layer0_outputs[3132];
    assign outputs[1597] = ~((layer0_outputs[388]) ^ (layer0_outputs[60]));
    assign outputs[1598] = layer0_outputs[3009];
    assign outputs[1599] = ~(layer0_outputs[5080]);
    assign outputs[1600] = (layer0_outputs[3423]) & ~(layer0_outputs[706]);
    assign outputs[1601] = ~(layer0_outputs[4089]) | (layer0_outputs[2577]);
    assign outputs[1602] = ~(layer0_outputs[4671]) | (layer0_outputs[4932]);
    assign outputs[1603] = layer0_outputs[3705];
    assign outputs[1604] = ~((layer0_outputs[868]) | (layer0_outputs[4809]));
    assign outputs[1605] = ~(layer0_outputs[3895]) | (layer0_outputs[4906]);
    assign outputs[1606] = ~(layer0_outputs[1584]);
    assign outputs[1607] = ~((layer0_outputs[2563]) ^ (layer0_outputs[259]));
    assign outputs[1608] = ~(layer0_outputs[1721]);
    assign outputs[1609] = ~(layer0_outputs[2202]) | (layer0_outputs[4499]);
    assign outputs[1610] = ~((layer0_outputs[4300]) ^ (layer0_outputs[2167]));
    assign outputs[1611] = (layer0_outputs[4347]) ^ (layer0_outputs[4454]);
    assign outputs[1612] = layer0_outputs[2660];
    assign outputs[1613] = ~((layer0_outputs[4022]) ^ (layer0_outputs[2927]));
    assign outputs[1614] = ~((layer0_outputs[1852]) ^ (layer0_outputs[2381]));
    assign outputs[1615] = (layer0_outputs[4676]) | (layer0_outputs[4917]);
    assign outputs[1616] = (layer0_outputs[4073]) & ~(layer0_outputs[144]);
    assign outputs[1617] = ~(layer0_outputs[2325]);
    assign outputs[1618] = (layer0_outputs[4366]) ^ (layer0_outputs[963]);
    assign outputs[1619] = layer0_outputs[1328];
    assign outputs[1620] = layer0_outputs[2090];
    assign outputs[1621] = layer0_outputs[3242];
    assign outputs[1622] = ~(layer0_outputs[2998]) | (layer0_outputs[2656]);
    assign outputs[1623] = layer0_outputs[2425];
    assign outputs[1624] = (layer0_outputs[5023]) ^ (layer0_outputs[4243]);
    assign outputs[1625] = ~(layer0_outputs[440]);
    assign outputs[1626] = ~(layer0_outputs[1740]);
    assign outputs[1627] = layer0_outputs[4776];
    assign outputs[1628] = ~(layer0_outputs[3147]);
    assign outputs[1629] = ~(layer0_outputs[1953]);
    assign outputs[1630] = ~(layer0_outputs[2279]);
    assign outputs[1631] = ~(layer0_outputs[3306]);
    assign outputs[1632] = (layer0_outputs[1132]) & (layer0_outputs[1201]);
    assign outputs[1633] = ~(layer0_outputs[2152]);
    assign outputs[1634] = ~(layer0_outputs[1138]);
    assign outputs[1635] = ~((layer0_outputs[2890]) & (layer0_outputs[2183]));
    assign outputs[1636] = ~(layer0_outputs[2549]) | (layer0_outputs[541]);
    assign outputs[1637] = (layer0_outputs[960]) & (layer0_outputs[1957]);
    assign outputs[1638] = (layer0_outputs[322]) & (layer0_outputs[50]);
    assign outputs[1639] = ~(layer0_outputs[1165]);
    assign outputs[1640] = ~(layer0_outputs[4432]) | (layer0_outputs[3601]);
    assign outputs[1641] = layer0_outputs[3754];
    assign outputs[1642] = ~((layer0_outputs[1041]) | (layer0_outputs[4423]));
    assign outputs[1643] = (layer0_outputs[2122]) & ~(layer0_outputs[2420]);
    assign outputs[1644] = ~(layer0_outputs[2862]) | (layer0_outputs[2386]);
    assign outputs[1645] = ~(layer0_outputs[3129]) | (layer0_outputs[3822]);
    assign outputs[1646] = ~(layer0_outputs[164]);
    assign outputs[1647] = ~((layer0_outputs[2437]) | (layer0_outputs[5014]));
    assign outputs[1648] = (layer0_outputs[332]) & (layer0_outputs[3551]);
    assign outputs[1649] = (layer0_outputs[3140]) | (layer0_outputs[2810]);
    assign outputs[1650] = ~(layer0_outputs[3466]);
    assign outputs[1651] = ~(layer0_outputs[3085]);
    assign outputs[1652] = layer0_outputs[1465];
    assign outputs[1653] = (layer0_outputs[1520]) & ~(layer0_outputs[3728]);
    assign outputs[1654] = layer0_outputs[4499];
    assign outputs[1655] = layer0_outputs[1649];
    assign outputs[1656] = (layer0_outputs[1109]) ^ (layer0_outputs[3301]);
    assign outputs[1657] = ~((layer0_outputs[3558]) | (layer0_outputs[1131]));
    assign outputs[1658] = ~((layer0_outputs[3106]) & (layer0_outputs[4672]));
    assign outputs[1659] = layer0_outputs[5087];
    assign outputs[1660] = ~(layer0_outputs[2575]);
    assign outputs[1661] = ~((layer0_outputs[2327]) & (layer0_outputs[2186]));
    assign outputs[1662] = (layer0_outputs[246]) & ~(layer0_outputs[1772]);
    assign outputs[1663] = layer0_outputs[1320];
    assign outputs[1664] = ~((layer0_outputs[3912]) & (layer0_outputs[1275]));
    assign outputs[1665] = ~((layer0_outputs[1176]) ^ (layer0_outputs[447]));
    assign outputs[1666] = ~(layer0_outputs[321]);
    assign outputs[1667] = (layer0_outputs[2430]) | (layer0_outputs[3677]);
    assign outputs[1668] = layer0_outputs[235];
    assign outputs[1669] = layer0_outputs[120];
    assign outputs[1670] = layer0_outputs[853];
    assign outputs[1671] = ~((layer0_outputs[1277]) & (layer0_outputs[4762]));
    assign outputs[1672] = ~(layer0_outputs[501]) | (layer0_outputs[3776]);
    assign outputs[1673] = ~(layer0_outputs[891]);
    assign outputs[1674] = ~(layer0_outputs[4947]);
    assign outputs[1675] = ~(layer0_outputs[1676]);
    assign outputs[1676] = (layer0_outputs[1679]) | (layer0_outputs[3220]);
    assign outputs[1677] = ~((layer0_outputs[1350]) & (layer0_outputs[2867]));
    assign outputs[1678] = (layer0_outputs[849]) & (layer0_outputs[4891]);
    assign outputs[1679] = 1'b1;
    assign outputs[1680] = (layer0_outputs[3947]) & ~(layer0_outputs[65]);
    assign outputs[1681] = (layer0_outputs[1230]) & (layer0_outputs[1968]);
    assign outputs[1682] = (layer0_outputs[3471]) ^ (layer0_outputs[4886]);
    assign outputs[1683] = (layer0_outputs[3180]) & ~(layer0_outputs[812]);
    assign outputs[1684] = ~(layer0_outputs[769]);
    assign outputs[1685] = (layer0_outputs[2727]) & (layer0_outputs[1959]);
    assign outputs[1686] = ~(layer0_outputs[297]);
    assign outputs[1687] = ~(layer0_outputs[2273]);
    assign outputs[1688] = ~((layer0_outputs[679]) ^ (layer0_outputs[4006]));
    assign outputs[1689] = ~((layer0_outputs[3178]) | (layer0_outputs[117]));
    assign outputs[1690] = ~(layer0_outputs[6]);
    assign outputs[1691] = (layer0_outputs[1459]) ^ (layer0_outputs[3145]);
    assign outputs[1692] = ~((layer0_outputs[2370]) ^ (layer0_outputs[2910]));
    assign outputs[1693] = (layer0_outputs[167]) & (layer0_outputs[4804]);
    assign outputs[1694] = ~(layer0_outputs[4610]);
    assign outputs[1695] = layer0_outputs[184];
    assign outputs[1696] = ~((layer0_outputs[5070]) ^ (layer0_outputs[3137]));
    assign outputs[1697] = (layer0_outputs[83]) ^ (layer0_outputs[49]);
    assign outputs[1698] = (layer0_outputs[406]) & ~(layer0_outputs[293]);
    assign outputs[1699] = layer0_outputs[1295];
    assign outputs[1700] = ~(layer0_outputs[1549]);
    assign outputs[1701] = ~((layer0_outputs[259]) | (layer0_outputs[3947]));
    assign outputs[1702] = ~(layer0_outputs[3272]);
    assign outputs[1703] = (layer0_outputs[1971]) & (layer0_outputs[2573]);
    assign outputs[1704] = ~(layer0_outputs[674]);
    assign outputs[1705] = ~((layer0_outputs[3663]) | (layer0_outputs[1927]));
    assign outputs[1706] = ~(layer0_outputs[1893]);
    assign outputs[1707] = ~(layer0_outputs[831]);
    assign outputs[1708] = (layer0_outputs[2853]) & (layer0_outputs[4815]);
    assign outputs[1709] = layer0_outputs[3964];
    assign outputs[1710] = ~((layer0_outputs[2918]) | (layer0_outputs[5050]));
    assign outputs[1711] = layer0_outputs[3069];
    assign outputs[1712] = ~((layer0_outputs[4665]) | (layer0_outputs[3477]));
    assign outputs[1713] = layer0_outputs[4906];
    assign outputs[1714] = (layer0_outputs[619]) ^ (layer0_outputs[784]);
    assign outputs[1715] = ~(layer0_outputs[4141]);
    assign outputs[1716] = (layer0_outputs[3269]) & (layer0_outputs[2024]);
    assign outputs[1717] = (layer0_outputs[1948]) | (layer0_outputs[2744]);
    assign outputs[1718] = (layer0_outputs[95]) & ~(layer0_outputs[2822]);
    assign outputs[1719] = (layer0_outputs[1851]) & ~(layer0_outputs[2336]);
    assign outputs[1720] = layer0_outputs[4831];
    assign outputs[1721] = ~((layer0_outputs[4620]) & (layer0_outputs[3977]));
    assign outputs[1722] = layer0_outputs[3825];
    assign outputs[1723] = ~((layer0_outputs[1436]) ^ (layer0_outputs[2329]));
    assign outputs[1724] = (layer0_outputs[1188]) & (layer0_outputs[2977]);
    assign outputs[1725] = layer0_outputs[3985];
    assign outputs[1726] = ~(layer0_outputs[3030]);
    assign outputs[1727] = (layer0_outputs[4744]) & (layer0_outputs[3438]);
    assign outputs[1728] = ~(layer0_outputs[4034]) | (layer0_outputs[404]);
    assign outputs[1729] = layer0_outputs[3709];
    assign outputs[1730] = ~(layer0_outputs[1790]) | (layer0_outputs[455]);
    assign outputs[1731] = layer0_outputs[689];
    assign outputs[1732] = ~(layer0_outputs[802]);
    assign outputs[1733] = layer0_outputs[3717];
    assign outputs[1734] = ~((layer0_outputs[3005]) | (layer0_outputs[2200]));
    assign outputs[1735] = layer0_outputs[3239];
    assign outputs[1736] = ~(layer0_outputs[1531]);
    assign outputs[1737] = ~((layer0_outputs[333]) ^ (layer0_outputs[4186]));
    assign outputs[1738] = ~(layer0_outputs[1020]);
    assign outputs[1739] = ~(layer0_outputs[3998]) | (layer0_outputs[2238]);
    assign outputs[1740] = layer0_outputs[2971];
    assign outputs[1741] = (layer0_outputs[1927]) ^ (layer0_outputs[2538]);
    assign outputs[1742] = ~(layer0_outputs[4276]);
    assign outputs[1743] = (layer0_outputs[761]) & ~(layer0_outputs[2460]);
    assign outputs[1744] = layer0_outputs[35];
    assign outputs[1745] = layer0_outputs[3327];
    assign outputs[1746] = (layer0_outputs[3900]) & ~(layer0_outputs[4530]);
    assign outputs[1747] = ~(layer0_outputs[1482]);
    assign outputs[1748] = (layer0_outputs[2042]) & ~(layer0_outputs[673]);
    assign outputs[1749] = (layer0_outputs[3300]) ^ (layer0_outputs[1597]);
    assign outputs[1750] = layer0_outputs[4339];
    assign outputs[1751] = layer0_outputs[3948];
    assign outputs[1752] = (layer0_outputs[4753]) ^ (layer0_outputs[2801]);
    assign outputs[1753] = layer0_outputs[1338];
    assign outputs[1754] = layer0_outputs[1420];
    assign outputs[1755] = ~((layer0_outputs[161]) ^ (layer0_outputs[2155]));
    assign outputs[1756] = ~(layer0_outputs[2167]);
    assign outputs[1757] = ~(layer0_outputs[4685]);
    assign outputs[1758] = ~(layer0_outputs[4258]);
    assign outputs[1759] = layer0_outputs[176];
    assign outputs[1760] = layer0_outputs[455];
    assign outputs[1761] = ~(layer0_outputs[4000]);
    assign outputs[1762] = layer0_outputs[4521];
    assign outputs[1763] = ~(layer0_outputs[1345]);
    assign outputs[1764] = ~((layer0_outputs[4763]) ^ (layer0_outputs[101]));
    assign outputs[1765] = layer0_outputs[2779];
    assign outputs[1766] = ~((layer0_outputs[4291]) ^ (layer0_outputs[3530]));
    assign outputs[1767] = (layer0_outputs[2307]) & ~(layer0_outputs[2839]);
    assign outputs[1768] = layer0_outputs[4795];
    assign outputs[1769] = ~((layer0_outputs[2836]) ^ (layer0_outputs[3588]));
    assign outputs[1770] = (layer0_outputs[4726]) & ~(layer0_outputs[4601]);
    assign outputs[1771] = layer0_outputs[4503];
    assign outputs[1772] = ~((layer0_outputs[3648]) ^ (layer0_outputs[3352]));
    assign outputs[1773] = ~((layer0_outputs[4567]) ^ (layer0_outputs[691]));
    assign outputs[1774] = ~(layer0_outputs[4796]) | (layer0_outputs[1354]);
    assign outputs[1775] = layer0_outputs[3469];
    assign outputs[1776] = layer0_outputs[4335];
    assign outputs[1777] = ~(layer0_outputs[1408]);
    assign outputs[1778] = 1'b1;
    assign outputs[1779] = (layer0_outputs[1692]) ^ (layer0_outputs[826]);
    assign outputs[1780] = ~(layer0_outputs[3383]);
    assign outputs[1781] = (layer0_outputs[1723]) ^ (layer0_outputs[1974]);
    assign outputs[1782] = ~(layer0_outputs[4692]);
    assign outputs[1783] = ~((layer0_outputs[1633]) & (layer0_outputs[5038]));
    assign outputs[1784] = (layer0_outputs[135]) & ~(layer0_outputs[4136]);
    assign outputs[1785] = ~(layer0_outputs[4433]);
    assign outputs[1786] = ~(layer0_outputs[493]) | (layer0_outputs[2053]);
    assign outputs[1787] = ~(layer0_outputs[323]);
    assign outputs[1788] = ~((layer0_outputs[2076]) & (layer0_outputs[619]));
    assign outputs[1789] = ~(layer0_outputs[2683]);
    assign outputs[1790] = ~((layer0_outputs[1833]) ^ (layer0_outputs[2886]));
    assign outputs[1791] = (layer0_outputs[4125]) & ~(layer0_outputs[709]);
    assign outputs[1792] = ~(layer0_outputs[4927]);
    assign outputs[1793] = ~((layer0_outputs[2714]) ^ (layer0_outputs[3297]));
    assign outputs[1794] = ~((layer0_outputs[3818]) & (layer0_outputs[4373]));
    assign outputs[1795] = ~(layer0_outputs[752]) | (layer0_outputs[541]);
    assign outputs[1796] = (layer0_outputs[1505]) ^ (layer0_outputs[3973]);
    assign outputs[1797] = ~(layer0_outputs[864]) | (layer0_outputs[1416]);
    assign outputs[1798] = ~(layer0_outputs[2343]);
    assign outputs[1799] = (layer0_outputs[1512]) | (layer0_outputs[4720]);
    assign outputs[1800] = (layer0_outputs[1254]) & (layer0_outputs[330]);
    assign outputs[1801] = (layer0_outputs[4202]) ^ (layer0_outputs[3247]);
    assign outputs[1802] = (layer0_outputs[1276]) & ~(layer0_outputs[5039]);
    assign outputs[1803] = ~(layer0_outputs[968]);
    assign outputs[1804] = ~((layer0_outputs[2732]) ^ (layer0_outputs[2173]));
    assign outputs[1805] = ~((layer0_outputs[2401]) ^ (layer0_outputs[4754]));
    assign outputs[1806] = layer0_outputs[3122];
    assign outputs[1807] = ~(layer0_outputs[2855]);
    assign outputs[1808] = (layer0_outputs[3612]) & ~(layer0_outputs[4256]);
    assign outputs[1809] = ~((layer0_outputs[239]) | (layer0_outputs[1488]));
    assign outputs[1810] = ~(layer0_outputs[2028]);
    assign outputs[1811] = ~(layer0_outputs[2903]) | (layer0_outputs[1401]);
    assign outputs[1812] = layer0_outputs[360];
    assign outputs[1813] = (layer0_outputs[2530]) & ~(layer0_outputs[3727]);
    assign outputs[1814] = (layer0_outputs[2915]) ^ (layer0_outputs[667]);
    assign outputs[1815] = ~((layer0_outputs[857]) ^ (layer0_outputs[358]));
    assign outputs[1816] = (layer0_outputs[3884]) & (layer0_outputs[3148]);
    assign outputs[1817] = ~((layer0_outputs[3047]) | (layer0_outputs[1107]));
    assign outputs[1818] = (layer0_outputs[2939]) | (layer0_outputs[3153]);
    assign outputs[1819] = ~((layer0_outputs[1169]) ^ (layer0_outputs[3139]));
    assign outputs[1820] = ~((layer0_outputs[2489]) ^ (layer0_outputs[5091]));
    assign outputs[1821] = ~(layer0_outputs[2109]) | (layer0_outputs[844]);
    assign outputs[1822] = (layer0_outputs[2324]) & (layer0_outputs[4451]);
    assign outputs[1823] = ~(layer0_outputs[1933]) | (layer0_outputs[697]);
    assign outputs[1824] = ~(layer0_outputs[4936]);
    assign outputs[1825] = ~(layer0_outputs[470]) | (layer0_outputs[431]);
    assign outputs[1826] = ~((layer0_outputs[5049]) | (layer0_outputs[775]));
    assign outputs[1827] = layer0_outputs[3000];
    assign outputs[1828] = (layer0_outputs[4224]) ^ (layer0_outputs[2678]);
    assign outputs[1829] = ~(layer0_outputs[1377]);
    assign outputs[1830] = (layer0_outputs[3894]) ^ (layer0_outputs[1900]);
    assign outputs[1831] = ~((layer0_outputs[1068]) ^ (layer0_outputs[4616]));
    assign outputs[1832] = ~((layer0_outputs[4866]) ^ (layer0_outputs[3698]));
    assign outputs[1833] = ~((layer0_outputs[2075]) | (layer0_outputs[4109]));
    assign outputs[1834] = (layer0_outputs[1333]) ^ (layer0_outputs[4871]);
    assign outputs[1835] = ~(layer0_outputs[177]) | (layer0_outputs[107]);
    assign outputs[1836] = ~((layer0_outputs[4885]) ^ (layer0_outputs[5066]));
    assign outputs[1837] = ~(layer0_outputs[2672]);
    assign outputs[1838] = ~(layer0_outputs[437]) | (layer0_outputs[2447]);
    assign outputs[1839] = ~(layer0_outputs[1808]) | (layer0_outputs[1895]);
    assign outputs[1840] = layer0_outputs[3733];
    assign outputs[1841] = ~(layer0_outputs[1059]) | (layer0_outputs[2142]);
    assign outputs[1842] = (layer0_outputs[703]) ^ (layer0_outputs[1902]);
    assign outputs[1843] = (layer0_outputs[3345]) ^ (layer0_outputs[2861]);
    assign outputs[1844] = ~((layer0_outputs[2071]) ^ (layer0_outputs[2378]));
    assign outputs[1845] = layer0_outputs[2005];
    assign outputs[1846] = (layer0_outputs[4571]) ^ (layer0_outputs[708]);
    assign outputs[1847] = ~(layer0_outputs[2102]) | (layer0_outputs[3122]);
    assign outputs[1848] = ~(layer0_outputs[4274]);
    assign outputs[1849] = ~(layer0_outputs[1924]);
    assign outputs[1850] = layer0_outputs[1401];
    assign outputs[1851] = ~(layer0_outputs[432]);
    assign outputs[1852] = ~((layer0_outputs[313]) & (layer0_outputs[1746]));
    assign outputs[1853] = ~((layer0_outputs[514]) ^ (layer0_outputs[3998]));
    assign outputs[1854] = (layer0_outputs[5113]) & (layer0_outputs[3625]);
    assign outputs[1855] = (layer0_outputs[3266]) ^ (layer0_outputs[1539]);
    assign outputs[1856] = layer0_outputs[1328];
    assign outputs[1857] = layer0_outputs[3257];
    assign outputs[1858] = (layer0_outputs[2788]) & (layer0_outputs[3613]);
    assign outputs[1859] = ~((layer0_outputs[223]) ^ (layer0_outputs[4695]));
    assign outputs[1860] = 1'b1;
    assign outputs[1861] = ~(layer0_outputs[2125]);
    assign outputs[1862] = layer0_outputs[4930];
    assign outputs[1863] = ~(layer0_outputs[2002]);
    assign outputs[1864] = ~(layer0_outputs[3216]);
    assign outputs[1865] = (layer0_outputs[2007]) | (layer0_outputs[1082]);
    assign outputs[1866] = layer0_outputs[2936];
    assign outputs[1867] = layer0_outputs[1497];
    assign outputs[1868] = 1'b1;
    assign outputs[1869] = ~(layer0_outputs[3813]);
    assign outputs[1870] = ~((layer0_outputs[2433]) & (layer0_outputs[836]));
    assign outputs[1871] = (layer0_outputs[2380]) & ~(layer0_outputs[736]);
    assign outputs[1872] = ~(layer0_outputs[2132]);
    assign outputs[1873] = ~((layer0_outputs[130]) ^ (layer0_outputs[3864]));
    assign outputs[1874] = (layer0_outputs[1207]) & ~(layer0_outputs[4724]);
    assign outputs[1875] = ~((layer0_outputs[503]) | (layer0_outputs[4858]));
    assign outputs[1876] = layer0_outputs[1678];
    assign outputs[1877] = ~(layer0_outputs[1508]);
    assign outputs[1878] = (layer0_outputs[2889]) & (layer0_outputs[2806]);
    assign outputs[1879] = (layer0_outputs[2307]) & ~(layer0_outputs[1425]);
    assign outputs[1880] = (layer0_outputs[356]) | (layer0_outputs[910]);
    assign outputs[1881] = ~(layer0_outputs[4274]);
    assign outputs[1882] = ~((layer0_outputs[1381]) ^ (layer0_outputs[1441]));
    assign outputs[1883] = ~((layer0_outputs[2017]) & (layer0_outputs[4395]));
    assign outputs[1884] = ~((layer0_outputs[586]) ^ (layer0_outputs[3164]));
    assign outputs[1885] = (layer0_outputs[3991]) | (layer0_outputs[5011]);
    assign outputs[1886] = ~((layer0_outputs[813]) ^ (layer0_outputs[4244]));
    assign outputs[1887] = ~((layer0_outputs[3719]) & (layer0_outputs[4022]));
    assign outputs[1888] = ~(layer0_outputs[940]);
    assign outputs[1889] = (layer0_outputs[4638]) & (layer0_outputs[388]);
    assign outputs[1890] = ~(layer0_outputs[2109]);
    assign outputs[1891] = layer0_outputs[587];
    assign outputs[1892] = layer0_outputs[2373];
    assign outputs[1893] = ~(layer0_outputs[1273]);
    assign outputs[1894] = ~(layer0_outputs[1604]);
    assign outputs[1895] = layer0_outputs[4989];
    assign outputs[1896] = layer0_outputs[746];
    assign outputs[1897] = layer0_outputs[4515];
    assign outputs[1898] = layer0_outputs[901];
    assign outputs[1899] = ~(layer0_outputs[5066]) | (layer0_outputs[1159]);
    assign outputs[1900] = (layer0_outputs[3224]) & (layer0_outputs[4148]);
    assign outputs[1901] = (layer0_outputs[4851]) & (layer0_outputs[1217]);
    assign outputs[1902] = ~(layer0_outputs[980]);
    assign outputs[1903] = layer0_outputs[3660];
    assign outputs[1904] = layer0_outputs[3312];
    assign outputs[1905] = ~(layer0_outputs[4209]) | (layer0_outputs[4648]);
    assign outputs[1906] = layer0_outputs[1615];
    assign outputs[1907] = layer0_outputs[4949];
    assign outputs[1908] = ~((layer0_outputs[876]) | (layer0_outputs[748]));
    assign outputs[1909] = ~(layer0_outputs[4249]);
    assign outputs[1910] = ~(layer0_outputs[4079]) | (layer0_outputs[5119]);
    assign outputs[1911] = layer0_outputs[3175];
    assign outputs[1912] = ~(layer0_outputs[2674]) | (layer0_outputs[4767]);
    assign outputs[1913] = ~(layer0_outputs[5084]);
    assign outputs[1914] = (layer0_outputs[4649]) & (layer0_outputs[3952]);
    assign outputs[1915] = layer0_outputs[2439];
    assign outputs[1916] = layer0_outputs[3566];
    assign outputs[1917] = (layer0_outputs[2506]) & ~(layer0_outputs[4283]);
    assign outputs[1918] = ~(layer0_outputs[3371]);
    assign outputs[1919] = (layer0_outputs[1734]) ^ (layer0_outputs[3814]);
    assign outputs[1920] = (layer0_outputs[3682]) | (layer0_outputs[2270]);
    assign outputs[1921] = ~(layer0_outputs[4402]);
    assign outputs[1922] = (layer0_outputs[3031]) | (layer0_outputs[1089]);
    assign outputs[1923] = layer0_outputs[3700];
    assign outputs[1924] = layer0_outputs[896];
    assign outputs[1925] = layer0_outputs[5114];
    assign outputs[1926] = ~(layer0_outputs[592]);
    assign outputs[1927] = ~((layer0_outputs[1070]) & (layer0_outputs[1332]));
    assign outputs[1928] = ~(layer0_outputs[3526]);
    assign outputs[1929] = layer0_outputs[791];
    assign outputs[1930] = (layer0_outputs[2136]) & ~(layer0_outputs[3003]);
    assign outputs[1931] = layer0_outputs[1744];
    assign outputs[1932] = (layer0_outputs[4118]) & ~(layer0_outputs[4350]);
    assign outputs[1933] = layer0_outputs[5046];
    assign outputs[1934] = ~((layer0_outputs[4028]) | (layer0_outputs[276]));
    assign outputs[1935] = layer0_outputs[1027];
    assign outputs[1936] = ~((layer0_outputs[1749]) ^ (layer0_outputs[432]));
    assign outputs[1937] = ~(layer0_outputs[3226]) | (layer0_outputs[4830]);
    assign outputs[1938] = layer0_outputs[1507];
    assign outputs[1939] = ~(layer0_outputs[4996]) | (layer0_outputs[3019]);
    assign outputs[1940] = layer0_outputs[1814];
    assign outputs[1941] = ~(layer0_outputs[3267]);
    assign outputs[1942] = ~(layer0_outputs[2652]);
    assign outputs[1943] = ~(layer0_outputs[4013]);
    assign outputs[1944] = (layer0_outputs[1888]) ^ (layer0_outputs[2457]);
    assign outputs[1945] = layer0_outputs[3741];
    assign outputs[1946] = layer0_outputs[4107];
    assign outputs[1947] = ~(layer0_outputs[4526]);
    assign outputs[1948] = layer0_outputs[1762];
    assign outputs[1949] = layer0_outputs[3148];
    assign outputs[1950] = (layer0_outputs[1005]) ^ (layer0_outputs[4349]);
    assign outputs[1951] = (layer0_outputs[4654]) & (layer0_outputs[2530]);
    assign outputs[1952] = (layer0_outputs[2168]) ^ (layer0_outputs[703]);
    assign outputs[1953] = ~(layer0_outputs[2844]);
    assign outputs[1954] = ~((layer0_outputs[3360]) & (layer0_outputs[2453]));
    assign outputs[1955] = ~(layer0_outputs[1034]);
    assign outputs[1956] = ~((layer0_outputs[1272]) | (layer0_outputs[428]));
    assign outputs[1957] = layer0_outputs[4911];
    assign outputs[1958] = ~(layer0_outputs[362]) | (layer0_outputs[278]);
    assign outputs[1959] = ~(layer0_outputs[4023]);
    assign outputs[1960] = (layer0_outputs[2238]) | (layer0_outputs[301]);
    assign outputs[1961] = (layer0_outputs[3268]) & ~(layer0_outputs[780]);
    assign outputs[1962] = layer0_outputs[2910];
    assign outputs[1963] = ~(layer0_outputs[2418]);
    assign outputs[1964] = ~((layer0_outputs[4571]) ^ (layer0_outputs[3615]));
    assign outputs[1965] = ~(layer0_outputs[5090]);
    assign outputs[1966] = ~((layer0_outputs[1955]) & (layer0_outputs[918]));
    assign outputs[1967] = ~(layer0_outputs[108]);
    assign outputs[1968] = layer0_outputs[2458];
    assign outputs[1969] = (layer0_outputs[2567]) | (layer0_outputs[2693]);
    assign outputs[1970] = layer0_outputs[2254];
    assign outputs[1971] = ~(layer0_outputs[3687]) | (layer0_outputs[2308]);
    assign outputs[1972] = ~((layer0_outputs[102]) ^ (layer0_outputs[977]));
    assign outputs[1973] = ~((layer0_outputs[1389]) ^ (layer0_outputs[2714]));
    assign outputs[1974] = 1'b1;
    assign outputs[1975] = (layer0_outputs[1398]) ^ (layer0_outputs[2825]);
    assign outputs[1976] = ~((layer0_outputs[2527]) & (layer0_outputs[3694]));
    assign outputs[1977] = (layer0_outputs[2576]) & ~(layer0_outputs[338]);
    assign outputs[1978] = ~(layer0_outputs[4166]) | (layer0_outputs[2765]);
    assign outputs[1979] = 1'b1;
    assign outputs[1980] = ~((layer0_outputs[2999]) | (layer0_outputs[1342]));
    assign outputs[1981] = ~((layer0_outputs[4707]) | (layer0_outputs[1211]));
    assign outputs[1982] = (layer0_outputs[970]) & ~(layer0_outputs[2892]);
    assign outputs[1983] = ~(layer0_outputs[556]);
    assign outputs[1984] = layer0_outputs[3811];
    assign outputs[1985] = ~(layer0_outputs[491]);
    assign outputs[1986] = ~(layer0_outputs[483]);
    assign outputs[1987] = ~(layer0_outputs[704]);
    assign outputs[1988] = ~((layer0_outputs[1938]) ^ (layer0_outputs[2229]));
    assign outputs[1989] = (layer0_outputs[4468]) & ~(layer0_outputs[4801]);
    assign outputs[1990] = (layer0_outputs[4427]) ^ (layer0_outputs[4488]);
    assign outputs[1991] = (layer0_outputs[3095]) & ~(layer0_outputs[3442]);
    assign outputs[1992] = ~((layer0_outputs[3595]) ^ (layer0_outputs[4249]));
    assign outputs[1993] = ~((layer0_outputs[1119]) & (layer0_outputs[1911]));
    assign outputs[1994] = ~(layer0_outputs[2868]) | (layer0_outputs[2763]);
    assign outputs[1995] = ~((layer0_outputs[3563]) & (layer0_outputs[2994]));
    assign outputs[1996] = layer0_outputs[4750];
    assign outputs[1997] = ~(layer0_outputs[2596]);
    assign outputs[1998] = ~((layer0_outputs[4244]) ^ (layer0_outputs[3282]));
    assign outputs[1999] = (layer0_outputs[40]) & ~(layer0_outputs[215]);
    assign outputs[2000] = (layer0_outputs[2352]) & ~(layer0_outputs[1650]);
    assign outputs[2001] = ~((layer0_outputs[835]) & (layer0_outputs[2948]));
    assign outputs[2002] = (layer0_outputs[738]) ^ (layer0_outputs[4422]);
    assign outputs[2003] = (layer0_outputs[4314]) & ~(layer0_outputs[3595]);
    assign outputs[2004] = (layer0_outputs[3520]) ^ (layer0_outputs[4150]);
    assign outputs[2005] = layer0_outputs[1480];
    assign outputs[2006] = layer0_outputs[4272];
    assign outputs[2007] = ~((layer0_outputs[2377]) ^ (layer0_outputs[1125]));
    assign outputs[2008] = (layer0_outputs[3303]) & ~(layer0_outputs[2952]);
    assign outputs[2009] = ~((layer0_outputs[281]) & (layer0_outputs[1275]));
    assign outputs[2010] = (layer0_outputs[3454]) & (layer0_outputs[1390]);
    assign outputs[2011] = (layer0_outputs[2427]) | (layer0_outputs[1496]);
    assign outputs[2012] = ~(layer0_outputs[3477]);
    assign outputs[2013] = ~((layer0_outputs[3396]) ^ (layer0_outputs[1454]));
    assign outputs[2014] = ~(layer0_outputs[4362]) | (layer0_outputs[5072]);
    assign outputs[2015] = layer0_outputs[1478];
    assign outputs[2016] = ~(layer0_outputs[4117]);
    assign outputs[2017] = ~((layer0_outputs[3829]) ^ (layer0_outputs[385]));
    assign outputs[2018] = (layer0_outputs[1685]) & ~(layer0_outputs[1915]);
    assign outputs[2019] = layer0_outputs[3898];
    assign outputs[2020] = (layer0_outputs[268]) | (layer0_outputs[3843]);
    assign outputs[2021] = ~((layer0_outputs[1602]) ^ (layer0_outputs[918]));
    assign outputs[2022] = (layer0_outputs[1011]) & ~(layer0_outputs[3051]);
    assign outputs[2023] = layer0_outputs[1708];
    assign outputs[2024] = layer0_outputs[153];
    assign outputs[2025] = layer0_outputs[4789];
    assign outputs[2026] = layer0_outputs[1940];
    assign outputs[2027] = layer0_outputs[2316];
    assign outputs[2028] = ~(layer0_outputs[1900]);
    assign outputs[2029] = ~((layer0_outputs[340]) | (layer0_outputs[555]));
    assign outputs[2030] = ~(layer0_outputs[1515]);
    assign outputs[2031] = ~((layer0_outputs[2699]) & (layer0_outputs[2578]));
    assign outputs[2032] = ~(layer0_outputs[4465]);
    assign outputs[2033] = ~(layer0_outputs[1491]);
    assign outputs[2034] = ~((layer0_outputs[728]) ^ (layer0_outputs[4346]));
    assign outputs[2035] = (layer0_outputs[4029]) & (layer0_outputs[5051]);
    assign outputs[2036] = (layer0_outputs[1954]) & (layer0_outputs[5003]);
    assign outputs[2037] = ~(layer0_outputs[3504]) | (layer0_outputs[3608]);
    assign outputs[2038] = ~(layer0_outputs[2240]);
    assign outputs[2039] = ~(layer0_outputs[4203]);
    assign outputs[2040] = ~((layer0_outputs[3006]) | (layer0_outputs[3868]));
    assign outputs[2041] = ~(layer0_outputs[2250]);
    assign outputs[2042] = layer0_outputs[3010];
    assign outputs[2043] = 1'b1;
    assign outputs[2044] = (layer0_outputs[2955]) | (layer0_outputs[3464]);
    assign outputs[2045] = layer0_outputs[3440];
    assign outputs[2046] = ~(layer0_outputs[4199]) | (layer0_outputs[474]);
    assign outputs[2047] = (layer0_outputs[3281]) | (layer0_outputs[2188]);
    assign outputs[2048] = layer0_outputs[2013];
    assign outputs[2049] = ~(layer0_outputs[3891]) | (layer0_outputs[4157]);
    assign outputs[2050] = layer0_outputs[4178];
    assign outputs[2051] = (layer0_outputs[1654]) & ~(layer0_outputs[3337]);
    assign outputs[2052] = layer0_outputs[3662];
    assign outputs[2053] = ~((layer0_outputs[1978]) | (layer0_outputs[995]));
    assign outputs[2054] = ~(layer0_outputs[1524]) | (layer0_outputs[1864]);
    assign outputs[2055] = ~((layer0_outputs[2794]) ^ (layer0_outputs[2796]));
    assign outputs[2056] = layer0_outputs[4816];
    assign outputs[2057] = (layer0_outputs[436]) & ~(layer0_outputs[3354]);
    assign outputs[2058] = layer0_outputs[2736];
    assign outputs[2059] = ~(layer0_outputs[791]);
    assign outputs[2060] = ~((layer0_outputs[271]) | (layer0_outputs[4722]));
    assign outputs[2061] = (layer0_outputs[4168]) & ~(layer0_outputs[633]);
    assign outputs[2062] = ~((layer0_outputs[1822]) ^ (layer0_outputs[3090]));
    assign outputs[2063] = (layer0_outputs[476]) & (layer0_outputs[449]);
    assign outputs[2064] = ~((layer0_outputs[4026]) | (layer0_outputs[1242]));
    assign outputs[2065] = ~((layer0_outputs[4647]) ^ (layer0_outputs[4737]));
    assign outputs[2066] = ~((layer0_outputs[4672]) & (layer0_outputs[1298]));
    assign outputs[2067] = (layer0_outputs[3365]) & ~(layer0_outputs[2383]);
    assign outputs[2068] = ~(layer0_outputs[4231]);
    assign outputs[2069] = layer0_outputs[2187];
    assign outputs[2070] = (layer0_outputs[4694]) & ~(layer0_outputs[658]);
    assign outputs[2071] = (layer0_outputs[1494]) | (layer0_outputs[754]);
    assign outputs[2072] = ~(layer0_outputs[546]);
    assign outputs[2073] = ~(layer0_outputs[613]) | (layer0_outputs[3231]);
    assign outputs[2074] = (layer0_outputs[2916]) ^ (layer0_outputs[500]);
    assign outputs[2075] = ~((layer0_outputs[4782]) ^ (layer0_outputs[1327]));
    assign outputs[2076] = (layer0_outputs[4949]) & ~(layer0_outputs[4069]);
    assign outputs[2077] = (layer0_outputs[3855]) ^ (layer0_outputs[3535]);
    assign outputs[2078] = (layer0_outputs[1716]) & ~(layer0_outputs[3353]);
    assign outputs[2079] = ~(layer0_outputs[1811]);
    assign outputs[2080] = (layer0_outputs[2499]) ^ (layer0_outputs[1351]);
    assign outputs[2081] = (layer0_outputs[4881]) & ~(layer0_outputs[2677]);
    assign outputs[2082] = ~(layer0_outputs[1410]) | (layer0_outputs[3527]);
    assign outputs[2083] = ~(layer0_outputs[866]);
    assign outputs[2084] = ~(layer0_outputs[4411]);
    assign outputs[2085] = layer0_outputs[671];
    assign outputs[2086] = (layer0_outputs[277]) & (layer0_outputs[4718]);
    assign outputs[2087] = ~((layer0_outputs[2406]) | (layer0_outputs[3131]));
    assign outputs[2088] = ~(layer0_outputs[3175]);
    assign outputs[2089] = layer0_outputs[2796];
    assign outputs[2090] = ~((layer0_outputs[3770]) & (layer0_outputs[3389]));
    assign outputs[2091] = (layer0_outputs[2961]) & ~(layer0_outputs[1378]);
    assign outputs[2092] = (layer0_outputs[2684]) & ~(layer0_outputs[4861]);
    assign outputs[2093] = ~(layer0_outputs[3133]);
    assign outputs[2094] = (layer0_outputs[635]) ^ (layer0_outputs[2704]);
    assign outputs[2095] = ~((layer0_outputs[225]) | (layer0_outputs[3862]));
    assign outputs[2096] = (layer0_outputs[882]) & (layer0_outputs[4404]);
    assign outputs[2097] = (layer0_outputs[3863]) ^ (layer0_outputs[4655]);
    assign outputs[2098] = ~((layer0_outputs[2206]) | (layer0_outputs[2231]));
    assign outputs[2099] = ~(layer0_outputs[4887]);
    assign outputs[2100] = ~(layer0_outputs[810]);
    assign outputs[2101] = (layer0_outputs[3363]) & ~(layer0_outputs[473]);
    assign outputs[2102] = ~(layer0_outputs[4098]) | (layer0_outputs[761]);
    assign outputs[2103] = layer0_outputs[530];
    assign outputs[2104] = ~(layer0_outputs[182]);
    assign outputs[2105] = layer0_outputs[2098];
    assign outputs[2106] = layer0_outputs[1128];
    assign outputs[2107] = ~(layer0_outputs[1498]);
    assign outputs[2108] = (layer0_outputs[1982]) & ~(layer0_outputs[201]);
    assign outputs[2109] = ~(layer0_outputs[431]);
    assign outputs[2110] = (layer0_outputs[4266]) & ~(layer0_outputs[2449]);
    assign outputs[2111] = ~(layer0_outputs[3126]);
    assign outputs[2112] = (layer0_outputs[1907]) & (layer0_outputs[3443]);
    assign outputs[2113] = layer0_outputs[794];
    assign outputs[2114] = (layer0_outputs[691]) & ~(layer0_outputs[4494]);
    assign outputs[2115] = (layer0_outputs[171]) & (layer0_outputs[4915]);
    assign outputs[2116] = ~((layer0_outputs[2452]) ^ (layer0_outputs[4745]));
    assign outputs[2117] = layer0_outputs[1121];
    assign outputs[2118] = (layer0_outputs[1540]) & ~(layer0_outputs[2735]);
    assign outputs[2119] = (layer0_outputs[1424]) & (layer0_outputs[3161]);
    assign outputs[2120] = (layer0_outputs[2341]) & ~(layer0_outputs[4994]);
    assign outputs[2121] = layer0_outputs[1844];
    assign outputs[2122] = ~(layer0_outputs[4384]) | (layer0_outputs[5024]);
    assign outputs[2123] = layer0_outputs[3641];
    assign outputs[2124] = (layer0_outputs[2511]) ^ (layer0_outputs[2474]);
    assign outputs[2125] = layer0_outputs[3679];
    assign outputs[2126] = (layer0_outputs[3713]) ^ (layer0_outputs[4514]);
    assign outputs[2127] = ~((layer0_outputs[4763]) ^ (layer0_outputs[2]));
    assign outputs[2128] = ~(layer0_outputs[2795]);
    assign outputs[2129] = ~(layer0_outputs[822]);
    assign outputs[2130] = layer0_outputs[2303];
    assign outputs[2131] = (layer0_outputs[2112]) & ~(layer0_outputs[3597]);
    assign outputs[2132] = ~((layer0_outputs[459]) ^ (layer0_outputs[4769]));
    assign outputs[2133] = ~((layer0_outputs[2691]) & (layer0_outputs[1813]));
    assign outputs[2134] = layer0_outputs[4188];
    assign outputs[2135] = layer0_outputs[5115];
    assign outputs[2136] = layer0_outputs[4615];
    assign outputs[2137] = (layer0_outputs[2232]) ^ (layer0_outputs[1606]);
    assign outputs[2138] = layer0_outputs[1663];
    assign outputs[2139] = (layer0_outputs[2088]) ^ (layer0_outputs[394]);
    assign outputs[2140] = ~((layer0_outputs[3870]) ^ (layer0_outputs[990]));
    assign outputs[2141] = layer0_outputs[1511];
    assign outputs[2142] = (layer0_outputs[1394]) & ~(layer0_outputs[2771]);
    assign outputs[2143] = ~(layer0_outputs[2129]);
    assign outputs[2144] = ~((layer0_outputs[4632]) ^ (layer0_outputs[1979]));
    assign outputs[2145] = layer0_outputs[4964];
    assign outputs[2146] = (layer0_outputs[2591]) | (layer0_outputs[1567]);
    assign outputs[2147] = (layer0_outputs[1990]) & ~(layer0_outputs[3316]);
    assign outputs[2148] = (layer0_outputs[15]) ^ (layer0_outputs[1228]);
    assign outputs[2149] = (layer0_outputs[4583]) & (layer0_outputs[3017]);
    assign outputs[2150] = (layer0_outputs[3149]) & (layer0_outputs[3341]);
    assign outputs[2151] = (layer0_outputs[4895]) ^ (layer0_outputs[1965]);
    assign outputs[2152] = (layer0_outputs[1244]) & (layer0_outputs[3478]);
    assign outputs[2153] = ~((layer0_outputs[3093]) ^ (layer0_outputs[3164]));
    assign outputs[2154] = (layer0_outputs[4738]) & (layer0_outputs[4492]);
    assign outputs[2155] = ~(layer0_outputs[1322]) | (layer0_outputs[419]);
    assign outputs[2156] = ~((layer0_outputs[1996]) ^ (layer0_outputs[5025]));
    assign outputs[2157] = ~(layer0_outputs[3934]) | (layer0_outputs[4821]);
    assign outputs[2158] = (layer0_outputs[3158]) ^ (layer0_outputs[138]);
    assign outputs[2159] = (layer0_outputs[90]) & ~(layer0_outputs[2639]);
    assign outputs[2160] = layer0_outputs[2662];
    assign outputs[2161] = ~((layer0_outputs[5076]) ^ (layer0_outputs[1274]));
    assign outputs[2162] = ~((layer0_outputs[2997]) ^ (layer0_outputs[2407]));
    assign outputs[2163] = layer0_outputs[1849];
    assign outputs[2164] = layer0_outputs[3953];
    assign outputs[2165] = layer0_outputs[2857];
    assign outputs[2166] = layer0_outputs[1781];
    assign outputs[2167] = ~((layer0_outputs[2296]) | (layer0_outputs[2041]));
    assign outputs[2168] = layer0_outputs[2439];
    assign outputs[2169] = ~((layer0_outputs[3537]) ^ (layer0_outputs[1995]));
    assign outputs[2170] = (layer0_outputs[1554]) & ~(layer0_outputs[1260]);
    assign outputs[2171] = ~((layer0_outputs[3655]) & (layer0_outputs[3561]));
    assign outputs[2172] = ~((layer0_outputs[2783]) | (layer0_outputs[499]));
    assign outputs[2173] = ~(layer0_outputs[4412]);
    assign outputs[2174] = ~(layer0_outputs[4154]);
    assign outputs[2175] = (layer0_outputs[1740]) & (layer0_outputs[4894]);
    assign outputs[2176] = ~(layer0_outputs[3173]) | (layer0_outputs[3932]);
    assign outputs[2177] = ~(layer0_outputs[1902]);
    assign outputs[2178] = (layer0_outputs[3563]) & ~(layer0_outputs[575]);
    assign outputs[2179] = (layer0_outputs[266]) & ~(layer0_outputs[2503]);
    assign outputs[2180] = ~(layer0_outputs[162]) | (layer0_outputs[1484]);
    assign outputs[2181] = (layer0_outputs[4519]) | (layer0_outputs[1823]);
    assign outputs[2182] = ~((layer0_outputs[1100]) ^ (layer0_outputs[4354]));
    assign outputs[2183] = ~((layer0_outputs[2249]) & (layer0_outputs[655]));
    assign outputs[2184] = layer0_outputs[3432];
    assign outputs[2185] = ~((layer0_outputs[1651]) ^ (layer0_outputs[2963]));
    assign outputs[2186] = ~((layer0_outputs[2918]) ^ (layer0_outputs[2820]));
    assign outputs[2187] = (layer0_outputs[4855]) & ~(layer0_outputs[2969]);
    assign outputs[2188] = layer0_outputs[445];
    assign outputs[2189] = (layer0_outputs[4284]) & (layer0_outputs[4027]);
    assign outputs[2190] = ~(layer0_outputs[3043]);
    assign outputs[2191] = layer0_outputs[5104];
    assign outputs[2192] = ~(layer0_outputs[4334]);
    assign outputs[2193] = layer0_outputs[3866];
    assign outputs[2194] = ~((layer0_outputs[1443]) & (layer0_outputs[2178]));
    assign outputs[2195] = (layer0_outputs[2703]) & ~(layer0_outputs[4942]);
    assign outputs[2196] = (layer0_outputs[1288]) & ~(layer0_outputs[3086]);
    assign outputs[2197] = layer0_outputs[3431];
    assign outputs[2198] = ~(layer0_outputs[1685]);
    assign outputs[2199] = ~(layer0_outputs[3494]);
    assign outputs[2200] = (layer0_outputs[923]) & ~(layer0_outputs[4418]);
    assign outputs[2201] = layer0_outputs[3824];
    assign outputs[2202] = (layer0_outputs[1110]) ^ (layer0_outputs[4528]);
    assign outputs[2203] = (layer0_outputs[4725]) ^ (layer0_outputs[2582]);
    assign outputs[2204] = ~(layer0_outputs[3451]);
    assign outputs[2205] = ~(layer0_outputs[926]);
    assign outputs[2206] = ~(layer0_outputs[310]);
    assign outputs[2207] = layer0_outputs[2207];
    assign outputs[2208] = (layer0_outputs[1960]) & ~(layer0_outputs[1590]);
    assign outputs[2209] = ~(layer0_outputs[5012]);
    assign outputs[2210] = layer0_outputs[4650];
    assign outputs[2211] = ~((layer0_outputs[3106]) ^ (layer0_outputs[3575]));
    assign outputs[2212] = ~((layer0_outputs[3187]) | (layer0_outputs[3832]));
    assign outputs[2213] = ~((layer0_outputs[3125]) ^ (layer0_outputs[1009]));
    assign outputs[2214] = (layer0_outputs[1277]) & (layer0_outputs[1035]);
    assign outputs[2215] = ~(layer0_outputs[1448]);
    assign outputs[2216] = (layer0_outputs[2283]) & (layer0_outputs[1825]);
    assign outputs[2217] = layer0_outputs[3457];
    assign outputs[2218] = ~((layer0_outputs[1733]) ^ (layer0_outputs[4017]));
    assign outputs[2219] = layer0_outputs[1174];
    assign outputs[2220] = layer0_outputs[1024];
    assign outputs[2221] = ~((layer0_outputs[2467]) ^ (layer0_outputs[3842]));
    assign outputs[2222] = layer0_outputs[1611];
    assign outputs[2223] = (layer0_outputs[471]) & (layer0_outputs[4978]);
    assign outputs[2224] = layer0_outputs[979];
    assign outputs[2225] = ~((layer0_outputs[546]) ^ (layer0_outputs[3992]));
    assign outputs[2226] = ~((layer0_outputs[3515]) ^ (layer0_outputs[3994]));
    assign outputs[2227] = ~(layer0_outputs[1465]);
    assign outputs[2228] = (layer0_outputs[1892]) & ~(layer0_outputs[4544]);
    assign outputs[2229] = ~((layer0_outputs[2204]) ^ (layer0_outputs[3635]));
    assign outputs[2230] = (layer0_outputs[4680]) & (layer0_outputs[1607]);
    assign outputs[2231] = layer0_outputs[596];
    assign outputs[2232] = layer0_outputs[5064];
    assign outputs[2233] = layer0_outputs[4281];
    assign outputs[2234] = ~((layer0_outputs[341]) ^ (layer0_outputs[1397]));
    assign outputs[2235] = ~(layer0_outputs[479]);
    assign outputs[2236] = ~(layer0_outputs[1347]);
    assign outputs[2237] = (layer0_outputs[5068]) ^ (layer0_outputs[3867]);
    assign outputs[2238] = (layer0_outputs[2298]) & ~(layer0_outputs[5001]);
    assign outputs[2239] = layer0_outputs[4000];
    assign outputs[2240] = ~(layer0_outputs[3825]);
    assign outputs[2241] = (layer0_outputs[1922]) & (layer0_outputs[4572]);
    assign outputs[2242] = ~(layer0_outputs[3566]);
    assign outputs[2243] = (layer0_outputs[3517]) & (layer0_outputs[979]);
    assign outputs[2244] = ~((layer0_outputs[1220]) ^ (layer0_outputs[1160]));
    assign outputs[2245] = layer0_outputs[2547];
    assign outputs[2246] = ~((layer0_outputs[2708]) ^ (layer0_outputs[4730]));
    assign outputs[2247] = (layer0_outputs[2156]) ^ (layer0_outputs[2497]);
    assign outputs[2248] = (layer0_outputs[1697]) ^ (layer0_outputs[2093]);
    assign outputs[2249] = ~(layer0_outputs[3946]);
    assign outputs[2250] = 1'b0;
    assign outputs[2251] = (layer0_outputs[1793]) ^ (layer0_outputs[2131]);
    assign outputs[2252] = (layer0_outputs[4971]) ^ (layer0_outputs[2509]);
    assign outputs[2253] = layer0_outputs[4214];
    assign outputs[2254] = ~((layer0_outputs[537]) ^ (layer0_outputs[161]));
    assign outputs[2255] = ~((layer0_outputs[1317]) | (layer0_outputs[87]));
    assign outputs[2256] = (layer0_outputs[1262]) ^ (layer0_outputs[2813]);
    assign outputs[2257] = (layer0_outputs[4212]) & (layer0_outputs[2550]);
    assign outputs[2258] = layer0_outputs[1245];
    assign outputs[2259] = ~(layer0_outputs[4817]);
    assign outputs[2260] = ~((layer0_outputs[3470]) | (layer0_outputs[2312]));
    assign outputs[2261] = (layer0_outputs[3317]) ^ (layer0_outputs[2601]);
    assign outputs[2262] = ~((layer0_outputs[2854]) ^ (layer0_outputs[4104]));
    assign outputs[2263] = ~(layer0_outputs[1287]);
    assign outputs[2264] = ~(layer0_outputs[3787]) | (layer0_outputs[1953]);
    assign outputs[2265] = ~(layer0_outputs[2110]);
    assign outputs[2266] = ~((layer0_outputs[1815]) ^ (layer0_outputs[4393]));
    assign outputs[2267] = (layer0_outputs[1573]) & (layer0_outputs[1516]);
    assign outputs[2268] = ~(layer0_outputs[4513]);
    assign outputs[2269] = ~((layer0_outputs[4297]) | (layer0_outputs[1146]));
    assign outputs[2270] = ~((layer0_outputs[714]) & (layer0_outputs[1753]));
    assign outputs[2271] = ~(layer0_outputs[1349]);
    assign outputs[2272] = (layer0_outputs[89]) & ~(layer0_outputs[1757]);
    assign outputs[2273] = ~((layer0_outputs[4258]) ^ (layer0_outputs[3649]));
    assign outputs[2274] = (layer0_outputs[2495]) & (layer0_outputs[874]);
    assign outputs[2275] = ~(layer0_outputs[2959]);
    assign outputs[2276] = ~((layer0_outputs[3221]) | (layer0_outputs[994]));
    assign outputs[2277] = ~(layer0_outputs[2707]);
    assign outputs[2278] = (layer0_outputs[129]) ^ (layer0_outputs[3867]);
    assign outputs[2279] = ~(layer0_outputs[4961]);
    assign outputs[2280] = layer0_outputs[3668];
    assign outputs[2281] = ~(layer0_outputs[3898]);
    assign outputs[2282] = (layer0_outputs[4813]) & ~(layer0_outputs[4099]);
    assign outputs[2283] = ~(layer0_outputs[5033]);
    assign outputs[2284] = (layer0_outputs[2874]) & ~(layer0_outputs[218]);
    assign outputs[2285] = (layer0_outputs[4743]) & (layer0_outputs[4322]);
    assign outputs[2286] = (layer0_outputs[4761]) & (layer0_outputs[195]);
    assign outputs[2287] = ~((layer0_outputs[4213]) | (layer0_outputs[1804]));
    assign outputs[2288] = layer0_outputs[4100];
    assign outputs[2289] = 1'b1;
    assign outputs[2290] = (layer0_outputs[3621]) & ~(layer0_outputs[991]);
    assign outputs[2291] = ~((layer0_outputs[920]) ^ (layer0_outputs[1404]));
    assign outputs[2292] = layer0_outputs[4918];
    assign outputs[2293] = (layer0_outputs[233]) & ~(layer0_outputs[830]);
    assign outputs[2294] = layer0_outputs[1726];
    assign outputs[2295] = layer0_outputs[1700];
    assign outputs[2296] = ~((layer0_outputs[616]) ^ (layer0_outputs[2771]));
    assign outputs[2297] = ~(layer0_outputs[191]);
    assign outputs[2298] = layer0_outputs[4770];
    assign outputs[2299] = layer0_outputs[1047];
    assign outputs[2300] = (layer0_outputs[2574]) ^ (layer0_outputs[4848]);
    assign outputs[2301] = ~(layer0_outputs[1497]);
    assign outputs[2302] = layer0_outputs[4583];
    assign outputs[2303] = layer0_outputs[1706];
    assign outputs[2304] = ~(layer0_outputs[4716]) | (layer0_outputs[3198]);
    assign outputs[2305] = (layer0_outputs[1527]) & ~(layer0_outputs[1255]);
    assign outputs[2306] = (layer0_outputs[84]) & ~(layer0_outputs[1217]);
    assign outputs[2307] = ~((layer0_outputs[859]) ^ (layer0_outputs[2742]));
    assign outputs[2308] = ~(layer0_outputs[1282]);
    assign outputs[2309] = (layer0_outputs[4500]) & (layer0_outputs[4142]);
    assign outputs[2310] = ~(layer0_outputs[4998]) | (layer0_outputs[2413]);
    assign outputs[2311] = ~((layer0_outputs[849]) ^ (layer0_outputs[786]));
    assign outputs[2312] = layer0_outputs[1490];
    assign outputs[2313] = (layer0_outputs[2726]) & (layer0_outputs[2681]);
    assign outputs[2314] = (layer0_outputs[3581]) ^ (layer0_outputs[4130]);
    assign outputs[2315] = ~(layer0_outputs[3337]);
    assign outputs[2316] = ~(layer0_outputs[3778]);
    assign outputs[2317] = ~(layer0_outputs[3101]);
    assign outputs[2318] = (layer0_outputs[4883]) & ~(layer0_outputs[4611]);
    assign outputs[2319] = (layer0_outputs[1886]) & ~(layer0_outputs[3971]);
    assign outputs[2320] = (layer0_outputs[2646]) & (layer0_outputs[4034]);
    assign outputs[2321] = ~((layer0_outputs[441]) | (layer0_outputs[3538]));
    assign outputs[2322] = layer0_outputs[1399];
    assign outputs[2323] = ~((layer0_outputs[3369]) ^ (layer0_outputs[3026]));
    assign outputs[2324] = layer0_outputs[2925];
    assign outputs[2325] = ~((layer0_outputs[3670]) | (layer0_outputs[537]));
    assign outputs[2326] = layer0_outputs[771];
    assign outputs[2327] = (layer0_outputs[1031]) ^ (layer0_outputs[3112]);
    assign outputs[2328] = (layer0_outputs[3571]) & ~(layer0_outputs[4445]);
    assign outputs[2329] = ~(layer0_outputs[1021]);
    assign outputs[2330] = ~(layer0_outputs[1866]);
    assign outputs[2331] = (layer0_outputs[2580]) & ~(layer0_outputs[1341]);
    assign outputs[2332] = layer0_outputs[353];
    assign outputs[2333] = (layer0_outputs[2991]) & ~(layer0_outputs[1962]);
    assign outputs[2334] = layer0_outputs[1007];
    assign outputs[2335] = layer0_outputs[4396];
    assign outputs[2336] = layer0_outputs[4200];
    assign outputs[2337] = layer0_outputs[839];
    assign outputs[2338] = ~(layer0_outputs[4481]);
    assign outputs[2339] = layer0_outputs[1960];
    assign outputs[2340] = layer0_outputs[1617];
    assign outputs[2341] = ~(layer0_outputs[933]);
    assign outputs[2342] = ~((layer0_outputs[2904]) | (layer0_outputs[2342]));
    assign outputs[2343] = ~(layer0_outputs[2727]);
    assign outputs[2344] = ~((layer0_outputs[4518]) & (layer0_outputs[491]));
    assign outputs[2345] = ~(layer0_outputs[4804]);
    assign outputs[2346] = layer0_outputs[1000];
    assign outputs[2347] = ~((layer0_outputs[2712]) ^ (layer0_outputs[826]));
    assign outputs[2348] = (layer0_outputs[2395]) ^ (layer0_outputs[4138]);
    assign outputs[2349] = ~((layer0_outputs[3234]) ^ (layer0_outputs[2900]));
    assign outputs[2350] = ~((layer0_outputs[49]) ^ (layer0_outputs[545]));
    assign outputs[2351] = (layer0_outputs[2808]) ^ (layer0_outputs[2981]);
    assign outputs[2352] = (layer0_outputs[855]) | (layer0_outputs[3322]);
    assign outputs[2353] = layer0_outputs[1846];
    assign outputs[2354] = ~(layer0_outputs[1030]);
    assign outputs[2355] = ~(layer0_outputs[4507]);
    assign outputs[2356] = ~((layer0_outputs[3753]) ^ (layer0_outputs[1157]));
    assign outputs[2357] = (layer0_outputs[2032]) & ~(layer0_outputs[4368]);
    assign outputs[2358] = (layer0_outputs[3560]) & ~(layer0_outputs[1728]);
    assign outputs[2359] = layer0_outputs[1575];
    assign outputs[2360] = ~((layer0_outputs[2223]) ^ (layer0_outputs[4680]));
    assign outputs[2361] = 1'b0;
    assign outputs[2362] = ~(layer0_outputs[3174]);
    assign outputs[2363] = ~((layer0_outputs[3506]) ^ (layer0_outputs[4844]));
    assign outputs[2364] = (layer0_outputs[281]) & ~(layer0_outputs[3798]);
    assign outputs[2365] = (layer0_outputs[609]) & ~(layer0_outputs[261]);
    assign outputs[2366] = ~(layer0_outputs[1001]);
    assign outputs[2367] = ~((layer0_outputs[2684]) | (layer0_outputs[809]));
    assign outputs[2368] = ~(layer0_outputs[3280]);
    assign outputs[2369] = (layer0_outputs[2699]) & ~(layer0_outputs[1471]);
    assign outputs[2370] = (layer0_outputs[1047]) & ~(layer0_outputs[965]);
    assign outputs[2371] = ~((layer0_outputs[5012]) | (layer0_outputs[1748]));
    assign outputs[2372] = ~((layer0_outputs[3329]) ^ (layer0_outputs[2339]));
    assign outputs[2373] = layer0_outputs[2056];
    assign outputs[2374] = ~(layer0_outputs[3979]) | (layer0_outputs[1660]);
    assign outputs[2375] = ~((layer0_outputs[951]) & (layer0_outputs[549]));
    assign outputs[2376] = layer0_outputs[1550];
    assign outputs[2377] = layer0_outputs[5020];
    assign outputs[2378] = ~((layer0_outputs[4667]) ^ (layer0_outputs[2831]));
    assign outputs[2379] = layer0_outputs[239];
    assign outputs[2380] = ~(layer0_outputs[2162]);
    assign outputs[2381] = ~((layer0_outputs[937]) ^ (layer0_outputs[843]));
    assign outputs[2382] = layer0_outputs[1646];
    assign outputs[2383] = layer0_outputs[1198];
    assign outputs[2384] = (layer0_outputs[1678]) & ~(layer0_outputs[2321]);
    assign outputs[2385] = (layer0_outputs[2069]) ^ (layer0_outputs[4646]);
    assign outputs[2386] = ~((layer0_outputs[1707]) ^ (layer0_outputs[28]));
    assign outputs[2387] = ~((layer0_outputs[4609]) ^ (layer0_outputs[1951]));
    assign outputs[2388] = (layer0_outputs[2030]) & ~(layer0_outputs[392]);
    assign outputs[2389] = ~((layer0_outputs[4730]) ^ (layer0_outputs[1836]));
    assign outputs[2390] = ~((layer0_outputs[591]) & (layer0_outputs[832]));
    assign outputs[2391] = (layer0_outputs[4743]) & (layer0_outputs[3837]);
    assign outputs[2392] = ~(layer0_outputs[1193]) | (layer0_outputs[1156]);
    assign outputs[2393] = (layer0_outputs[5048]) & ~(layer0_outputs[123]);
    assign outputs[2394] = (layer0_outputs[4558]) & ~(layer0_outputs[641]);
    assign outputs[2395] = layer0_outputs[2409];
    assign outputs[2396] = ~((layer0_outputs[920]) ^ (layer0_outputs[4330]));
    assign outputs[2397] = layer0_outputs[1406];
    assign outputs[2398] = layer0_outputs[1726];
    assign outputs[2399] = ~(layer0_outputs[1259]);
    assign outputs[2400] = ~((layer0_outputs[630]) ^ (layer0_outputs[48]));
    assign outputs[2401] = (layer0_outputs[734]) ^ (layer0_outputs[5022]);
    assign outputs[2402] = ~(layer0_outputs[5054]);
    assign outputs[2403] = ~(layer0_outputs[2291]);
    assign outputs[2404] = (layer0_outputs[1445]) & ~(layer0_outputs[2960]);
    assign outputs[2405] = layer0_outputs[2320];
    assign outputs[2406] = layer0_outputs[1398];
    assign outputs[2407] = layer0_outputs[4109];
    assign outputs[2408] = (layer0_outputs[2040]) ^ (layer0_outputs[701]);
    assign outputs[2409] = 1'b1;
    assign outputs[2410] = ~((layer0_outputs[3685]) | (layer0_outputs[2561]));
    assign outputs[2411] = (layer0_outputs[4014]) ^ (layer0_outputs[1935]);
    assign outputs[2412] = (layer0_outputs[2197]) & ~(layer0_outputs[3277]);
    assign outputs[2413] = (layer0_outputs[355]) & ~(layer0_outputs[5081]);
    assign outputs[2414] = ~((layer0_outputs[3441]) | (layer0_outputs[1707]));
    assign outputs[2415] = layer0_outputs[1367];
    assign outputs[2416] = ~((layer0_outputs[5026]) ^ (layer0_outputs[3156]));
    assign outputs[2417] = (layer0_outputs[4958]) & ~(layer0_outputs[1409]);
    assign outputs[2418] = (layer0_outputs[1017]) & ~(layer0_outputs[2127]);
    assign outputs[2419] = (layer0_outputs[4593]) & (layer0_outputs[710]);
    assign outputs[2420] = ~(layer0_outputs[469]);
    assign outputs[2421] = (layer0_outputs[4447]) ^ (layer0_outputs[3579]);
    assign outputs[2422] = (layer0_outputs[304]) & ~(layer0_outputs[4201]);
    assign outputs[2423] = ~((layer0_outputs[2089]) | (layer0_outputs[1640]));
    assign outputs[2424] = layer0_outputs[260];
    assign outputs[2425] = (layer0_outputs[3729]) ^ (layer0_outputs[1826]);
    assign outputs[2426] = (layer0_outputs[2083]) ^ (layer0_outputs[11]);
    assign outputs[2427] = layer0_outputs[183];
    assign outputs[2428] = ~((layer0_outputs[1260]) | (layer0_outputs[3238]));
    assign outputs[2429] = ~((layer0_outputs[835]) | (layer0_outputs[1334]));
    assign outputs[2430] = (layer0_outputs[2389]) & (layer0_outputs[2446]);
    assign outputs[2431] = layer0_outputs[2012];
    assign outputs[2432] = layer0_outputs[2297];
    assign outputs[2433] = (layer0_outputs[1313]) | (layer0_outputs[2203]);
    assign outputs[2434] = (layer0_outputs[3858]) ^ (layer0_outputs[5024]);
    assign outputs[2435] = (layer0_outputs[811]) & ~(layer0_outputs[1521]);
    assign outputs[2436] = ~(layer0_outputs[4941]);
    assign outputs[2437] = (layer0_outputs[4878]) | (layer0_outputs[462]);
    assign outputs[2438] = (layer0_outputs[3096]) & (layer0_outputs[1393]);
    assign outputs[2439] = (layer0_outputs[3138]) & (layer0_outputs[3839]);
    assign outputs[2440] = ~((layer0_outputs[267]) & (layer0_outputs[2637]));
    assign outputs[2441] = ~((layer0_outputs[4729]) ^ (layer0_outputs[3021]));
    assign outputs[2442] = ~((layer0_outputs[4753]) | (layer0_outputs[1702]));
    assign outputs[2443] = ~(layer0_outputs[3492]) | (layer0_outputs[4420]);
    assign outputs[2444] = ~(layer0_outputs[1820]);
    assign outputs[2445] = ~(layer0_outputs[610]);
    assign outputs[2446] = ~((layer0_outputs[1589]) | (layer0_outputs[747]));
    assign outputs[2447] = ~(layer0_outputs[2332]);
    assign outputs[2448] = ~(layer0_outputs[1339]);
    assign outputs[2449] = ~(layer0_outputs[2157]);
    assign outputs[2450] = ~(layer0_outputs[2027]);
    assign outputs[2451] = (layer0_outputs[2315]) & ~(layer0_outputs[2488]);
    assign outputs[2452] = (layer0_outputs[5065]) ^ (layer0_outputs[3136]);
    assign outputs[2453] = (layer0_outputs[5030]) & ~(layer0_outputs[3510]);
    assign outputs[2454] = (layer0_outputs[3357]) & ~(layer0_outputs[4385]);
    assign outputs[2455] = (layer0_outputs[3115]) & ~(layer0_outputs[67]);
    assign outputs[2456] = ~(layer0_outputs[1029]);
    assign outputs[2457] = (layer0_outputs[787]) ^ (layer0_outputs[4547]);
    assign outputs[2458] = (layer0_outputs[39]) & ~(layer0_outputs[3332]);
    assign outputs[2459] = (layer0_outputs[4678]) | (layer0_outputs[2262]);
    assign outputs[2460] = (layer0_outputs[4882]) & ~(layer0_outputs[486]);
    assign outputs[2461] = layer0_outputs[678];
    assign outputs[2462] = ~(layer0_outputs[2899]);
    assign outputs[2463] = (layer0_outputs[1101]) ^ (layer0_outputs[1880]);
    assign outputs[2464] = ~((layer0_outputs[1247]) | (layer0_outputs[3702]));
    assign outputs[2465] = layer0_outputs[690];
    assign outputs[2466] = (layer0_outputs[1512]) ^ (layer0_outputs[1203]);
    assign outputs[2467] = ~(layer0_outputs[3118]);
    assign outputs[2468] = ~(layer0_outputs[3693]) | (layer0_outputs[2330]);
    assign outputs[2469] = ~((layer0_outputs[3958]) & (layer0_outputs[4061]));
    assign outputs[2470] = ~(layer0_outputs[3390]);
    assign outputs[2471] = layer0_outputs[2521];
    assign outputs[2472] = (layer0_outputs[4802]) & ~(layer0_outputs[1761]);
    assign outputs[2473] = ~((layer0_outputs[1360]) & (layer0_outputs[2968]));
    assign outputs[2474] = layer0_outputs[3593];
    assign outputs[2475] = (layer0_outputs[1438]) & (layer0_outputs[928]);
    assign outputs[2476] = layer0_outputs[5103];
    assign outputs[2477] = (layer0_outputs[171]) ^ (layer0_outputs[1440]);
    assign outputs[2478] = ~((layer0_outputs[4919]) ^ (layer0_outputs[3305]));
    assign outputs[2479] = ~(layer0_outputs[4143]) | (layer0_outputs[3681]);
    assign outputs[2480] = ~((layer0_outputs[4457]) ^ (layer0_outputs[2776]));
    assign outputs[2481] = ~((layer0_outputs[4124]) | (layer0_outputs[3905]));
    assign outputs[2482] = layer0_outputs[2767];
    assign outputs[2483] = (layer0_outputs[4896]) & ~(layer0_outputs[3674]);
    assign outputs[2484] = (layer0_outputs[631]) & ~(layer0_outputs[160]);
    assign outputs[2485] = ~(layer0_outputs[3981]);
    assign outputs[2486] = (layer0_outputs[2956]) & ~(layer0_outputs[4797]);
    assign outputs[2487] = layer0_outputs[4060];
    assign outputs[2488] = layer0_outputs[2762];
    assign outputs[2489] = (layer0_outputs[3134]) & ~(layer0_outputs[4156]);
    assign outputs[2490] = (layer0_outputs[4321]) & ~(layer0_outputs[2617]);
    assign outputs[2491] = (layer0_outputs[1386]) & ~(layer0_outputs[2148]);
    assign outputs[2492] = ~(layer0_outputs[2696]);
    assign outputs[2493] = ~((layer0_outputs[69]) | (layer0_outputs[2818]));
    assign outputs[2494] = 1'b0;
    assign outputs[2495] = (layer0_outputs[2977]) & (layer0_outputs[2097]);
    assign outputs[2496] = (layer0_outputs[2120]) & (layer0_outputs[3387]);
    assign outputs[2497] = (layer0_outputs[2030]) & (layer0_outputs[4872]);
    assign outputs[2498] = ~((layer0_outputs[3750]) | (layer0_outputs[5084]));
    assign outputs[2499] = layer0_outputs[4234];
    assign outputs[2500] = (layer0_outputs[427]) ^ (layer0_outputs[2851]);
    assign outputs[2501] = ~(layer0_outputs[2698]);
    assign outputs[2502] = 1'b0;
    assign outputs[2503] = (layer0_outputs[932]) ^ (layer0_outputs[2251]);
    assign outputs[2504] = layer0_outputs[2063];
    assign outputs[2505] = layer0_outputs[4836];
    assign outputs[2506] = ~(layer0_outputs[4528]);
    assign outputs[2507] = ~(layer0_outputs[4952]);
    assign outputs[2508] = ~((layer0_outputs[4935]) ^ (layer0_outputs[3131]));
    assign outputs[2509] = layer0_outputs[3945];
    assign outputs[2510] = ~((layer0_outputs[3931]) ^ (layer0_outputs[1458]));
    assign outputs[2511] = (layer0_outputs[732]) & ~(layer0_outputs[22]);
    assign outputs[2512] = (layer0_outputs[4186]) ^ (layer0_outputs[3760]);
    assign outputs[2513] = layer0_outputs[4211];
    assign outputs[2514] = (layer0_outputs[1851]) & ~(layer0_outputs[2891]);
    assign outputs[2515] = ~((layer0_outputs[4684]) ^ (layer0_outputs[2149]));
    assign outputs[2516] = (layer0_outputs[4396]) & ~(layer0_outputs[2512]);
    assign outputs[2517] = layer0_outputs[4237];
    assign outputs[2518] = ~((layer0_outputs[2632]) ^ (layer0_outputs[509]));
    assign outputs[2519] = ~(layer0_outputs[5042]);
    assign outputs[2520] = ~(layer0_outputs[2768]);
    assign outputs[2521] = ~(layer0_outputs[3770]);
    assign outputs[2522] = layer0_outputs[3258];
    assign outputs[2523] = ~((layer0_outputs[4440]) ^ (layer0_outputs[727]));
    assign outputs[2524] = (layer0_outputs[1226]) ^ (layer0_outputs[1144]);
    assign outputs[2525] = ~(layer0_outputs[3638]);
    assign outputs[2526] = (layer0_outputs[2139]) ^ (layer0_outputs[3576]);
    assign outputs[2527] = ~((layer0_outputs[3515]) ^ (layer0_outputs[514]));
    assign outputs[2528] = ~(layer0_outputs[4016]);
    assign outputs[2529] = ~((layer0_outputs[1197]) ^ (layer0_outputs[1185]));
    assign outputs[2530] = layer0_outputs[3022];
    assign outputs[2531] = ~((layer0_outputs[2045]) & (layer0_outputs[4786]));
    assign outputs[2532] = (layer0_outputs[4108]) & ~(layer0_outputs[1448]);
    assign outputs[2533] = (layer0_outputs[3792]) & (layer0_outputs[2817]);
    assign outputs[2534] = ~(layer0_outputs[3280]);
    assign outputs[2535] = ~(layer0_outputs[1562]);
    assign outputs[2536] = layer0_outputs[1972];
    assign outputs[2537] = (layer0_outputs[1528]) & ~(layer0_outputs[2471]);
    assign outputs[2538] = ~(layer0_outputs[3020]);
    assign outputs[2539] = layer0_outputs[743];
    assign outputs[2540] = (layer0_outputs[3288]) & ~(layer0_outputs[3927]);
    assign outputs[2541] = ~((layer0_outputs[1899]) ^ (layer0_outputs[3505]));
    assign outputs[2542] = layer0_outputs[4043];
    assign outputs[2543] = layer0_outputs[366];
    assign outputs[2544] = (layer0_outputs[3837]) ^ (layer0_outputs[1526]);
    assign outputs[2545] = ~(layer0_outputs[1447]);
    assign outputs[2546] = ~(layer0_outputs[4574]);
    assign outputs[2547] = ~((layer0_outputs[3135]) & (layer0_outputs[1218]));
    assign outputs[2548] = layer0_outputs[956];
    assign outputs[2549] = (layer0_outputs[1747]) & ~(layer0_outputs[3265]);
    assign outputs[2550] = (layer0_outputs[41]) ^ (layer0_outputs[3581]);
    assign outputs[2551] = ~((layer0_outputs[3385]) ^ (layer0_outputs[579]));
    assign outputs[2552] = 1'b0;
    assign outputs[2553] = ~((layer0_outputs[3167]) ^ (layer0_outputs[3057]));
    assign outputs[2554] = ~((layer0_outputs[126]) | (layer0_outputs[4962]));
    assign outputs[2555] = ~(layer0_outputs[229]);
    assign outputs[2556] = ~(layer0_outputs[4225]);
    assign outputs[2557] = (layer0_outputs[4640]) ^ (layer0_outputs[3620]);
    assign outputs[2558] = layer0_outputs[4341];
    assign outputs[2559] = (layer0_outputs[3632]) & (layer0_outputs[227]);
    assign outputs[2560] = (layer0_outputs[3083]) | (layer0_outputs[545]);
    assign outputs[2561] = (layer0_outputs[3484]) & ~(layer0_outputs[1185]);
    assign outputs[2562] = ~((layer0_outputs[4733]) ^ (layer0_outputs[1705]));
    assign outputs[2563] = layer0_outputs[4627];
    assign outputs[2564] = ~((layer0_outputs[621]) ^ (layer0_outputs[1928]));
    assign outputs[2565] = ~((layer0_outputs[4177]) & (layer0_outputs[4130]));
    assign outputs[2566] = (layer0_outputs[4105]) ^ (layer0_outputs[68]);
    assign outputs[2567] = ~((layer0_outputs[940]) ^ (layer0_outputs[443]));
    assign outputs[2568] = layer0_outputs[208];
    assign outputs[2569] = ~(layer0_outputs[1004]);
    assign outputs[2570] = layer0_outputs[4428];
    assign outputs[2571] = layer0_outputs[3925];
    assign outputs[2572] = ~((layer0_outputs[4603]) | (layer0_outputs[3531]));
    assign outputs[2573] = layer0_outputs[4005];
    assign outputs[2574] = layer0_outputs[3150];
    assign outputs[2575] = layer0_outputs[3669];
    assign outputs[2576] = ~(layer0_outputs[2288]);
    assign outputs[2577] = layer0_outputs[4178];
    assign outputs[2578] = ~((layer0_outputs[626]) | (layer0_outputs[2729]));
    assign outputs[2579] = (layer0_outputs[4683]) & ~(layer0_outputs[5010]);
    assign outputs[2580] = ~((layer0_outputs[1634]) | (layer0_outputs[3358]));
    assign outputs[2581] = layer0_outputs[3087];
    assign outputs[2582] = ~(layer0_outputs[958]);
    assign outputs[2583] = ~((layer0_outputs[2325]) | (layer0_outputs[904]));
    assign outputs[2584] = (layer0_outputs[3968]) & ~(layer0_outputs[4241]);
    assign outputs[2585] = ~((layer0_outputs[2103]) | (layer0_outputs[508]));
    assign outputs[2586] = (layer0_outputs[4165]) & (layer0_outputs[4768]);
    assign outputs[2587] = layer0_outputs[3260];
    assign outputs[2588] = (layer0_outputs[3576]) & (layer0_outputs[583]);
    assign outputs[2589] = ~(layer0_outputs[3653]) | (layer0_outputs[2344]);
    assign outputs[2590] = ~(layer0_outputs[310]) | (layer0_outputs[2134]);
    assign outputs[2591] = ~(layer0_outputs[2242]);
    assign outputs[2592] = (layer0_outputs[2534]) & (layer0_outputs[2324]);
    assign outputs[2593] = ~(layer0_outputs[349]);
    assign outputs[2594] = ~(layer0_outputs[1532]);
    assign outputs[2595] = ~(layer0_outputs[360]);
    assign outputs[2596] = layer0_outputs[3503];
    assign outputs[2597] = ~((layer0_outputs[1609]) ^ (layer0_outputs[4342]));
    assign outputs[2598] = ~((layer0_outputs[1898]) ^ (layer0_outputs[233]));
    assign outputs[2599] = (layer0_outputs[1025]) & ~(layer0_outputs[4127]);
    assign outputs[2600] = ~(layer0_outputs[1378]);
    assign outputs[2601] = (layer0_outputs[3697]) & ~(layer0_outputs[254]);
    assign outputs[2602] = layer0_outputs[3182];
    assign outputs[2603] = layer0_outputs[1904];
    assign outputs[2604] = ~(layer0_outputs[1088]);
    assign outputs[2605] = ~(layer0_outputs[3990]);
    assign outputs[2606] = ~((layer0_outputs[3293]) ^ (layer0_outputs[4092]));
    assign outputs[2607] = ~(layer0_outputs[926]);
    assign outputs[2608] = ~(layer0_outputs[598]);
    assign outputs[2609] = ~(layer0_outputs[783]) | (layer0_outputs[3568]);
    assign outputs[2610] = ~(layer0_outputs[1600]);
    assign outputs[2611] = ~((layer0_outputs[3189]) ^ (layer0_outputs[529]));
    assign outputs[2612] = ~((layer0_outputs[2838]) | (layer0_outputs[503]));
    assign outputs[2613] = ~((layer0_outputs[79]) & (layer0_outputs[1447]));
    assign outputs[2614] = layer0_outputs[4004];
    assign outputs[2615] = ~(layer0_outputs[2345]);
    assign outputs[2616] = (layer0_outputs[4261]) & ~(layer0_outputs[4197]);
    assign outputs[2617] = ~(layer0_outputs[2320]) | (layer0_outputs[1756]);
    assign outputs[2618] = (layer0_outputs[4811]) ^ (layer0_outputs[1468]);
    assign outputs[2619] = (layer0_outputs[620]) | (layer0_outputs[2273]);
    assign outputs[2620] = ~(layer0_outputs[1283]) | (layer0_outputs[4937]);
    assign outputs[2621] = ~(layer0_outputs[3104]);
    assign outputs[2622] = ~((layer0_outputs[1803]) ^ (layer0_outputs[3176]));
    assign outputs[2623] = (layer0_outputs[2697]) | (layer0_outputs[1587]);
    assign outputs[2624] = ~(layer0_outputs[57]) | (layer0_outputs[2480]);
    assign outputs[2625] = ~(layer0_outputs[1425]);
    assign outputs[2626] = ~((layer0_outputs[385]) ^ (layer0_outputs[520]));
    assign outputs[2627] = (layer0_outputs[4985]) & ~(layer0_outputs[2347]);
    assign outputs[2628] = ~((layer0_outputs[471]) ^ (layer0_outputs[4599]));
    assign outputs[2629] = (layer0_outputs[1816]) & (layer0_outputs[1906]);
    assign outputs[2630] = ~(layer0_outputs[3457]);
    assign outputs[2631] = (layer0_outputs[3322]) | (layer0_outputs[1021]);
    assign outputs[2632] = ~((layer0_outputs[3296]) | (layer0_outputs[414]));
    assign outputs[2633] = (layer0_outputs[1411]) ^ (layer0_outputs[3143]);
    assign outputs[2634] = ~((layer0_outputs[24]) | (layer0_outputs[2738]));
    assign outputs[2635] = ~((layer0_outputs[3540]) ^ (layer0_outputs[4225]));
    assign outputs[2636] = ~(layer0_outputs[3997]) | (layer0_outputs[1346]);
    assign outputs[2637] = ~((layer0_outputs[737]) ^ (layer0_outputs[1879]));
    assign outputs[2638] = ~((layer0_outputs[4491]) ^ (layer0_outputs[1478]));
    assign outputs[2639] = ~(layer0_outputs[4315]);
    assign outputs[2640] = ~(layer0_outputs[47]);
    assign outputs[2641] = layer0_outputs[2929];
    assign outputs[2642] = ~(layer0_outputs[262]) | (layer0_outputs[2322]);
    assign outputs[2643] = (layer0_outputs[1636]) & (layer0_outputs[2357]);
    assign outputs[2644] = 1'b0;
    assign outputs[2645] = ~(layer0_outputs[3745]) | (layer0_outputs[1131]);
    assign outputs[2646] = ~(layer0_outputs[1789]) | (layer0_outputs[4044]);
    assign outputs[2647] = (layer0_outputs[234]) & ~(layer0_outputs[2967]);
    assign outputs[2648] = (layer0_outputs[401]) ^ (layer0_outputs[2780]);
    assign outputs[2649] = ~(layer0_outputs[2435]);
    assign outputs[2650] = ~(layer0_outputs[3502]) | (layer0_outputs[3726]);
    assign outputs[2651] = layer0_outputs[2781];
    assign outputs[2652] = 1'b1;
    assign outputs[2653] = layer0_outputs[1208];
    assign outputs[2654] = ~((layer0_outputs[4684]) ^ (layer0_outputs[2114]));
    assign outputs[2655] = ~((layer0_outputs[139]) | (layer0_outputs[4778]));
    assign outputs[2656] = ~((layer0_outputs[4125]) ^ (layer0_outputs[880]));
    assign outputs[2657] = layer0_outputs[442];
    assign outputs[2658] = layer0_outputs[1709];
    assign outputs[2659] = layer0_outputs[3034];
    assign outputs[2660] = (layer0_outputs[4862]) & (layer0_outputs[3973]);
    assign outputs[2661] = layer0_outputs[1134];
    assign outputs[2662] = ~(layer0_outputs[3041]) | (layer0_outputs[2408]);
    assign outputs[2663] = layer0_outputs[4536];
    assign outputs[2664] = ~(layer0_outputs[4912]);
    assign outputs[2665] = layer0_outputs[3881];
    assign outputs[2666] = ~(layer0_outputs[1206]);
    assign outputs[2667] = ~((layer0_outputs[4024]) | (layer0_outputs[563]));
    assign outputs[2668] = ~((layer0_outputs[4678]) & (layer0_outputs[1111]));
    assign outputs[2669] = ~(layer0_outputs[1184]) | (layer0_outputs[2668]);
    assign outputs[2670] = layer0_outputs[4727];
    assign outputs[2671] = layer0_outputs[1149];
    assign outputs[2672] = ~(layer0_outputs[2937]);
    assign outputs[2673] = layer0_outputs[3682];
    assign outputs[2674] = ~((layer0_outputs[1567]) | (layer0_outputs[5007]));
    assign outputs[2675] = (layer0_outputs[1257]) & ~(layer0_outputs[3883]);
    assign outputs[2676] = (layer0_outputs[2842]) ^ (layer0_outputs[4487]);
    assign outputs[2677] = layer0_outputs[4698];
    assign outputs[2678] = (layer0_outputs[4478]) & (layer0_outputs[1568]);
    assign outputs[2679] = (layer0_outputs[3129]) & (layer0_outputs[4974]);
    assign outputs[2680] = (layer0_outputs[2617]) ^ (layer0_outputs[4990]);
    assign outputs[2681] = (layer0_outputs[4214]) & ~(layer0_outputs[2732]);
    assign outputs[2682] = (layer0_outputs[2098]) & ~(layer0_outputs[5009]);
    assign outputs[2683] = ~(layer0_outputs[101]);
    assign outputs[2684] = ~(layer0_outputs[1312]);
    assign outputs[2685] = (layer0_outputs[4261]) ^ (layer0_outputs[3358]);
    assign outputs[2686] = ~((layer0_outputs[3235]) & (layer0_outputs[4959]));
    assign outputs[2687] = ~((layer0_outputs[306]) | (layer0_outputs[2586]));
    assign outputs[2688] = ~(layer0_outputs[1225]);
    assign outputs[2689] = (layer0_outputs[4756]) & ~(layer0_outputs[4563]);
    assign outputs[2690] = layer0_outputs[3264];
    assign outputs[2691] = ~(layer0_outputs[1224]) | (layer0_outputs[3756]);
    assign outputs[2692] = (layer0_outputs[1426]) & (layer0_outputs[3134]);
    assign outputs[2693] = (layer0_outputs[1235]) | (layer0_outputs[3749]);
    assign outputs[2694] = ~(layer0_outputs[561]);
    assign outputs[2695] = layer0_outputs[1290];
    assign outputs[2696] = (layer0_outputs[608]) ^ (layer0_outputs[1637]);
    assign outputs[2697] = ~((layer0_outputs[3541]) ^ (layer0_outputs[686]));
    assign outputs[2698] = (layer0_outputs[152]) ^ (layer0_outputs[2743]);
    assign outputs[2699] = (layer0_outputs[327]) ^ (layer0_outputs[2913]);
    assign outputs[2700] = layer0_outputs[1671];
    assign outputs[2701] = ~((layer0_outputs[2494]) ^ (layer0_outputs[3377]));
    assign outputs[2702] = (layer0_outputs[3549]) ^ (layer0_outputs[4303]);
    assign outputs[2703] = ~(layer0_outputs[2297]) | (layer0_outputs[4981]);
    assign outputs[2704] = ~(layer0_outputs[4230]);
    assign outputs[2705] = layer0_outputs[5063];
    assign outputs[2706] = layer0_outputs[3183];
    assign outputs[2707] = ~(layer0_outputs[4625]);
    assign outputs[2708] = ~((layer0_outputs[3195]) ^ (layer0_outputs[3503]));
    assign outputs[2709] = ~((layer0_outputs[3508]) ^ (layer0_outputs[2366]));
    assign outputs[2710] = ~((layer0_outputs[4550]) & (layer0_outputs[2430]));
    assign outputs[2711] = ~(layer0_outputs[1729]);
    assign outputs[2712] = (layer0_outputs[2932]) | (layer0_outputs[3765]);
    assign outputs[2713] = ~(layer0_outputs[2368]);
    assign outputs[2714] = (layer0_outputs[62]) | (layer0_outputs[226]);
    assign outputs[2715] = (layer0_outputs[220]) & (layer0_outputs[2371]);
    assign outputs[2716] = ~((layer0_outputs[1684]) ^ (layer0_outputs[1292]));
    assign outputs[2717] = (layer0_outputs[2392]) ^ (layer0_outputs[1020]);
    assign outputs[2718] = ~(layer0_outputs[4714]);
    assign outputs[2719] = (layer0_outputs[1518]) & ~(layer0_outputs[391]);
    assign outputs[2720] = ~((layer0_outputs[3467]) ^ (layer0_outputs[2827]));
    assign outputs[2721] = (layer0_outputs[660]) ^ (layer0_outputs[4675]);
    assign outputs[2722] = layer0_outputs[4820];
    assign outputs[2723] = ~(layer0_outputs[3920]) | (layer0_outputs[3569]);
    assign outputs[2724] = ~(layer0_outputs[4527]);
    assign outputs[2725] = (layer0_outputs[4395]) ^ (layer0_outputs[3957]);
    assign outputs[2726] = (layer0_outputs[374]) & ~(layer0_outputs[4344]);
    assign outputs[2727] = (layer0_outputs[1819]) & ~(layer0_outputs[1555]);
    assign outputs[2728] = ~(layer0_outputs[4111]);
    assign outputs[2729] = ~((layer0_outputs[4407]) ^ (layer0_outputs[1159]));
    assign outputs[2730] = ~(layer0_outputs[2686]);
    assign outputs[2731] = (layer0_outputs[4796]) ^ (layer0_outputs[3491]);
    assign outputs[2732] = layer0_outputs[86];
    assign outputs[2733] = ~(layer0_outputs[4449]);
    assign outputs[2734] = ~(layer0_outputs[3324]);
    assign outputs[2735] = (layer0_outputs[2208]) | (layer0_outputs[1147]);
    assign outputs[2736] = layer0_outputs[4517];
    assign outputs[2737] = layer0_outputs[3200];
    assign outputs[2738] = ~((layer0_outputs[1931]) & (layer0_outputs[3899]));
    assign outputs[2739] = ~((layer0_outputs[976]) | (layer0_outputs[638]));
    assign outputs[2740] = ~((layer0_outputs[3137]) & (layer0_outputs[5017]));
    assign outputs[2741] = layer0_outputs[8];
    assign outputs[2742] = ~(layer0_outputs[4847]);
    assign outputs[2743] = ~((layer0_outputs[315]) ^ (layer0_outputs[456]));
    assign outputs[2744] = (layer0_outputs[2854]) & ~(layer0_outputs[3098]);
    assign outputs[2745] = ~(layer0_outputs[91]);
    assign outputs[2746] = (layer0_outputs[4579]) & ~(layer0_outputs[1428]);
    assign outputs[2747] = ~(layer0_outputs[713]) | (layer0_outputs[3449]);
    assign outputs[2748] = ~(layer0_outputs[3686]) | (layer0_outputs[416]);
    assign outputs[2749] = (layer0_outputs[4718]) & (layer0_outputs[4165]);
    assign outputs[2750] = layer0_outputs[1172];
    assign outputs[2751] = ~((layer0_outputs[2722]) | (layer0_outputs[1939]));
    assign outputs[2752] = layer0_outputs[4426];
    assign outputs[2753] = (layer0_outputs[5045]) ^ (layer0_outputs[3960]);
    assign outputs[2754] = ~((layer0_outputs[134]) | (layer0_outputs[4828]));
    assign outputs[2755] = layer0_outputs[1143];
    assign outputs[2756] = ~(layer0_outputs[3660]);
    assign outputs[2757] = layer0_outputs[1348];
    assign outputs[2758] = layer0_outputs[5038];
    assign outputs[2759] = (layer0_outputs[4254]) & ~(layer0_outputs[1528]);
    assign outputs[2760] = (layer0_outputs[4649]) & ~(layer0_outputs[1375]);
    assign outputs[2761] = (layer0_outputs[4591]) ^ (layer0_outputs[4976]);
    assign outputs[2762] = (layer0_outputs[4992]) | (layer0_outputs[2399]);
    assign outputs[2763] = ~(layer0_outputs[3893]);
    assign outputs[2764] = (layer0_outputs[2078]) ^ (layer0_outputs[1574]);
    assign outputs[2765] = layer0_outputs[3754];
    assign outputs[2766] = ~(layer0_outputs[3793]);
    assign outputs[2767] = ~(layer0_outputs[842]);
    assign outputs[2768] = ~((layer0_outputs[2107]) ^ (layer0_outputs[1928]));
    assign outputs[2769] = layer0_outputs[2894];
    assign outputs[2770] = ~((layer0_outputs[3921]) ^ (layer0_outputs[4783]));
    assign outputs[2771] = layer0_outputs[1003];
    assign outputs[2772] = ~((layer0_outputs[4351]) ^ (layer0_outputs[4231]));
    assign outputs[2773] = ~(layer0_outputs[2990]);
    assign outputs[2774] = layer0_outputs[381];
    assign outputs[2775] = ~(layer0_outputs[3684]);
    assign outputs[2776] = ~((layer0_outputs[3420]) & (layer0_outputs[29]));
    assign outputs[2777] = (layer0_outputs[4397]) & (layer0_outputs[2141]);
    assign outputs[2778] = ~(layer0_outputs[4115]) | (layer0_outputs[4741]);
    assign outputs[2779] = ~((layer0_outputs[4582]) & (layer0_outputs[4929]));
    assign outputs[2780] = ~(layer0_outputs[556]);
    assign outputs[2781] = ~((layer0_outputs[467]) & (layer0_outputs[2798]));
    assign outputs[2782] = layer0_outputs[4833];
    assign outputs[2783] = ~(layer0_outputs[644]);
    assign outputs[2784] = layer0_outputs[4748];
    assign outputs[2785] = layer0_outputs[217];
    assign outputs[2786] = ~((layer0_outputs[2932]) | (layer0_outputs[3738]));
    assign outputs[2787] = layer0_outputs[2615];
    assign outputs[2788] = (layer0_outputs[5057]) | (layer0_outputs[1449]);
    assign outputs[2789] = ~(layer0_outputs[2709]) | (layer0_outputs[2902]);
    assign outputs[2790] = ~(layer0_outputs[576]);
    assign outputs[2791] = ~((layer0_outputs[4047]) & (layer0_outputs[1165]));
    assign outputs[2792] = (layer0_outputs[50]) & ~(layer0_outputs[4849]);
    assign outputs[2793] = ~(layer0_outputs[3431]) | (layer0_outputs[4532]);
    assign outputs[2794] = (layer0_outputs[4524]) & ~(layer0_outputs[1004]);
    assign outputs[2795] = ~(layer0_outputs[2585]);
    assign outputs[2796] = ~((layer0_outputs[3663]) ^ (layer0_outputs[2531]));
    assign outputs[2797] = ~(layer0_outputs[4279]);
    assign outputs[2798] = ~(layer0_outputs[373]) | (layer0_outputs[1392]);
    assign outputs[2799] = ~(layer0_outputs[4915]);
    assign outputs[2800] = layer0_outputs[4599];
    assign outputs[2801] = layer0_outputs[108];
    assign outputs[2802] = ~((layer0_outputs[2076]) ^ (layer0_outputs[2600]));
    assign outputs[2803] = ~((layer0_outputs[4549]) ^ (layer0_outputs[41]));
    assign outputs[2804] = (layer0_outputs[3119]) ^ (layer0_outputs[867]);
    assign outputs[2805] = (layer0_outputs[2634]) & (layer0_outputs[5117]);
    assign outputs[2806] = ~((layer0_outputs[4629]) ^ (layer0_outputs[3513]));
    assign outputs[2807] = ~(layer0_outputs[4747]);
    assign outputs[2808] = ~((layer0_outputs[2881]) ^ (layer0_outputs[1745]));
    assign outputs[2809] = ~((layer0_outputs[997]) ^ (layer0_outputs[4559]));
    assign outputs[2810] = layer0_outputs[3952];
    assign outputs[2811] = ~(layer0_outputs[82]);
    assign outputs[2812] = ~((layer0_outputs[204]) ^ (layer0_outputs[1367]));
    assign outputs[2813] = ~((layer0_outputs[2382]) | (layer0_outputs[2899]));
    assign outputs[2814] = ~(layer0_outputs[143]) | (layer0_outputs[4681]);
    assign outputs[2815] = layer0_outputs[1880];
    assign outputs[2816] = ~(layer0_outputs[3587]);
    assign outputs[2817] = layer0_outputs[2943];
    assign outputs[2818] = ~(layer0_outputs[4266]);
    assign outputs[2819] = ~(layer0_outputs[599]) | (layer0_outputs[3475]);
    assign outputs[2820] = layer0_outputs[1983];
    assign outputs[2821] = ~((layer0_outputs[3687]) ^ (layer0_outputs[3969]));
    assign outputs[2822] = layer0_outputs[3336];
    assign outputs[2823] = (layer0_outputs[323]) & (layer0_outputs[2669]);
    assign outputs[2824] = (layer0_outputs[2934]) & ~(layer0_outputs[2022]);
    assign outputs[2825] = (layer0_outputs[3232]) & (layer0_outputs[1561]);
    assign outputs[2826] = ~((layer0_outputs[2046]) ^ (layer0_outputs[4850]));
    assign outputs[2827] = layer0_outputs[567];
    assign outputs[2828] = (layer0_outputs[4912]) & ~(layer0_outputs[51]);
    assign outputs[2829] = ~(layer0_outputs[4810]);
    assign outputs[2830] = layer0_outputs[2023];
    assign outputs[2831] = layer0_outputs[283];
    assign outputs[2832] = layer0_outputs[796];
    assign outputs[2833] = (layer0_outputs[1730]) & ~(layer0_outputs[1442]);
    assign outputs[2834] = (layer0_outputs[3291]) ^ (layer0_outputs[4374]);
    assign outputs[2835] = (layer0_outputs[1994]) & ~(layer0_outputs[128]);
    assign outputs[2836] = (layer0_outputs[2569]) & (layer0_outputs[1091]);
    assign outputs[2837] = (layer0_outputs[518]) & (layer0_outputs[150]);
    assign outputs[2838] = ~((layer0_outputs[4944]) | (layer0_outputs[1657]));
    assign outputs[2839] = (layer0_outputs[5063]) & ~(layer0_outputs[1800]);
    assign outputs[2840] = layer0_outputs[1453];
    assign outputs[2841] = layer0_outputs[216];
    assign outputs[2842] = layer0_outputs[4842];
    assign outputs[2843] = layer0_outputs[3010];
    assign outputs[2844] = (layer0_outputs[739]) ^ (layer0_outputs[680]);
    assign outputs[2845] = ~((layer0_outputs[2521]) ^ (layer0_outputs[1481]));
    assign outputs[2846] = ~((layer0_outputs[3718]) ^ (layer0_outputs[1577]));
    assign outputs[2847] = ~(layer0_outputs[955]);
    assign outputs[2848] = ~((layer0_outputs[3542]) | (layer0_outputs[3589]));
    assign outputs[2849] = ~(layer0_outputs[228]);
    assign outputs[2850] = ~(layer0_outputs[1524]);
    assign outputs[2851] = (layer0_outputs[1129]) & ~(layer0_outputs[3926]);
    assign outputs[2852] = (layer0_outputs[758]) ^ (layer0_outputs[1566]);
    assign outputs[2853] = ~((layer0_outputs[1683]) ^ (layer0_outputs[3600]));
    assign outputs[2854] = ~(layer0_outputs[56]) | (layer0_outputs[2905]);
    assign outputs[2855] = ~((layer0_outputs[185]) ^ (layer0_outputs[573]));
    assign outputs[2856] = ~(layer0_outputs[4939]);
    assign outputs[2857] = ~(layer0_outputs[454]);
    assign outputs[2858] = ~((layer0_outputs[2185]) | (layer0_outputs[1243]));
    assign outputs[2859] = layer0_outputs[3892];
    assign outputs[2860] = ~((layer0_outputs[2579]) ^ (layer0_outputs[2837]));
    assign outputs[2861] = layer0_outputs[3402];
    assign outputs[2862] = (layer0_outputs[890]) ^ (layer0_outputs[1104]);
    assign outputs[2863] = (layer0_outputs[1645]) ^ (layer0_outputs[1883]);
    assign outputs[2864] = ~(layer0_outputs[2741]) | (layer0_outputs[3415]);
    assign outputs[2865] = ~((layer0_outputs[1945]) & (layer0_outputs[4713]));
    assign outputs[2866] = ~(layer0_outputs[3704]) | (layer0_outputs[3529]);
    assign outputs[2867] = ~((layer0_outputs[2644]) | (layer0_outputs[2126]));
    assign outputs[2868] = ~((layer0_outputs[3820]) ^ (layer0_outputs[4468]));
    assign outputs[2869] = layer0_outputs[3510];
    assign outputs[2870] = layer0_outputs[63];
    assign outputs[2871] = layer0_outputs[364];
    assign outputs[2872] = ~(layer0_outputs[148]);
    assign outputs[2873] = (layer0_outputs[513]) & ~(layer0_outputs[1107]);
    assign outputs[2874] = 1'b1;
    assign outputs[2875] = (layer0_outputs[1671]) & (layer0_outputs[1857]);
    assign outputs[2876] = ~((layer0_outputs[1427]) | (layer0_outputs[3192]));
    assign outputs[2877] = (layer0_outputs[3409]) & ~(layer0_outputs[125]);
    assign outputs[2878] = ~((layer0_outputs[140]) | (layer0_outputs[1910]));
    assign outputs[2879] = ~((layer0_outputs[3794]) ^ (layer0_outputs[3422]));
    assign outputs[2880] = ~((layer0_outputs[1583]) & (layer0_outputs[648]));
    assign outputs[2881] = ~(layer0_outputs[1817]);
    assign outputs[2882] = (layer0_outputs[1372]) ^ (layer0_outputs[481]);
    assign outputs[2883] = ~((layer0_outputs[116]) ^ (layer0_outputs[2333]));
    assign outputs[2884] = layer0_outputs[89];
    assign outputs[2885] = ~((layer0_outputs[3804]) ^ (layer0_outputs[301]));
    assign outputs[2886] = ~(layer0_outputs[4140]) | (layer0_outputs[4609]);
    assign outputs[2887] = (layer0_outputs[156]) & ~(layer0_outputs[174]);
    assign outputs[2888] = ~(layer0_outputs[2373]);
    assign outputs[2889] = layer0_outputs[3089];
    assign outputs[2890] = layer0_outputs[584];
    assign outputs[2891] = ~(layer0_outputs[871]);
    assign outputs[2892] = layer0_outputs[4180];
    assign outputs[2893] = ~((layer0_outputs[4383]) ^ (layer0_outputs[1416]));
    assign outputs[2894] = ~(layer0_outputs[3312]);
    assign outputs[2895] = layer0_outputs[1321];
    assign outputs[2896] = (layer0_outputs[1405]) | (layer0_outputs[4853]);
    assign outputs[2897] = layer0_outputs[2928];
    assign outputs[2898] = layer0_outputs[4984];
    assign outputs[2899] = ~((layer0_outputs[1698]) | (layer0_outputs[3939]));
    assign outputs[2900] = layer0_outputs[753];
    assign outputs[2901] = ~((layer0_outputs[26]) | (layer0_outputs[2276]));
    assign outputs[2902] = ~((layer0_outputs[3052]) & (layer0_outputs[4343]));
    assign outputs[2903] = ~(layer0_outputs[1543]) | (layer0_outputs[899]);
    assign outputs[2904] = ~((layer0_outputs[504]) ^ (layer0_outputs[2661]));
    assign outputs[2905] = ~((layer0_outputs[2548]) | (layer0_outputs[2385]));
    assign outputs[2906] = ~((layer0_outputs[288]) & (layer0_outputs[4617]));
    assign outputs[2907] = ~(layer0_outputs[2747]);
    assign outputs[2908] = (layer0_outputs[3940]) & ~(layer0_outputs[3278]);
    assign outputs[2909] = ~(layer0_outputs[2429]);
    assign outputs[2910] = ~((layer0_outputs[1855]) & (layer0_outputs[553]));
    assign outputs[2911] = ~(layer0_outputs[2560]);
    assign outputs[2912] = layer0_outputs[1510];
    assign outputs[2913] = layer0_outputs[4175];
    assign outputs[2914] = ~((layer0_outputs[4696]) ^ (layer0_outputs[4215]));
    assign outputs[2915] = ~(layer0_outputs[3840]);
    assign outputs[2916] = ~((layer0_outputs[382]) ^ (layer0_outputs[2442]));
    assign outputs[2917] = (layer0_outputs[528]) ^ (layer0_outputs[3971]);
    assign outputs[2918] = ~((layer0_outputs[3472]) & (layer0_outputs[3212]));
    assign outputs[2919] = ~(layer0_outputs[3012]) | (layer0_outputs[4587]);
    assign outputs[2920] = layer0_outputs[2881];
    assign outputs[2921] = ~(layer0_outputs[2219]);
    assign outputs[2922] = ~(layer0_outputs[3652]) | (layer0_outputs[377]);
    assign outputs[2923] = layer0_outputs[1431];
    assign outputs[2924] = layer0_outputs[3945];
    assign outputs[2925] = ~(layer0_outputs[2826]);
    assign outputs[2926] = (layer0_outputs[4876]) | (layer0_outputs[3788]);
    assign outputs[2927] = ~(layer0_outputs[1753]);
    assign outputs[2928] = layer0_outputs[3603];
    assign outputs[2929] = (layer0_outputs[710]) ^ (layer0_outputs[2441]);
    assign outputs[2930] = ~(layer0_outputs[3915]);
    assign outputs[2931] = (layer0_outputs[2972]) ^ (layer0_outputs[1314]);
    assign outputs[2932] = (layer0_outputs[1826]) ^ (layer0_outputs[3276]);
    assign outputs[2933] = ~((layer0_outputs[2346]) ^ (layer0_outputs[2581]));
    assign outputs[2934] = (layer0_outputs[1879]) ^ (layer0_outputs[4256]);
    assign outputs[2935] = layer0_outputs[4577];
    assign outputs[2936] = ~(layer0_outputs[1798]);
    assign outputs[2937] = ~(layer0_outputs[3805]) | (layer0_outputs[4981]);
    assign outputs[2938] = ~((layer0_outputs[2210]) | (layer0_outputs[3499]));
    assign outputs[2939] = (layer0_outputs[2911]) & ~(layer0_outputs[1530]);
    assign outputs[2940] = (layer0_outputs[4779]) & ~(layer0_outputs[3844]);
    assign outputs[2941] = (layer0_outputs[1290]) & (layer0_outputs[2628]);
    assign outputs[2942] = (layer0_outputs[3247]) & (layer0_outputs[4293]);
    assign outputs[2943] = ~((layer0_outputs[682]) ^ (layer0_outputs[1419]));
    assign outputs[2944] = (layer0_outputs[4827]) ^ (layer0_outputs[900]);
    assign outputs[2945] = ~(layer0_outputs[1630]);
    assign outputs[2946] = ~((layer0_outputs[896]) & (layer0_outputs[94]));
    assign outputs[2947] = (layer0_outputs[2803]) & ~(layer0_outputs[0]);
    assign outputs[2948] = ~(layer0_outputs[3330]);
    assign outputs[2949] = ~(layer0_outputs[4210]) | (layer0_outputs[2867]);
    assign outputs[2950] = ~(layer0_outputs[3552]);
    assign outputs[2951] = ~(layer0_outputs[1218]);
    assign outputs[2952] = ~((layer0_outputs[4630]) ^ (layer0_outputs[2349]));
    assign outputs[2953] = ~(layer0_outputs[4476]);
    assign outputs[2954] = ~(layer0_outputs[4968]);
    assign outputs[2955] = layer0_outputs[779];
    assign outputs[2956] = (layer0_outputs[4582]) ^ (layer0_outputs[1070]);
    assign outputs[2957] = (layer0_outputs[3631]) & ~(layer0_outputs[1582]);
    assign outputs[2958] = layer0_outputs[160];
    assign outputs[2959] = ~(layer0_outputs[523]);
    assign outputs[2960] = (layer0_outputs[808]) ^ (layer0_outputs[3812]);
    assign outputs[2961] = layer0_outputs[612];
    assign outputs[2962] = ~(layer0_outputs[2150]);
    assign outputs[2963] = ~(layer0_outputs[1838]);
    assign outputs[2964] = ~(layer0_outputs[3871]);
    assign outputs[2965] = (layer0_outputs[287]) | (layer0_outputs[4263]);
    assign outputs[2966] = ~((layer0_outputs[1166]) ^ (layer0_outputs[4212]));
    assign outputs[2967] = ~(layer0_outputs[1081]);
    assign outputs[2968] = ~(layer0_outputs[3261]);
    assign outputs[2969] = (layer0_outputs[4843]) & (layer0_outputs[283]);
    assign outputs[2970] = layer0_outputs[4820];
    assign outputs[2971] = layer0_outputs[612];
    assign outputs[2972] = ~(layer0_outputs[1387]) | (layer0_outputs[452]);
    assign outputs[2973] = ~((layer0_outputs[3661]) ^ (layer0_outputs[3275]));
    assign outputs[2974] = ~((layer0_outputs[1215]) & (layer0_outputs[2281]));
    assign outputs[2975] = (layer0_outputs[5101]) & ~(layer0_outputs[1872]);
    assign outputs[2976] = ~((layer0_outputs[24]) | (layer0_outputs[2180]));
    assign outputs[2977] = ~(layer0_outputs[4893]) | (layer0_outputs[997]);
    assign outputs[2978] = ~((layer0_outputs[3060]) ^ (layer0_outputs[224]));
    assign outputs[2979] = (layer0_outputs[4893]) | (layer0_outputs[336]);
    assign outputs[2980] = layer0_outputs[4122];
    assign outputs[2981] = layer0_outputs[119];
    assign outputs[2982] = (layer0_outputs[4788]) & ~(layer0_outputs[4350]);
    assign outputs[2983] = ~(layer0_outputs[4854]);
    assign outputs[2984] = (layer0_outputs[2788]) & (layer0_outputs[3554]);
    assign outputs[2985] = layer0_outputs[4135];
    assign outputs[2986] = ~((layer0_outputs[1584]) & (layer0_outputs[3372]));
    assign outputs[2987] = (layer0_outputs[2863]) & ~(layer0_outputs[2180]);
    assign outputs[2988] = (layer0_outputs[4564]) & (layer0_outputs[1941]);
    assign outputs[2989] = (layer0_outputs[1983]) ^ (layer0_outputs[3903]);
    assign outputs[2990] = layer0_outputs[3572];
    assign outputs[2991] = ~((layer0_outputs[3544]) ^ (layer0_outputs[4839]));
    assign outputs[2992] = layer0_outputs[4805];
    assign outputs[2993] = ~(layer0_outputs[1667]) | (layer0_outputs[1344]);
    assign outputs[2994] = (layer0_outputs[656]) & ~(layer0_outputs[607]);
    assign outputs[2995] = (layer0_outputs[2157]) & ~(layer0_outputs[4139]);
    assign outputs[2996] = ~((layer0_outputs[3594]) ^ (layer0_outputs[3887]));
    assign outputs[2997] = ~(layer0_outputs[988]) | (layer0_outputs[4205]);
    assign outputs[2998] = layer0_outputs[2784];
    assign outputs[2999] = layer0_outputs[1703];
    assign outputs[3000] = ~((layer0_outputs[1412]) | (layer0_outputs[1695]));
    assign outputs[3001] = (layer0_outputs[1108]) ^ (layer0_outputs[3624]);
    assign outputs[3002] = ~(layer0_outputs[3410]) | (layer0_outputs[4515]);
    assign outputs[3003] = (layer0_outputs[662]) | (layer0_outputs[4466]);
    assign outputs[3004] = layer0_outputs[3988];
    assign outputs[3005] = ~(layer0_outputs[3093]) | (layer0_outputs[2018]);
    assign outputs[3006] = ~((layer0_outputs[17]) ^ (layer0_outputs[600]));
    assign outputs[3007] = ~((layer0_outputs[4482]) & (layer0_outputs[3587]));
    assign outputs[3008] = ~(layer0_outputs[1461]);
    assign outputs[3009] = layer0_outputs[3610];
    assign outputs[3010] = ~((layer0_outputs[3854]) ^ (layer0_outputs[3826]));
    assign outputs[3011] = ~((layer0_outputs[883]) | (layer0_outputs[2912]));
    assign outputs[3012] = layer0_outputs[1238];
    assign outputs[3013] = ~(layer0_outputs[2504]);
    assign outputs[3014] = ~(layer0_outputs[3616]);
    assign outputs[3015] = ~(layer0_outputs[2453]) | (layer0_outputs[196]);
    assign outputs[3016] = layer0_outputs[942];
    assign outputs[3017] = (layer0_outputs[2338]) & (layer0_outputs[129]);
    assign outputs[3018] = (layer0_outputs[4055]) ^ (layer0_outputs[724]);
    assign outputs[3019] = (layer0_outputs[1399]) & ~(layer0_outputs[4552]);
    assign outputs[3020] = (layer0_outputs[3270]) & (layer0_outputs[3343]);
    assign outputs[3021] = ~((layer0_outputs[1711]) | (layer0_outputs[4828]));
    assign outputs[3022] = (layer0_outputs[4934]) | (layer0_outputs[2418]);
    assign outputs[3023] = (layer0_outputs[642]) & ~(layer0_outputs[4811]);
    assign outputs[3024] = (layer0_outputs[4126]) ^ (layer0_outputs[924]);
    assign outputs[3025] = layer0_outputs[1326];
    assign outputs[3026] = layer0_outputs[540];
    assign outputs[3027] = ~(layer0_outputs[3848]);
    assign outputs[3028] = ~(layer0_outputs[3042]) | (layer0_outputs[999]);
    assign outputs[3029] = (layer0_outputs[3528]) ^ (layer0_outputs[4129]);
    assign outputs[3030] = layer0_outputs[4461];
    assign outputs[3031] = ~(layer0_outputs[2469]);
    assign outputs[3032] = ~(layer0_outputs[2314]) | (layer0_outputs[2713]);
    assign outputs[3033] = layer0_outputs[4161];
    assign outputs[3034] = (layer0_outputs[2394]) & (layer0_outputs[2946]);
    assign outputs[3035] = 1'b0;
    assign outputs[3036] = ~((layer0_outputs[2984]) ^ (layer0_outputs[2715]));
    assign outputs[3037] = (layer0_outputs[4508]) ^ (layer0_outputs[473]);
    assign outputs[3038] = ~(layer0_outputs[2865]) | (layer0_outputs[4858]);
    assign outputs[3039] = ~(layer0_outputs[1995]);
    assign outputs[3040] = ~(layer0_outputs[4894]);
    assign outputs[3041] = layer0_outputs[944];
    assign outputs[3042] = ~((layer0_outputs[1583]) ^ (layer0_outputs[650]));
    assign outputs[3043] = ~(layer0_outputs[911]);
    assign outputs[3044] = layer0_outputs[3922];
    assign outputs[3045] = ~(layer0_outputs[140]) | (layer0_outputs[3494]);
    assign outputs[3046] = (layer0_outputs[1449]) | (layer0_outputs[1246]);
    assign outputs[3047] = layer0_outputs[4171];
    assign outputs[3048] = layer0_outputs[5032];
    assign outputs[3049] = ~(layer0_outputs[4527]);
    assign outputs[3050] = ~((layer0_outputs[1908]) ^ (layer0_outputs[1305]));
    assign outputs[3051] = layer0_outputs[366];
    assign outputs[3052] = ~(layer0_outputs[2266]);
    assign outputs[3053] = layer0_outputs[670];
    assign outputs[3054] = layer0_outputs[3929];
    assign outputs[3055] = layer0_outputs[4410];
    assign outputs[3056] = (layer0_outputs[4768]) ^ (layer0_outputs[5116]);
    assign outputs[3057] = ~(layer0_outputs[3948]);
    assign outputs[3058] = (layer0_outputs[4051]) ^ (layer0_outputs[1144]);
    assign outputs[3059] = ~(layer0_outputs[3849]);
    assign outputs[3060] = ~(layer0_outputs[2444]);
    assign outputs[3061] = ~(layer0_outputs[1690]) | (layer0_outputs[3512]);
    assign outputs[3062] = ~(layer0_outputs[4509]);
    assign outputs[3063] = layer0_outputs[447];
    assign outputs[3064] = (layer0_outputs[3154]) ^ (layer0_outputs[642]);
    assign outputs[3065] = ~((layer0_outputs[1357]) ^ (layer0_outputs[3703]));
    assign outputs[3066] = layer0_outputs[3875];
    assign outputs[3067] = ~((layer0_outputs[4096]) ^ (layer0_outputs[4523]));
    assign outputs[3068] = ~(layer0_outputs[3919]) | (layer0_outputs[3597]);
    assign outputs[3069] = ~(layer0_outputs[1018]) | (layer0_outputs[3263]);
    assign outputs[3070] = layer0_outputs[538];
    assign outputs[3071] = ~(layer0_outputs[599]);
    assign outputs[3072] = ~((layer0_outputs[1017]) & (layer0_outputs[1523]));
    assign outputs[3073] = (layer0_outputs[253]) & ~(layer0_outputs[1122]);
    assign outputs[3074] = ~(layer0_outputs[325]);
    assign outputs[3075] = ~((layer0_outputs[3555]) | (layer0_outputs[2302]));
    assign outputs[3076] = (layer0_outputs[4511]) & ~(layer0_outputs[38]);
    assign outputs[3077] = ~((layer0_outputs[1321]) | (layer0_outputs[2975]));
    assign outputs[3078] = layer0_outputs[2356];
    assign outputs[3079] = layer0_outputs[931];
    assign outputs[3080] = layer0_outputs[1252];
    assign outputs[3081] = (layer0_outputs[242]) ^ (layer0_outputs[268]);
    assign outputs[3082] = ~((layer0_outputs[1456]) & (layer0_outputs[1035]));
    assign outputs[3083] = layer0_outputs[374];
    assign outputs[3084] = ~((layer0_outputs[20]) ^ (layer0_outputs[526]));
    assign outputs[3085] = layer0_outputs[5082];
    assign outputs[3086] = ~((layer0_outputs[73]) & (layer0_outputs[3263]));
    assign outputs[3087] = layer0_outputs[2087];
    assign outputs[3088] = ~((layer0_outputs[291]) ^ (layer0_outputs[1429]));
    assign outputs[3089] = ~((layer0_outputs[3014]) ^ (layer0_outputs[207]));
    assign outputs[3090] = (layer0_outputs[3716]) & ~(layer0_outputs[3230]);
    assign outputs[3091] = (layer0_outputs[1992]) ^ (layer0_outputs[1015]);
    assign outputs[3092] = ~(layer0_outputs[5010]) | (layer0_outputs[4410]);
    assign outputs[3093] = (layer0_outputs[4123]) ^ (layer0_outputs[2315]);
    assign outputs[3094] = ~(layer0_outputs[238]);
    assign outputs[3095] = layer0_outputs[3917];
    assign outputs[3096] = (layer0_outputs[3121]) & (layer0_outputs[5018]);
    assign outputs[3097] = (layer0_outputs[3619]) ^ (layer0_outputs[1812]);
    assign outputs[3098] = (layer0_outputs[423]) | (layer0_outputs[2124]);
    assign outputs[3099] = (layer0_outputs[3301]) ^ (layer0_outputs[4588]);
    assign outputs[3100] = ~((layer0_outputs[903]) ^ (layer0_outputs[1024]));
    assign outputs[3101] = (layer0_outputs[2641]) & ~(layer0_outputs[824]);
    assign outputs[3102] = ~(layer0_outputs[873]);
    assign outputs[3103] = (layer0_outputs[2915]) & ~(layer0_outputs[2496]);
    assign outputs[3104] = ~((layer0_outputs[5061]) ^ (layer0_outputs[553]));
    assign outputs[3105] = (layer0_outputs[1265]) & ~(layer0_outputs[1920]);
    assign outputs[3106] = layer0_outputs[4520];
    assign outputs[3107] = (layer0_outputs[1997]) & (layer0_outputs[2104]);
    assign outputs[3108] = ~((layer0_outputs[1919]) & (layer0_outputs[2701]));
    assign outputs[3109] = (layer0_outputs[1689]) | (layer0_outputs[3962]);
    assign outputs[3110] = ~((layer0_outputs[2917]) | (layer0_outputs[146]));
    assign outputs[3111] = (layer0_outputs[19]) & ~(layer0_outputs[1]);
    assign outputs[3112] = ~(layer0_outputs[4613]);
    assign outputs[3113] = ~((layer0_outputs[572]) & (layer0_outputs[2221]));
    assign outputs[3114] = ~(layer0_outputs[3391]);
    assign outputs[3115] = ~(layer0_outputs[4238]);
    assign outputs[3116] = ~(layer0_outputs[1142]);
    assign outputs[3117] = (layer0_outputs[1216]) & ~(layer0_outputs[1342]);
    assign outputs[3118] = ~((layer0_outputs[4685]) ^ (layer0_outputs[2976]));
    assign outputs[3119] = layer0_outputs[2216];
    assign outputs[3120] = ~((layer0_outputs[677]) & (layer0_outputs[2259]));
    assign outputs[3121] = ~(layer0_outputs[365]);
    assign outputs[3122] = (layer0_outputs[4012]) & ~(layer0_outputs[4123]);
    assign outputs[3123] = ~(layer0_outputs[3638]);
    assign outputs[3124] = ~(layer0_outputs[4953]);
    assign outputs[3125] = ~(layer0_outputs[4611]);
    assign outputs[3126] = layer0_outputs[4816];
    assign outputs[3127] = ~(layer0_outputs[4479]);
    assign outputs[3128] = ~((layer0_outputs[4948]) | (layer0_outputs[10]));
    assign outputs[3129] = (layer0_outputs[3000]) | (layer0_outputs[1697]);
    assign outputs[3130] = ~(layer0_outputs[32]) | (layer0_outputs[1245]);
    assign outputs[3131] = ~((layer0_outputs[2994]) & (layer0_outputs[1139]));
    assign outputs[3132] = ~(layer0_outputs[4631]);
    assign outputs[3133] = ~((layer0_outputs[104]) ^ (layer0_outputs[5044]));
    assign outputs[3134] = ~(layer0_outputs[2101]);
    assign outputs[3135] = (layer0_outputs[4655]) ^ (layer0_outputs[254]);
    assign outputs[3136] = ~((layer0_outputs[2728]) ^ (layer0_outputs[3360]));
    assign outputs[3137] = ~((layer0_outputs[2636]) ^ (layer0_outputs[945]));
    assign outputs[3138] = layer0_outputs[1236];
    assign outputs[3139] = ~(layer0_outputs[4557]);
    assign outputs[3140] = (layer0_outputs[1745]) & ~(layer0_outputs[457]);
    assign outputs[3141] = ~(layer0_outputs[4146]);
    assign outputs[3142] = (layer0_outputs[4879]) & ~(layer0_outputs[3637]);
    assign outputs[3143] = ~(layer0_outputs[1552]);
    assign outputs[3144] = ~(layer0_outputs[308]);
    assign outputs[3145] = (layer0_outputs[4659]) & ~(layer0_outputs[380]);
    assign outputs[3146] = ~(layer0_outputs[569]);
    assign outputs[3147] = ~(layer0_outputs[1578]);
    assign outputs[3148] = (layer0_outputs[4614]) & (layer0_outputs[4703]);
    assign outputs[3149] = (layer0_outputs[3199]) & (layer0_outputs[4852]);
    assign outputs[3150] = layer0_outputs[399];
    assign outputs[3151] = layer0_outputs[2664];
    assign outputs[3152] = ~(layer0_outputs[986]);
    assign outputs[3153] = layer0_outputs[1551];
    assign outputs[3154] = ~(layer0_outputs[476]);
    assign outputs[3155] = ~((layer0_outputs[3716]) & (layer0_outputs[240]));
    assign outputs[3156] = ~(layer0_outputs[4719]);
    assign outputs[3157] = (layer0_outputs[3270]) ^ (layer0_outputs[4849]);
    assign outputs[3158] = ~(layer0_outputs[3780]);
    assign outputs[3159] = layer0_outputs[4078];
    assign outputs[3160] = ~(layer0_outputs[718]);
    assign outputs[3161] = ~(layer0_outputs[2671]);
    assign outputs[3162] = layer0_outputs[2913];
    assign outputs[3163] = ~((layer0_outputs[3249]) | (layer0_outputs[4113]));
    assign outputs[3164] = (layer0_outputs[2995]) ^ (layer0_outputs[1664]);
    assign outputs[3165] = ~((layer0_outputs[4623]) ^ (layer0_outputs[1064]));
    assign outputs[3166] = ~(layer0_outputs[3117]);
    assign outputs[3167] = layer0_outputs[2925];
    assign outputs[3168] = (layer0_outputs[2728]) & ~(layer0_outputs[4039]);
    assign outputs[3169] = ~(layer0_outputs[2688]);
    assign outputs[3170] = ~(layer0_outputs[4905]);
    assign outputs[3171] = layer0_outputs[236];
    assign outputs[3172] = ~(layer0_outputs[4204]) | (layer0_outputs[3712]);
    assign outputs[3173] = (layer0_outputs[3388]) & (layer0_outputs[4237]);
    assign outputs[3174] = ~(layer0_outputs[4605]);
    assign outputs[3175] = layer0_outputs[46];
    assign outputs[3176] = layer0_outputs[3459];
    assign outputs[3177] = ~(layer0_outputs[4742]);
    assign outputs[3178] = ~(layer0_outputs[3847]);
    assign outputs[3179] = (layer0_outputs[1180]) ^ (layer0_outputs[3349]);
    assign outputs[3180] = ~((layer0_outputs[1075]) ^ (layer0_outputs[209]));
    assign outputs[3181] = ~((layer0_outputs[4587]) ^ (layer0_outputs[421]));
    assign outputs[3182] = layer0_outputs[782];
    assign outputs[3183] = ~(layer0_outputs[983]);
    assign outputs[3184] = ~(layer0_outputs[492]);
    assign outputs[3185] = ~(layer0_outputs[1203]);
    assign outputs[3186] = (layer0_outputs[317]) & (layer0_outputs[4290]);
    assign outputs[3187] = ~(layer0_outputs[616]);
    assign outputs[3188] = layer0_outputs[2816];
    assign outputs[3189] = ~((layer0_outputs[4785]) & (layer0_outputs[298]));
    assign outputs[3190] = (layer0_outputs[4089]) & ~(layer0_outputs[1670]);
    assign outputs[3191] = (layer0_outputs[350]) ^ (layer0_outputs[4650]);
    assign outputs[3192] = ~((layer0_outputs[3896]) ^ (layer0_outputs[4459]));
    assign outputs[3193] = (layer0_outputs[4218]) & ~(layer0_outputs[271]);
    assign outputs[3194] = ~(layer0_outputs[3088]) | (layer0_outputs[337]);
    assign outputs[3195] = (layer0_outputs[542]) ^ (layer0_outputs[4512]);
    assign outputs[3196] = ~((layer0_outputs[4602]) ^ (layer0_outputs[2717]));
    assign outputs[3197] = (layer0_outputs[3382]) & (layer0_outputs[3805]);
    assign outputs[3198] = ~(layer0_outputs[2145]) | (layer0_outputs[3027]);
    assign outputs[3199] = (layer0_outputs[3138]) ^ (layer0_outputs[368]);
    assign outputs[3200] = ~(layer0_outputs[1451]);
    assign outputs[3201] = ~(layer0_outputs[4513]);
    assign outputs[3202] = (layer0_outputs[4927]) & ~(layer0_outputs[700]);
    assign outputs[3203] = layer0_outputs[1026];
    assign outputs[3204] = (layer0_outputs[1012]) & ~(layer0_outputs[100]);
    assign outputs[3205] = (layer0_outputs[224]) & ~(layer0_outputs[3146]);
    assign outputs[3206] = ~(layer0_outputs[1214]);
    assign outputs[3207] = layer0_outputs[4640];
    assign outputs[3208] = layer0_outputs[1981];
    assign outputs[3209] = layer0_outputs[741];
    assign outputs[3210] = ~((layer0_outputs[3607]) | (layer0_outputs[4952]));
    assign outputs[3211] = (layer0_outputs[3703]) | (layer0_outputs[4224]);
    assign outputs[3212] = (layer0_outputs[3407]) ^ (layer0_outputs[424]);
    assign outputs[3213] = ~(layer0_outputs[773]) | (layer0_outputs[756]);
    assign outputs[3214] = ~((layer0_outputs[2308]) | (layer0_outputs[2791]));
    assign outputs[3215] = layer0_outputs[1049];
    assign outputs[3216] = (layer0_outputs[1464]) & ~(layer0_outputs[83]);
    assign outputs[3217] = ~(layer0_outputs[3936]) | (layer0_outputs[4108]);
    assign outputs[3218] = ~((layer0_outputs[4391]) | (layer0_outputs[2513]));
    assign outputs[3219] = (layer0_outputs[582]) & ~(layer0_outputs[2753]);
    assign outputs[3220] = layer0_outputs[1770];
    assign outputs[3221] = layer0_outputs[3592];
    assign outputs[3222] = layer0_outputs[2084];
    assign outputs[3223] = layer0_outputs[818];
    assign outputs[3224] = (layer0_outputs[3747]) & ~(layer0_outputs[2843]);
    assign outputs[3225] = layer0_outputs[622];
    assign outputs[3226] = ~(layer0_outputs[3225]);
    assign outputs[3227] = ~((layer0_outputs[2711]) | (layer0_outputs[4600]));
    assign outputs[3228] = ~((layer0_outputs[3517]) ^ (layer0_outputs[2677]));
    assign outputs[3229] = ~(layer0_outputs[4580]) | (layer0_outputs[837]);
    assign outputs[3230] = (layer0_outputs[4082]) & (layer0_outputs[1767]);
    assign outputs[3231] = ~(layer0_outputs[4381]);
    assign outputs[3232] = (layer0_outputs[2175]) & ~(layer0_outputs[4233]);
    assign outputs[3233] = (layer0_outputs[1961]) | (layer0_outputs[895]);
    assign outputs[3234] = layer0_outputs[2652];
    assign outputs[3235] = layer0_outputs[3250];
    assign outputs[3236] = ~((layer0_outputs[790]) & (layer0_outputs[3940]));
    assign outputs[3237] = ~((layer0_outputs[2391]) | (layer0_outputs[523]));
    assign outputs[3238] = ~(layer0_outputs[2477]) | (layer0_outputs[4293]);
    assign outputs[3239] = (layer0_outputs[3857]) ^ (layer0_outputs[5073]);
    assign outputs[3240] = (layer0_outputs[2182]) & ~(layer0_outputs[2594]);
    assign outputs[3241] = ~(layer0_outputs[173]);
    assign outputs[3242] = layer0_outputs[3388];
    assign outputs[3243] = (layer0_outputs[3808]) & (layer0_outputs[5039]);
    assign outputs[3244] = ~(layer0_outputs[3946]) | (layer0_outputs[72]);
    assign outputs[3245] = ~(layer0_outputs[1500]);
    assign outputs[3246] = ~(layer0_outputs[2468]);
    assign outputs[3247] = layer0_outputs[174];
    assign outputs[3248] = ~((layer0_outputs[1337]) | (layer0_outputs[679]));
    assign outputs[3249] = ~((layer0_outputs[628]) ^ (layer0_outputs[4887]));
    assign outputs[3250] = (layer0_outputs[167]) & (layer0_outputs[2793]);
    assign outputs[3251] = (layer0_outputs[5095]) ^ (layer0_outputs[5105]);
    assign outputs[3252] = ~(layer0_outputs[3541]);
    assign outputs[3253] = ~(layer0_outputs[446]);
    assign outputs[3254] = ~((layer0_outputs[4375]) ^ (layer0_outputs[3794]));
    assign outputs[3255] = (layer0_outputs[3961]) ^ (layer0_outputs[1118]);
    assign outputs[3256] = (layer0_outputs[4347]) ^ (layer0_outputs[1438]);
    assign outputs[3257] = ~(layer0_outputs[2983]);
    assign outputs[3258] = ~(layer0_outputs[1595]);
    assign outputs[3259] = ~(layer0_outputs[5027]);
    assign outputs[3260] = ~((layer0_outputs[380]) | (layer0_outputs[3198]));
    assign outputs[3261] = ~(layer0_outputs[1575]) | (layer0_outputs[4173]);
    assign outputs[3262] = ~(layer0_outputs[1785]);
    assign outputs[3263] = layer0_outputs[2014];
    assign outputs[3264] = (layer0_outputs[4370]) & ~(layer0_outputs[1455]);
    assign outputs[3265] = ~((layer0_outputs[3523]) & (layer0_outputs[1533]));
    assign outputs[3266] = (layer0_outputs[478]) ^ (layer0_outputs[2613]);
    assign outputs[3267] = layer0_outputs[509];
    assign outputs[3268] = layer0_outputs[709];
    assign outputs[3269] = (layer0_outputs[56]) & ~(layer0_outputs[2532]);
    assign outputs[3270] = ~(layer0_outputs[2277]) | (layer0_outputs[26]);
    assign outputs[3271] = (layer0_outputs[2546]) ^ (layer0_outputs[158]);
    assign outputs[3272] = layer0_outputs[4254];
    assign outputs[3273] = layer0_outputs[2330];
    assign outputs[3274] = (layer0_outputs[2942]) & ~(layer0_outputs[907]);
    assign outputs[3275] = ~((layer0_outputs[418]) | (layer0_outputs[2691]));
    assign outputs[3276] = layer0_outputs[1732];
    assign outputs[3277] = ~((layer0_outputs[4152]) | (layer0_outputs[4895]));
    assign outputs[3278] = ~((layer0_outputs[2876]) | (layer0_outputs[1160]));
    assign outputs[3279] = ~((layer0_outputs[2249]) ^ (layer0_outputs[3058]));
    assign outputs[3280] = (layer0_outputs[2945]) | (layer0_outputs[3493]);
    assign outputs[3281] = (layer0_outputs[2725]) ^ (layer0_outputs[1742]);
    assign outputs[3282] = (layer0_outputs[2515]) & (layer0_outputs[4983]);
    assign outputs[3283] = ~((layer0_outputs[1947]) | (layer0_outputs[800]));
    assign outputs[3284] = (layer0_outputs[2237]) & ~(layer0_outputs[1461]);
    assign outputs[3285] = layer0_outputs[4965];
    assign outputs[3286] = ~((layer0_outputs[1982]) ^ (layer0_outputs[3573]));
    assign outputs[3287] = ~((layer0_outputs[4791]) ^ (layer0_outputs[2318]));
    assign outputs[3288] = ~((layer0_outputs[2398]) & (layer0_outputs[2720]));
    assign outputs[3289] = ~((layer0_outputs[2537]) ^ (layer0_outputs[88]));
    assign outputs[3290] = ~((layer0_outputs[4207]) & (layer0_outputs[3553]));
    assign outputs[3291] = ~(layer0_outputs[2870]);
    assign outputs[3292] = ~((layer0_outputs[5030]) ^ (layer0_outputs[236]));
    assign outputs[3293] = (layer0_outputs[2522]) & ~(layer0_outputs[4464]);
    assign outputs[3294] = ~(layer0_outputs[1172]);
    assign outputs[3295] = ~((layer0_outputs[1591]) & (layer0_outputs[3083]));
    assign outputs[3296] = (layer0_outputs[488]) & (layer0_outputs[3562]);
    assign outputs[3297] = ~((layer0_outputs[3181]) & (layer0_outputs[435]));
    assign outputs[3298] = (layer0_outputs[60]) ^ (layer0_outputs[3412]);
    assign outputs[3299] = (layer0_outputs[3368]) ^ (layer0_outputs[2033]);
    assign outputs[3300] = (layer0_outputs[3342]) ^ (layer0_outputs[626]);
    assign outputs[3301] = (layer0_outputs[3199]) ^ (layer0_outputs[3299]);
    assign outputs[3302] = ~(layer0_outputs[4533]);
    assign outputs[3303] = ~((layer0_outputs[3490]) & (layer0_outputs[3404]));
    assign outputs[3304] = ~(layer0_outputs[1999]);
    assign outputs[3305] = layer0_outputs[1369];
    assign outputs[3306] = layer0_outputs[1333];
    assign outputs[3307] = ~((layer0_outputs[715]) & (layer0_outputs[3767]));
    assign outputs[3308] = layer0_outputs[3594];
    assign outputs[3309] = (layer0_outputs[3667]) | (layer0_outputs[3757]);
    assign outputs[3310] = ~((layer0_outputs[162]) & (layer0_outputs[3161]));
    assign outputs[3311] = (layer0_outputs[4555]) & ~(layer0_outputs[263]);
    assign outputs[3312] = (layer0_outputs[3913]) ^ (layer0_outputs[3339]);
    assign outputs[3313] = (layer0_outputs[786]) & ~(layer0_outputs[4771]);
    assign outputs[3314] = (layer0_outputs[1069]) & ~(layer0_outputs[1092]);
    assign outputs[3315] = (layer0_outputs[2072]) ^ (layer0_outputs[511]);
    assign outputs[3316] = (layer0_outputs[4642]) & (layer0_outputs[2003]);
    assign outputs[3317] = layer0_outputs[879];
    assign outputs[3318] = ~((layer0_outputs[4015]) | (layer0_outputs[452]));
    assign outputs[3319] = ~((layer0_outputs[554]) ^ (layer0_outputs[3205]));
    assign outputs[3320] = ~(layer0_outputs[2176]);
    assign outputs[3321] = layer0_outputs[1096];
    assign outputs[3322] = ~((layer0_outputs[457]) ^ (layer0_outputs[462]));
    assign outputs[3323] = ~((layer0_outputs[1011]) | (layer0_outputs[2678]));
    assign outputs[3324] = layer0_outputs[669];
    assign outputs[3325] = ~(layer0_outputs[3540]) | (layer0_outputs[3711]);
    assign outputs[3326] = ~((layer0_outputs[3741]) ^ (layer0_outputs[602]));
    assign outputs[3327] = layer0_outputs[3180];
    assign outputs[3328] = (layer0_outputs[810]) & ~(layer0_outputs[2972]);
    assign outputs[3329] = ~((layer0_outputs[106]) ^ (layer0_outputs[1744]));
    assign outputs[3330] = ~(layer0_outputs[2929]);
    assign outputs[3331] = ~((layer0_outputs[852]) | (layer0_outputs[3104]));
    assign outputs[3332] = (layer0_outputs[3874]) & (layer0_outputs[1018]);
    assign outputs[3333] = ~(layer0_outputs[1797]) | (layer0_outputs[1864]);
    assign outputs[3334] = ~((layer0_outputs[2964]) ^ (layer0_outputs[1059]));
    assign outputs[3335] = ~(layer0_outputs[1576]);
    assign outputs[3336] = layer0_outputs[2473];
    assign outputs[3337] = ~(layer0_outputs[5104]);
    assign outputs[3338] = layer0_outputs[3534];
    assign outputs[3339] = (layer0_outputs[4990]) ^ (layer0_outputs[3951]);
    assign outputs[3340] = layer0_outputs[5014];
    assign outputs[3341] = (layer0_outputs[4577]) ^ (layer0_outputs[4483]);
    assign outputs[3342] = ~(layer0_outputs[3295]) | (layer0_outputs[2950]);
    assign outputs[3343] = ~((layer0_outputs[4962]) ^ (layer0_outputs[4466]));
    assign outputs[3344] = layer0_outputs[2922];
    assign outputs[3345] = (layer0_outputs[4941]) & (layer0_outputs[1151]);
    assign outputs[3346] = ~(layer0_outputs[4750]);
    assign outputs[3347] = layer0_outputs[5100];
    assign outputs[3348] = ~(layer0_outputs[917]) | (layer0_outputs[2542]);
    assign outputs[3349] = ~((layer0_outputs[4424]) ^ (layer0_outputs[2184]));
    assign outputs[3350] = layer0_outputs[4210];
    assign outputs[3351] = ~(layer0_outputs[2067]) | (layer0_outputs[4657]);
    assign outputs[3352] = (layer0_outputs[909]) & ~(layer0_outputs[2554]);
    assign outputs[3353] = ~((layer0_outputs[2676]) ^ (layer0_outputs[1201]));
    assign outputs[3354] = layer0_outputs[4729];
    assign outputs[3355] = ~((layer0_outputs[3861]) | (layer0_outputs[4064]));
    assign outputs[3356] = layer0_outputs[618];
    assign outputs[3357] = layer0_outputs[2354];
    assign outputs[3358] = ~(layer0_outputs[159]) | (layer0_outputs[177]);
    assign outputs[3359] = layer0_outputs[3668];
    assign outputs[3360] = (layer0_outputs[5106]) ^ (layer0_outputs[2106]);
    assign outputs[3361] = ~(layer0_outputs[467]) | (layer0_outputs[1330]);
    assign outputs[3362] = layer0_outputs[3376];
    assign outputs[3363] = (layer0_outputs[1499]) ^ (layer0_outputs[3362]);
    assign outputs[3364] = ~(layer0_outputs[340]);
    assign outputs[3365] = layer0_outputs[4879];
    assign outputs[3366] = layer0_outputs[2963];
    assign outputs[3367] = (layer0_outputs[1324]) ^ (layer0_outputs[4413]);
    assign outputs[3368] = ~(layer0_outputs[1871]);
    assign outputs[3369] = layer0_outputs[3201];
    assign outputs[3370] = (layer0_outputs[801]) & ~(layer0_outputs[296]);
    assign outputs[3371] = ~((layer0_outputs[92]) ^ (layer0_outputs[348]));
    assign outputs[3372] = (layer0_outputs[2830]) & (layer0_outputs[4590]);
    assign outputs[3373] = ~((layer0_outputs[520]) | (layer0_outputs[4779]));
    assign outputs[3374] = layer0_outputs[91];
    assign outputs[3375] = layer0_outputs[1073];
    assign outputs[3376] = ~(layer0_outputs[4874]) | (layer0_outputs[2265]);
    assign outputs[3377] = layer0_outputs[2205];
    assign outputs[3378] = ~(layer0_outputs[25]) | (layer0_outputs[3169]);
    assign outputs[3379] = layer0_outputs[3283];
    assign outputs[3380] = layer0_outputs[2610];
    assign outputs[3381] = ~((layer0_outputs[151]) | (layer0_outputs[865]));
    assign outputs[3382] = ~(layer0_outputs[2209]);
    assign outputs[3383] = ~(layer0_outputs[1561]);
    assign outputs[3384] = layer0_outputs[3437];
    assign outputs[3385] = layer0_outputs[1633];
    assign outputs[3386] = (layer0_outputs[4145]) ^ (layer0_outputs[4024]);
    assign outputs[3387] = layer0_outputs[5004];
    assign outputs[3388] = ~(layer0_outputs[3233]);
    assign outputs[3389] = ~(layer0_outputs[2657]);
    assign outputs[3390] = layer0_outputs[3826];
    assign outputs[3391] = (layer0_outputs[3883]) & ~(layer0_outputs[1659]);
    assign outputs[3392] = (layer0_outputs[3980]) ^ (layer0_outputs[1485]);
    assign outputs[3393] = layer0_outputs[1508];
    assign outputs[3394] = ~((layer0_outputs[3468]) ^ (layer0_outputs[4148]));
    assign outputs[3395] = ~((layer0_outputs[3298]) & (layer0_outputs[1246]));
    assign outputs[3396] = ~(layer0_outputs[4250]);
    assign outputs[3397] = (layer0_outputs[2415]) & ~(layer0_outputs[3929]);
    assign outputs[3398] = layer0_outputs[3866];
    assign outputs[3399] = ~(layer0_outputs[5041]);
    assign outputs[3400] = ~((layer0_outputs[4153]) ^ (layer0_outputs[205]));
    assign outputs[3401] = layer0_outputs[3194];
    assign outputs[3402] = ~((layer0_outputs[4003]) ^ (layer0_outputs[3943]));
    assign outputs[3403] = ~(layer0_outputs[1716]) | (layer0_outputs[1647]);
    assign outputs[3404] = ~(layer0_outputs[1229]);
    assign outputs[3405] = ~((layer0_outputs[2194]) ^ (layer0_outputs[3043]));
    assign outputs[3406] = layer0_outputs[4267];
    assign outputs[3407] = (layer0_outputs[3317]) ^ (layer0_outputs[3889]);
    assign outputs[3408] = layer0_outputs[723];
    assign outputs[3409] = layer0_outputs[1760];
    assign outputs[3410] = ~((layer0_outputs[2166]) ^ (layer0_outputs[2015]));
    assign outputs[3411] = layer0_outputs[3949];
    assign outputs[3412] = layer0_outputs[4404];
    assign outputs[3413] = ~(layer0_outputs[31]);
    assign outputs[3414] = ~(layer0_outputs[2726]);
    assign outputs[3415] = (layer0_outputs[934]) & ~(layer0_outputs[1302]);
    assign outputs[3416] = (layer0_outputs[2539]) ^ (layer0_outputs[2472]);
    assign outputs[3417] = layer0_outputs[3836];
    assign outputs[3418] = ~(layer0_outputs[4666]);
    assign outputs[3419] = ~((layer0_outputs[4197]) ^ (layer0_outputs[4221]));
    assign outputs[3420] = layer0_outputs[868];
    assign outputs[3421] = ~(layer0_outputs[2361]);
    assign outputs[3422] = ~(layer0_outputs[427]);
    assign outputs[3423] = (layer0_outputs[1315]) | (layer0_outputs[4525]);
    assign outputs[3424] = ~((layer0_outputs[2170]) ^ (layer0_outputs[3956]));
    assign outputs[3425] = ~(layer0_outputs[4917]);
    assign outputs[3426] = ~((layer0_outputs[2513]) ^ (layer0_outputs[2955]));
    assign outputs[3427] = (layer0_outputs[5003]) & ~(layer0_outputs[4102]);
    assign outputs[3428] = (layer0_outputs[1727]) ^ (layer0_outputs[1930]);
    assign outputs[3429] = (layer0_outputs[1426]) ^ (layer0_outputs[2745]);
    assign outputs[3430] = ~(layer0_outputs[4516]) | (layer0_outputs[2198]);
    assign outputs[3431] = ~((layer0_outputs[3245]) ^ (layer0_outputs[4826]));
    assign outputs[3432] = layer0_outputs[3029];
    assign outputs[3433] = layer0_outputs[2258];
    assign outputs[3434] = ~((layer0_outputs[883]) ^ (layer0_outputs[5053]));
    assign outputs[3435] = layer0_outputs[1115];
    assign outputs[3436] = ~((layer0_outputs[3262]) | (layer0_outputs[1602]));
    assign outputs[3437] = ~((layer0_outputs[3089]) ^ (layer0_outputs[3352]));
    assign outputs[3438] = ~(layer0_outputs[4409]) | (layer0_outputs[4749]);
    assign outputs[3439] = (layer0_outputs[2052]) & ~(layer0_outputs[2121]);
    assign outputs[3440] = ~(layer0_outputs[2622]);
    assign outputs[3441] = layer0_outputs[2639];
    assign outputs[3442] = layer0_outputs[2435];
    assign outputs[3443] = (layer0_outputs[948]) & ~(layer0_outputs[3448]);
    assign outputs[3444] = ~(layer0_outputs[4926]);
    assign outputs[3445] = layer0_outputs[2673];
    assign outputs[3446] = ~((layer0_outputs[4660]) ^ (layer0_outputs[3319]));
    assign outputs[3447] = ~(layer0_outputs[3536]) | (layer0_outputs[961]);
    assign outputs[3448] = ~(layer0_outputs[2909]);
    assign outputs[3449] = ~(layer0_outputs[2983]);
    assign outputs[3450] = layer0_outputs[4007];
    assign outputs[3451] = ~((layer0_outputs[351]) | (layer0_outputs[4938]));
    assign outputs[3452] = ~((layer0_outputs[2592]) | (layer0_outputs[566]));
    assign outputs[3453] = (layer0_outputs[2560]) & ~(layer0_outputs[4297]);
    assign outputs[3454] = ~(layer0_outputs[2209]);
    assign outputs[3455] = (layer0_outputs[4495]) ^ (layer0_outputs[2820]);
    assign outputs[3456] = ~((layer0_outputs[4406]) ^ (layer0_outputs[182]));
    assign outputs[3457] = (layer0_outputs[4543]) & ~(layer0_outputs[4954]);
    assign outputs[3458] = (layer0_outputs[3427]) & ~(layer0_outputs[1869]);
    assign outputs[3459] = ~(layer0_outputs[2067]);
    assign outputs[3460] = ~(layer0_outputs[487]);
    assign outputs[3461] = layer0_outputs[3398];
    assign outputs[3462] = (layer0_outputs[4101]) ^ (layer0_outputs[895]);
    assign outputs[3463] = (layer0_outputs[4918]) ^ (layer0_outputs[1453]);
    assign outputs[3464] = layer0_outputs[795];
    assign outputs[3465] = layer0_outputs[1285];
    assign outputs[3466] = ~((layer0_outputs[2917]) | (layer0_outputs[3982]));
    assign outputs[3467] = ~((layer0_outputs[2391]) | (layer0_outputs[1477]));
    assign outputs[3468] = ~((layer0_outputs[478]) ^ (layer0_outputs[1659]));
    assign outputs[3469] = ~((layer0_outputs[4776]) & (layer0_outputs[2285]));
    assign outputs[3470] = layer0_outputs[3965];
    assign outputs[3471] = (layer0_outputs[5023]) ^ (layer0_outputs[133]);
    assign outputs[3472] = (layer0_outputs[4471]) & ~(layer0_outputs[4182]);
    assign outputs[3473] = ~((layer0_outputs[4690]) | (layer0_outputs[4606]));
    assign outputs[3474] = ~((layer0_outputs[1097]) ^ (layer0_outputs[4832]));
    assign outputs[3475] = (layer0_outputs[617]) & ~(layer0_outputs[2443]);
    assign outputs[3476] = (layer0_outputs[1658]) & (layer0_outputs[2581]);
    assign outputs[3477] = ~(layer0_outputs[1901]);
    assign outputs[3478] = (layer0_outputs[1194]) & ~(layer0_outputs[4472]);
    assign outputs[3479] = ~(layer0_outputs[3982]);
    assign outputs[3480] = ~((layer0_outputs[1196]) ^ (layer0_outputs[1799]));
    assign outputs[3481] = ~((layer0_outputs[4020]) ^ (layer0_outputs[2715]));
    assign outputs[3482] = layer0_outputs[657];
    assign outputs[3483] = ~(layer0_outputs[3251]);
    assign outputs[3484] = ~(layer0_outputs[3392]);
    assign outputs[3485] = layer0_outputs[1846];
    assign outputs[3486] = ~((layer0_outputs[672]) & (layer0_outputs[1782]));
    assign outputs[3487] = ~(layer0_outputs[2653]);
    assign outputs[3488] = (layer0_outputs[1894]) & (layer0_outputs[1958]);
    assign outputs[3489] = ~(layer0_outputs[3823]);
    assign outputs[3490] = ~((layer0_outputs[3206]) | (layer0_outputs[3181]));
    assign outputs[3491] = (layer0_outputs[357]) ^ (layer0_outputs[4097]);
    assign outputs[3492] = ~((layer0_outputs[2590]) | (layer0_outputs[1691]));
    assign outputs[3493] = layer0_outputs[5081];
    assign outputs[3494] = layer0_outputs[4065];
    assign outputs[3495] = layer0_outputs[3978];
    assign outputs[3496] = ~(layer0_outputs[4313]);
    assign outputs[3497] = layer0_outputs[1295];
    assign outputs[3498] = ~(layer0_outputs[1234]);
    assign outputs[3499] = ~(layer0_outputs[2305]);
    assign outputs[3500] = layer0_outputs[1514];
    assign outputs[3501] = ~(layer0_outputs[318]);
    assign outputs[3502] = layer0_outputs[900];
    assign outputs[3503] = layer0_outputs[1751];
    assign outputs[3504] = ~(layer0_outputs[4076]);
    assign outputs[3505] = ~(layer0_outputs[1266]);
    assign outputs[3506] = (layer0_outputs[1728]) ^ (layer0_outputs[4253]);
    assign outputs[3507] = layer0_outputs[948];
    assign outputs[3508] = layer0_outputs[211];
    assign outputs[3509] = ~(layer0_outputs[2584]);
    assign outputs[3510] = (layer0_outputs[461]) & ~(layer0_outputs[1409]);
    assign outputs[3511] = layer0_outputs[1262];
    assign outputs[3512] = (layer0_outputs[1874]) & ~(layer0_outputs[3550]);
    assign outputs[3513] = (layer0_outputs[4283]) & ~(layer0_outputs[2973]);
    assign outputs[3514] = (layer0_outputs[2104]) & ~(layer0_outputs[3657]);
    assign outputs[3515] = (layer0_outputs[1681]) & ~(layer0_outputs[2647]);
    assign outputs[3516] = (layer0_outputs[2222]) | (layer0_outputs[4263]);
    assign outputs[3517] = (layer0_outputs[915]) | (layer0_outputs[1057]);
    assign outputs[3518] = layer0_outputs[3622];
    assign outputs[3519] = layer0_outputs[3545];
    assign outputs[3520] = (layer0_outputs[2456]) & ~(layer0_outputs[4664]);
    assign outputs[3521] = layer0_outputs[3279];
    assign outputs[3522] = layer0_outputs[1861];
    assign outputs[3523] = layer0_outputs[3123];
    assign outputs[3524] = (layer0_outputs[4397]) ^ (layer0_outputs[3891]);
    assign outputs[3525] = layer0_outputs[3040];
    assign outputs[3526] = (layer0_outputs[2336]) | (layer0_outputs[3711]);
    assign outputs[3527] = layer0_outputs[4094];
    assign outputs[3528] = layer0_outputs[3236];
    assign outputs[3529] = ~(layer0_outputs[4103]) | (layer0_outputs[3789]);
    assign outputs[3530] = layer0_outputs[2859];
    assign outputs[3531] = (layer0_outputs[195]) ^ (layer0_outputs[1990]);
    assign outputs[3532] = ~((layer0_outputs[4867]) | (layer0_outputs[4464]));
    assign outputs[3533] = layer0_outputs[3763];
    assign outputs[3534] = (layer0_outputs[4850]) ^ (layer0_outputs[1153]);
    assign outputs[3535] = (layer0_outputs[4282]) & (layer0_outputs[45]);
    assign outputs[3536] = layer0_outputs[4840];
    assign outputs[3537] = ~((layer0_outputs[4403]) ^ (layer0_outputs[4829]));
    assign outputs[3538] = (layer0_outputs[3074]) & (layer0_outputs[2110]);
    assign outputs[3539] = ~(layer0_outputs[3113]);
    assign outputs[3540] = ~(layer0_outputs[4097]);
    assign outputs[3541] = ~(layer0_outputs[4260]);
    assign outputs[3542] = (layer0_outputs[111]) ^ (layer0_outputs[2013]);
    assign outputs[3543] = ~((layer0_outputs[947]) ^ (layer0_outputs[2719]));
    assign outputs[3544] = (layer0_outputs[1666]) | (layer0_outputs[3279]);
    assign outputs[3545] = ~((layer0_outputs[3001]) & (layer0_outputs[4265]));
    assign outputs[3546] = ~(layer0_outputs[1913]);
    assign outputs[3547] = layer0_outputs[4830];
    assign outputs[3548] = ~(layer0_outputs[519]);
    assign outputs[3549] = ~(layer0_outputs[894]);
    assign outputs[3550] = layer0_outputs[3267];
    assign outputs[3551] = ~(layer0_outputs[1128]);
    assign outputs[3552] = ~((layer0_outputs[1988]) ^ (layer0_outputs[1391]));
    assign outputs[3553] = ~(layer0_outputs[1440]);
    assign outputs[3554] = layer0_outputs[1806];
    assign outputs[3555] = ~(layer0_outputs[4963]) | (layer0_outputs[1227]);
    assign outputs[3556] = layer0_outputs[2924];
    assign outputs[3557] = (layer0_outputs[4687]) & ~(layer0_outputs[1998]);
    assign outputs[3558] = (layer0_outputs[4386]) ^ (layer0_outputs[1043]);
    assign outputs[3559] = ~((layer0_outputs[2656]) | (layer0_outputs[4014]));
    assign outputs[3560] = ~((layer0_outputs[2172]) ^ (layer0_outputs[3444]));
    assign outputs[3561] = layer0_outputs[428];
    assign outputs[3562] = ~(layer0_outputs[3523]) | (layer0_outputs[3849]);
    assign outputs[3563] = ~(layer0_outputs[4546]);
    assign outputs[3564] = ~(layer0_outputs[3]);
    assign outputs[3565] = (layer0_outputs[4309]) & (layer0_outputs[1974]);
    assign outputs[3566] = ~(layer0_outputs[1037]);
    assign outputs[3567] = (layer0_outputs[4018]) & ~(layer0_outputs[2776]);
    assign outputs[3568] = (layer0_outputs[1209]) & (layer0_outputs[2402]);
    assign outputs[3569] = (layer0_outputs[3461]) & ~(layer0_outputs[2933]);
    assign outputs[3570] = ~(layer0_outputs[3208]);
    assign outputs[3571] = ~(layer0_outputs[2221]);
    assign outputs[3572] = ~(layer0_outputs[3602]);
    assign outputs[3573] = ~(layer0_outputs[2486]) | (layer0_outputs[3831]);
    assign outputs[3574] = ~(layer0_outputs[480]) | (layer0_outputs[1450]);
    assign outputs[3575] = 1'b0;
    assign outputs[3576] = (layer0_outputs[4708]) ^ (layer0_outputs[3693]);
    assign outputs[3577] = ~(layer0_outputs[30]);
    assign outputs[3578] = ~((layer0_outputs[4617]) ^ (layer0_outputs[4]));
    assign outputs[3579] = (layer0_outputs[2230]) | (layer0_outputs[1779]);
    assign outputs[3580] = layer0_outputs[273];
    assign outputs[3581] = ~(layer0_outputs[2554]);
    assign outputs[3582] = ~((layer0_outputs[1189]) | (layer0_outputs[4028]));
    assign outputs[3583] = ~((layer0_outputs[217]) ^ (layer0_outputs[1852]));
    assign outputs[3584] = (layer0_outputs[1407]) | (layer0_outputs[3953]);
    assign outputs[3585] = ~((layer0_outputs[4361]) & (layer0_outputs[4402]));
    assign outputs[3586] = ~(layer0_outputs[3534]);
    assign outputs[3587] = ~(layer0_outputs[3506]) | (layer0_outputs[4799]);
    assign outputs[3588] = ~((layer0_outputs[3782]) ^ (layer0_outputs[4384]));
    assign outputs[3589] = (layer0_outputs[512]) & ~(layer0_outputs[1115]);
    assign outputs[3590] = ~(layer0_outputs[2822]) | (layer0_outputs[2897]);
    assign outputs[3591] = ~(layer0_outputs[4644]);
    assign outputs[3592] = ~(layer0_outputs[2128]);
    assign outputs[3593] = ~((layer0_outputs[4644]) | (layer0_outputs[915]));
    assign outputs[3594] = ~(layer0_outputs[4739]);
    assign outputs[3595] = ~((layer0_outputs[4436]) ^ (layer0_outputs[4160]));
    assign outputs[3596] = ~((layer0_outputs[762]) ^ (layer0_outputs[4063]));
    assign outputs[3597] = (layer0_outputs[4074]) & ~(layer0_outputs[1831]);
    assign outputs[3598] = ~((layer0_outputs[4841]) ^ (layer0_outputs[1993]));
    assign outputs[3599] = ~((layer0_outputs[2978]) ^ (layer0_outputs[2269]));
    assign outputs[3600] = layer0_outputs[2673];
    assign outputs[3601] = ~((layer0_outputs[4493]) | (layer0_outputs[494]));
    assign outputs[3602] = layer0_outputs[3868];
    assign outputs[3603] = layer0_outputs[3133];
    assign outputs[3604] = ~(layer0_outputs[1044]);
    assign outputs[3605] = (layer0_outputs[1250]) ^ (layer0_outputs[861]);
    assign outputs[3606] = ~((layer0_outputs[4029]) & (layer0_outputs[4265]));
    assign outputs[3607] = ~((layer0_outputs[200]) ^ (layer0_outputs[2605]));
    assign outputs[3608] = (layer0_outputs[2058]) & ~(layer0_outputs[1544]);
    assign outputs[3609] = (layer0_outputs[3762]) ^ (layer0_outputs[4867]);
    assign outputs[3610] = (layer0_outputs[1178]) & ~(layer0_outputs[2538]);
    assign outputs[3611] = (layer0_outputs[4802]) & ~(layer0_outputs[1415]);
    assign outputs[3612] = layer0_outputs[1662];
    assign outputs[3613] = (layer0_outputs[3612]) & ~(layer0_outputs[3578]);
    assign outputs[3614] = ~(layer0_outputs[1709]);
    assign outputs[3615] = layer0_outputs[905];
    assign outputs[3616] = ~(layer0_outputs[2608]);
    assign outputs[3617] = ~(layer0_outputs[1349]);
    assign outputs[3618] = (layer0_outputs[361]) ^ (layer0_outputs[2018]);
    assign outputs[3619] = ~((layer0_outputs[1876]) ^ (layer0_outputs[1388]));
    assign outputs[3620] = (layer0_outputs[2133]) & ~(layer0_outputs[3547]);
    assign outputs[3621] = (layer0_outputs[58]) ^ (layer0_outputs[4463]);
    assign outputs[3622] = (layer0_outputs[85]) & (layer0_outputs[3723]);
    assign outputs[3623] = (layer0_outputs[4260]) & ~(layer0_outputs[2071]);
    assign outputs[3624] = ~(layer0_outputs[2380]) | (layer0_outputs[3465]);
    assign outputs[3625] = layer0_outputs[4490];
    assign outputs[3626] = (layer0_outputs[1279]) & ~(layer0_outputs[699]);
    assign outputs[3627] = layer0_outputs[993];
    assign outputs[3628] = (layer0_outputs[3686]) & ~(layer0_outputs[4021]);
    assign outputs[3629] = layer0_outputs[4379];
    assign outputs[3630] = ~(layer0_outputs[2431]) | (layer0_outputs[3058]);
    assign outputs[3631] = (layer0_outputs[3235]) & (layer0_outputs[4339]);
    assign outputs[3632] = (layer0_outputs[53]) & ~(layer0_outputs[3100]);
    assign outputs[3633] = (layer0_outputs[429]) & ~(layer0_outputs[912]);
    assign outputs[3634] = (layer0_outputs[4819]) ^ (layer0_outputs[2392]);
    assign outputs[3635] = layer0_outputs[987];
    assign outputs[3636] = ~((layer0_outputs[4310]) ^ (layer0_outputs[2502]));
    assign outputs[3637] = layer0_outputs[4345];
    assign outputs[3638] = (layer0_outputs[787]) & (layer0_outputs[5110]);
    assign outputs[3639] = layer0_outputs[3041];
    assign outputs[3640] = (layer0_outputs[486]) ^ (layer0_outputs[3356]);
    assign outputs[3641] = (layer0_outputs[4082]) & ~(layer0_outputs[2041]);
    assign outputs[3642] = (layer0_outputs[1792]) & (layer0_outputs[4842]);
    assign outputs[3643] = (layer0_outputs[2316]) ^ (layer0_outputs[45]);
    assign outputs[3644] = ~((layer0_outputs[2484]) ^ (layer0_outputs[3785]));
    assign outputs[3645] = layer0_outputs[1873];
    assign outputs[3646] = ~(layer0_outputs[3852]);
    assign outputs[3647] = (layer0_outputs[2779]) & (layer0_outputs[1101]);
    assign outputs[3648] = layer0_outputs[4327];
    assign outputs[3649] = (layer0_outputs[2365]) & ~(layer0_outputs[4267]);
    assign outputs[3650] = layer0_outputs[4700];
    assign outputs[3651] = layer0_outputs[4967];
    assign outputs[3652] = ~(layer0_outputs[2236]);
    assign outputs[3653] = layer0_outputs[2589];
    assign outputs[3654] = ~((layer0_outputs[3488]) | (layer0_outputs[4390]));
    assign outputs[3655] = layer0_outputs[3434];
    assign outputs[3656] = ~(layer0_outputs[4835]);
    assign outputs[3657] = ~((layer0_outputs[3022]) ^ (layer0_outputs[4985]));
    assign outputs[3658] = (layer0_outputs[3019]) & ~(layer0_outputs[248]);
    assign outputs[3659] = ~((layer0_outputs[5043]) ^ (layer0_outputs[134]));
    assign outputs[3660] = ~(layer0_outputs[1124]);
    assign outputs[3661] = ~(layer0_outputs[2687]);
    assign outputs[3662] = (layer0_outputs[3643]) & (layer0_outputs[4326]);
    assign outputs[3663] = ~(layer0_outputs[4364]);
    assign outputs[3664] = ~((layer0_outputs[664]) | (layer0_outputs[3409]));
    assign outputs[3665] = ~((layer0_outputs[1358]) | (layer0_outputs[4434]));
    assign outputs[3666] = ~(layer0_outputs[1483]);
    assign outputs[3667] = (layer0_outputs[863]) ^ (layer0_outputs[2311]);
    assign outputs[3668] = ~((layer0_outputs[1052]) & (layer0_outputs[2057]));
    assign outputs[3669] = layer0_outputs[2289];
    assign outputs[3670] = (layer0_outputs[4377]) & ~(layer0_outputs[398]);
    assign outputs[3671] = ~(layer0_outputs[1824]);
    assign outputs[3672] = ~(layer0_outputs[942]);
    assign outputs[3673] = ~(layer0_outputs[219]);
    assign outputs[3674] = (layer0_outputs[4025]) & ~(layer0_outputs[4898]);
    assign outputs[3675] = (layer0_outputs[1060]) & ~(layer0_outputs[717]);
    assign outputs[3676] = ~(layer0_outputs[2956]);
    assign outputs[3677] = (layer0_outputs[3634]) & ~(layer0_outputs[1929]);
    assign outputs[3678] = ~((layer0_outputs[2003]) ^ (layer0_outputs[1343]));
    assign outputs[3679] = (layer0_outputs[966]) & ~(layer0_outputs[4361]);
    assign outputs[3680] = (layer0_outputs[1935]) & ~(layer0_outputs[3009]);
    assign outputs[3681] = ~((layer0_outputs[1242]) ^ (layer0_outputs[954]));
    assign outputs[3682] = ~(layer0_outputs[331]);
    assign outputs[3683] = layer0_outputs[4570];
    assign outputs[3684] = ~(layer0_outputs[2000]);
    assign outputs[3685] = layer0_outputs[450];
    assign outputs[3686] = (layer0_outputs[2093]) & ~(layer0_outputs[2986]);
    assign outputs[3687] = ~((layer0_outputs[3063]) ^ (layer0_outputs[1599]));
    assign outputs[3688] = (layer0_outputs[1247]) ^ (layer0_outputs[2358]);
    assign outputs[3689] = (layer0_outputs[9]) ^ (layer0_outputs[1289]);
    assign outputs[3690] = ~((layer0_outputs[1981]) ^ (layer0_outputs[551]));
    assign outputs[3691] = (layer0_outputs[4559]) ^ (layer0_outputs[500]);
    assign outputs[3692] = (layer0_outputs[1627]) ^ (layer0_outputs[3240]);
    assign outputs[3693] = (layer0_outputs[614]) & (layer0_outputs[1344]);
    assign outputs[3694] = ~((layer0_outputs[3165]) | (layer0_outputs[3888]));
    assign outputs[3695] = layer0_outputs[2722];
    assign outputs[3696] = layer0_outputs[2246];
    assign outputs[3697] = ~(layer0_outputs[3471]);
    assign outputs[3698] = (layer0_outputs[2809]) & ~(layer0_outputs[2566]);
    assign outputs[3699] = layer0_outputs[1368];
    assign outputs[3700] = (layer0_outputs[3511]) & (layer0_outputs[90]);
    assign outputs[3701] = (layer0_outputs[2815]) & ~(layer0_outputs[1624]);
    assign outputs[3702] = layer0_outputs[2723];
    assign outputs[3703] = (layer0_outputs[4509]) & ~(layer0_outputs[126]);
    assign outputs[3704] = ~(layer0_outputs[98]);
    assign outputs[3705] = (layer0_outputs[3096]) & (layer0_outputs[656]);
    assign outputs[3706] = ~((layer0_outputs[3742]) | (layer0_outputs[1148]));
    assign outputs[3707] = ~((layer0_outputs[674]) ^ (layer0_outputs[4485]));
    assign outputs[3708] = (layer0_outputs[4896]) & ~(layer0_outputs[2354]);
    assign outputs[3709] = layer0_outputs[665];
    assign outputs[3710] = (layer0_outputs[4576]) & (layer0_outputs[270]);
    assign outputs[3711] = (layer0_outputs[4686]) | (layer0_outputs[3838]);
    assign outputs[3712] = layer0_outputs[1608];
    assign outputs[3713] = (layer0_outputs[4376]) & ~(layer0_outputs[2816]);
    assign outputs[3714] = 1'b0;
    assign outputs[3715] = layer0_outputs[3979];
    assign outputs[3716] = ~((layer0_outputs[2408]) | (layer0_outputs[5060]));
    assign outputs[3717] = (layer0_outputs[2387]) & ~(layer0_outputs[3323]);
    assign outputs[3718] = (layer0_outputs[3684]) & ~(layer0_outputs[4124]);
    assign outputs[3719] = layer0_outputs[2343];
    assign outputs[3720] = ~(layer0_outputs[4199]);
    assign outputs[3721] = ~(layer0_outputs[1433]);
    assign outputs[3722] = layer0_outputs[3857];
    assign outputs[3723] = ~(layer0_outputs[3044]);
    assign outputs[3724] = (layer0_outputs[3379]) & (layer0_outputs[294]);
    assign outputs[3725] = (layer0_outputs[1371]) & ~(layer0_outputs[1705]);
    assign outputs[3726] = ~(layer0_outputs[3397]) | (layer0_outputs[420]);
    assign outputs[3727] = layer0_outputs[2156];
    assign outputs[3728] = layer0_outputs[1006];
    assign outputs[3729] = ~(layer0_outputs[3557]);
    assign outputs[3730] = (layer0_outputs[884]) & ~(layer0_outputs[4633]);
    assign outputs[3731] = layer0_outputs[637];
    assign outputs[3732] = ~((layer0_outputs[4916]) | (layer0_outputs[1221]));
    assign outputs[3733] = ~(layer0_outputs[180]) | (layer0_outputs[58]);
    assign outputs[3734] = layer0_outputs[4621];
    assign outputs[3735] = ~(layer0_outputs[2295]);
    assign outputs[3736] = (layer0_outputs[1519]) ^ (layer0_outputs[4453]);
    assign outputs[3737] = ~(layer0_outputs[4812]);
    assign outputs[3738] = (layer0_outputs[4315]) & ~(layer0_outputs[4668]);
    assign outputs[3739] = ~(layer0_outputs[7]);
    assign outputs[3740] = ~((layer0_outputs[4332]) ^ (layer0_outputs[4821]));
    assign outputs[3741] = layer0_outputs[2998];
    assign outputs[3742] = layer0_outputs[2696];
    assign outputs[3743] = ~(layer0_outputs[4614]);
    assign outputs[3744] = ~(layer0_outputs[875]);
    assign outputs[3745] = layer0_outputs[344];
    assign outputs[3746] = ~((layer0_outputs[3645]) ^ (layer0_outputs[4400]));
    assign outputs[3747] = ~(layer0_outputs[375]) | (layer0_outputs[2138]);
    assign outputs[3748] = (layer0_outputs[559]) & ~(layer0_outputs[856]);
    assign outputs[3749] = (layer0_outputs[3996]) ^ (layer0_outputs[2540]);
    assign outputs[3750] = (layer0_outputs[3323]) ^ (layer0_outputs[1533]);
    assign outputs[3751] = ~((layer0_outputs[4217]) ^ (layer0_outputs[1477]));
    assign outputs[3752] = (layer0_outputs[4181]) ^ (layer0_outputs[1007]);
    assign outputs[3753] = (layer0_outputs[4544]) | (layer0_outputs[346]);
    assign outputs[3754] = (layer0_outputs[1992]) & ~(layer0_outputs[2333]);
    assign outputs[3755] = (layer0_outputs[4531]) & (layer0_outputs[3412]);
    assign outputs[3756] = layer0_outputs[4389];
    assign outputs[3757] = ~((layer0_outputs[1289]) & (layer0_outputs[1394]));
    assign outputs[3758] = 1'b0;
    assign outputs[3759] = layer0_outputs[4565];
    assign outputs[3760] = ~(layer0_outputs[4385]);
    assign outputs[3761] = (layer0_outputs[1580]) & (layer0_outputs[5069]);
    assign outputs[3762] = ~((layer0_outputs[618]) ^ (layer0_outputs[3941]));
    assign outputs[3763] = (layer0_outputs[247]) & ~(layer0_outputs[1267]);
    assign outputs[3764] = (layer0_outputs[2754]) ^ (layer0_outputs[3524]);
    assign outputs[3765] = layer0_outputs[4132];
    assign outputs[3766] = (layer0_outputs[4251]) & (layer0_outputs[575]);
    assign outputs[3767] = (layer0_outputs[1150]) & ~(layer0_outputs[498]);
    assign outputs[3768] = ~(layer0_outputs[2459]);
    assign outputs[3769] = layer0_outputs[788];
    assign outputs[3770] = layer0_outputs[973];
    assign outputs[3771] = ~((layer0_outputs[2670]) ^ (layer0_outputs[4345]));
    assign outputs[3772] = (layer0_outputs[4588]) | (layer0_outputs[2331]);
    assign outputs[3773] = ~((layer0_outputs[4608]) | (layer0_outputs[2841]));
    assign outputs[3774] = ~((layer0_outputs[1613]) | (layer0_outputs[100]));
    assign outputs[3775] = ~(layer0_outputs[2369]);
    assign outputs[3776] = layer0_outputs[451];
    assign outputs[3777] = ~((layer0_outputs[2433]) | (layer0_outputs[2794]));
    assign outputs[3778] = ~(layer0_outputs[3039]);
    assign outputs[3779] = ~((layer0_outputs[3385]) | (layer0_outputs[4613]));
    assign outputs[3780] = layer0_outputs[4184];
    assign outputs[3781] = (layer0_outputs[4340]) & (layer0_outputs[2952]);
    assign outputs[3782] = (layer0_outputs[2425]) & (layer0_outputs[3840]);
    assign outputs[3783] = ~(layer0_outputs[4474]) | (layer0_outputs[2334]);
    assign outputs[3784] = ~(layer0_outputs[2888]);
    assign outputs[3785] = ~(layer0_outputs[4253]);
    assign outputs[3786] = (layer0_outputs[1600]) & ~(layer0_outputs[1326]);
    assign outputs[3787] = (layer0_outputs[4598]) ^ (layer0_outputs[2969]);
    assign outputs[3788] = layer0_outputs[4735];
    assign outputs[3789] = (layer0_outputs[138]) ^ (layer0_outputs[2946]);
    assign outputs[3790] = (layer0_outputs[1083]) & (layer0_outputs[2021]);
    assign outputs[3791] = (layer0_outputs[256]) & ~(layer0_outputs[2275]);
    assign outputs[3792] = (layer0_outputs[2578]) ^ (layer0_outputs[4688]);
    assign outputs[3793] = ~((layer0_outputs[376]) | (layer0_outputs[2411]));
    assign outputs[3794] = layer0_outputs[685];
    assign outputs[3795] = ~(layer0_outputs[3145]);
    assign outputs[3796] = ~(layer0_outputs[1996]) | (layer0_outputs[407]);
    assign outputs[3797] = (layer0_outputs[264]) & ~(layer0_outputs[4167]);
    assign outputs[3798] = (layer0_outputs[510]) & ~(layer0_outputs[2695]);
    assign outputs[3799] = ~(layer0_outputs[147]);
    assign outputs[3800] = ~((layer0_outputs[1708]) ^ (layer0_outputs[4738]));
    assign outputs[3801] = ~(layer0_outputs[3160]);
    assign outputs[3802] = ~((layer0_outputs[2597]) | (layer0_outputs[4835]));
    assign outputs[3803] = layer0_outputs[4792];
    assign outputs[3804] = ~(layer0_outputs[2350]);
    assign outputs[3805] = ~(layer0_outputs[4388]);
    assign outputs[3806] = ~(layer0_outputs[640]) | (layer0_outputs[114]);
    assign outputs[3807] = (layer0_outputs[251]) & ~(layer0_outputs[1704]);
    assign outputs[3808] = ~(layer0_outputs[4561]);
    assign outputs[3809] = (layer0_outputs[964]) & (layer0_outputs[934]);
    assign outputs[3810] = layer0_outputs[1258];
    assign outputs[3811] = ~((layer0_outputs[1923]) ^ (layer0_outputs[3619]));
    assign outputs[3812] = (layer0_outputs[2421]) & ~(layer0_outputs[5076]);
    assign outputs[3813] = (layer0_outputs[3271]) & (layer0_outputs[892]);
    assign outputs[3814] = ~((layer0_outputs[2123]) ^ (layer0_outputs[832]));
    assign outputs[3815] = ~((layer0_outputs[3797]) ^ (layer0_outputs[1763]));
    assign outputs[3816] = ~((layer0_outputs[2376]) ^ (layer0_outputs[2426]));
    assign outputs[3817] = ~((layer0_outputs[4189]) ^ (layer0_outputs[3981]));
    assign outputs[3818] = (layer0_outputs[4064]) ^ (layer0_outputs[4298]);
    assign outputs[3819] = ~(layer0_outputs[1056]);
    assign outputs[3820] = layer0_outputs[3584];
    assign outputs[3821] = (layer0_outputs[1064]) & (layer0_outputs[4421]);
    assign outputs[3822] = ~((layer0_outputs[2680]) ^ (layer0_outputs[474]));
    assign outputs[3823] = ~(layer0_outputs[3357]);
    assign outputs[3824] = (layer0_outputs[3673]) & (layer0_outputs[4357]);
    assign outputs[3825] = ~((layer0_outputs[3965]) | (layer0_outputs[3556]));
    assign outputs[3826] = (layer0_outputs[1713]) ^ (layer0_outputs[4643]);
    assign outputs[3827] = (layer0_outputs[3755]) ^ (layer0_outputs[3413]);
    assign outputs[3828] = (layer0_outputs[2774]) & ~(layer0_outputs[3664]);
    assign outputs[3829] = (layer0_outputs[2606]) & ~(layer0_outputs[3321]);
    assign outputs[3830] = (layer0_outputs[4085]) ^ (layer0_outputs[3443]);
    assign outputs[3831] = ~((layer0_outputs[4445]) | (layer0_outputs[3722]));
    assign outputs[3832] = ~(layer0_outputs[4931]);
    assign outputs[3833] = (layer0_outputs[2410]) ^ (layer0_outputs[3378]);
    assign outputs[3834] = layer0_outputs[451];
    assign outputs[3835] = layer0_outputs[420];
    assign outputs[3836] = ~(layer0_outputs[1764]);
    assign outputs[3837] = (layer0_outputs[4626]) ^ (layer0_outputs[3823]);
    assign outputs[3838] = (layer0_outputs[527]) ^ (layer0_outputs[2184]);
    assign outputs[3839] = ~(layer0_outputs[1899]) | (layer0_outputs[3378]);
    assign outputs[3840] = (layer0_outputs[561]) | (layer0_outputs[3692]);
    assign outputs[3841] = layer0_outputs[3498];
    assign outputs[3842] = layer0_outputs[2359];
    assign outputs[3843] = ~((layer0_outputs[1966]) ^ (layer0_outputs[1094]));
    assign outputs[3844] = ~(layer0_outputs[749]);
    assign outputs[3845] = (layer0_outputs[2007]) ^ (layer0_outputs[4181]);
    assign outputs[3846] = layer0_outputs[1126];
    assign outputs[3847] = layer0_outputs[800];
    assign outputs[3848] = ~((layer0_outputs[495]) & (layer0_outputs[4325]));
    assign outputs[3849] = (layer0_outputs[365]) & (layer0_outputs[1114]);
    assign outputs[3850] = (layer0_outputs[4823]) ^ (layer0_outputs[4993]);
    assign outputs[3851] = (layer0_outputs[4362]) & ~(layer0_outputs[3853]);
    assign outputs[3852] = ~(layer0_outputs[3036]);
    assign outputs[3853] = ~(layer0_outputs[701]);
    assign outputs[3854] = (layer0_outputs[3766]) & ~(layer0_outputs[244]);
    assign outputs[3855] = ~((layer0_outputs[4566]) | (layer0_outputs[2293]));
    assign outputs[3856] = (layer0_outputs[66]) | (layer0_outputs[4951]);
    assign outputs[3857] = (layer0_outputs[3197]) & ~(layer0_outputs[574]);
    assign outputs[3858] = layer0_outputs[218];
    assign outputs[3859] = layer0_outputs[933];
    assign outputs[3860] = ~((layer0_outputs[3496]) ^ (layer0_outputs[74]));
    assign outputs[3861] = ~((layer0_outputs[4252]) ^ (layer0_outputs[4975]));
    assign outputs[3862] = (layer0_outputs[3127]) | (layer0_outputs[2196]);
    assign outputs[3863] = (layer0_outputs[1040]) ^ (layer0_outputs[2850]);
    assign outputs[3864] = ~((layer0_outputs[3707]) | (layer0_outputs[870]));
    assign outputs[3865] = (layer0_outputs[692]) & ~(layer0_outputs[4921]);
    assign outputs[3866] = layer0_outputs[3071];
    assign outputs[3867] = ~(layer0_outputs[2716]);
    assign outputs[3868] = (layer0_outputs[4697]) & (layer0_outputs[4251]);
    assign outputs[3869] = ~(layer0_outputs[2549]);
    assign outputs[3870] = layer0_outputs[1808];
    assign outputs[3871] = layer0_outputs[3779];
    assign outputs[3872] = (layer0_outputs[265]) & ~(layer0_outputs[412]);
    assign outputs[3873] = ~(layer0_outputs[3726]);
    assign outputs[3874] = (layer0_outputs[4117]) & ~(layer0_outputs[2485]);
    assign outputs[3875] = ~(layer0_outputs[1184]) | (layer0_outputs[502]);
    assign outputs[3876] = (layer0_outputs[4279]) & ~(layer0_outputs[1648]);
    assign outputs[3877] = ~((layer0_outputs[4393]) | (layer0_outputs[27]));
    assign outputs[3878] = ~(layer0_outputs[3456]) | (layer0_outputs[2089]);
    assign outputs[3879] = (layer0_outputs[1298]) ^ (layer0_outputs[2462]);
    assign outputs[3880] = ~((layer0_outputs[4987]) ^ (layer0_outputs[1414]));
    assign outputs[3881] = ~(layer0_outputs[3256]);
    assign outputs[3882] = ~((layer0_outputs[1741]) ^ (layer0_outputs[71]));
    assign outputs[3883] = ~(layer0_outputs[4174]);
    assign outputs[3884] = layer0_outputs[2629];
    assign outputs[3885] = (layer0_outputs[5058]) ^ (layer0_outputs[4031]);
    assign outputs[3886] = ~((layer0_outputs[1782]) ^ (layer0_outputs[1523]));
    assign outputs[3887] = layer0_outputs[409];
    assign outputs[3888] = (layer0_outputs[2627]) & ~(layer0_outputs[2718]);
    assign outputs[3889] = (layer0_outputs[123]) ^ (layer0_outputs[2594]);
    assign outputs[3890] = layer0_outputs[1355];
    assign outputs[3891] = ~(layer0_outputs[1597]);
    assign outputs[3892] = (layer0_outputs[382]) & (layer0_outputs[2811]);
    assign outputs[3893] = layer0_outputs[1997];
    assign outputs[3894] = ~((layer0_outputs[904]) | (layer0_outputs[1192]));
    assign outputs[3895] = layer0_outputs[4511];
    assign outputs[3896] = ~((layer0_outputs[2413]) | (layer0_outputs[3529]));
    assign outputs[3897] = (layer0_outputs[4869]) & (layer0_outputs[265]);
    assign outputs[3898] = (layer0_outputs[5028]) ^ (layer0_outputs[3447]);
    assign outputs[3899] = ~(layer0_outputs[155]);
    assign outputs[3900] = ~(layer0_outputs[1334]);
    assign outputs[3901] = (layer0_outputs[1993]) ^ (layer0_outputs[2060]);
    assign outputs[3902] = layer0_outputs[261];
    assign outputs[3903] = layer0_outputs[2266];
    assign outputs[3904] = ~((layer0_outputs[4236]) | (layer0_outputs[4102]));
    assign outputs[3905] = ~(layer0_outputs[1985]) | (layer0_outputs[3873]);
    assign outputs[3906] = ~(layer0_outputs[4890]);
    assign outputs[3907] = layer0_outputs[3304];
    assign outputs[3908] = (layer0_outputs[1890]) ^ (layer0_outputs[4187]);
    assign outputs[3909] = layer0_outputs[40];
    assign outputs[3910] = layer0_outputs[3449];
    assign outputs[3911] = layer0_outputs[4333];
    assign outputs[3912] = (layer0_outputs[3218]) & ~(layer0_outputs[3885]);
    assign outputs[3913] = layer0_outputs[2101];
    assign outputs[3914] = (layer0_outputs[5015]) & ~(layer0_outputs[2676]);
    assign outputs[3915] = (layer0_outputs[755]) & ~(layer0_outputs[4845]);
    assign outputs[3916] = ~(layer0_outputs[1717]);
    assign outputs[3917] = layer0_outputs[2647];
    assign outputs[3918] = (layer0_outputs[4926]) & (layer0_outputs[413]);
    assign outputs[3919] = layer0_outputs[2396];
    assign outputs[3920] = layer0_outputs[1934];
    assign outputs[3921] = ~(layer0_outputs[2215]);
    assign outputs[3922] = (layer0_outputs[1863]) ^ (layer0_outputs[1008]);
    assign outputs[3923] = ~(layer0_outputs[3783]);
    assign outputs[3924] = (layer0_outputs[1560]) & ~(layer0_outputs[2587]);
    assign outputs[3925] = ~(layer0_outputs[2172]) | (layer0_outputs[4070]);
    assign outputs[3926] = (layer0_outputs[4752]) & ~(layer0_outputs[389]);
    assign outputs[3927] = (layer0_outputs[4320]) & ~(layer0_outputs[2503]);
    assign outputs[3928] = ~(layer0_outputs[4408]);
    assign outputs[3929] = ~(layer0_outputs[215]);
    assign outputs[3930] = (layer0_outputs[2196]) | (layer0_outputs[4810]);
    assign outputs[3931] = (layer0_outputs[2518]) & (layer0_outputs[3975]);
    assign outputs[3932] = (layer0_outputs[3630]) & ~(layer0_outputs[3038]);
    assign outputs[3933] = ~(layer0_outputs[4081]) | (layer0_outputs[2010]);
    assign outputs[3934] = (layer0_outputs[3689]) ^ (layer0_outputs[4575]);
    assign outputs[3935] = layer0_outputs[4195];
    assign outputs[3936] = ~((layer0_outputs[535]) ^ (layer0_outputs[959]));
    assign outputs[3937] = ~(layer0_outputs[781]);
    assign outputs[3938] = ~((layer0_outputs[3015]) | (layer0_outputs[2469]));
    assign outputs[3939] = (layer0_outputs[1555]) ^ (layer0_outputs[3309]);
    assign outputs[3940] = ~((layer0_outputs[2524]) | (layer0_outputs[76]));
    assign outputs[3941] = (layer0_outputs[1207]) & ~(layer0_outputs[3207]);
    assign outputs[3942] = ~((layer0_outputs[2179]) | (layer0_outputs[780]));
    assign outputs[3943] = ~((layer0_outputs[3168]) ^ (layer0_outputs[1026]));
    assign outputs[3944] = (layer0_outputs[1629]) ^ (layer0_outputs[2085]);
    assign outputs[3945] = layer0_outputs[4242];
    assign outputs[3946] = (layer0_outputs[3495]) & ~(layer0_outputs[4194]);
    assign outputs[3947] = (layer0_outputs[1257]) ^ (layer0_outputs[1196]);
    assign outputs[3948] = (layer0_outputs[2533]) & (layer0_outputs[2926]);
    assign outputs[3949] = layer0_outputs[4947];
    assign outputs[3950] = (layer0_outputs[3603]) & ~(layer0_outputs[4174]);
    assign outputs[3951] = (layer0_outputs[395]) & (layer0_outputs[4522]);
    assign outputs[3952] = ~((layer0_outputs[3459]) ^ (layer0_outputs[3255]));
    assign outputs[3953] = (layer0_outputs[3630]) ^ (layer0_outputs[2137]);
    assign outputs[3954] = (layer0_outputs[3458]) & ~(layer0_outputs[415]);
    assign outputs[3955] = (layer0_outputs[4216]) & ~(layer0_outputs[5114]);
    assign outputs[3956] = ~(layer0_outputs[913]);
    assign outputs[3957] = 1'b0;
    assign outputs[3958] = ~(layer0_outputs[3688]);
    assign outputs[3959] = layer0_outputs[1861];
    assign outputs[3960] = (layer0_outputs[3835]) & (layer0_outputs[4235]);
    assign outputs[3961] = ~((layer0_outputs[3242]) ^ (layer0_outputs[2821]));
    assign outputs[3962] = ~((layer0_outputs[3048]) ^ (layer0_outputs[2470]));
    assign outputs[3963] = ~(layer0_outputs[2634]);
    assign outputs[3964] = ~((layer0_outputs[2248]) ^ (layer0_outputs[4564]));
    assign outputs[3965] = (layer0_outputs[4192]) ^ (layer0_outputs[2443]);
    assign outputs[3966] = layer0_outputs[3618];
    assign outputs[3967] = layer0_outputs[2975];
    assign outputs[3968] = ~((layer0_outputs[2032]) ^ (layer0_outputs[3739]));
    assign outputs[3969] = ~(layer0_outputs[2292]);
    assign outputs[3970] = layer0_outputs[93];
    assign outputs[3971] = ~((layer0_outputs[625]) ^ (layer0_outputs[1205]));
    assign outputs[3972] = (layer0_outputs[4777]) & (layer0_outputs[1303]);
    assign outputs[3973] = ~((layer0_outputs[3162]) ^ (layer0_outputs[4026]));
    assign outputs[3974] = ~(layer0_outputs[1912]);
    assign outputs[3975] = layer0_outputs[744];
    assign outputs[3976] = ~(layer0_outputs[4058]);
    assign outputs[3977] = (layer0_outputs[1222]) & ~(layer0_outputs[5071]);
    assign outputs[3978] = ~(layer0_outputs[3578]) | (layer0_outputs[2590]);
    assign outputs[3979] = ~(layer0_outputs[4942]);
    assign outputs[3980] = ~(layer0_outputs[540]);
    assign outputs[3981] = layer0_outputs[1758];
    assign outputs[3982] = ~((layer0_outputs[1652]) & (layer0_outputs[1193]));
    assign outputs[3983] = ~(layer0_outputs[5033]);
    assign outputs[3984] = ~((layer0_outputs[2287]) ^ (layer0_outputs[3159]));
    assign outputs[3985] = ~(layer0_outputs[1268]) | (layer0_outputs[70]);
    assign outputs[3986] = (layer0_outputs[1682]) ^ (layer0_outputs[320]);
    assign outputs[3987] = layer0_outputs[3796];
    assign outputs[3988] = ~(layer0_outputs[1565]);
    assign outputs[3989] = ~(layer0_outputs[4434]);
    assign outputs[3990] = layer0_outputs[3079];
    assign outputs[3991] = (layer0_outputs[3943]) & ~(layer0_outputs[5032]);
    assign outputs[3992] = ~(layer0_outputs[4168]);
    assign outputs[3993] = (layer0_outputs[5009]) & (layer0_outputs[232]);
    assign outputs[3994] = layer0_outputs[2675];
    assign outputs[3995] = (layer0_outputs[4446]) & ~(layer0_outputs[2335]);
    assign outputs[3996] = ~((layer0_outputs[543]) ^ (layer0_outputs[5028]));
    assign outputs[3997] = ~(layer0_outputs[3268]);
    assign outputs[3998] = layer0_outputs[1698];
    assign outputs[3999] = (layer0_outputs[2496]) ^ (layer0_outputs[3738]);
    assign outputs[4000] = layer0_outputs[1282];
    assign outputs[4001] = ~((layer0_outputs[4377]) ^ (layer0_outputs[3438]));
    assign outputs[4002] = (layer0_outputs[2808]) & (layer0_outputs[4373]);
    assign outputs[4003] = (layer0_outputs[2255]) & ~(layer0_outputs[4966]);
    assign outputs[4004] = layer0_outputs[299];
    assign outputs[4005] = ~(layer0_outputs[901]);
    assign outputs[4006] = ~(layer0_outputs[2105]);
    assign outputs[4007] = (layer0_outputs[3839]) ^ (layer0_outputs[2384]);
    assign outputs[4008] = (layer0_outputs[3804]) ^ (layer0_outputs[1291]);
    assign outputs[4009] = (layer0_outputs[3356]) ^ (layer0_outputs[3833]);
    assign outputs[4010] = ~((layer0_outputs[1304]) | (layer0_outputs[4155]));
    assign outputs[4011] = ~((layer0_outputs[2092]) | (layer0_outputs[1359]));
    assign outputs[4012] = (layer0_outputs[4442]) & ~(layer0_outputs[2039]);
    assign outputs[4013] = ~(layer0_outputs[458]);
    assign outputs[4014] = ~((layer0_outputs[4709]) ^ (layer0_outputs[1412]));
    assign outputs[4015] = (layer0_outputs[3274]) & ~(layer0_outputs[1702]);
    assign outputs[4016] = ~(layer0_outputs[1022]);
    assign outputs[4017] = (layer0_outputs[4281]) & ~(layer0_outputs[955]);
    assign outputs[4018] = layer0_outputs[4379];
    assign outputs[4019] = (layer0_outputs[2243]) ^ (layer0_outputs[2065]);
    assign outputs[4020] = ~(layer0_outputs[4594]);
    assign outputs[4021] = ~(layer0_outputs[2612]);
    assign outputs[4022] = ~(layer0_outputs[862]);
    assign outputs[4023] = (layer0_outputs[4960]) & ~(layer0_outputs[5098]);
    assign outputs[4024] = ~((layer0_outputs[513]) & (layer0_outputs[5073]));
    assign outputs[4025] = layer0_outputs[3656];
    assign outputs[4026] = (layer0_outputs[4221]) ^ (layer0_outputs[1593]);
    assign outputs[4027] = (layer0_outputs[923]) & (layer0_outputs[2119]);
    assign outputs[4028] = (layer0_outputs[2217]) & (layer0_outputs[4222]);
    assign outputs[4029] = ~(layer0_outputs[4461]);
    assign outputs[4030] = ~((layer0_outputs[1670]) | (layer0_outputs[3516]));
    assign outputs[4031] = ~(layer0_outputs[2515]) | (layer0_outputs[2904]);
    assign outputs[4032] = layer0_outputs[2210];
    assign outputs[4033] = layer0_outputs[1424];
    assign outputs[4034] = ~((layer0_outputs[4688]) ^ (layer0_outputs[4674]));
    assign outputs[4035] = layer0_outputs[1361];
    assign outputs[4036] = layer0_outputs[80];
    assign outputs[4037] = (layer0_outputs[1692]) & ~(layer0_outputs[3208]);
    assign outputs[4038] = ~(layer0_outputs[5099]);
    assign outputs[4039] = (layer0_outputs[1010]) & ~(layer0_outputs[1750]);
    assign outputs[4040] = 1'b0;
    assign outputs[4041] = ~(layer0_outputs[1511]);
    assign outputs[4042] = layer0_outputs[5103];
    assign outputs[4043] = ~((layer0_outputs[4770]) | (layer0_outputs[2799]));
    assign outputs[4044] = ~((layer0_outputs[2967]) ^ (layer0_outputs[1192]));
    assign outputs[4045] = (layer0_outputs[1658]) & ~(layer0_outputs[4633]);
    assign outputs[4046] = layer0_outputs[3386];
    assign outputs[4047] = ~(layer0_outputs[1855]);
    assign outputs[4048] = ~(layer0_outputs[4190]);
    assign outputs[4049] = ~(layer0_outputs[2710]) | (layer0_outputs[653]);
    assign outputs[4050] = (layer0_outputs[744]) & (layer0_outputs[3972]);
    assign outputs[4051] = (layer0_outputs[4619]) & (layer0_outputs[4593]);
    assign outputs[4052] = layer0_outputs[4467];
    assign outputs[4053] = ~(layer0_outputs[1541]);
    assign outputs[4054] = ~(layer0_outputs[3328]);
    assign outputs[4055] = ~((layer0_outputs[797]) ^ (layer0_outputs[2933]));
    assign outputs[4056] = 1'b0;
    assign outputs[4057] = layer0_outputs[1510];
    assign outputs[4058] = (layer0_outputs[1759]) | (layer0_outputs[1632]);
    assign outputs[4059] = layer0_outputs[3807];
    assign outputs[4060] = (layer0_outputs[1601]) & ~(layer0_outputs[1322]);
    assign outputs[4061] = ~(layer0_outputs[778]);
    assign outputs[4062] = (layer0_outputs[3013]) & ~(layer0_outputs[3107]);
    assign outputs[4063] = ~(layer0_outputs[3817]);
    assign outputs[4064] = layer0_outputs[2887];
    assign outputs[4065] = (layer0_outputs[731]) ^ (layer0_outputs[1778]);
    assign outputs[4066] = ~(layer0_outputs[2599]);
    assign outputs[4067] = ~((layer0_outputs[4973]) & (layer0_outputs[5000]));
    assign outputs[4068] = (layer0_outputs[1547]) ^ (layer0_outputs[4995]);
    assign outputs[4069] = (layer0_outputs[2158]) & ~(layer0_outputs[250]);
    assign outputs[4070] = ~((layer0_outputs[280]) ^ (layer0_outputs[2940]));
    assign outputs[4071] = layer0_outputs[1570];
    assign outputs[4072] = layer0_outputs[1145];
    assign outputs[4073] = (layer0_outputs[4950]) & (layer0_outputs[2142]);
    assign outputs[4074] = ~(layer0_outputs[521]);
    assign outputs[4075] = ~(layer0_outputs[3368]);
    assign outputs[4076] = ~(layer0_outputs[1069]);
    assign outputs[4077] = ~((layer0_outputs[4542]) | (layer0_outputs[3785]));
    assign outputs[4078] = ~((layer0_outputs[2786]) | (layer0_outputs[4270]));
    assign outputs[4079] = layer0_outputs[2396];
    assign outputs[4080] = (layer0_outputs[3059]) & ~(layer0_outputs[2660]);
    assign outputs[4081] = ~(layer0_outputs[252]);
    assign outputs[4082] = ~((layer0_outputs[1434]) | (layer0_outputs[1013]));
    assign outputs[4083] = ~(layer0_outputs[3896]) | (layer0_outputs[4999]);
    assign outputs[4084] = ~(layer0_outputs[329]);
    assign outputs[4085] = layer0_outputs[3906];
    assign outputs[4086] = (layer0_outputs[13]) ^ (layer0_outputs[2285]);
    assign outputs[4087] = ~((layer0_outputs[4540]) ^ (layer0_outputs[116]));
    assign outputs[4088] = layer0_outputs[163];
    assign outputs[4089] = (layer0_outputs[3580]) & ~(layer0_outputs[147]);
    assign outputs[4090] = (layer0_outputs[506]) | (layer0_outputs[1545]);
    assign outputs[4091] = ~((layer0_outputs[411]) | (layer0_outputs[3519]));
    assign outputs[4092] = (layer0_outputs[2244]) & (layer0_outputs[3956]);
    assign outputs[4093] = layer0_outputs[1630];
    assign outputs[4094] = ~((layer0_outputs[4010]) | (layer0_outputs[4023]));
    assign outputs[4095] = (layer0_outputs[4963]) & (layer0_outputs[1585]);
    assign outputs[4096] = ~((layer0_outputs[5067]) | (layer0_outputs[3829]));
    assign outputs[4097] = ~(layer0_outputs[1134]);
    assign outputs[4098] = (layer0_outputs[5]) & ~(layer0_outputs[481]);
    assign outputs[4099] = ~(layer0_outputs[954]);
    assign outputs[4100] = layer0_outputs[351];
    assign outputs[4101] = ~(layer0_outputs[4825]);
    assign outputs[4102] = layer0_outputs[2488];
    assign outputs[4103] = (layer0_outputs[4905]) ^ (layer0_outputs[1889]);
    assign outputs[4104] = ~(layer0_outputs[3950]);
    assign outputs[4105] = ~((layer0_outputs[4294]) ^ (layer0_outputs[1309]));
    assign outputs[4106] = layer0_outputs[2073];
    assign outputs[4107] = (layer0_outputs[2979]) & ~(layer0_outputs[752]);
    assign outputs[4108] = ~((layer0_outputs[1914]) ^ (layer0_outputs[4533]));
    assign outputs[4109] = (layer0_outputs[3654]) | (layer0_outputs[1680]);
    assign outputs[4110] = (layer0_outputs[229]) & ~(layer0_outputs[2386]);
    assign outputs[4111] = ~(layer0_outputs[4543]) | (layer0_outputs[3789]);
    assign outputs[4112] = ~(layer0_outputs[4438]) | (layer0_outputs[3319]);
    assign outputs[4113] = (layer0_outputs[2085]) & ~(layer0_outputs[4405]);
    assign outputs[4114] = ~(layer0_outputs[4933]) | (layer0_outputs[3078]);
    assign outputs[4115] = ~(layer0_outputs[4247]);
    assign outputs[4116] = (layer0_outputs[1346]) | (layer0_outputs[3635]);
    assign outputs[4117] = ~(layer0_outputs[3983]);
    assign outputs[4118] = (layer0_outputs[3874]) & ~(layer0_outputs[870]);
    assign outputs[4119] = (layer0_outputs[4338]) & (layer0_outputs[3340]);
    assign outputs[4120] = layer0_outputs[2006];
    assign outputs[4121] = ~(layer0_outputs[4534]);
    assign outputs[4122] = ~(layer0_outputs[707]);
    assign outputs[4123] = (layer0_outputs[4694]) ^ (layer0_outputs[4463]);
    assign outputs[4124] = (layer0_outputs[3452]) | (layer0_outputs[3143]);
    assign outputs[4125] = (layer0_outputs[1765]) & (layer0_outputs[2507]);
    assign outputs[4126] = ~((layer0_outputs[3120]) ^ (layer0_outputs[1435]));
    assign outputs[4127] = ~(layer0_outputs[4712]);
    assign outputs[4128] = (layer0_outputs[2784]) & (layer0_outputs[1012]);
    assign outputs[4129] = ~(layer0_outputs[646]);
    assign outputs[4130] = layer0_outputs[421];
    assign outputs[4131] = ~(layer0_outputs[2668]);
    assign outputs[4132] = (layer0_outputs[1804]) ^ (layer0_outputs[1677]);
    assign outputs[4133] = ~(layer0_outputs[981]) | (layer0_outputs[1986]);
    assign outputs[4134] = (layer0_outputs[71]) | (layer0_outputs[2875]);
    assign outputs[4135] = 1'b1;
    assign outputs[4136] = layer0_outputs[3469];
    assign outputs[4137] = ~(layer0_outputs[1352]);
    assign outputs[4138] = ~(layer0_outputs[881]) | (layer0_outputs[2970]);
    assign outputs[4139] = ~((layer0_outputs[396]) & (layer0_outputs[1677]));
    assign outputs[4140] = (layer0_outputs[644]) | (layer0_outputs[3911]);
    assign outputs[4141] = ~(layer0_outputs[815]);
    assign outputs[4142] = (layer0_outputs[1204]) & ~(layer0_outputs[4323]);
    assign outputs[4143] = layer0_outputs[4607];
    assign outputs[4144] = ~(layer0_outputs[4853]) | (layer0_outputs[3651]);
    assign outputs[4145] = ~(layer0_outputs[638]);
    assign outputs[4146] = layer0_outputs[1266];
    assign outputs[4147] = ~((layer0_outputs[1916]) ^ (layer0_outputs[3959]));
    assign outputs[4148] = ~(layer0_outputs[4961]);
    assign outputs[4149] = layer0_outputs[4331];
    assign outputs[4150] = layer0_outputs[443];
    assign outputs[4151] = 1'b1;
    assign outputs[4152] = layer0_outputs[2909];
    assign outputs[4153] = (layer0_outputs[33]) & (layer0_outputs[1091]);
    assign outputs[4154] = ~(layer0_outputs[1840]) | (layer0_outputs[3275]);
    assign outputs[4155] = ~(layer0_outputs[2951]) | (layer0_outputs[2000]);
    assign outputs[4156] = ~(layer0_outputs[5088]) | (layer0_outputs[680]);
    assign outputs[4157] = ~((layer0_outputs[634]) | (layer0_outputs[1830]));
    assign outputs[4158] = ~((layer0_outputs[4606]) ^ (layer0_outputs[4997]));
    assign outputs[4159] = ~(layer0_outputs[3374]) | (layer0_outputs[2475]);
    assign outputs[4160] = layer0_outputs[2415];
    assign outputs[4161] = ~(layer0_outputs[2287]);
    assign outputs[4162] = ~(layer0_outputs[2629]);
    assign outputs[4163] = (layer0_outputs[4156]) & ~(layer0_outputs[202]);
    assign outputs[4164] = ~((layer0_outputs[3047]) | (layer0_outputs[391]));
    assign outputs[4165] = ~(layer0_outputs[1501]) | (layer0_outputs[2733]);
    assign outputs[4166] = (layer0_outputs[695]) ^ (layer0_outputs[5098]);
    assign outputs[4167] = ~((layer0_outputs[3228]) | (layer0_outputs[2290]));
    assign outputs[4168] = (layer0_outputs[924]) | (layer0_outputs[2768]);
    assign outputs[4169] = ~(layer0_outputs[305]);
    assign outputs[4170] = (layer0_outputs[2432]) & ~(layer0_outputs[1434]);
    assign outputs[4171] = layer0_outputs[2749];
    assign outputs[4172] = (layer0_outputs[1564]) & (layer0_outputs[1542]);
    assign outputs[4173] = layer0_outputs[1116];
    assign outputs[4174] = (layer0_outputs[4741]) ^ (layer0_outputs[3364]);
    assign outputs[4175] = (layer0_outputs[1866]) & (layer0_outputs[1395]);
    assign outputs[4176] = ~((layer0_outputs[3217]) ^ (layer0_outputs[3399]));
    assign outputs[4177] = layer0_outputs[4766];
    assign outputs[4178] = ~((layer0_outputs[891]) ^ (layer0_outputs[4791]));
    assign outputs[4179] = ~(layer0_outputs[3004]);
    assign outputs[4180] = ~((layer0_outputs[735]) ^ (layer0_outputs[1977]));
    assign outputs[4181] = (layer0_outputs[2573]) & ~(layer0_outputs[4062]);
    assign outputs[4182] = ~((layer0_outputs[4715]) | (layer0_outputs[419]));
    assign outputs[4183] = (layer0_outputs[1868]) ^ (layer0_outputs[4534]);
    assign outputs[4184] = layer0_outputs[1714];
    assign outputs[4185] = layer0_outputs[4353];
    assign outputs[4186] = ~((layer0_outputs[4149]) | (layer0_outputs[4203]));
    assign outputs[4187] = (layer0_outputs[2964]) | (layer0_outputs[276]);
    assign outputs[4188] = layer0_outputs[289];
    assign outputs[4189] = layer0_outputs[3055];
    assign outputs[4190] = (layer0_outputs[768]) & ~(layer0_outputs[4275]);
    assign outputs[4191] = (layer0_outputs[2100]) ^ (layer0_outputs[16]);
    assign outputs[4192] = ~((layer0_outputs[1767]) ^ (layer0_outputs[2604]));
    assign outputs[4193] = layer0_outputs[1432];
    assign outputs[4194] = layer0_outputs[142];
    assign outputs[4195] = ~(layer0_outputs[2792]);
    assign outputs[4196] = layer0_outputs[4336];
    assign outputs[4197] = layer0_outputs[378];
    assign outputs[4198] = ~(layer0_outputs[2871]);
    assign outputs[4199] = ~(layer0_outputs[3051]) | (layer0_outputs[194]);
    assign outputs[4200] = ~((layer0_outputs[911]) & (layer0_outputs[5074]));
    assign outputs[4201] = (layer0_outputs[2807]) & ~(layer0_outputs[3361]);
    assign outputs[4202] = layer0_outputs[10];
    assign outputs[4203] = ~(layer0_outputs[647]);
    assign outputs[4204] = ~(layer0_outputs[2504]) | (layer0_outputs[3441]);
    assign outputs[4205] = ~(layer0_outputs[4140]) | (layer0_outputs[2702]);
    assign outputs[4206] = layer0_outputs[3855];
    assign outputs[4207] = ~(layer0_outputs[5113]);
    assign outputs[4208] = layer0_outputs[2075];
    assign outputs[4209] = (layer0_outputs[1964]) & (layer0_outputs[150]);
    assign outputs[4210] = (layer0_outputs[1296]) ^ (layer0_outputs[2292]);
    assign outputs[4211] = (layer0_outputs[1620]) & ~(layer0_outputs[4601]);
    assign outputs[4212] = (layer0_outputs[2936]) ^ (layer0_outputs[4371]);
    assign outputs[4213] = layer0_outputs[115];
    assign outputs[4214] = ~((layer0_outputs[1265]) & (layer0_outputs[3513]));
    assign outputs[4215] = layer0_outputs[3795];
    assign outputs[4216] = ~(layer0_outputs[2789]);
    assign outputs[4217] = (layer0_outputs[5094]) ^ (layer0_outputs[3454]);
    assign outputs[4218] = ~((layer0_outputs[4019]) & (layer0_outputs[442]));
    assign outputs[4219] = ~(layer0_outputs[865]);
    assign outputs[4220] = (layer0_outputs[2593]) | (layer0_outputs[3624]);
    assign outputs[4221] = layer0_outputs[1155];
    assign outputs[4222] = ~((layer0_outputs[2450]) & (layer0_outputs[991]));
    assign outputs[4223] = ~((layer0_outputs[2229]) ^ (layer0_outputs[2339]));
    assign outputs[4224] = ~(layer0_outputs[2492]) | (layer0_outputs[4737]);
    assign outputs[4225] = ~(layer0_outputs[2505]);
    assign outputs[4226] = layer0_outputs[2596];
    assign outputs[4227] = ~(layer0_outputs[4575]);
    assign outputs[4228] = ~(layer0_outputs[112]) | (layer0_outputs[1922]);
    assign outputs[4229] = (layer0_outputs[1863]) | (layer0_outputs[4415]);
    assign outputs[4230] = ~(layer0_outputs[2107]);
    assign outputs[4231] = layer0_outputs[55];
    assign outputs[4232] = layer0_outputs[1097];
    assign outputs[4233] = layer0_outputs[198];
    assign outputs[4234] = ~(layer0_outputs[4152]);
    assign outputs[4235] = layer0_outputs[3732];
    assign outputs[4236] = layer0_outputs[4984];
    assign outputs[4237] = ~(layer0_outputs[2606]);
    assign outputs[4238] = layer0_outputs[273];
    assign outputs[4239] = layer0_outputs[4477];
    assign outputs[4240] = layer0_outputs[789];
    assign outputs[4241] = ~((layer0_outputs[4004]) & (layer0_outputs[1942]));
    assign outputs[4242] = ~(layer0_outputs[166]);
    assign outputs[4243] = ~(layer0_outputs[3264]);
    assign outputs[4244] = ~((layer0_outputs[2603]) & (layer0_outputs[3558]));
    assign outputs[4245] = ~(layer0_outputs[783]);
    assign outputs[4246] = ~(layer0_outputs[1873]);
    assign outputs[4247] = ~(layer0_outputs[3248]);
    assign outputs[4248] = (layer0_outputs[3053]) ^ (layer0_outputs[1609]);
    assign outputs[4249] = ~((layer0_outputs[4634]) | (layer0_outputs[3501]));
    assign outputs[4250] = (layer0_outputs[2667]) ^ (layer0_outputs[33]);
    assign outputs[4251] = ~(layer0_outputs[1027]);
    assign outputs[4252] = ~(layer0_outputs[889]) | (layer0_outputs[3414]);
    assign outputs[4253] = (layer0_outputs[2851]) | (layer0_outputs[1579]);
    assign outputs[4254] = ~((layer0_outputs[594]) | (layer0_outputs[458]));
    assign outputs[4255] = ~((layer0_outputs[2136]) & (layer0_outputs[932]));
    assign outputs[4256] = layer0_outputs[1122];
    assign outputs[4257] = layer0_outputs[1940];
    assign outputs[4258] = ~((layer0_outputs[3314]) ^ (layer0_outputs[4700]));
    assign outputs[4259] = layer0_outputs[5093];
    assign outputs[4260] = layer0_outputs[3272];
    assign outputs[4261] = layer0_outputs[4084];
    assign outputs[4262] = (layer0_outputs[1504]) & ~(layer0_outputs[4957]);
    assign outputs[4263] = layer0_outputs[183];
    assign outputs[4264] = (layer0_outputs[3909]) ^ (layer0_outputs[389]);
    assign outputs[4265] = ~((layer0_outputs[122]) ^ (layer0_outputs[2848]));
    assign outputs[4266] = layer0_outputs[4934];
    assign outputs[4267] = ~(layer0_outputs[245]) | (layer0_outputs[5096]);
    assign outputs[4268] = ~(layer0_outputs[2294]);
    assign outputs[4269] = layer0_outputs[3172];
    assign outputs[4270] = (layer0_outputs[3278]) ^ (layer0_outputs[4480]);
    assign outputs[4271] = ~(layer0_outputs[577]);
    assign outputs[4272] = (layer0_outputs[345]) ^ (layer0_outputs[3689]);
    assign outputs[4273] = ~(layer0_outputs[3622]) | (layer0_outputs[1370]);
    assign outputs[4274] = (layer0_outputs[3966]) & ~(layer0_outputs[4086]);
    assign outputs[4275] = layer0_outputs[4215];
    assign outputs[4276] = (layer0_outputs[4067]) ^ (layer0_outputs[3146]);
    assign outputs[4277] = (layer0_outputs[331]) & (layer0_outputs[1972]);
    assign outputs[4278] = ~(layer0_outputs[640]);
    assign outputs[4279] = layer0_outputs[828];
    assign outputs[4280] = (layer0_outputs[34]) ^ (layer0_outputs[1038]);
    assign outputs[4281] = ~((layer0_outputs[3405]) & (layer0_outputs[2966]));
    assign outputs[4282] = ~(layer0_outputs[2870]);
    assign outputs[4283] = ~(layer0_outputs[3347]);
    assign outputs[4284] = layer0_outputs[3646];
    assign outputs[4285] = (layer0_outputs[4095]) ^ (layer0_outputs[2244]);
    assign outputs[4286] = (layer0_outputs[4629]) | (layer0_outputs[4272]);
    assign outputs[4287] = layer0_outputs[59];
    assign outputs[4288] = ~(layer0_outputs[262]) | (layer0_outputs[3233]);
    assign outputs[4289] = ~(layer0_outputs[3639]);
    assign outputs[4290] = ~(layer0_outputs[4444]);
    assign outputs[4291] = ~((layer0_outputs[1377]) ^ (layer0_outputs[1747]));
    assign outputs[4292] = layer0_outputs[789];
    assign outputs[4293] = layer0_outputs[1433];
    assign outputs[4294] = (layer0_outputs[953]) | (layer0_outputs[3187]);
    assign outputs[4295] = (layer0_outputs[4309]) ^ (layer0_outputs[4316]);
    assign outputs[4296] = (layer0_outputs[2126]) ^ (layer0_outputs[2016]);
    assign outputs[4297] = layer0_outputs[1284];
    assign outputs[4298] = ~(layer0_outputs[4717]);
    assign outputs[4299] = layer0_outputs[5083];
    assign outputs[4300] = ~(layer0_outputs[4486]);
    assign outputs[4301] = ~((layer0_outputs[903]) ^ (layer0_outputs[1727]));
    assign outputs[4302] = (layer0_outputs[3508]) & ~(layer0_outputs[3032]);
    assign outputs[4303] = (layer0_outputs[3872]) | (layer0_outputs[2194]);
    assign outputs[4304] = ~((layer0_outputs[1269]) ^ (layer0_outputs[622]));
    assign outputs[4305] = ~(layer0_outputs[22]);
    assign outputs[4306] = (layer0_outputs[1226]) ^ (layer0_outputs[2034]);
    assign outputs[4307] = ~(layer0_outputs[846]);
    assign outputs[4308] = (layer0_outputs[3909]) & ~(layer0_outputs[2133]);
    assign outputs[4309] = (layer0_outputs[2274]) | (layer0_outputs[4866]);
    assign outputs[4310] = layer0_outputs[3411];
    assign outputs[4311] = ~((layer0_outputs[4875]) & (layer0_outputs[439]));
    assign outputs[4312] = layer0_outputs[3802];
    assign outputs[4313] = ~(layer0_outputs[2821]) | (layer0_outputs[1556]);
    assign outputs[4314] = (layer0_outputs[4094]) & ~(layer0_outputs[1785]);
    assign outputs[4315] = (layer0_outputs[4788]) & ~(layer0_outputs[4716]);
    assign outputs[4316] = (layer0_outputs[967]) & ~(layer0_outputs[423]);
    assign outputs[4317] = ~(layer0_outputs[4677]);
    assign outputs[4318] = ~((layer0_outputs[3918]) ^ (layer0_outputs[4041]));
    assign outputs[4319] = layer0_outputs[4107];
    assign outputs[4320] = ~((layer0_outputs[1563]) | (layer0_outputs[2544]));
    assign outputs[4321] = ~((layer0_outputs[1839]) ^ (layer0_outputs[3786]));
    assign outputs[4322] = layer0_outputs[1179];
    assign outputs[4323] = (layer0_outputs[362]) & ~(layer0_outputs[4360]);
    assign outputs[4324] = ~((layer0_outputs[2068]) & (layer0_outputs[3838]));
    assign outputs[4325] = ~(layer0_outputs[3462]) | (layer0_outputs[1340]);
    assign outputs[4326] = layer0_outputs[2814];
    assign outputs[4327] = (layer0_outputs[3775]) & (layer0_outputs[2291]);
    assign outputs[4328] = ~(layer0_outputs[1498]);
    assign outputs[4329] = ~(layer0_outputs[4489]);
    assign outputs[4330] = layer0_outputs[4465];
    assign outputs[4331] = layer0_outputs[3567];
    assign outputs[4332] = ~(layer0_outputs[4504]) | (layer0_outputs[890]);
    assign outputs[4333] = 1'b1;
    assign outputs[4334] = ~(layer0_outputs[303]);
    assign outputs[4335] = (layer0_outputs[2029]) ^ (layer0_outputs[929]);
    assign outputs[4336] = ~(layer0_outputs[1347]);
    assign outputs[4337] = (layer0_outputs[4924]) | (layer0_outputs[4128]);
    assign outputs[4338] = ~(layer0_outputs[4888]);
    assign outputs[4339] = (layer0_outputs[3393]) | (layer0_outputs[4877]);
    assign outputs[4340] = layer0_outputs[131];
    assign outputs[4341] = layer0_outputs[755];
    assign outputs[4342] = ~((layer0_outputs[4068]) ^ (layer0_outputs[2690]));
    assign outputs[4343] = ~(layer0_outputs[4271]);
    assign outputs[4344] = (layer0_outputs[1644]) & ~(layer0_outputs[3353]);
    assign outputs[4345] = ~((layer0_outputs[2466]) ^ (layer0_outputs[2805]));
    assign outputs[4346] = ~(layer0_outputs[2571]);
    assign outputs[4347] = (layer0_outputs[2848]) ^ (layer0_outputs[1096]);
    assign outputs[4348] = ~(layer0_outputs[4032]) | (layer0_outputs[2127]);
    assign outputs[4349] = layer0_outputs[1473];
    assign outputs[4350] = ~(layer0_outputs[2697]) | (layer0_outputs[2417]);
    assign outputs[4351] = ~(layer0_outputs[1756]) | (layer0_outputs[2651]);
    assign outputs[4352] = (layer0_outputs[2499]) & ~(layer0_outputs[726]);
    assign outputs[4353] = ~(layer0_outputs[2729]);
    assign outputs[4354] = layer0_outputs[1095];
    assign outputs[4355] = ~((layer0_outputs[4053]) | (layer0_outputs[864]));
    assign outputs[4356] = (layer0_outputs[1865]) ^ (layer0_outputs[4311]);
    assign outputs[4357] = ~(layer0_outputs[3758]);
    assign outputs[4358] = layer0_outputs[4484];
    assign outputs[4359] = (layer0_outputs[4755]) ^ (layer0_outputs[2637]);
    assign outputs[4360] = ~((layer0_outputs[797]) & (layer0_outputs[1643]));
    assign outputs[4361] = (layer0_outputs[5013]) ^ (layer0_outputs[4270]);
    assign outputs[4362] = ~(layer0_outputs[2208]);
    assign outputs[4363] = (layer0_outputs[3803]) & ~(layer0_outputs[191]);
    assign outputs[4364] = layer0_outputs[1095];
    assign outputs[4365] = ~(layer0_outputs[4073]);
    assign outputs[4366] = layer0_outputs[1969];
    assign outputs[4367] = (layer0_outputs[1984]) & (layer0_outputs[1868]);
    assign outputs[4368] = ~(layer0_outputs[3132]) | (layer0_outputs[3318]);
    assign outputs[4369] = ~((layer0_outputs[2921]) | (layer0_outputs[4728]));
    assign outputs[4370] = (layer0_outputs[3930]) | (layer0_outputs[4430]);
    assign outputs[4371] = ~(layer0_outputs[2845]);
    assign outputs[4372] = ~(layer0_outputs[4970]) | (layer0_outputs[3016]);
    assign outputs[4373] = ~((layer0_outputs[4623]) ^ (layer0_outputs[3330]));
    assign outputs[4374] = (layer0_outputs[3254]) | (layer0_outputs[1738]);
    assign outputs[4375] = layer0_outputs[1641];
    assign outputs[4376] = layer0_outputs[54];
    assign outputs[4377] = ~((layer0_outputs[497]) | (layer0_outputs[996]));
    assign outputs[4378] = (layer0_outputs[192]) & (layer0_outputs[4909]);
    assign outputs[4379] = ~((layer0_outputs[4708]) & (layer0_outputs[3536]));
    assign outputs[4380] = ~((layer0_outputs[2871]) ^ (layer0_outputs[3325]));
    assign outputs[4381] = ~((layer0_outputs[3922]) ^ (layer0_outputs[1300]));
    assign outputs[4382] = layer0_outputs[1044];
    assign outputs[4383] = layer0_outputs[785];
    assign outputs[4384] = ~(layer0_outputs[1973]);
    assign outputs[4385] = layer0_outputs[4886];
    assign outputs[4386] = ~(layer0_outputs[2390]);
    assign outputs[4387] = layer0_outputs[3648];
    assign outputs[4388] = ~(layer0_outputs[2111]) | (layer0_outputs[3895]);
    assign outputs[4389] = ~(layer0_outputs[384]) | (layer0_outputs[2823]);
    assign outputs[4390] = ~(layer0_outputs[2357]) | (layer0_outputs[1506]);
    assign outputs[4391] = (layer0_outputs[1015]) & ~(layer0_outputs[558]);
    assign outputs[4392] = ~(layer0_outputs[3097]);
    assign outputs[4393] = (layer0_outputs[4501]) | (layer0_outputs[4653]);
    assign outputs[4394] = 1'b1;
    assign outputs[4395] = (layer0_outputs[2532]) & (layer0_outputs[3713]);
    assign outputs[4396] = layer0_outputs[2879];
    assign outputs[4397] = ~((layer0_outputs[946]) ^ (layer0_outputs[854]));
    assign outputs[4398] = ~(layer0_outputs[172]);
    assign outputs[4399] = layer0_outputs[235];
    assign outputs[4400] = ~(layer0_outputs[2304]);
    assign outputs[4401] = layer0_outputs[1881];
    assign outputs[4402] = (layer0_outputs[5086]) & (layer0_outputs[3730]);
    assign outputs[4403] = layer0_outputs[729];
    assign outputs[4404] = (layer0_outputs[3787]) ^ (layer0_outputs[326]);
    assign outputs[4405] = ~(layer0_outputs[4320]) | (layer0_outputs[3306]);
    assign outputs[4406] = layer0_outputs[4335];
    assign outputs[4407] = ~(layer0_outputs[4053]);
    assign outputs[4408] = layer0_outputs[2793];
    assign outputs[4409] = (layer0_outputs[2432]) & (layer0_outputs[3546]);
    assign outputs[4410] = ~(layer0_outputs[1034]);
    assign outputs[4411] = (layer0_outputs[472]) & ~(layer0_outputs[2461]);
    assign outputs[4412] = ~((layer0_outputs[1686]) & (layer0_outputs[688]));
    assign outputs[4413] = layer0_outputs[2424];
    assign outputs[4414] = layer0_outputs[86];
    assign outputs[4415] = (layer0_outputs[3331]) & ~(layer0_outputs[4191]);
    assign outputs[4416] = ~(layer0_outputs[2379]) | (layer0_outputs[1142]);
    assign outputs[4417] = (layer0_outputs[2623]) | (layer0_outputs[1952]);
    assign outputs[4418] = layer0_outputs[4187];
    assign outputs[4419] = (layer0_outputs[3044]) ^ (layer0_outputs[580]);
    assign outputs[4420] = ~(layer0_outputs[3282]) | (layer0_outputs[1975]);
    assign outputs[4421] = (layer0_outputs[4189]) & ~(layer0_outputs[3475]);
    assign outputs[4422] = layer0_outputs[105];
    assign outputs[4423] = layer0_outputs[3117];
    assign outputs[4424] = ~(layer0_outputs[1302]);
    assign outputs[4425] = ~((layer0_outputs[975]) ^ (layer0_outputs[1943]));
    assign outputs[4426] = layer0_outputs[1443];
    assign outputs[4427] = (layer0_outputs[1601]) ^ (layer0_outputs[3290]);
    assign outputs[4428] = ~((layer0_outputs[3919]) ^ (layer0_outputs[1475]));
    assign outputs[4429] = ~(layer0_outputs[2445]);
    assign outputs[4430] = (layer0_outputs[2236]) ^ (layer0_outputs[929]);
    assign outputs[4431] = (layer0_outputs[4863]) | (layer0_outputs[4668]);
    assign outputs[4432] = (layer0_outputs[4976]) & (layer0_outputs[2170]);
    assign outputs[4433] = ~(layer0_outputs[2930]);
    assign outputs[4434] = ~((layer0_outputs[2240]) & (layer0_outputs[935]));
    assign outputs[4435] = layer0_outputs[712];
    assign outputs[4436] = ~(layer0_outputs[3425]);
    assign outputs[4437] = (layer0_outputs[3346]) ^ (layer0_outputs[1243]);
    assign outputs[4438] = ~((layer0_outputs[2367]) ^ (layer0_outputs[448]));
    assign outputs[4439] = (layer0_outputs[490]) ^ (layer0_outputs[4363]);
    assign outputs[4440] = layer0_outputs[4353];
    assign outputs[4441] = ~(layer0_outputs[4035]);
    assign outputs[4442] = ~((layer0_outputs[3389]) & (layer0_outputs[1114]));
    assign outputs[4443] = (layer0_outputs[4376]) & ~(layer0_outputs[722]);
    assign outputs[4444] = ~(layer0_outputs[4940]);
    assign outputs[4445] = layer0_outputs[4113];
    assign outputs[4446] = ~(layer0_outputs[396]);
    assign outputs[4447] = ~(layer0_outputs[2319]);
    assign outputs[4448] = layer0_outputs[2992];
    assign outputs[4449] = ~(layer0_outputs[2565]) | (layer0_outputs[547]);
    assign outputs[4450] = ~((layer0_outputs[2037]) ^ (layer0_outputs[2490]));
    assign outputs[4451] = (layer0_outputs[4285]) ^ (layer0_outputs[3141]);
    assign outputs[4452] = (layer0_outputs[1612]) & ~(layer0_outputs[1286]);
    assign outputs[4453] = ~((layer0_outputs[1791]) ^ (layer0_outputs[880]));
    assign outputs[4454] = (layer0_outputs[1787]) & (layer0_outputs[3886]);
    assign outputs[4455] = ~(layer0_outputs[2928]);
    assign outputs[4456] = ~(layer0_outputs[3710]);
    assign outputs[4457] = (layer0_outputs[1825]) & ~(layer0_outputs[4288]);
    assign outputs[4458] = layer0_outputs[4429];
    assign outputs[4459] = layer0_outputs[3308];
    assign outputs[4460] = (layer0_outputs[4824]) & (layer0_outputs[1787]);
    assign outputs[4461] = ~(layer0_outputs[3472]);
    assign outputs[4462] = (layer0_outputs[1010]) & (layer0_outputs[1908]);
    assign outputs[4463] = layer0_outputs[3869];
    assign outputs[4464] = layer0_outputs[2362];
    assign outputs[4465] = layer0_outputs[828];
    assign outputs[4466] = ~(layer0_outputs[4996]);
    assign outputs[4467] = (layer0_outputs[1558]) ^ (layer0_outputs[4657]);
    assign outputs[4468] = (layer0_outputs[1968]) & (layer0_outputs[1251]);
    assign outputs[4469] = layer0_outputs[587];
    assign outputs[4470] = ~(layer0_outputs[309]) | (layer0_outputs[3772]);
    assign outputs[4471] = ~((layer0_outputs[3918]) ^ (layer0_outputs[2082]));
    assign outputs[4472] = ~(layer0_outputs[1687]) | (layer0_outputs[3157]);
    assign outputs[4473] = ~(layer0_outputs[1176]);
    assign outputs[4474] = (layer0_outputs[535]) ^ (layer0_outputs[2517]);
    assign outputs[4475] = ~((layer0_outputs[3683]) | (layer0_outputs[3257]));
    assign outputs[4476] = ~(layer0_outputs[3695]);
    assign outputs[4477] = layer0_outputs[609];
    assign outputs[4478] = ~(layer0_outputs[139]);
    assign outputs[4479] = layer0_outputs[3764];
    assign outputs[4480] = layer0_outputs[4805];
    assign outputs[4481] = ~((layer0_outputs[202]) | (layer0_outputs[1276]));
    assign outputs[4482] = layer0_outputs[578];
    assign outputs[4483] = ~(layer0_outputs[5044]) | (layer0_outputs[3478]);
    assign outputs[4484] = ~(layer0_outputs[5008]);
    assign outputs[4485] = ~(layer0_outputs[4213]);
    assign outputs[4486] = (layer0_outputs[4683]) & ~(layer0_outputs[3006]);
    assign outputs[4487] = (layer0_outputs[2006]) | (layer0_outputs[3115]);
    assign outputs[4488] = ~((layer0_outputs[1571]) ^ (layer0_outputs[1387]));
    assign outputs[4489] = layer0_outputs[3803];
    assign outputs[4490] = (layer0_outputs[985]) ^ (layer0_outputs[1721]);
    assign outputs[4491] = (layer0_outputs[2847]) & (layer0_outputs[601]);
    assign outputs[4492] = layer0_outputs[1970];
    assign outputs[4493] = (layer0_outputs[1205]) ^ (layer0_outputs[856]);
    assign outputs[4494] = ~(layer0_outputs[2158]);
    assign outputs[4495] = (layer0_outputs[4011]) ^ (layer0_outputs[1318]);
    assign outputs[4496] = ~(layer0_outputs[3763]) | (layer0_outputs[408]);
    assign outputs[4497] = layer0_outputs[1392];
    assign outputs[4498] = ~((layer0_outputs[850]) ^ (layer0_outputs[1976]));
    assign outputs[4499] = ~(layer0_outputs[2873]);
    assign outputs[4500] = ~(layer0_outputs[2192]) | (layer0_outputs[99]);
    assign outputs[4501] = ~(layer0_outputs[3370]);
    assign outputs[4502] = (layer0_outputs[1297]) & ~(layer0_outputs[4656]);
    assign outputs[4503] = (layer0_outputs[4545]) | (layer0_outputs[2493]);
    assign outputs[4504] = (layer0_outputs[4705]) | (layer0_outputs[1834]);
    assign outputs[4505] = (layer0_outputs[4732]) ^ (layer0_outputs[2280]);
    assign outputs[4506] = (layer0_outputs[2756]) | (layer0_outputs[3320]);
    assign outputs[4507] = (layer0_outputs[1746]) & (layer0_outputs[3380]);
    assign outputs[4508] = layer0_outputs[1639];
    assign outputs[4509] = (layer0_outputs[3308]) & ~(layer0_outputs[2902]);
    assign outputs[4510] = (layer0_outputs[4095]) | (layer0_outputs[1489]);
    assign outputs[4511] = ~(layer0_outputs[2164]);
    assign outputs[4512] = ~(layer0_outputs[1190]);
    assign outputs[4513] = (layer0_outputs[1681]) & (layer0_outputs[1431]);
    assign outputs[4514] = (layer0_outputs[5083]) & ~(layer0_outputs[3349]);
    assign outputs[4515] = ~(layer0_outputs[3376]);
    assign outputs[4516] = 1'b1;
    assign outputs[4517] = layer0_outputs[370];
    assign outputs[4518] = ~((layer0_outputs[4437]) ^ (layer0_outputs[4744]));
    assign outputs[4519] = layer0_outputs[3260];
    assign outputs[4520] = ~((layer0_outputs[4904]) ^ (layer0_outputs[484]));
    assign outputs[4521] = ~(layer0_outputs[1903]);
    assign outputs[4522] = ~(layer0_outputs[4136]);
    assign outputs[4523] = (layer0_outputs[2182]) | (layer0_outputs[3486]);
    assign outputs[4524] = ~((layer0_outputs[4596]) | (layer0_outputs[1446]));
    assign outputs[4525] = ~(layer0_outputs[470]);
    assign outputs[4526] = ~(layer0_outputs[2643]);
    assign outputs[4527] = ~((layer0_outputs[2467]) & (layer0_outputs[555]));
    assign outputs[4528] = (layer0_outputs[3509]) ^ (layer0_outputs[3913]);
    assign outputs[4529] = layer0_outputs[2353];
    assign outputs[4530] = ~(layer0_outputs[2643]);
    assign outputs[4531] = layer0_outputs[3144];
    assign outputs[4532] = (layer0_outputs[2195]) & (layer0_outputs[1239]);
    assign outputs[4533] = layer0_outputs[3737];
    assign outputs[4534] = ~((layer0_outputs[718]) ^ (layer0_outputs[816]));
    assign outputs[4535] = ~(layer0_outputs[4573]);
    assign outputs[4536] = ~((layer0_outputs[3546]) ^ (layer0_outputs[3933]));
    assign outputs[4537] = (layer0_outputs[4669]) ^ (layer0_outputs[1656]);
    assign outputs[4538] = layer0_outputs[3391];
    assign outputs[4539] = ~(layer0_outputs[2563]);
    assign outputs[4540] = (layer0_outputs[3252]) & (layer0_outputs[4554]);
    assign outputs[4541] = ~((layer0_outputs[1492]) ^ (layer0_outputs[697]));
    assign outputs[4542] = ~((layer0_outputs[1669]) ^ (layer0_outputs[4545]));
    assign outputs[4543] = ~(layer0_outputs[559]);
    assign outputs[4544] = ~(layer0_outputs[4945]) | (layer0_outputs[4808]);
    assign outputs[4545] = ~(layer0_outputs[1757]);
    assign outputs[4546] = (layer0_outputs[2736]) & ~(layer0_outputs[4597]);
    assign outputs[4547] = ~((layer0_outputs[1562]) | (layer0_outputs[722]));
    assign outputs[4548] = layer0_outputs[3605];
    assign outputs[4549] = (layer0_outputs[971]) & ~(layer0_outputs[3862]);
    assign outputs[4550] = ~((layer0_outputs[1080]) ^ (layer0_outputs[1045]));
    assign outputs[4551] = ~((layer0_outputs[2914]) ^ (layer0_outputs[2949]));
    assign outputs[4552] = ~((layer0_outputs[3520]) ^ (layer0_outputs[643]));
    assign outputs[4553] = layer0_outputs[2317];
    assign outputs[4554] = (layer0_outputs[4085]) & (layer0_outputs[2394]);
    assign outputs[4555] = layer0_outputs[1077];
    assign outputs[4556] = ~((layer0_outputs[4504]) & (layer0_outputs[2337]));
    assign outputs[4557] = ~((layer0_outputs[2042]) ^ (layer0_outputs[2803]));
    assign outputs[4558] = ~((layer0_outputs[3474]) ^ (layer0_outputs[4093]));
    assign outputs[4559] = layer0_outputs[1212];
    assign outputs[4560] = ~(layer0_outputs[4892]) | (layer0_outputs[4948]);
    assign outputs[4561] = ~(layer0_outputs[193]);
    assign outputs[4562] = ~(layer0_outputs[2564]);
    assign outputs[4563] = (layer0_outputs[1456]) ^ (layer0_outputs[1317]);
    assign outputs[4564] = (layer0_outputs[517]) ^ (layer0_outputs[3525]);
    assign outputs[4565] = layer0_outputs[5034];
    assign outputs[4566] = layer0_outputs[2597];
    assign outputs[4567] = (layer0_outputs[525]) & ~(layer0_outputs[5021]);
    assign outputs[4568] = ~(layer0_outputs[1487]) | (layer0_outputs[739]);
    assign outputs[4569] = ~(layer0_outputs[3212]);
    assign outputs[4570] = ~(layer0_outputs[3584]);
    assign outputs[4571] = (layer0_outputs[2033]) & ~(layer0_outputs[320]);
    assign outputs[4572] = layer0_outputs[2974];
    assign outputs[4573] = ~(layer0_outputs[4435]);
    assign outputs[4574] = ~(layer0_outputs[104]) | (layer0_outputs[2545]);
    assign outputs[4575] = ~((layer0_outputs[2705]) ^ (layer0_outputs[5102]));
    assign outputs[4576] = ~((layer0_outputs[272]) ^ (layer0_outputs[2859]));
    assign outputs[4577] = (layer0_outputs[211]) ^ (layer0_outputs[1415]);
    assign outputs[4578] = layer0_outputs[1694];
    assign outputs[4579] = (layer0_outputs[4843]) & ~(layer0_outputs[4087]);
    assign outputs[4580] = (layer0_outputs[1383]) | (layer0_outputs[321]);
    assign outputs[4581] = ~((layer0_outputs[3318]) & (layer0_outputs[118]));
    assign outputs[4582] = layer0_outputs[3942];
    assign outputs[4583] = ~(layer0_outputs[1830]);
    assign outputs[4584] = (layer0_outputs[2416]) | (layer0_outputs[3881]);
    assign outputs[4585] = (layer0_outputs[4009]) ^ (layer0_outputs[792]);
    assign outputs[4586] = ~(layer0_outputs[314]);
    assign outputs[4587] = layer0_outputs[4319];
    assign outputs[4588] = ~(layer0_outputs[3615]);
    assign outputs[4589] = (layer0_outputs[2252]) ^ (layer0_outputs[3522]);
    assign outputs[4590] = layer0_outputs[3708];
    assign outputs[4591] = layer0_outputs[1223];
    assign outputs[4592] = layer0_outputs[2502];
    assign outputs[4593] = ~(layer0_outputs[4765]);
    assign outputs[4594] = ~(layer0_outputs[1072]);
    assign outputs[4595] = ~(layer0_outputs[606]);
    assign outputs[4596] = ~(layer0_outputs[373]);
    assign outputs[4597] = ~(layer0_outputs[4367]);
    assign outputs[4598] = ~(layer0_outputs[3397]) | (layer0_outputs[2375]);
    assign outputs[4599] = ~(layer0_outputs[2971]);
    assign outputs[4600] = (layer0_outputs[5077]) | (layer0_outputs[3302]);
    assign outputs[4601] = (layer0_outputs[1163]) & (layer0_outputs[2809]);
    assign outputs[4602] = ~(layer0_outputs[433]);
    assign outputs[4603] = ~(layer0_outputs[4047]);
    assign outputs[4604] = ~(layer0_outputs[4183]);
    assign outputs[4605] = ~((layer0_outputs[1057]) & (layer0_outputs[3025]));
    assign outputs[4606] = ~(layer0_outputs[647]);
    assign outputs[4607] = layer0_outputs[2612];
    assign outputs[4608] = ~((layer0_outputs[4143]) ^ (layer0_outputs[969]));
    assign outputs[4609] = (layer0_outputs[3524]) ^ (layer0_outputs[1906]);
    assign outputs[4610] = (layer0_outputs[1506]) ^ (layer0_outputs[2062]);
    assign outputs[4611] = (layer0_outputs[3975]) & (layer0_outputs[4516]);
    assign outputs[4612] = ~(layer0_outputs[1675]) | (layer0_outputs[1944]);
    assign outputs[4613] = (layer0_outputs[3001]) & (layer0_outputs[1325]);
    assign outputs[4614] = (layer0_outputs[4417]) ^ (layer0_outputs[4859]);
    assign outputs[4615] = ~((layer0_outputs[446]) ^ (layer0_outputs[3543]));
    assign outputs[4616] = ~(layer0_outputs[2615]);
    assign outputs[4617] = layer0_outputs[4195];
    assign outputs[4618] = ~((layer0_outputs[1616]) ^ (layer0_outputs[4439]));
    assign outputs[4619] = (layer0_outputs[288]) & ~(layer0_outputs[3447]);
    assign outputs[4620] = ~((layer0_outputs[5056]) ^ (layer0_outputs[4562]));
    assign outputs[4621] = ~((layer0_outputs[749]) & (layer0_outputs[4340]));
    assign outputs[4622] = (layer0_outputs[539]) & ~(layer0_outputs[871]);
    assign outputs[4623] = (layer0_outputs[3582]) ^ (layer0_outputs[2837]);
    assign outputs[4624] = (layer0_outputs[922]) & ~(layer0_outputs[1292]);
    assign outputs[4625] = ~(layer0_outputs[257]) | (layer0_outputs[2301]);
    assign outputs[4626] = layer0_outputs[1849];
    assign outputs[4627] = ~(layer0_outputs[3479]);
    assign outputs[4628] = (layer0_outputs[3092]) & ~(layer0_outputs[1043]);
    assign outputs[4629] = 1'b0;
    assign outputs[4630] = ~((layer0_outputs[1835]) ^ (layer0_outputs[339]));
    assign outputs[4631] = layer0_outputs[2117];
    assign outputs[4632] = ~((layer0_outputs[308]) | (layer0_outputs[334]));
    assign outputs[4633] = ~((layer0_outputs[2449]) ^ (layer0_outputs[605]));
    assign outputs[4634] = (layer0_outputs[1878]) & ~(layer0_outputs[1036]);
    assign outputs[4635] = (layer0_outputs[4411]) & ~(layer0_outputs[343]);
    assign outputs[4636] = (layer0_outputs[5047]) ^ (layer0_outputs[222]);
    assign outputs[4637] = ~(layer0_outputs[2465]);
    assign outputs[4638] = (layer0_outputs[4160]) & ~(layer0_outputs[2350]);
    assign outputs[4639] = layer0_outputs[2501];
    assign outputs[4640] = ~((layer0_outputs[3374]) ^ (layer0_outputs[1220]));
    assign outputs[4641] = ~(layer0_outputs[765]);
    assign outputs[4642] = (layer0_outputs[4016]) & ~(layer0_outputs[1487]);
    assign outputs[4643] = ~(layer0_outputs[4975]);
    assign outputs[4644] = layer0_outputs[413];
    assign outputs[4645] = layer0_outputs[1722];
    assign outputs[4646] = layer0_outputs[4079];
    assign outputs[4647] = ~((layer0_outputs[1280]) | (layer0_outputs[4144]));
    assign outputs[4648] = ~(layer0_outputs[848]);
    assign outputs[4649] = (layer0_outputs[2954]) & ~(layer0_outputs[2002]);
    assign outputs[4650] = ~(layer0_outputs[78]);
    assign outputs[4651] = ~(layer0_outputs[604]);
    assign outputs[4652] = ~((layer0_outputs[1046]) | (layer0_outputs[426]));
    assign outputs[4653] = (layer0_outputs[740]) | (layer0_outputs[1299]);
    assign outputs[4654] = (layer0_outputs[2177]) ^ (layer0_outputs[110]);
    assign outputs[4655] = (layer0_outputs[1559]) & ~(layer0_outputs[4992]);
    assign outputs[4656] = layer0_outputs[3193];
    assign outputs[4657] = (layer0_outputs[4495]) & (layer0_outputs[3768]);
    assign outputs[4658] = ~((layer0_outputs[197]) | (layer0_outputs[910]));
    assign outputs[4659] = layer0_outputs[4837];
    assign outputs[4660] = ~(layer0_outputs[2868]);
    assign outputs[4661] = (layer0_outputs[231]) & ~(layer0_outputs[2645]);
    assign outputs[4662] = (layer0_outputs[192]) ^ (layer0_outputs[2791]);
    assign outputs[4663] = (layer0_outputs[3963]) & ~(layer0_outputs[3944]);
    assign outputs[4664] = ~((layer0_outputs[2383]) ^ (layer0_outputs[3422]));
    assign outputs[4665] = (layer0_outputs[3646]) & (layer0_outputs[4620]);
    assign outputs[4666] = (layer0_outputs[3241]) ^ (layer0_outputs[3421]);
    assign outputs[4667] = (layer0_outputs[641]) | (layer0_outputs[2965]);
    assign outputs[4668] = (layer0_outputs[1374]) & ~(layer0_outputs[595]);
    assign outputs[4669] = layer0_outputs[581];
    assign outputs[4670] = ~((layer0_outputs[124]) | (layer0_outputs[3426]));
    assign outputs[4671] = ~(layer0_outputs[3463]) | (layer0_outputs[803]);
    assign outputs[4672] = ~(layer0_outputs[4058]);
    assign outputs[4673] = ~(layer0_outputs[2125]);
    assign outputs[4674] = ~(layer0_outputs[1495]) | (layer0_outputs[2262]);
    assign outputs[4675] = (layer0_outputs[4712]) | (layer0_outputs[4704]);
    assign outputs[4676] = (layer0_outputs[4401]) & ~(layer0_outputs[4011]);
    assign outputs[4677] = (layer0_outputs[5078]) ^ (layer0_outputs[4938]);
    assign outputs[4678] = layer0_outputs[352];
    assign outputs[4679] = ~(layer0_outputs[4013]);
    assign outputs[4680] = (layer0_outputs[2989]) & ~(layer0_outputs[3565]);
    assign outputs[4681] = ~((layer0_outputs[3018]) ^ (layer0_outputs[1130]));
    assign outputs[4682] = (layer0_outputs[379]) & ~(layer0_outputs[3865]);
    assign outputs[4683] = ~(layer0_outputs[1281]);
    assign outputs[4684] = ~(layer0_outputs[2850]) | (layer0_outputs[2642]);
    assign outputs[4685] = (layer0_outputs[342]) ^ (layer0_outputs[143]);
    assign outputs[4686] = (layer0_outputs[330]) & ~(layer0_outputs[3227]);
    assign outputs[4687] = layer0_outputs[3683];
    assign outputs[4688] = 1'b1;
    assign outputs[4689] = (layer0_outputs[2393]) & (layer0_outputs[4164]);
    assign outputs[4690] = ~(layer0_outputs[2082]);
    assign outputs[4691] = (layer0_outputs[3362]) ^ (layer0_outputs[3099]);
    assign outputs[4692] = (layer0_outputs[3657]) ^ (layer0_outputs[2387]);
    assign outputs[4693] = (layer0_outputs[4171]) & (layer0_outputs[3714]);
    assign outputs[4694] = ~(layer0_outputs[3954]);
    assign outputs[4695] = (layer0_outputs[2241]) & ~(layer0_outputs[3142]);
    assign outputs[4696] = ~((layer0_outputs[1493]) | (layer0_outputs[1820]));
    assign outputs[4697] = (layer0_outputs[2724]) & ~(layer0_outputs[1252]);
    assign outputs[4698] = ~(layer0_outputs[3677]);
    assign outputs[4699] = ~(layer0_outputs[4369]);
    assign outputs[4700] = (layer0_outputs[1754]) ^ (layer0_outputs[1568]);
    assign outputs[4701] = layer0_outputs[3396];
    assign outputs[4702] = ~(layer0_outputs[4530]);
    assign outputs[4703] = ~(layer0_outputs[4078]);
    assign outputs[4704] = layer0_outputs[1867];
    assign outputs[4705] = (layer0_outputs[623]) ^ (layer0_outputs[3710]);
    assign outputs[4706] = (layer0_outputs[845]) & ~(layer0_outputs[5111]);
    assign outputs[4707] = ~((layer0_outputs[1084]) | (layer0_outputs[4706]));
    assign outputs[4708] = ~((layer0_outputs[1503]) | (layer0_outputs[1080]));
    assign outputs[4709] = ~(layer0_outputs[1042]);
    assign outputs[4710] = layer0_outputs[1363];
    assign outputs[4711] = (layer0_outputs[2774]) & ~(layer0_outputs[1140]);
    assign outputs[4712] = (layer0_outputs[4689]) & ~(layer0_outputs[3589]);
    assign outputs[4713] = layer0_outputs[3433];
    assign outputs[4714] = layer0_outputs[2052];
    assign outputs[4715] = ~(layer0_outputs[371]);
    assign outputs[4716] = layer0_outputs[169];
    assign outputs[4717] = layer0_outputs[3593];
    assign outputs[4718] = (layer0_outputs[928]) & (layer0_outputs[3694]);
    assign outputs[4719] = layer0_outputs[4413];
    assign outputs[4720] = layer0_outputs[2012];
    assign outputs[4721] = layer0_outputs[121];
    assign outputs[4722] = (layer0_outputs[1739]) & ~(layer0_outputs[2692]);
    assign outputs[4723] = ~((layer0_outputs[2481]) ^ (layer0_outputs[3223]));
    assign outputs[4724] = (layer0_outputs[5106]) & (layer0_outputs[5043]);
    assign outputs[4725] = layer0_outputs[2907];
    assign outputs[4726] = (layer0_outputs[3870]) & ~(layer0_outputs[2500]);
    assign outputs[4727] = (layer0_outputs[3570]) & ~(layer0_outputs[4502]);
    assign outputs[4728] = (layer0_outputs[1045]) ^ (layer0_outputs[2759]);
    assign outputs[4729] = layer0_outputs[468];
    assign outputs[4730] = ~(layer0_outputs[998]);
    assign outputs[4731] = (layer0_outputs[82]) & ~(layer0_outputs[4663]);
    assign outputs[4732] = (layer0_outputs[3735]) ^ (layer0_outputs[3230]);
    assign outputs[4733] = (layer0_outputs[4819]) ^ (layer0_outputs[4114]);
    assign outputs[4734] = (layer0_outputs[3827]) ^ (layer0_outputs[4910]);
    assign outputs[4735] = (layer0_outputs[1382]) & ~(layer0_outputs[3717]);
    assign outputs[4736] = layer0_outputs[4247];
    assign outputs[4737] = ~(layer0_outputs[2078]);
    assign outputs[4738] = (layer0_outputs[4979]) & ~(layer0_outputs[4833]);
    assign outputs[4739] = (layer0_outputs[916]) & ~(layer0_outputs[1576]);
    assign outputs[4740] = ~((layer0_outputs[2410]) | (layer0_outputs[1050]));
    assign outputs[4741] = ~(layer0_outputs[3937]) | (layer0_outputs[2961]);
    assign outputs[4742] = (layer0_outputs[1918]) & ~(layer0_outputs[3210]);
    assign outputs[4743] = layer0_outputs[3028];
    assign outputs[4744] = layer0_outputs[52];
    assign outputs[4745] = ~(layer0_outputs[4008]);
    assign outputs[4746] = (layer0_outputs[1989]) ^ (layer0_outputs[260]);
    assign outputs[4747] = layer0_outputs[1152];
    assign outputs[4748] = (layer0_outputs[5101]) & ~(layer0_outputs[1223]);
    assign outputs[4749] = ~(layer0_outputs[4059]);
    assign outputs[4750] = ~((layer0_outputs[1087]) | (layer0_outputs[4348]));
    assign outputs[4751] = (layer0_outputs[3650]) ^ (layer0_outputs[3338]);
    assign outputs[4752] = (layer0_outputs[1827]) ^ (layer0_outputs[4046]);
    assign outputs[4753] = (layer0_outputs[536]) & (layer0_outputs[223]);
    assign outputs[4754] = (layer0_outputs[4172]) & ~(layer0_outputs[3903]);
    assign outputs[4755] = (layer0_outputs[4812]) ^ (layer0_outputs[633]);
    assign outputs[4756] = ~((layer0_outputs[4510]) | (layer0_outputs[3326]));
    assign outputs[4757] = ~(layer0_outputs[4786]);
    assign outputs[4758] = ~(layer0_outputs[1850]);
    assign outputs[4759] = layer0_outputs[1234];
    assign outputs[4760] = ~((layer0_outputs[1383]) ^ (layer0_outputs[1238]));
    assign outputs[4761] = ~((layer0_outputs[1954]) & (layer0_outputs[4163]));
    assign outputs[4762] = (layer0_outputs[2570]) ^ (layer0_outputs[3814]);
    assign outputs[4763] = layer0_outputs[3037];
    assign outputs[4764] = layer0_outputs[2016];
    assign outputs[4765] = ~((layer0_outputs[3833]) ^ (layer0_outputs[3675]));
    assign outputs[4766] = layer0_outputs[314];
    assign outputs[4767] = (layer0_outputs[3244]) ^ (layer0_outputs[1877]);
    assign outputs[4768] = ~((layer0_outputs[2962]) ^ (layer0_outputs[1773]));
    assign outputs[4769] = (layer0_outputs[1862]) | (layer0_outputs[1848]);
    assign outputs[4770] = ~((layer0_outputs[2160]) | (layer0_outputs[199]));
    assign outputs[4771] = ~(layer0_outputs[2066]);
    assign outputs[4772] = (layer0_outputs[1117]) & ~(layer0_outputs[1466]);
    assign outputs[4773] = (layer0_outputs[1853]) ^ (layer0_outputs[1074]);
    assign outputs[4774] = layer0_outputs[4002];
    assign outputs[4775] = ~((layer0_outputs[4711]) ^ (layer0_outputs[3759]));
    assign outputs[4776] = layer0_outputs[5045];
    assign outputs[4777] = (layer0_outputs[1722]) & ~(layer0_outputs[4486]);
    assign outputs[4778] = layer0_outputs[1563];
    assign outputs[4779] = (layer0_outputs[1187]) & ~(layer0_outputs[170]);
    assign outputs[4780] = ~(layer0_outputs[4916]);
    assign outputs[4781] = ~((layer0_outputs[4175]) | (layer0_outputs[2064]));
    assign outputs[4782] = layer0_outputs[851];
    assign outputs[4783] = layer0_outputs[3274];
    assign outputs[4784] = ~((layer0_outputs[1949]) ^ (layer0_outputs[1137]));
    assign outputs[4785] = layer0_outputs[3105];
    assign outputs[4786] = ~(layer0_outputs[921]) | (layer0_outputs[1635]);
    assign outputs[4787] = layer0_outputs[962];
    assign outputs[4788] = layer0_outputs[3777];
    assign outputs[4789] = ~(layer0_outputs[2348]);
    assign outputs[4790] = ~(layer0_outputs[1952]);
    assign outputs[4791] = ~((layer0_outputs[3229]) ^ (layer0_outputs[3367]));
    assign outputs[4792] = ~(layer0_outputs[3163]);
    assign outputs[4793] = ~(layer0_outputs[3516]);
    assign outputs[4794] = ~(layer0_outputs[2099]) | (layer0_outputs[237]);
    assign outputs[4795] = ~(layer0_outputs[1046]);
    assign outputs[4796] = ~(layer0_outputs[246]);
    assign outputs[4797] = layer0_outputs[1946];
    assign outputs[4798] = layer0_outputs[1368];
    assign outputs[4799] = ~(layer0_outputs[4328]);
    assign outputs[4800] = ~(layer0_outputs[3902]);
    assign outputs[4801] = (layer0_outputs[1739]) & ~(layer0_outputs[6]);
    assign outputs[4802] = layer0_outputs[3950];
    assign outputs[4803] = ~((layer0_outputs[3712]) & (layer0_outputs[3551]));
    assign outputs[4804] = ~((layer0_outputs[4399]) ^ (layer0_outputs[4711]));
    assign outputs[4805] = (layer0_outputs[731]) | (layer0_outputs[3015]);
    assign outputs[4806] = layer0_outputs[4307];
    assign outputs[4807] = (layer0_outputs[1371]) & (layer0_outputs[2135]);
    assign outputs[4808] = layer0_outputs[4298];
    assign outputs[4809] = (layer0_outputs[2829]) & (layer0_outputs[1717]);
    assign outputs[4810] = layer0_outputs[4913];
    assign outputs[4811] = (layer0_outputs[4356]) & ~(layer0_outputs[822]);
    assign outputs[4812] = ~((layer0_outputs[2555]) | (layer0_outputs[1147]));
    assign outputs[4813] = (layer0_outputs[2010]) | (layer0_outputs[3004]);
    assign outputs[4814] = ~((layer0_outputs[527]) | (layer0_outputs[2833]));
    assign outputs[4815] = (layer0_outputs[4727]) & ~(layer0_outputs[770]);
    assign outputs[4816] = layer0_outputs[1548];
    assign outputs[4817] = ~(layer0_outputs[3375]) | (layer0_outputs[2858]);
    assign outputs[4818] = ~((layer0_outputs[1444]) | (layer0_outputs[2795]));
    assign outputs[4819] = layer0_outputs[115];
    assign outputs[4820] = layer0_outputs[2665];
    assign outputs[4821] = ~(layer0_outputs[3774]);
    assign outputs[4822] = layer0_outputs[1358];
    assign outputs[4823] = (layer0_outputs[3678]) ^ (layer0_outputs[3821]);
    assign outputs[4824] = (layer0_outputs[2787]) & (layer0_outputs[2589]);
    assign outputs[4825] = ~(layer0_outputs[3548]);
    assign outputs[4826] = layer0_outputs[2205];
    assign outputs[4827] = (layer0_outputs[721]) & (layer0_outputs[1980]);
    assign outputs[4828] = layer0_outputs[4367];
    assign outputs[4829] = (layer0_outputs[2701]) & (layer0_outputs[684]);
    assign outputs[4830] = layer0_outputs[3124];
    assign outputs[4831] = (layer0_outputs[768]) & ~(layer0_outputs[978]);
    assign outputs[4832] = layer0_outputs[3255];
    assign outputs[4833] = layer0_outputs[154];
    assign outputs[4834] = ~(layer0_outputs[3614]);
    assign outputs[4835] = (layer0_outputs[1149]) ^ (layer0_outputs[2876]);
    assign outputs[4836] = (layer0_outputs[1882]) & ~(layer0_outputs[799]);
    assign outputs[4837] = (layer0_outputs[3024]) & ~(layer0_outputs[4419]);
    assign outputs[4838] = layer0_outputs[4607];
    assign outputs[4839] = (layer0_outputs[1225]) & (layer0_outputs[166]);
    assign outputs[4840] = layer0_outputs[695];
    assign outputs[4841] = (layer0_outputs[1991]) & ~(layer0_outputs[3479]);
    assign outputs[4842] = ~(layer0_outputs[2849]);
    assign outputs[4843] = ~((layer0_outputs[2965]) | (layer0_outputs[2843]));
    assign outputs[4844] = ~((layer0_outputs[568]) | (layer0_outputs[562]));
    assign outputs[4845] = ~(layer0_outputs[4922]);
    assign outputs[4846] = (layer0_outputs[5019]) ^ (layer0_outputs[1763]);
    assign outputs[4847] = layer0_outputs[3582];
    assign outputs[4848] = (layer0_outputs[1943]) & ~(layer0_outputs[996]);
    assign outputs[4849] = (layer0_outputs[1556]) ^ (layer0_outputs[3586]);
    assign outputs[4850] = layer0_outputs[2653];
    assign outputs[4851] = ~(layer0_outputs[4572]);
    assign outputs[4852] = (layer0_outputs[3453]) & ~(layer0_outputs[538]);
    assign outputs[4853] = ~((layer0_outputs[426]) ^ (layer0_outputs[2947]));
    assign outputs[4854] = (layer0_outputs[57]) ^ (layer0_outputs[2103]);
    assign outputs[4855] = ~(layer0_outputs[8]);
    assign outputs[4856] = (layer0_outputs[4045]) & ~(layer0_outputs[1592]);
    assign outputs[4857] = (layer0_outputs[4852]) & (layer0_outputs[5075]);
    assign outputs[4858] = ~(layer0_outputs[146]);
    assign outputs[4859] = ~(layer0_outputs[3497]);
    assign outputs[4860] = (layer0_outputs[909]) & (layer0_outputs[1913]);
    assign outputs[4861] = ~(layer0_outputs[813]);
    assign outputs[4862] = (layer0_outputs[2454]) & (layer0_outputs[2852]);
    assign outputs[4863] = (layer0_outputs[1083]) & ~(layer0_outputs[2422]);
    assign outputs[4864] = (layer0_outputs[4074]) & (layer0_outputs[3470]);
    assign outputs[4865] = ~(layer0_outputs[4551]);
    assign outputs[4866] = ~((layer0_outputs[4973]) ^ (layer0_outputs[1540]));
    assign outputs[4867] = layer0_outputs[3751];
    assign outputs[4868] = layer0_outputs[4409];
    assign outputs[4869] = ~((layer0_outputs[1618]) | (layer0_outputs[3747]));
    assign outputs[4870] = ~((layer0_outputs[4691]) ^ (layer0_outputs[3542]));
    assign outputs[4871] = (layer0_outputs[2253]) & ~(layer0_outputs[3556]);
    assign outputs[4872] = (layer0_outputs[1553]) & ~(layer0_outputs[408]);
    assign outputs[4873] = (layer0_outputs[2631]) & (layer0_outputs[2746]);
    assign outputs[4874] = (layer0_outputs[1723]) ^ (layer0_outputs[1270]);
    assign outputs[4875] = ~((layer0_outputs[952]) | (layer0_outputs[1874]));
    assign outputs[4876] = (layer0_outputs[771]) & ~(layer0_outputs[1200]);
    assign outputs[4877] = (layer0_outputs[2704]) ^ (layer0_outputs[3151]);
    assign outputs[4878] = ~((layer0_outputs[3996]) | (layer0_outputs[490]));
    assign outputs[4879] = (layer0_outputs[1620]) ^ (layer0_outputs[4664]);
    assign outputs[4880] = ~(layer0_outputs[657]);
    assign outputs[4881] = (layer0_outputs[318]) & ~(layer0_outputs[1194]);
    assign outputs[4882] = layer0_outputs[2251];
    assign outputs[4883] = (layer0_outputs[620]) ^ (layer0_outputs[1250]);
    assign outputs[4884] = layer0_outputs[1656];
    assign outputs[4885] = (layer0_outputs[3204]) | (layer0_outputs[5080]);
    assign outputs[4886] = (layer0_outputs[1543]) & (layer0_outputs[2159]);
    assign outputs[4887] = (layer0_outputs[2511]) & (layer0_outputs[845]);
    assign outputs[4888] = (layer0_outputs[5013]) | (layer0_outputs[3836]);
    assign outputs[4889] = ~((layer0_outputs[1112]) | (layer0_outputs[28]));
    assign outputs[4890] = ~(layer0_outputs[1699]);
    assign outputs[4891] = layer0_outputs[3033];
    assign outputs[4892] = layer0_outputs[4943];
    assign outputs[4893] = ~((layer0_outputs[3991]) | (layer0_outputs[571]));
    assign outputs[4894] = layer0_outputs[3037];
    assign outputs[4895] = ~((layer0_outputs[145]) ^ (layer0_outputs[1312]));
    assign outputs[4896] = ~(layer0_outputs[1356]) | (layer0_outputs[3664]);
    assign outputs[4897] = (layer0_outputs[4273]) & ~(layer0_outputs[2760]);
    assign outputs[4898] = (layer0_outputs[1278]) ^ (layer0_outputs[2981]);
    assign outputs[4899] = ~(layer0_outputs[1307]) | (layer0_outputs[4881]);
    assign outputs[4900] = (layer0_outputs[1570]) & (layer0_outputs[1871]);
    assign outputs[4901] = (layer0_outputs[1088]) & (layer0_outputs[1306]);
    assign outputs[4902] = ~(layer0_outputs[4929]);
    assign outputs[4903] = (layer0_outputs[3743]) ^ (layer0_outputs[1856]);
    assign outputs[4904] = layer0_outputs[1884];
    assign outputs[4905] = (layer0_outputs[4658]) & (layer0_outputs[3865]);
    assign outputs[4906] = layer0_outputs[1865];
    assign outputs[4907] = (layer0_outputs[3416]) & ~(layer0_outputs[927]);
    assign outputs[4908] = ~(layer0_outputs[806]);
    assign outputs[4909] = ~(layer0_outputs[269]);
    assign outputs[4910] = (layer0_outputs[1256]) ^ (layer0_outputs[4920]);
    assign outputs[4911] = layer0_outputs[930];
    assign outputs[4912] = layer0_outputs[1230];
    assign outputs[4913] = ~((layer0_outputs[4065]) | (layer0_outputs[1537]));
    assign outputs[4914] = (layer0_outputs[2935]) ^ (layer0_outputs[3736]);
    assign outputs[4915] = ~(layer0_outputs[4856]) | (layer0_outputs[2583]);
    assign outputs[4916] = ~(layer0_outputs[2300]);
    assign outputs[4917] = ~(layer0_outputs[3987]);
    assign outputs[4918] = (layer0_outputs[2872]) & ~(layer0_outputs[4538]);
    assign outputs[4919] = layer0_outputs[189];
    assign outputs[4920] = (layer0_outputs[4162]) ^ (layer0_outputs[4661]);
    assign outputs[4921] = ~(layer0_outputs[3406]);
    assign outputs[4922] = ~(layer0_outputs[2050]);
    assign outputs[4923] = layer0_outputs[2420];
    assign outputs[4924] = layer0_outputs[4803];
    assign outputs[4925] = ~(layer0_outputs[719]) | (layer0_outputs[4690]);
    assign outputs[4926] = ~(layer0_outputs[3567]);
    assign outputs[4927] = (layer0_outputs[1393]) & (layer0_outputs[23]);
    assign outputs[4928] = (layer0_outputs[916]) & (layer0_outputs[5062]);
    assign outputs[4929] = layer0_outputs[3050];
    assign outputs[4930] = ~((layer0_outputs[2942]) | (layer0_outputs[1039]));
    assign outputs[4931] = ~((layer0_outputs[3243]) & (layer0_outputs[1350]));
    assign outputs[4932] = ~(layer0_outputs[4517]);
    assign outputs[4933] = ~((layer0_outputs[2990]) & (layer0_outputs[4974]));
    assign outputs[4934] = ~((layer0_outputs[2888]) | (layer0_outputs[3911]));
    assign outputs[4935] = ~((layer0_outputs[4389]) ^ (layer0_outputs[2611]));
    assign outputs[4936] = ~(layer0_outputs[1158]);
    assign outputs[4937] = ~(layer0_outputs[919]);
    assign outputs[4938] = (layer0_outputs[1732]) ^ (layer0_outputs[190]);
    assign outputs[4939] = layer0_outputs[4560];
    assign outputs[4940] = ~((layer0_outputs[2250]) | (layer0_outputs[972]));
    assign outputs[4941] = ~(layer0_outputs[3328]);
    assign outputs[4942] = (layer0_outputs[5016]) & (layer0_outputs[2351]);
    assign outputs[4943] = (layer0_outputs[1950]) & ~(layer0_outputs[3347]);
    assign outputs[4944] = ~((layer0_outputs[1486]) | (layer0_outputs[3531]));
    assign outputs[4945] = layer0_outputs[1883];
    assign outputs[4946] = ~((layer0_outputs[3900]) & (layer0_outputs[2278]));
    assign outputs[4947] = ~((layer0_outputs[4088]) & (layer0_outputs[2953]));
    assign outputs[4948] = layer0_outputs[1987];
    assign outputs[4949] = layer0_outputs[31];
    assign outputs[4950] = (layer0_outputs[5082]) & (layer0_outputs[1673]);
    assign outputs[4951] = layer0_outputs[51];
    assign outputs[4952] = ~(layer0_outputs[4365]);
    assign outputs[4953] = (layer0_outputs[2811]) & ~(layer0_outputs[3885]);
    assign outputs[4954] = ~(layer0_outputs[819]);
    assign outputs[4955] = (layer0_outputs[1674]) ^ (layer0_outputs[682]);
    assign outputs[4956] = ~((layer0_outputs[3954]) | (layer0_outputs[1807]));
    assign outputs[4957] = (layer0_outputs[3853]) ^ (layer0_outputs[3986]);
    assign outputs[4958] = ~(layer0_outputs[2310]);
    assign outputs[4959] = ~(layer0_outputs[3062]);
    assign outputs[4960] = (layer0_outputs[847]) ^ (layer0_outputs[132]);
    assign outputs[4961] = ~((layer0_outputs[3969]) ^ (layer0_outputs[740]));
    assign outputs[4962] = layer0_outputs[4355];
    assign outputs[4963] = layer0_outputs[1674];
    assign outputs[4964] = ~(layer0_outputs[2801]);
    assign outputs[4965] = layer0_outputs[3050];
    assign outputs[4966] = (layer0_outputs[234]) & ~(layer0_outputs[1734]);
    assign outputs[4967] = ~((layer0_outputs[1696]) | (layer0_outputs[547]));
    assign outputs[4968] = layer0_outputs[4722];
    assign outputs[4969] = layer0_outputs[877];
    assign outputs[4970] = (layer0_outputs[1263]) & ~(layer0_outputs[2476]);
    assign outputs[4971] = (layer0_outputs[2077]) ^ (layer0_outputs[4070]);
    assign outputs[4972] = layer0_outputs[4505];
    assign outputs[4973] = layer0_outputs[4387];
    assign outputs[4974] = ~((layer0_outputs[3970]) ^ (layer0_outputs[4008]));
    assign outputs[4975] = layer0_outputs[1033];
    assign outputs[4976] = ~(layer0_outputs[3743]);
    assign outputs[4977] = (layer0_outputs[1887]) & ~(layer0_outputs[4033]);
    assign outputs[4978] = (layer0_outputs[1699]) ^ (layer0_outputs[2213]);
    assign outputs[4979] = ~((layer0_outputs[2381]) & (layer0_outputs[3830]));
    assign outputs[4980] = (layer0_outputs[2376]) & ~(layer0_outputs[149]);
    assign outputs[4981] = (layer0_outputs[821]) & ~(layer0_outputs[4153]);
    assign outputs[4982] = (layer0_outputs[4869]) & ~(layer0_outputs[1446]);
    assign outputs[4983] = ~(layer0_outputs[2329]);
    assign outputs[4984] = ~((layer0_outputs[1104]) | (layer0_outputs[369]));
    assign outputs[4985] = (layer0_outputs[210]) ^ (layer0_outputs[4204]);
    assign outputs[4986] = (layer0_outputs[3873]) & ~(layer0_outputs[2256]);
    assign outputs[4987] = ~(layer0_outputs[124]);
    assign outputs[4988] = ~(layer0_outputs[4304]);
    assign outputs[4989] = (layer0_outputs[1072]) ^ (layer0_outputs[142]);
    assign outputs[4990] = ~((layer0_outputs[2883]) ^ (layer0_outputs[2980]));
    assign outputs[4991] = (layer0_outputs[2]) & (layer0_outputs[4448]);
    assign outputs[4992] = ~(layer0_outputs[2687]);
    assign outputs[4993] = ~((layer0_outputs[681]) ^ (layer0_outputs[1645]));
    assign outputs[4994] = (layer0_outputs[302]) & ~(layer0_outputs[3769]);
    assign outputs[4995] = (layer0_outputs[732]) & ~(layer0_outputs[3907]);
    assign outputs[4996] = layer0_outputs[1686];
    assign outputs[4997] = layer0_outputs[1463];
    assign outputs[4998] = (layer0_outputs[4747]) & (layer0_outputs[1857]);
    assign outputs[4999] = ~(layer0_outputs[96]) | (layer0_outputs[3386]);
    assign outputs[5000] = ~(layer0_outputs[333]);
    assign outputs[5001] = (layer0_outputs[2671]) & (layer0_outputs[4546]);
    assign outputs[5002] = ~((layer0_outputs[713]) ^ (layer0_outputs[3928]));
    assign outputs[5003] = ~(layer0_outputs[1649]);
    assign outputs[5004] = (layer0_outputs[2582]) & ~(layer0_outputs[2951]);
    assign outputs[5005] = (layer0_outputs[592]) & ~(layer0_outputs[5027]);
    assign outputs[5006] = ~(layer0_outputs[4352]);
    assign outputs[5007] = (layer0_outputs[425]) ^ (layer0_outputs[936]);
    assign outputs[5008] = ~(layer0_outputs[4365]);
    assign outputs[5009] = (layer0_outputs[1956]) & (layer0_outputs[2407]);
    assign outputs[5010] = (layer0_outputs[1213]) ^ (layer0_outputs[4096]);
    assign outputs[5011] = layer0_outputs[3105];
    assign outputs[5012] = ~(layer0_outputs[2814]);
    assign outputs[5013] = (layer0_outputs[3771]) & ~(layer0_outputs[2492]);
    assign outputs[5014] = (layer0_outputs[1626]) & ~(layer0_outputs[564]);
    assign outputs[5015] = (layer0_outputs[1762]) ^ (layer0_outputs[4863]);
    assign outputs[5016] = ~(layer0_outputs[4900]);
    assign outputs[5017] = ~(layer0_outputs[1917]) | (layer0_outputs[4245]);
    assign outputs[5018] = ~(layer0_outputs[3210]);
    assign outputs[5019] = ~((layer0_outputs[4112]) | (layer0_outputs[3856]));
    assign outputs[5020] = ~(layer0_outputs[1793]) | (layer0_outputs[2224]);
    assign outputs[5021] = (layer0_outputs[4431]) & ~(layer0_outputs[3177]);
    assign outputs[5022] = (layer0_outputs[1019]) & ~(layer0_outputs[2500]);
    assign outputs[5023] = ~((layer0_outputs[949]) & (layer0_outputs[2422]));
    assign outputs[5024] = ~(layer0_outputs[2459]);
    assign outputs[5025] = (layer0_outputs[824]) ^ (layer0_outputs[2235]);
    assign outputs[5026] = ~((layer0_outputs[941]) & (layer0_outputs[4972]));
    assign outputs[5027] = (layer0_outputs[2197]) & (layer0_outputs[3780]);
    assign outputs[5028] = (layer0_outputs[667]) | (layer0_outputs[4764]);
    assign outputs[5029] = layer0_outputs[4638];
    assign outputs[5030] = (layer0_outputs[1798]) & ~(layer0_outputs[899]);
    assign outputs[5031] = (layer0_outputs[672]) & ~(layer0_outputs[629]);
    assign outputs[5032] = ~((layer0_outputs[5096]) | (layer0_outputs[1249]));
    assign outputs[5033] = ~(layer0_outputs[2775]);
    assign outputs[5034] = (layer0_outputs[1669]) & (layer0_outputs[4051]);
    assign outputs[5035] = (layer0_outputs[2037]) ^ (layer0_outputs[767]);
    assign outputs[5036] = ~(layer0_outputs[557]);
    assign outputs[5037] = ~((layer0_outputs[2303]) ^ (layer0_outputs[885]));
    assign outputs[5038] = layer0_outputs[2907];
    assign outputs[5039] = (layer0_outputs[4878]) | (layer0_outputs[2294]);
    assign outputs[5040] = layer0_outputs[2533];
    assign outputs[5041] = (layer0_outputs[4208]) & ~(layer0_outputs[1419]);
    assign outputs[5042] = ~((layer0_outputs[4781]) ^ (layer0_outputs[994]));
    assign outputs[5043] = (layer0_outputs[2048]) & (layer0_outputs[1090]);
    assign outputs[5044] = ~((layer0_outputs[422]) | (layer0_outputs[1116]));
    assign outputs[5045] = (layer0_outputs[4625]) & ~(layer0_outputs[136]);
    assign outputs[5046] = (layer0_outputs[1255]) | (layer0_outputs[1737]);
    assign outputs[5047] = ~((layer0_outputs[1578]) | (layer0_outputs[1068]));
    assign outputs[5048] = ~(layer0_outputs[2620]);
    assign outputs[5049] = (layer0_outputs[3305]) & (layer0_outputs[3064]);
    assign outputs[5050] = (layer0_outputs[2941]) & ~(layer0_outputs[1359]);
    assign outputs[5051] = layer0_outputs[460];
    assign outputs[5052] = (layer0_outputs[4897]) & (layer0_outputs[2777]);
    assign outputs[5053] = layer0_outputs[4721];
    assign outputs[5054] = (layer0_outputs[3364]) & ~(layer0_outputs[75]);
    assign outputs[5055] = layer0_outputs[4557];
    assign outputs[5056] = ~((layer0_outputs[2345]) ^ (layer0_outputs[3880]));
    assign outputs[5057] = ~((layer0_outputs[5049]) | (layer0_outputs[2174]));
    assign outputs[5058] = ~((layer0_outputs[597]) ^ (layer0_outputs[4897]));
    assign outputs[5059] = ~(layer0_outputs[1353]);
    assign outputs[5060] = ~((layer0_outputs[4311]) | (layer0_outputs[861]));
    assign outputs[5061] = (layer0_outputs[646]) & ~(layer0_outputs[1274]);
    assign outputs[5062] = (layer0_outputs[831]) & ~(layer0_outputs[3902]);
    assign outputs[5063] = ~(layer0_outputs[4581]) | (layer0_outputs[1183]);
    assign outputs[5064] = (layer0_outputs[2945]) & ~(layer0_outputs[3462]);
    assign outputs[5065] = layer0_outputs[2412];
    assign outputs[5066] = (layer0_outputs[917]) & ~(layer0_outputs[1859]);
    assign outputs[5067] = ~((layer0_outputs[1796]) | (layer0_outputs[482]));
    assign outputs[5068] = ~((layer0_outputs[2165]) & (layer0_outputs[3070]));
    assign outputs[5069] = ~(layer0_outputs[4077]) | (layer0_outputs[3269]);
    assign outputs[5070] = (layer0_outputs[2864]) & (layer0_outputs[3023]);
    assign outputs[5071] = (layer0_outputs[1911]) & ~(layer0_outputs[1376]);
    assign outputs[5072] = (layer0_outputs[1155]) & (layer0_outputs[4330]);
    assign outputs[5073] = (layer0_outputs[3751]) & (layer0_outputs[4978]);
    assign outputs[5074] = (layer0_outputs[2609]) ^ (layer0_outputs[1485]);
    assign outputs[5075] = layer0_outputs[2970];
    assign outputs[5076] = ~((layer0_outputs[2833]) | (layer0_outputs[4473]));
    assign outputs[5077] = layer0_outputs[4438];
    assign outputs[5078] = layer0_outputs[4986];
    assign outputs[5079] = ~((layer0_outputs[4861]) & (layer0_outputs[3121]));
    assign outputs[5080] = ~((layer0_outputs[4675]) ^ (layer0_outputs[2181]));
    assign outputs[5081] = layer0_outputs[2164];
    assign outputs[5082] = layer0_outputs[3183];
    assign outputs[5083] = ~(layer0_outputs[605]);
    assign outputs[5084] = (layer0_outputs[2255]) & ~(layer0_outputs[4616]);
    assign outputs[5085] = layer0_outputs[874];
    assign outputs[5086] = (layer0_outputs[809]) ^ (layer0_outputs[2626]);
    assign outputs[5087] = (layer0_outputs[3066]) ^ (layer0_outputs[3166]);
    assign outputs[5088] = ~((layer0_outputs[3616]) | (layer0_outputs[334]));
    assign outputs[5089] = layer0_outputs[530];
    assign outputs[5090] = layer0_outputs[84];
    assign outputs[5091] = ~((layer0_outputs[1539]) & (layer0_outputs[3070]));
    assign outputs[5092] = ~((layer0_outputs[5046]) ^ (layer0_outputs[372]));
    assign outputs[5093] = (layer0_outputs[4269]) & ~(layer0_outputs[4469]);
    assign outputs[5094] = ~((layer0_outputs[3191]) ^ (layer0_outputs[681]));
    assign outputs[5095] = layer0_outputs[2288];
    assign outputs[5096] = (layer0_outputs[4220]) & ~(layer0_outputs[3768]);
    assign outputs[5097] = (layer0_outputs[1181]) & ~(layer0_outputs[4603]);
    assign outputs[5098] = (layer0_outputs[2553]) & ~(layer0_outputs[1310]);
    assign outputs[5099] = layer0_outputs[802];
    assign outputs[5100] = ~(layer0_outputs[3036]);
    assign outputs[5101] = layer0_outputs[2572];
    assign outputs[5102] = ~((layer0_outputs[2474]) ^ (layer0_outputs[1278]));
    assign outputs[5103] = (layer0_outputs[1315]) & (layer0_outputs[4296]);
    assign outputs[5104] = ~((layer0_outputs[908]) | (layer0_outputs[2832]));
    assign outputs[5105] = layer0_outputs[1653];
    assign outputs[5106] = layer0_outputs[2438];
    assign outputs[5107] = (layer0_outputs[3777]) ^ (layer0_outputs[581]);
    assign outputs[5108] = ~((layer0_outputs[3828]) ^ (layer0_outputs[4417]));
    assign outputs[5109] = ~((layer0_outputs[565]) | (layer0_outputs[1704]));
    assign outputs[5110] = (layer0_outputs[2755]) ^ (layer0_outputs[2118]);
    assign outputs[5111] = ~((layer0_outputs[2115]) & (layer0_outputs[4790]));
    assign outputs[5112] = (layer0_outputs[645]) ^ (layer0_outputs[4062]);
    assign outputs[5113] = 1'b0;
    assign outputs[5114] = ~((layer0_outputs[2537]) | (layer0_outputs[359]));
    assign outputs[5115] = layer0_outputs[2402];
    assign outputs[5116] = (layer0_outputs[4088]) & ~(layer0_outputs[3512]);
    assign outputs[5117] = (layer0_outputs[2497]) & ~(layer0_outputs[4928]);
    assign outputs[5118] = (layer0_outputs[1517]) & ~(layer0_outputs[4663]);
    assign outputs[5119] = (layer0_outputs[3017]) & ~(layer0_outputs[3599]);
endmodule
