library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(10239 downto 0);
    signal layer1_outputs: std_logic_vector(10239 downto 0);
    signal layer2_outputs: std_logic_vector(10239 downto 0);
    signal layer3_outputs: std_logic_vector(10239 downto 0);
    signal layer4_outputs: std_logic_vector(10239 downto 0);
    signal layer5_outputs: std_logic_vector(10239 downto 0);
    signal layer6_outputs: std_logic_vector(10239 downto 0);
    signal layer7_outputs: std_logic_vector(10239 downto 0);
    signal layer8_outputs: std_logic_vector(10239 downto 0);

begin
    layer0_outputs(0) <= not (a or b);
    layer0_outputs(1) <= 1'b1;
    layer0_outputs(2) <= not b;
    layer0_outputs(3) <= not b or a;
    layer0_outputs(4) <= a;
    layer0_outputs(5) <= not a;
    layer0_outputs(6) <= not (a or b);
    layer0_outputs(7) <= b and not a;
    layer0_outputs(8) <= not a;
    layer0_outputs(9) <= a and not b;
    layer0_outputs(10) <= not a;
    layer0_outputs(11) <= a;
    layer0_outputs(12) <= a and not b;
    layer0_outputs(13) <= 1'b1;
    layer0_outputs(14) <= not (a xor b);
    layer0_outputs(15) <= a or b;
    layer0_outputs(16) <= 1'b0;
    layer0_outputs(17) <= a and not b;
    layer0_outputs(18) <= b;
    layer0_outputs(19) <= b;
    layer0_outputs(20) <= not (a xor b);
    layer0_outputs(21) <= not (a and b);
    layer0_outputs(22) <= 1'b0;
    layer0_outputs(23) <= b;
    layer0_outputs(24) <= a or b;
    layer0_outputs(25) <= not (a xor b);
    layer0_outputs(26) <= a;
    layer0_outputs(27) <= b and not a;
    layer0_outputs(28) <= a;
    layer0_outputs(29) <= a and b;
    layer0_outputs(30) <= 1'b0;
    layer0_outputs(31) <= b and not a;
    layer0_outputs(32) <= not a;
    layer0_outputs(33) <= not b;
    layer0_outputs(34) <= not a;
    layer0_outputs(35) <= not (a xor b);
    layer0_outputs(36) <= a xor b;
    layer0_outputs(37) <= a or b;
    layer0_outputs(38) <= a or b;
    layer0_outputs(39) <= not (a and b);
    layer0_outputs(40) <= a and b;
    layer0_outputs(41) <= a and b;
    layer0_outputs(42) <= not a;
    layer0_outputs(43) <= not (a or b);
    layer0_outputs(44) <= b;
    layer0_outputs(45) <= 1'b1;
    layer0_outputs(46) <= 1'b1;
    layer0_outputs(47) <= not (a and b);
    layer0_outputs(48) <= a and b;
    layer0_outputs(49) <= 1'b1;
    layer0_outputs(50) <= 1'b0;
    layer0_outputs(51) <= b;
    layer0_outputs(52) <= not a;
    layer0_outputs(53) <= not a or b;
    layer0_outputs(54) <= a or b;
    layer0_outputs(55) <= not a or b;
    layer0_outputs(56) <= 1'b0;
    layer0_outputs(57) <= not (a or b);
    layer0_outputs(58) <= not b;
    layer0_outputs(59) <= not a or b;
    layer0_outputs(60) <= b;
    layer0_outputs(61) <= b and not a;
    layer0_outputs(62) <= not a;
    layer0_outputs(63) <= not b;
    layer0_outputs(64) <= a and b;
    layer0_outputs(65) <= 1'b0;
    layer0_outputs(66) <= not a;
    layer0_outputs(67) <= b;
    layer0_outputs(68) <= not (a or b);
    layer0_outputs(69) <= not a;
    layer0_outputs(70) <= 1'b0;
    layer0_outputs(71) <= not b or a;
    layer0_outputs(72) <= not a;
    layer0_outputs(73) <= 1'b0;
    layer0_outputs(74) <= not b;
    layer0_outputs(75) <= not (a or b);
    layer0_outputs(76) <= a;
    layer0_outputs(77) <= not a or b;
    layer0_outputs(78) <= b;
    layer0_outputs(79) <= a or b;
    layer0_outputs(80) <= a or b;
    layer0_outputs(81) <= not a;
    layer0_outputs(82) <= 1'b0;
    layer0_outputs(83) <= not (a or b);
    layer0_outputs(84) <= a or b;
    layer0_outputs(85) <= 1'b1;
    layer0_outputs(86) <= not a or b;
    layer0_outputs(87) <= not (a and b);
    layer0_outputs(88) <= a and not b;
    layer0_outputs(89) <= not (a xor b);
    layer0_outputs(90) <= not b or a;
    layer0_outputs(91) <= a;
    layer0_outputs(92) <= a;
    layer0_outputs(93) <= a;
    layer0_outputs(94) <= a and b;
    layer0_outputs(95) <= not (a and b);
    layer0_outputs(96) <= a and b;
    layer0_outputs(97) <= b;
    layer0_outputs(98) <= not (a and b);
    layer0_outputs(99) <= not a;
    layer0_outputs(100) <= not (a xor b);
    layer0_outputs(101) <= 1'b0;
    layer0_outputs(102) <= not (a or b);
    layer0_outputs(103) <= not (a and b);
    layer0_outputs(104) <= a and not b;
    layer0_outputs(105) <= a xor b;
    layer0_outputs(106) <= a;
    layer0_outputs(107) <= not b;
    layer0_outputs(108) <= not b;
    layer0_outputs(109) <= a and b;
    layer0_outputs(110) <= not (a xor b);
    layer0_outputs(111) <= not (a and b);
    layer0_outputs(112) <= not (a and b);
    layer0_outputs(113) <= a;
    layer0_outputs(114) <= not (a xor b);
    layer0_outputs(115) <= a or b;
    layer0_outputs(116) <= a xor b;
    layer0_outputs(117) <= b;
    layer0_outputs(118) <= not a or b;
    layer0_outputs(119) <= b;
    layer0_outputs(120) <= 1'b0;
    layer0_outputs(121) <= not (a xor b);
    layer0_outputs(122) <= b;
    layer0_outputs(123) <= 1'b0;
    layer0_outputs(124) <= not b or a;
    layer0_outputs(125) <= not (a or b);
    layer0_outputs(126) <= a;
    layer0_outputs(127) <= not b;
    layer0_outputs(128) <= not b or a;
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= not (a or b);
    layer0_outputs(131) <= not a;
    layer0_outputs(132) <= b;
    layer0_outputs(133) <= not b or a;
    layer0_outputs(134) <= not b or a;
    layer0_outputs(135) <= not (a and b);
    layer0_outputs(136) <= not a or b;
    layer0_outputs(137) <= 1'b1;
    layer0_outputs(138) <= b;
    layer0_outputs(139) <= a;
    layer0_outputs(140) <= not b or a;
    layer0_outputs(141) <= 1'b1;
    layer0_outputs(142) <= a;
    layer0_outputs(143) <= a and not b;
    layer0_outputs(144) <= a and not b;
    layer0_outputs(145) <= a and b;
    layer0_outputs(146) <= b;
    layer0_outputs(147) <= not (a or b);
    layer0_outputs(148) <= a and b;
    layer0_outputs(149) <= not a or b;
    layer0_outputs(150) <= a or b;
    layer0_outputs(151) <= not (a or b);
    layer0_outputs(152) <= a and not b;
    layer0_outputs(153) <= b;
    layer0_outputs(154) <= a or b;
    layer0_outputs(155) <= not a or b;
    layer0_outputs(156) <= not b or a;
    layer0_outputs(157) <= a and not b;
    layer0_outputs(158) <= 1'b0;
    layer0_outputs(159) <= a and b;
    layer0_outputs(160) <= a or b;
    layer0_outputs(161) <= a;
    layer0_outputs(162) <= a and b;
    layer0_outputs(163) <= 1'b0;
    layer0_outputs(164) <= b and not a;
    layer0_outputs(165) <= not (a and b);
    layer0_outputs(166) <= not b or a;
    layer0_outputs(167) <= not b;
    layer0_outputs(168) <= a;
    layer0_outputs(169) <= b;
    layer0_outputs(170) <= 1'b0;
    layer0_outputs(171) <= a and b;
    layer0_outputs(172) <= not (a and b);
    layer0_outputs(173) <= 1'b0;
    layer0_outputs(174) <= not b;
    layer0_outputs(175) <= a;
    layer0_outputs(176) <= not b or a;
    layer0_outputs(177) <= not a or b;
    layer0_outputs(178) <= 1'b0;
    layer0_outputs(179) <= a and b;
    layer0_outputs(180) <= not b or a;
    layer0_outputs(181) <= not a;
    layer0_outputs(182) <= a and not b;
    layer0_outputs(183) <= b and not a;
    layer0_outputs(184) <= 1'b1;
    layer0_outputs(185) <= not a or b;
    layer0_outputs(186) <= not (a and b);
    layer0_outputs(187) <= not (a and b);
    layer0_outputs(188) <= 1'b0;
    layer0_outputs(189) <= not (a or b);
    layer0_outputs(190) <= a and not b;
    layer0_outputs(191) <= b and not a;
    layer0_outputs(192) <= 1'b1;
    layer0_outputs(193) <= a;
    layer0_outputs(194) <= not b or a;
    layer0_outputs(195) <= not b or a;
    layer0_outputs(196) <= not (a xor b);
    layer0_outputs(197) <= 1'b1;
    layer0_outputs(198) <= not (a or b);
    layer0_outputs(199) <= not a or b;
    layer0_outputs(200) <= b;
    layer0_outputs(201) <= a and not b;
    layer0_outputs(202) <= a and b;
    layer0_outputs(203) <= b and not a;
    layer0_outputs(204) <= not a;
    layer0_outputs(205) <= b;
    layer0_outputs(206) <= 1'b1;
    layer0_outputs(207) <= not (a and b);
    layer0_outputs(208) <= a or b;
    layer0_outputs(209) <= 1'b0;
    layer0_outputs(210) <= a and b;
    layer0_outputs(211) <= a or b;
    layer0_outputs(212) <= not (a or b);
    layer0_outputs(213) <= a xor b;
    layer0_outputs(214) <= a and not b;
    layer0_outputs(215) <= a or b;
    layer0_outputs(216) <= a or b;
    layer0_outputs(217) <= 1'b1;
    layer0_outputs(218) <= a xor b;
    layer0_outputs(219) <= a and b;
    layer0_outputs(220) <= a and not b;
    layer0_outputs(221) <= not b;
    layer0_outputs(222) <= not b;
    layer0_outputs(223) <= b and not a;
    layer0_outputs(224) <= a xor b;
    layer0_outputs(225) <= b;
    layer0_outputs(226) <= b and not a;
    layer0_outputs(227) <= 1'b0;
    layer0_outputs(228) <= not (a and b);
    layer0_outputs(229) <= not b or a;
    layer0_outputs(230) <= not a or b;
    layer0_outputs(231) <= not (a or b);
    layer0_outputs(232) <= b;
    layer0_outputs(233) <= a;
    layer0_outputs(234) <= 1'b1;
    layer0_outputs(235) <= not a or b;
    layer0_outputs(236) <= a;
    layer0_outputs(237) <= 1'b1;
    layer0_outputs(238) <= not b or a;
    layer0_outputs(239) <= 1'b0;
    layer0_outputs(240) <= 1'b0;
    layer0_outputs(241) <= a or b;
    layer0_outputs(242) <= a and not b;
    layer0_outputs(243) <= not (a and b);
    layer0_outputs(244) <= not (a and b);
    layer0_outputs(245) <= not (a xor b);
    layer0_outputs(246) <= not a;
    layer0_outputs(247) <= a or b;
    layer0_outputs(248) <= b and not a;
    layer0_outputs(249) <= a;
    layer0_outputs(250) <= 1'b0;
    layer0_outputs(251) <= not a;
    layer0_outputs(252) <= not a or b;
    layer0_outputs(253) <= a or b;
    layer0_outputs(254) <= 1'b1;
    layer0_outputs(255) <= a and not b;
    layer0_outputs(256) <= a and not b;
    layer0_outputs(257) <= not a or b;
    layer0_outputs(258) <= a and not b;
    layer0_outputs(259) <= not a or b;
    layer0_outputs(260) <= 1'b1;
    layer0_outputs(261) <= not a or b;
    layer0_outputs(262) <= b;
    layer0_outputs(263) <= a and b;
    layer0_outputs(264) <= not (a or b);
    layer0_outputs(265) <= b;
    layer0_outputs(266) <= 1'b1;
    layer0_outputs(267) <= not (a or b);
    layer0_outputs(268) <= a and not b;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= 1'b1;
    layer0_outputs(271) <= a and not b;
    layer0_outputs(272) <= a;
    layer0_outputs(273) <= a and not b;
    layer0_outputs(274) <= b and not a;
    layer0_outputs(275) <= 1'b1;
    layer0_outputs(276) <= b;
    layer0_outputs(277) <= not (a or b);
    layer0_outputs(278) <= not a;
    layer0_outputs(279) <= a or b;
    layer0_outputs(280) <= not (a or b);
    layer0_outputs(281) <= a or b;
    layer0_outputs(282) <= not a or b;
    layer0_outputs(283) <= not (a and b);
    layer0_outputs(284) <= b;
    layer0_outputs(285) <= a xor b;
    layer0_outputs(286) <= a;
    layer0_outputs(287) <= b;
    layer0_outputs(288) <= not (a xor b);
    layer0_outputs(289) <= b;
    layer0_outputs(290) <= b;
    layer0_outputs(291) <= not (a xor b);
    layer0_outputs(292) <= a;
    layer0_outputs(293) <= 1'b1;
    layer0_outputs(294) <= not (a and b);
    layer0_outputs(295) <= a;
    layer0_outputs(296) <= not a or b;
    layer0_outputs(297) <= not a;
    layer0_outputs(298) <= a and b;
    layer0_outputs(299) <= not (a and b);
    layer0_outputs(300) <= not (a or b);
    layer0_outputs(301) <= a or b;
    layer0_outputs(302) <= b and not a;
    layer0_outputs(303) <= not a or b;
    layer0_outputs(304) <= a or b;
    layer0_outputs(305) <= b and not a;
    layer0_outputs(306) <= b;
    layer0_outputs(307) <= not (a and b);
    layer0_outputs(308) <= a;
    layer0_outputs(309) <= b and not a;
    layer0_outputs(310) <= 1'b1;
    layer0_outputs(311) <= not b or a;
    layer0_outputs(312) <= 1'b1;
    layer0_outputs(313) <= not (a or b);
    layer0_outputs(314) <= b and not a;
    layer0_outputs(315) <= not a or b;
    layer0_outputs(316) <= 1'b0;
    layer0_outputs(317) <= b and not a;
    layer0_outputs(318) <= not (a or b);
    layer0_outputs(319) <= a or b;
    layer0_outputs(320) <= a xor b;
    layer0_outputs(321) <= not a;
    layer0_outputs(322) <= b;
    layer0_outputs(323) <= not a;
    layer0_outputs(324) <= not (a and b);
    layer0_outputs(325) <= 1'b0;
    layer0_outputs(326) <= not b;
    layer0_outputs(327) <= not (a xor b);
    layer0_outputs(328) <= not (a and b);
    layer0_outputs(329) <= not (a or b);
    layer0_outputs(330) <= 1'b0;
    layer0_outputs(331) <= not b;
    layer0_outputs(332) <= a and not b;
    layer0_outputs(333) <= not a or b;
    layer0_outputs(334) <= a or b;
    layer0_outputs(335) <= b and not a;
    layer0_outputs(336) <= 1'b1;
    layer0_outputs(337) <= b;
    layer0_outputs(338) <= 1'b0;
    layer0_outputs(339) <= a or b;
    layer0_outputs(340) <= b and not a;
    layer0_outputs(341) <= a and b;
    layer0_outputs(342) <= a and not b;
    layer0_outputs(343) <= a and b;
    layer0_outputs(344) <= b;
    layer0_outputs(345) <= b;
    layer0_outputs(346) <= not (a xor b);
    layer0_outputs(347) <= not (a or b);
    layer0_outputs(348) <= a;
    layer0_outputs(349) <= a and not b;
    layer0_outputs(350) <= not (a xor b);
    layer0_outputs(351) <= not (a xor b);
    layer0_outputs(352) <= b and not a;
    layer0_outputs(353) <= 1'b1;
    layer0_outputs(354) <= not a or b;
    layer0_outputs(355) <= not a or b;
    layer0_outputs(356) <= not b;
    layer0_outputs(357) <= b and not a;
    layer0_outputs(358) <= a and not b;
    layer0_outputs(359) <= a;
    layer0_outputs(360) <= a and not b;
    layer0_outputs(361) <= not a;
    layer0_outputs(362) <= a;
    layer0_outputs(363) <= a;
    layer0_outputs(364) <= 1'b0;
    layer0_outputs(365) <= not (a and b);
    layer0_outputs(366) <= not b or a;
    layer0_outputs(367) <= 1'b1;
    layer0_outputs(368) <= not b or a;
    layer0_outputs(369) <= b and not a;
    layer0_outputs(370) <= a or b;
    layer0_outputs(371) <= 1'b0;
    layer0_outputs(372) <= a;
    layer0_outputs(373) <= not a;
    layer0_outputs(374) <= b;
    layer0_outputs(375) <= 1'b0;
    layer0_outputs(376) <= a and b;
    layer0_outputs(377) <= b;
    layer0_outputs(378) <= b and not a;
    layer0_outputs(379) <= not b or a;
    layer0_outputs(380) <= not b;
    layer0_outputs(381) <= not b;
    layer0_outputs(382) <= not b or a;
    layer0_outputs(383) <= not b;
    layer0_outputs(384) <= not (a or b);
    layer0_outputs(385) <= b;
    layer0_outputs(386) <= not (a or b);
    layer0_outputs(387) <= a or b;
    layer0_outputs(388) <= a and not b;
    layer0_outputs(389) <= not b;
    layer0_outputs(390) <= 1'b0;
    layer0_outputs(391) <= a xor b;
    layer0_outputs(392) <= 1'b0;
    layer0_outputs(393) <= not a or b;
    layer0_outputs(394) <= a xor b;
    layer0_outputs(395) <= 1'b1;
    layer0_outputs(396) <= not (a and b);
    layer0_outputs(397) <= not (a and b);
    layer0_outputs(398) <= not b;
    layer0_outputs(399) <= a and not b;
    layer0_outputs(400) <= not b;
    layer0_outputs(401) <= not (a and b);
    layer0_outputs(402) <= not b;
    layer0_outputs(403) <= a;
    layer0_outputs(404) <= not a or b;
    layer0_outputs(405) <= not a;
    layer0_outputs(406) <= not b or a;
    layer0_outputs(407) <= not b or a;
    layer0_outputs(408) <= a and b;
    layer0_outputs(409) <= not a;
    layer0_outputs(410) <= not a or b;
    layer0_outputs(411) <= not (a xor b);
    layer0_outputs(412) <= not (a and b);
    layer0_outputs(413) <= not (a or b);
    layer0_outputs(414) <= not (a or b);
    layer0_outputs(415) <= a xor b;
    layer0_outputs(416) <= 1'b1;
    layer0_outputs(417) <= a or b;
    layer0_outputs(418) <= not a;
    layer0_outputs(419) <= not (a xor b);
    layer0_outputs(420) <= 1'b0;
    layer0_outputs(421) <= a and b;
    layer0_outputs(422) <= not (a or b);
    layer0_outputs(423) <= a and not b;
    layer0_outputs(424) <= a;
    layer0_outputs(425) <= a and b;
    layer0_outputs(426) <= not (a xor b);
    layer0_outputs(427) <= a or b;
    layer0_outputs(428) <= not b or a;
    layer0_outputs(429) <= not b or a;
    layer0_outputs(430) <= not a or b;
    layer0_outputs(431) <= not b;
    layer0_outputs(432) <= not b;
    layer0_outputs(433) <= b and not a;
    layer0_outputs(434) <= b;
    layer0_outputs(435) <= not a;
    layer0_outputs(436) <= not (a or b);
    layer0_outputs(437) <= not a;
    layer0_outputs(438) <= a and b;
    layer0_outputs(439) <= not (a and b);
    layer0_outputs(440) <= not a or b;
    layer0_outputs(441) <= a and b;
    layer0_outputs(442) <= not (a or b);
    layer0_outputs(443) <= b and not a;
    layer0_outputs(444) <= b;
    layer0_outputs(445) <= a;
    layer0_outputs(446) <= b;
    layer0_outputs(447) <= not b;
    layer0_outputs(448) <= b;
    layer0_outputs(449) <= not (a and b);
    layer0_outputs(450) <= a and not b;
    layer0_outputs(451) <= not a;
    layer0_outputs(452) <= a and not b;
    layer0_outputs(453) <= not (a xor b);
    layer0_outputs(454) <= a xor b;
    layer0_outputs(455) <= not a;
    layer0_outputs(456) <= a;
    layer0_outputs(457) <= a;
    layer0_outputs(458) <= not b;
    layer0_outputs(459) <= 1'b1;
    layer0_outputs(460) <= 1'b0;
    layer0_outputs(461) <= b and not a;
    layer0_outputs(462) <= not a or b;
    layer0_outputs(463) <= 1'b0;
    layer0_outputs(464) <= a;
    layer0_outputs(465) <= not a or b;
    layer0_outputs(466) <= not (a and b);
    layer0_outputs(467) <= not (a and b);
    layer0_outputs(468) <= not b;
    layer0_outputs(469) <= not (a xor b);
    layer0_outputs(470) <= not a or b;
    layer0_outputs(471) <= not b or a;
    layer0_outputs(472) <= a;
    layer0_outputs(473) <= not b or a;
    layer0_outputs(474) <= a;
    layer0_outputs(475) <= a;
    layer0_outputs(476) <= b;
    layer0_outputs(477) <= a and b;
    layer0_outputs(478) <= a and b;
    layer0_outputs(479) <= b and not a;
    layer0_outputs(480) <= not (a xor b);
    layer0_outputs(481) <= not b;
    layer0_outputs(482) <= not (a and b);
    layer0_outputs(483) <= a xor b;
    layer0_outputs(484) <= 1'b1;
    layer0_outputs(485) <= 1'b1;
    layer0_outputs(486) <= a and b;
    layer0_outputs(487) <= a and not b;
    layer0_outputs(488) <= not (a or b);
    layer0_outputs(489) <= a and not b;
    layer0_outputs(490) <= not (a and b);
    layer0_outputs(491) <= a;
    layer0_outputs(492) <= a;
    layer0_outputs(493) <= 1'b0;
    layer0_outputs(494) <= not a or b;
    layer0_outputs(495) <= a and b;
    layer0_outputs(496) <= b and not a;
    layer0_outputs(497) <= not (a or b);
    layer0_outputs(498) <= not a or b;
    layer0_outputs(499) <= a or b;
    layer0_outputs(500) <= a and not b;
    layer0_outputs(501) <= not (a or b);
    layer0_outputs(502) <= not (a or b);
    layer0_outputs(503) <= not a or b;
    layer0_outputs(504) <= not (a and b);
    layer0_outputs(505) <= a and b;
    layer0_outputs(506) <= not b;
    layer0_outputs(507) <= not a or b;
    layer0_outputs(508) <= a and not b;
    layer0_outputs(509) <= a xor b;
    layer0_outputs(510) <= not a or b;
    layer0_outputs(511) <= b;
    layer0_outputs(512) <= a and not b;
    layer0_outputs(513) <= a and not b;
    layer0_outputs(514) <= b and not a;
    layer0_outputs(515) <= a or b;
    layer0_outputs(516) <= not b;
    layer0_outputs(517) <= not b or a;
    layer0_outputs(518) <= a and b;
    layer0_outputs(519) <= b;
    layer0_outputs(520) <= not (a and b);
    layer0_outputs(521) <= 1'b0;
    layer0_outputs(522) <= not b;
    layer0_outputs(523) <= b and not a;
    layer0_outputs(524) <= not b or a;
    layer0_outputs(525) <= not (a or b);
    layer0_outputs(526) <= a;
    layer0_outputs(527) <= a and b;
    layer0_outputs(528) <= not a or b;
    layer0_outputs(529) <= not b;
    layer0_outputs(530) <= not (a and b);
    layer0_outputs(531) <= b and not a;
    layer0_outputs(532) <= a and b;
    layer0_outputs(533) <= b;
    layer0_outputs(534) <= a xor b;
    layer0_outputs(535) <= not (a and b);
    layer0_outputs(536) <= not b;
    layer0_outputs(537) <= not a;
    layer0_outputs(538) <= not a;
    layer0_outputs(539) <= b and not a;
    layer0_outputs(540) <= not (a xor b);
    layer0_outputs(541) <= b and not a;
    layer0_outputs(542) <= a xor b;
    layer0_outputs(543) <= not (a or b);
    layer0_outputs(544) <= 1'b0;
    layer0_outputs(545) <= not b;
    layer0_outputs(546) <= not (a or b);
    layer0_outputs(547) <= not b;
    layer0_outputs(548) <= a and not b;
    layer0_outputs(549) <= not b or a;
    layer0_outputs(550) <= not a or b;
    layer0_outputs(551) <= a and b;
    layer0_outputs(552) <= a or b;
    layer0_outputs(553) <= b;
    layer0_outputs(554) <= a xor b;
    layer0_outputs(555) <= a or b;
    layer0_outputs(556) <= not b;
    layer0_outputs(557) <= not (a and b);
    layer0_outputs(558) <= a or b;
    layer0_outputs(559) <= not a or b;
    layer0_outputs(560) <= not b or a;
    layer0_outputs(561) <= b and not a;
    layer0_outputs(562) <= 1'b0;
    layer0_outputs(563) <= not (a or b);
    layer0_outputs(564) <= a xor b;
    layer0_outputs(565) <= not (a and b);
    layer0_outputs(566) <= not b;
    layer0_outputs(567) <= not b;
    layer0_outputs(568) <= not (a xor b);
    layer0_outputs(569) <= not (a xor b);
    layer0_outputs(570) <= b and not a;
    layer0_outputs(571) <= 1'b0;
    layer0_outputs(572) <= not b or a;
    layer0_outputs(573) <= not (a xor b);
    layer0_outputs(574) <= a or b;
    layer0_outputs(575) <= b and not a;
    layer0_outputs(576) <= a or b;
    layer0_outputs(577) <= not a or b;
    layer0_outputs(578) <= not a;
    layer0_outputs(579) <= b and not a;
    layer0_outputs(580) <= 1'b1;
    layer0_outputs(581) <= not b or a;
    layer0_outputs(582) <= a xor b;
    layer0_outputs(583) <= a and not b;
    layer0_outputs(584) <= not (a and b);
    layer0_outputs(585) <= b;
    layer0_outputs(586) <= a and not b;
    layer0_outputs(587) <= 1'b1;
    layer0_outputs(588) <= not (a xor b);
    layer0_outputs(589) <= 1'b1;
    layer0_outputs(590) <= not b;
    layer0_outputs(591) <= not b or a;
    layer0_outputs(592) <= a and b;
    layer0_outputs(593) <= not (a and b);
    layer0_outputs(594) <= a;
    layer0_outputs(595) <= 1'b1;
    layer0_outputs(596) <= not a or b;
    layer0_outputs(597) <= not (a xor b);
    layer0_outputs(598) <= b and not a;
    layer0_outputs(599) <= not a or b;
    layer0_outputs(600) <= b;
    layer0_outputs(601) <= a or b;
    layer0_outputs(602) <= a and b;
    layer0_outputs(603) <= b;
    layer0_outputs(604) <= b;
    layer0_outputs(605) <= not b;
    layer0_outputs(606) <= not (a xor b);
    layer0_outputs(607) <= b and not a;
    layer0_outputs(608) <= b;
    layer0_outputs(609) <= not a or b;
    layer0_outputs(610) <= not (a and b);
    layer0_outputs(611) <= a;
    layer0_outputs(612) <= b;
    layer0_outputs(613) <= not b or a;
    layer0_outputs(614) <= 1'b1;
    layer0_outputs(615) <= a;
    layer0_outputs(616) <= a and not b;
    layer0_outputs(617) <= a and not b;
    layer0_outputs(618) <= a and not b;
    layer0_outputs(619) <= not (a and b);
    layer0_outputs(620) <= not a;
    layer0_outputs(621) <= b;
    layer0_outputs(622) <= a xor b;
    layer0_outputs(623) <= a xor b;
    layer0_outputs(624) <= b;
    layer0_outputs(625) <= b and not a;
    layer0_outputs(626) <= b;
    layer0_outputs(627) <= a and not b;
    layer0_outputs(628) <= not (a xor b);
    layer0_outputs(629) <= a and b;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= 1'b1;
    layer0_outputs(632) <= 1'b0;
    layer0_outputs(633) <= not (a or b);
    layer0_outputs(634) <= a and b;
    layer0_outputs(635) <= not b;
    layer0_outputs(636) <= not (a xor b);
    layer0_outputs(637) <= 1'b1;
    layer0_outputs(638) <= not a or b;
    layer0_outputs(639) <= not (a xor b);
    layer0_outputs(640) <= a xor b;
    layer0_outputs(641) <= a;
    layer0_outputs(642) <= a and b;
    layer0_outputs(643) <= b;
    layer0_outputs(644) <= a and b;
    layer0_outputs(645) <= not b or a;
    layer0_outputs(646) <= 1'b0;
    layer0_outputs(647) <= not (a or b);
    layer0_outputs(648) <= 1'b1;
    layer0_outputs(649) <= not b or a;
    layer0_outputs(650) <= not a or b;
    layer0_outputs(651) <= 1'b0;
    layer0_outputs(652) <= not a;
    layer0_outputs(653) <= 1'b0;
    layer0_outputs(654) <= not (a and b);
    layer0_outputs(655) <= not (a or b);
    layer0_outputs(656) <= b;
    layer0_outputs(657) <= not b;
    layer0_outputs(658) <= a;
    layer0_outputs(659) <= not a;
    layer0_outputs(660) <= not b;
    layer0_outputs(661) <= 1'b0;
    layer0_outputs(662) <= not b;
    layer0_outputs(663) <= b and not a;
    layer0_outputs(664) <= a;
    layer0_outputs(665) <= not b;
    layer0_outputs(666) <= 1'b1;
    layer0_outputs(667) <= a and b;
    layer0_outputs(668) <= b and not a;
    layer0_outputs(669) <= a and not b;
    layer0_outputs(670) <= a;
    layer0_outputs(671) <= a;
    layer0_outputs(672) <= not (a or b);
    layer0_outputs(673) <= not a or b;
    layer0_outputs(674) <= not a;
    layer0_outputs(675) <= a or b;
    layer0_outputs(676) <= not (a or b);
    layer0_outputs(677) <= b;
    layer0_outputs(678) <= a;
    layer0_outputs(679) <= not (a or b);
    layer0_outputs(680) <= a;
    layer0_outputs(681) <= a and b;
    layer0_outputs(682) <= 1'b0;
    layer0_outputs(683) <= not (a or b);
    layer0_outputs(684) <= not (a or b);
    layer0_outputs(685) <= not a or b;
    layer0_outputs(686) <= a;
    layer0_outputs(687) <= not (a and b);
    layer0_outputs(688) <= b and not a;
    layer0_outputs(689) <= a;
    layer0_outputs(690) <= not b or a;
    layer0_outputs(691) <= not (a xor b);
    layer0_outputs(692) <= a;
    layer0_outputs(693) <= a;
    layer0_outputs(694) <= not a or b;
    layer0_outputs(695) <= not (a or b);
    layer0_outputs(696) <= not b;
    layer0_outputs(697) <= a xor b;
    layer0_outputs(698) <= a and b;
    layer0_outputs(699) <= not (a and b);
    layer0_outputs(700) <= not a or b;
    layer0_outputs(701) <= 1'b1;
    layer0_outputs(702) <= 1'b1;
    layer0_outputs(703) <= not a;
    layer0_outputs(704) <= 1'b1;
    layer0_outputs(705) <= not b or a;
    layer0_outputs(706) <= b and not a;
    layer0_outputs(707) <= a;
    layer0_outputs(708) <= b and not a;
    layer0_outputs(709) <= not b or a;
    layer0_outputs(710) <= b and not a;
    layer0_outputs(711) <= not a;
    layer0_outputs(712) <= a;
    layer0_outputs(713) <= b and not a;
    layer0_outputs(714) <= b;
    layer0_outputs(715) <= not a or b;
    layer0_outputs(716) <= not a or b;
    layer0_outputs(717) <= not (a and b);
    layer0_outputs(718) <= not b;
    layer0_outputs(719) <= not (a xor b);
    layer0_outputs(720) <= not b or a;
    layer0_outputs(721) <= a xor b;
    layer0_outputs(722) <= 1'b1;
    layer0_outputs(723) <= b and not a;
    layer0_outputs(724) <= not (a or b);
    layer0_outputs(725) <= not a;
    layer0_outputs(726) <= 1'b0;
    layer0_outputs(727) <= a;
    layer0_outputs(728) <= 1'b1;
    layer0_outputs(729) <= not a;
    layer0_outputs(730) <= a xor b;
    layer0_outputs(731) <= a or b;
    layer0_outputs(732) <= a and b;
    layer0_outputs(733) <= a xor b;
    layer0_outputs(734) <= not (a and b);
    layer0_outputs(735) <= not a;
    layer0_outputs(736) <= not (a or b);
    layer0_outputs(737) <= not b;
    layer0_outputs(738) <= not (a or b);
    layer0_outputs(739) <= not a or b;
    layer0_outputs(740) <= a or b;
    layer0_outputs(741) <= not (a or b);
    layer0_outputs(742) <= b;
    layer0_outputs(743) <= b;
    layer0_outputs(744) <= not b or a;
    layer0_outputs(745) <= not (a or b);
    layer0_outputs(746) <= 1'b1;
    layer0_outputs(747) <= not (a or b);
    layer0_outputs(748) <= not a or b;
    layer0_outputs(749) <= not a or b;
    layer0_outputs(750) <= a and not b;
    layer0_outputs(751) <= not b or a;
    layer0_outputs(752) <= 1'b0;
    layer0_outputs(753) <= not a;
    layer0_outputs(754) <= not a or b;
    layer0_outputs(755) <= not b;
    layer0_outputs(756) <= a and not b;
    layer0_outputs(757) <= not a or b;
    layer0_outputs(758) <= a xor b;
    layer0_outputs(759) <= a;
    layer0_outputs(760) <= b;
    layer0_outputs(761) <= 1'b1;
    layer0_outputs(762) <= not (a and b);
    layer0_outputs(763) <= 1'b0;
    layer0_outputs(764) <= 1'b1;
    layer0_outputs(765) <= a or b;
    layer0_outputs(766) <= a and not b;
    layer0_outputs(767) <= b and not a;
    layer0_outputs(768) <= a and not b;
    layer0_outputs(769) <= not (a and b);
    layer0_outputs(770) <= not a or b;
    layer0_outputs(771) <= b;
    layer0_outputs(772) <= not a;
    layer0_outputs(773) <= not a;
    layer0_outputs(774) <= not a;
    layer0_outputs(775) <= not b or a;
    layer0_outputs(776) <= a xor b;
    layer0_outputs(777) <= not (a and b);
    layer0_outputs(778) <= not (a xor b);
    layer0_outputs(779) <= not (a xor b);
    layer0_outputs(780) <= a;
    layer0_outputs(781) <= not (a or b);
    layer0_outputs(782) <= a;
    layer0_outputs(783) <= a or b;
    layer0_outputs(784) <= a and not b;
    layer0_outputs(785) <= b and not a;
    layer0_outputs(786) <= not a or b;
    layer0_outputs(787) <= not (a xor b);
    layer0_outputs(788) <= 1'b1;
    layer0_outputs(789) <= b;
    layer0_outputs(790) <= not a;
    layer0_outputs(791) <= not a or b;
    layer0_outputs(792) <= a and b;
    layer0_outputs(793) <= a or b;
    layer0_outputs(794) <= not b or a;
    layer0_outputs(795) <= a;
    layer0_outputs(796) <= not b;
    layer0_outputs(797) <= not (a and b);
    layer0_outputs(798) <= a and b;
    layer0_outputs(799) <= not a;
    layer0_outputs(800) <= a and not b;
    layer0_outputs(801) <= a xor b;
    layer0_outputs(802) <= 1'b1;
    layer0_outputs(803) <= b;
    layer0_outputs(804) <= b;
    layer0_outputs(805) <= a or b;
    layer0_outputs(806) <= b;
    layer0_outputs(807) <= not (a and b);
    layer0_outputs(808) <= b and not a;
    layer0_outputs(809) <= a or b;
    layer0_outputs(810) <= 1'b0;
    layer0_outputs(811) <= a or b;
    layer0_outputs(812) <= not a;
    layer0_outputs(813) <= not a;
    layer0_outputs(814) <= 1'b1;
    layer0_outputs(815) <= 1'b0;
    layer0_outputs(816) <= 1'b0;
    layer0_outputs(817) <= a;
    layer0_outputs(818) <= 1'b1;
    layer0_outputs(819) <= a and not b;
    layer0_outputs(820) <= a or b;
    layer0_outputs(821) <= a and not b;
    layer0_outputs(822) <= not a;
    layer0_outputs(823) <= a;
    layer0_outputs(824) <= a and b;
    layer0_outputs(825) <= not b or a;
    layer0_outputs(826) <= a and not b;
    layer0_outputs(827) <= 1'b0;
    layer0_outputs(828) <= not (a and b);
    layer0_outputs(829) <= not (a and b);
    layer0_outputs(830) <= b and not a;
    layer0_outputs(831) <= 1'b1;
    layer0_outputs(832) <= not b;
    layer0_outputs(833) <= not b or a;
    layer0_outputs(834) <= a;
    layer0_outputs(835) <= b;
    layer0_outputs(836) <= not (a xor b);
    layer0_outputs(837) <= 1'b0;
    layer0_outputs(838) <= a or b;
    layer0_outputs(839) <= not b or a;
    layer0_outputs(840) <= a and not b;
    layer0_outputs(841) <= not a or b;
    layer0_outputs(842) <= 1'b1;
    layer0_outputs(843) <= not b or a;
    layer0_outputs(844) <= not (a and b);
    layer0_outputs(845) <= 1'b1;
    layer0_outputs(846) <= a xor b;
    layer0_outputs(847) <= b and not a;
    layer0_outputs(848) <= a;
    layer0_outputs(849) <= a and b;
    layer0_outputs(850) <= a;
    layer0_outputs(851) <= a and b;
    layer0_outputs(852) <= 1'b0;
    layer0_outputs(853) <= a;
    layer0_outputs(854) <= a and b;
    layer0_outputs(855) <= a and not b;
    layer0_outputs(856) <= b and not a;
    layer0_outputs(857) <= not (a or b);
    layer0_outputs(858) <= 1'b1;
    layer0_outputs(859) <= b;
    layer0_outputs(860) <= not b;
    layer0_outputs(861) <= b;
    layer0_outputs(862) <= 1'b1;
    layer0_outputs(863) <= not b;
    layer0_outputs(864) <= 1'b1;
    layer0_outputs(865) <= not b or a;
    layer0_outputs(866) <= not b or a;
    layer0_outputs(867) <= a;
    layer0_outputs(868) <= 1'b1;
    layer0_outputs(869) <= 1'b1;
    layer0_outputs(870) <= a and not b;
    layer0_outputs(871) <= not b;
    layer0_outputs(872) <= a;
    layer0_outputs(873) <= not a or b;
    layer0_outputs(874) <= a and b;
    layer0_outputs(875) <= not b or a;
    layer0_outputs(876) <= not (a xor b);
    layer0_outputs(877) <= a xor b;
    layer0_outputs(878) <= 1'b0;
    layer0_outputs(879) <= not b or a;
    layer0_outputs(880) <= not a or b;
    layer0_outputs(881) <= not a;
    layer0_outputs(882) <= not (a or b);
    layer0_outputs(883) <= 1'b0;
    layer0_outputs(884) <= b and not a;
    layer0_outputs(885) <= not (a or b);
    layer0_outputs(886) <= not a;
    layer0_outputs(887) <= a and b;
    layer0_outputs(888) <= a xor b;
    layer0_outputs(889) <= not b or a;
    layer0_outputs(890) <= not a or b;
    layer0_outputs(891) <= not a;
    layer0_outputs(892) <= 1'b0;
    layer0_outputs(893) <= 1'b1;
    layer0_outputs(894) <= b;
    layer0_outputs(895) <= a xor b;
    layer0_outputs(896) <= b and not a;
    layer0_outputs(897) <= not b or a;
    layer0_outputs(898) <= a and not b;
    layer0_outputs(899) <= not b;
    layer0_outputs(900) <= 1'b0;
    layer0_outputs(901) <= a and not b;
    layer0_outputs(902) <= a xor b;
    layer0_outputs(903) <= 1'b0;
    layer0_outputs(904) <= 1'b1;
    layer0_outputs(905) <= a;
    layer0_outputs(906) <= not (a and b);
    layer0_outputs(907) <= a and b;
    layer0_outputs(908) <= not (a and b);
    layer0_outputs(909) <= not a or b;
    layer0_outputs(910) <= 1'b0;
    layer0_outputs(911) <= a;
    layer0_outputs(912) <= a and not b;
    layer0_outputs(913) <= not (a or b);
    layer0_outputs(914) <= a or b;
    layer0_outputs(915) <= b and not a;
    layer0_outputs(916) <= 1'b1;
    layer0_outputs(917) <= not (a and b);
    layer0_outputs(918) <= not a or b;
    layer0_outputs(919) <= not a or b;
    layer0_outputs(920) <= a;
    layer0_outputs(921) <= 1'b1;
    layer0_outputs(922) <= a and b;
    layer0_outputs(923) <= a;
    layer0_outputs(924) <= b and not a;
    layer0_outputs(925) <= not (a or b);
    layer0_outputs(926) <= not a;
    layer0_outputs(927) <= 1'b0;
    layer0_outputs(928) <= not (a xor b);
    layer0_outputs(929) <= a or b;
    layer0_outputs(930) <= 1'b1;
    layer0_outputs(931) <= not a or b;
    layer0_outputs(932) <= a and not b;
    layer0_outputs(933) <= b and not a;
    layer0_outputs(934) <= not (a xor b);
    layer0_outputs(935) <= b;
    layer0_outputs(936) <= b;
    layer0_outputs(937) <= not (a or b);
    layer0_outputs(938) <= not b or a;
    layer0_outputs(939) <= not b or a;
    layer0_outputs(940) <= 1'b1;
    layer0_outputs(941) <= not (a xor b);
    layer0_outputs(942) <= not b or a;
    layer0_outputs(943) <= b;
    layer0_outputs(944) <= not (a xor b);
    layer0_outputs(945) <= not b;
    layer0_outputs(946) <= 1'b0;
    layer0_outputs(947) <= a or b;
    layer0_outputs(948) <= not (a or b);
    layer0_outputs(949) <= b;
    layer0_outputs(950) <= 1'b0;
    layer0_outputs(951) <= a;
    layer0_outputs(952) <= 1'b0;
    layer0_outputs(953) <= b and not a;
    layer0_outputs(954) <= b and not a;
    layer0_outputs(955) <= a and b;
    layer0_outputs(956) <= not (a or b);
    layer0_outputs(957) <= a and not b;
    layer0_outputs(958) <= a;
    layer0_outputs(959) <= not (a and b);
    layer0_outputs(960) <= 1'b1;
    layer0_outputs(961) <= 1'b0;
    layer0_outputs(962) <= 1'b1;
    layer0_outputs(963) <= 1'b0;
    layer0_outputs(964) <= a xor b;
    layer0_outputs(965) <= 1'b0;
    layer0_outputs(966) <= not a or b;
    layer0_outputs(967) <= a;
    layer0_outputs(968) <= not (a and b);
    layer0_outputs(969) <= b;
    layer0_outputs(970) <= b and not a;
    layer0_outputs(971) <= a and b;
    layer0_outputs(972) <= not a;
    layer0_outputs(973) <= 1'b0;
    layer0_outputs(974) <= a xor b;
    layer0_outputs(975) <= not a or b;
    layer0_outputs(976) <= a;
    layer0_outputs(977) <= not a;
    layer0_outputs(978) <= a or b;
    layer0_outputs(979) <= not (a and b);
    layer0_outputs(980) <= not b or a;
    layer0_outputs(981) <= a xor b;
    layer0_outputs(982) <= b;
    layer0_outputs(983) <= not a;
    layer0_outputs(984) <= a and b;
    layer0_outputs(985) <= 1'b1;
    layer0_outputs(986) <= 1'b0;
    layer0_outputs(987) <= 1'b1;
    layer0_outputs(988) <= b;
    layer0_outputs(989) <= 1'b1;
    layer0_outputs(990) <= not a;
    layer0_outputs(991) <= a and not b;
    layer0_outputs(992) <= not b;
    layer0_outputs(993) <= not (a and b);
    layer0_outputs(994) <= a;
    layer0_outputs(995) <= not b;
    layer0_outputs(996) <= not (a xor b);
    layer0_outputs(997) <= 1'b1;
    layer0_outputs(998) <= not (a or b);
    layer0_outputs(999) <= a and not b;
    layer0_outputs(1000) <= b and not a;
    layer0_outputs(1001) <= b and not a;
    layer0_outputs(1002) <= not a;
    layer0_outputs(1003) <= a;
    layer0_outputs(1004) <= 1'b0;
    layer0_outputs(1005) <= b;
    layer0_outputs(1006) <= 1'b1;
    layer0_outputs(1007) <= a and b;
    layer0_outputs(1008) <= 1'b1;
    layer0_outputs(1009) <= a and not b;
    layer0_outputs(1010) <= a xor b;
    layer0_outputs(1011) <= not b or a;
    layer0_outputs(1012) <= 1'b1;
    layer0_outputs(1013) <= a;
    layer0_outputs(1014) <= a and not b;
    layer0_outputs(1015) <= 1'b0;
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= 1'b0;
    layer0_outputs(1018) <= not (a and b);
    layer0_outputs(1019) <= b and not a;
    layer0_outputs(1020) <= not (a or b);
    layer0_outputs(1021) <= a;
    layer0_outputs(1022) <= b and not a;
    layer0_outputs(1023) <= 1'b0;
    layer0_outputs(1024) <= a xor b;
    layer0_outputs(1025) <= a;
    layer0_outputs(1026) <= b and not a;
    layer0_outputs(1027) <= not b;
    layer0_outputs(1028) <= a or b;
    layer0_outputs(1029) <= a xor b;
    layer0_outputs(1030) <= a and not b;
    layer0_outputs(1031) <= 1'b1;
    layer0_outputs(1032) <= b and not a;
    layer0_outputs(1033) <= not (a xor b);
    layer0_outputs(1034) <= a;
    layer0_outputs(1035) <= a and b;
    layer0_outputs(1036) <= not a or b;
    layer0_outputs(1037) <= a and not b;
    layer0_outputs(1038) <= 1'b0;
    layer0_outputs(1039) <= a xor b;
    layer0_outputs(1040) <= b;
    layer0_outputs(1041) <= b;
    layer0_outputs(1042) <= a or b;
    layer0_outputs(1043) <= b;
    layer0_outputs(1044) <= not (a or b);
    layer0_outputs(1045) <= not b or a;
    layer0_outputs(1046) <= 1'b0;
    layer0_outputs(1047) <= a and b;
    layer0_outputs(1048) <= not (a and b);
    layer0_outputs(1049) <= b and not a;
    layer0_outputs(1050) <= b;
    layer0_outputs(1051) <= not b or a;
    layer0_outputs(1052) <= b;
    layer0_outputs(1053) <= a;
    layer0_outputs(1054) <= a and b;
    layer0_outputs(1055) <= not a;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= a or b;
    layer0_outputs(1058) <= not a;
    layer0_outputs(1059) <= 1'b1;
    layer0_outputs(1060) <= b and not a;
    layer0_outputs(1061) <= a or b;
    layer0_outputs(1062) <= a or b;
    layer0_outputs(1063) <= a and b;
    layer0_outputs(1064) <= b and not a;
    layer0_outputs(1065) <= not (a and b);
    layer0_outputs(1066) <= 1'b1;
    layer0_outputs(1067) <= not a or b;
    layer0_outputs(1068) <= a;
    layer0_outputs(1069) <= 1'b1;
    layer0_outputs(1070) <= a or b;
    layer0_outputs(1071) <= 1'b0;
    layer0_outputs(1072) <= a and not b;
    layer0_outputs(1073) <= b;
    layer0_outputs(1074) <= a and b;
    layer0_outputs(1075) <= not b or a;
    layer0_outputs(1076) <= not (a and b);
    layer0_outputs(1077) <= not (a xor b);
    layer0_outputs(1078) <= not a;
    layer0_outputs(1079) <= a and not b;
    layer0_outputs(1080) <= a or b;
    layer0_outputs(1081) <= a and b;
    layer0_outputs(1082) <= not a;
    layer0_outputs(1083) <= 1'b1;
    layer0_outputs(1084) <= not (a or b);
    layer0_outputs(1085) <= a;
    layer0_outputs(1086) <= not (a xor b);
    layer0_outputs(1087) <= 1'b0;
    layer0_outputs(1088) <= b and not a;
    layer0_outputs(1089) <= b and not a;
    layer0_outputs(1090) <= 1'b1;
    layer0_outputs(1091) <= not a or b;
    layer0_outputs(1092) <= a or b;
    layer0_outputs(1093) <= a;
    layer0_outputs(1094) <= a and not b;
    layer0_outputs(1095) <= a and not b;
    layer0_outputs(1096) <= a or b;
    layer0_outputs(1097) <= a;
    layer0_outputs(1098) <= not b or a;
    layer0_outputs(1099) <= a xor b;
    layer0_outputs(1100) <= not b or a;
    layer0_outputs(1101) <= 1'b0;
    layer0_outputs(1102) <= a or b;
    layer0_outputs(1103) <= a and not b;
    layer0_outputs(1104) <= not a;
    layer0_outputs(1105) <= b and not a;
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= a and b;
    layer0_outputs(1108) <= not a or b;
    layer0_outputs(1109) <= a xor b;
    layer0_outputs(1110) <= not (a or b);
    layer0_outputs(1111) <= not a;
    layer0_outputs(1112) <= not a or b;
    layer0_outputs(1113) <= not (a or b);
    layer0_outputs(1114) <= a and b;
    layer0_outputs(1115) <= not (a xor b);
    layer0_outputs(1116) <= not (a or b);
    layer0_outputs(1117) <= a and not b;
    layer0_outputs(1118) <= not a or b;
    layer0_outputs(1119) <= b and not a;
    layer0_outputs(1120) <= not (a and b);
    layer0_outputs(1121) <= b and not a;
    layer0_outputs(1122) <= a or b;
    layer0_outputs(1123) <= not a;
    layer0_outputs(1124) <= a;
    layer0_outputs(1125) <= a;
    layer0_outputs(1126) <= not a or b;
    layer0_outputs(1127) <= a or b;
    layer0_outputs(1128) <= b and not a;
    layer0_outputs(1129) <= not b or a;
    layer0_outputs(1130) <= a xor b;
    layer0_outputs(1131) <= not b;
    layer0_outputs(1132) <= b;
    layer0_outputs(1133) <= b and not a;
    layer0_outputs(1134) <= 1'b0;
    layer0_outputs(1135) <= not (a and b);
    layer0_outputs(1136) <= 1'b0;
    layer0_outputs(1137) <= not (a or b);
    layer0_outputs(1138) <= not a or b;
    layer0_outputs(1139) <= a;
    layer0_outputs(1140) <= not b;
    layer0_outputs(1141) <= not a or b;
    layer0_outputs(1142) <= not (a or b);
    layer0_outputs(1143) <= not b;
    layer0_outputs(1144) <= not (a and b);
    layer0_outputs(1145) <= a;
    layer0_outputs(1146) <= not b or a;
    layer0_outputs(1147) <= not (a or b);
    layer0_outputs(1148) <= not b;
    layer0_outputs(1149) <= not (a or b);
    layer0_outputs(1150) <= not (a or b);
    layer0_outputs(1151) <= a and not b;
    layer0_outputs(1152) <= a and b;
    layer0_outputs(1153) <= not b;
    layer0_outputs(1154) <= b;
    layer0_outputs(1155) <= a or b;
    layer0_outputs(1156) <= not b or a;
    layer0_outputs(1157) <= a and b;
    layer0_outputs(1158) <= b and not a;
    layer0_outputs(1159) <= b and not a;
    layer0_outputs(1160) <= 1'b0;
    layer0_outputs(1161) <= 1'b1;
    layer0_outputs(1162) <= a and b;
    layer0_outputs(1163) <= a xor b;
    layer0_outputs(1164) <= a xor b;
    layer0_outputs(1165) <= 1'b0;
    layer0_outputs(1166) <= not a;
    layer0_outputs(1167) <= a and not b;
    layer0_outputs(1168) <= a;
    layer0_outputs(1169) <= a or b;
    layer0_outputs(1170) <= not b;
    layer0_outputs(1171) <= 1'b0;
    layer0_outputs(1172) <= not b or a;
    layer0_outputs(1173) <= a and b;
    layer0_outputs(1174) <= a;
    layer0_outputs(1175) <= b;
    layer0_outputs(1176) <= not a;
    layer0_outputs(1177) <= b and not a;
    layer0_outputs(1178) <= b and not a;
    layer0_outputs(1179) <= not a or b;
    layer0_outputs(1180) <= not a or b;
    layer0_outputs(1181) <= not b;
    layer0_outputs(1182) <= a xor b;
    layer0_outputs(1183) <= 1'b0;
    layer0_outputs(1184) <= a or b;
    layer0_outputs(1185) <= not b or a;
    layer0_outputs(1186) <= 1'b1;
    layer0_outputs(1187) <= not a;
    layer0_outputs(1188) <= 1'b1;
    layer0_outputs(1189) <= not a or b;
    layer0_outputs(1190) <= a and b;
    layer0_outputs(1191) <= a xor b;
    layer0_outputs(1192) <= a and not b;
    layer0_outputs(1193) <= a;
    layer0_outputs(1194) <= not a or b;
    layer0_outputs(1195) <= a and not b;
    layer0_outputs(1196) <= not a;
    layer0_outputs(1197) <= not (a or b);
    layer0_outputs(1198) <= b and not a;
    layer0_outputs(1199) <= not (a and b);
    layer0_outputs(1200) <= not (a xor b);
    layer0_outputs(1201) <= not (a and b);
    layer0_outputs(1202) <= b;
    layer0_outputs(1203) <= b and not a;
    layer0_outputs(1204) <= a or b;
    layer0_outputs(1205) <= not b or a;
    layer0_outputs(1206) <= not (a or b);
    layer0_outputs(1207) <= 1'b0;
    layer0_outputs(1208) <= a and b;
    layer0_outputs(1209) <= a xor b;
    layer0_outputs(1210) <= not (a or b);
    layer0_outputs(1211) <= 1'b1;
    layer0_outputs(1212) <= a and b;
    layer0_outputs(1213) <= not a;
    layer0_outputs(1214) <= a;
    layer0_outputs(1215) <= not (a and b);
    layer0_outputs(1216) <= not (a or b);
    layer0_outputs(1217) <= not a;
    layer0_outputs(1218) <= a;
    layer0_outputs(1219) <= not b;
    layer0_outputs(1220) <= not a;
    layer0_outputs(1221) <= b;
    layer0_outputs(1222) <= a or b;
    layer0_outputs(1223) <= not a;
    layer0_outputs(1224) <= a and not b;
    layer0_outputs(1225) <= not b or a;
    layer0_outputs(1226) <= not a;
    layer0_outputs(1227) <= a xor b;
    layer0_outputs(1228) <= 1'b1;
    layer0_outputs(1229) <= a or b;
    layer0_outputs(1230) <= 1'b0;
    layer0_outputs(1231) <= a and not b;
    layer0_outputs(1232) <= 1'b0;
    layer0_outputs(1233) <= not a;
    layer0_outputs(1234) <= not b or a;
    layer0_outputs(1235) <= not a or b;
    layer0_outputs(1236) <= b and not a;
    layer0_outputs(1237) <= b;
    layer0_outputs(1238) <= a and not b;
    layer0_outputs(1239) <= a or b;
    layer0_outputs(1240) <= a xor b;
    layer0_outputs(1241) <= a xor b;
    layer0_outputs(1242) <= not (a xor b);
    layer0_outputs(1243) <= a or b;
    layer0_outputs(1244) <= not b or a;
    layer0_outputs(1245) <= a or b;
    layer0_outputs(1246) <= a and b;
    layer0_outputs(1247) <= 1'b1;
    layer0_outputs(1248) <= not a;
    layer0_outputs(1249) <= not (a or b);
    layer0_outputs(1250) <= a;
    layer0_outputs(1251) <= not b;
    layer0_outputs(1252) <= not (a xor b);
    layer0_outputs(1253) <= not b or a;
    layer0_outputs(1254) <= a and b;
    layer0_outputs(1255) <= 1'b1;
    layer0_outputs(1256) <= not (a and b);
    layer0_outputs(1257) <= not (a and b);
    layer0_outputs(1258) <= not (a or b);
    layer0_outputs(1259) <= b;
    layer0_outputs(1260) <= not b or a;
    layer0_outputs(1261) <= not (a xor b);
    layer0_outputs(1262) <= not a or b;
    layer0_outputs(1263) <= not b or a;
    layer0_outputs(1264) <= not a;
    layer0_outputs(1265) <= not b or a;
    layer0_outputs(1266) <= a;
    layer0_outputs(1267) <= a xor b;
    layer0_outputs(1268) <= b and not a;
    layer0_outputs(1269) <= 1'b1;
    layer0_outputs(1270) <= b and not a;
    layer0_outputs(1271) <= b;
    layer0_outputs(1272) <= not a or b;
    layer0_outputs(1273) <= not a;
    layer0_outputs(1274) <= not a or b;
    layer0_outputs(1275) <= not a;
    layer0_outputs(1276) <= not (a xor b);
    layer0_outputs(1277) <= not (a or b);
    layer0_outputs(1278) <= not (a or b);
    layer0_outputs(1279) <= not b;
    layer0_outputs(1280) <= a and not b;
    layer0_outputs(1281) <= b;
    layer0_outputs(1282) <= a and not b;
    layer0_outputs(1283) <= not b;
    layer0_outputs(1284) <= not (a xor b);
    layer0_outputs(1285) <= b;
    layer0_outputs(1286) <= not a or b;
    layer0_outputs(1287) <= 1'b0;
    layer0_outputs(1288) <= not a;
    layer0_outputs(1289) <= b and not a;
    layer0_outputs(1290) <= a and b;
    layer0_outputs(1291) <= a and b;
    layer0_outputs(1292) <= 1'b0;
    layer0_outputs(1293) <= b;
    layer0_outputs(1294) <= a or b;
    layer0_outputs(1295) <= not b or a;
    layer0_outputs(1296) <= not (a and b);
    layer0_outputs(1297) <= not a or b;
    layer0_outputs(1298) <= b;
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= 1'b0;
    layer0_outputs(1301) <= 1'b1;
    layer0_outputs(1302) <= a or b;
    layer0_outputs(1303) <= not a or b;
    layer0_outputs(1304) <= not (a and b);
    layer0_outputs(1305) <= not (a xor b);
    layer0_outputs(1306) <= not b or a;
    layer0_outputs(1307) <= not b;
    layer0_outputs(1308) <= a and b;
    layer0_outputs(1309) <= a or b;
    layer0_outputs(1310) <= 1'b0;
    layer0_outputs(1311) <= b;
    layer0_outputs(1312) <= not (a and b);
    layer0_outputs(1313) <= not a or b;
    layer0_outputs(1314) <= a or b;
    layer0_outputs(1315) <= b;
    layer0_outputs(1316) <= not a or b;
    layer0_outputs(1317) <= b;
    layer0_outputs(1318) <= b;
    layer0_outputs(1319) <= a and b;
    layer0_outputs(1320) <= b;
    layer0_outputs(1321) <= 1'b0;
    layer0_outputs(1322) <= a xor b;
    layer0_outputs(1323) <= 1'b1;
    layer0_outputs(1324) <= 1'b1;
    layer0_outputs(1325) <= 1'b1;
    layer0_outputs(1326) <= a or b;
    layer0_outputs(1327) <= not a;
    layer0_outputs(1328) <= not (a or b);
    layer0_outputs(1329) <= not (a or b);
    layer0_outputs(1330) <= b;
    layer0_outputs(1331) <= a and not b;
    layer0_outputs(1332) <= a and not b;
    layer0_outputs(1333) <= not b or a;
    layer0_outputs(1334) <= 1'b0;
    layer0_outputs(1335) <= 1'b0;
    layer0_outputs(1336) <= not b;
    layer0_outputs(1337) <= b;
    layer0_outputs(1338) <= a and b;
    layer0_outputs(1339) <= not b or a;
    layer0_outputs(1340) <= not (a xor b);
    layer0_outputs(1341) <= b and not a;
    layer0_outputs(1342) <= a and b;
    layer0_outputs(1343) <= not b or a;
    layer0_outputs(1344) <= b and not a;
    layer0_outputs(1345) <= not a;
    layer0_outputs(1346) <= not (a and b);
    layer0_outputs(1347) <= 1'b0;
    layer0_outputs(1348) <= not b or a;
    layer0_outputs(1349) <= b and not a;
    layer0_outputs(1350) <= not a or b;
    layer0_outputs(1351) <= b and not a;
    layer0_outputs(1352) <= not (a xor b);
    layer0_outputs(1353) <= not a;
    layer0_outputs(1354) <= not b;
    layer0_outputs(1355) <= 1'b0;
    layer0_outputs(1356) <= not a or b;
    layer0_outputs(1357) <= a or b;
    layer0_outputs(1358) <= not (a xor b);
    layer0_outputs(1359) <= not a;
    layer0_outputs(1360) <= not (a or b);
    layer0_outputs(1361) <= a and b;
    layer0_outputs(1362) <= a or b;
    layer0_outputs(1363) <= b and not a;
    layer0_outputs(1364) <= b;
    layer0_outputs(1365) <= not b;
    layer0_outputs(1366) <= not b;
    layer0_outputs(1367) <= b and not a;
    layer0_outputs(1368) <= not a;
    layer0_outputs(1369) <= a xor b;
    layer0_outputs(1370) <= not a or b;
    layer0_outputs(1371) <= b and not a;
    layer0_outputs(1372) <= a;
    layer0_outputs(1373) <= not (a or b);
    layer0_outputs(1374) <= a and b;
    layer0_outputs(1375) <= not b;
    layer0_outputs(1376) <= a or b;
    layer0_outputs(1377) <= not b;
    layer0_outputs(1378) <= a or b;
    layer0_outputs(1379) <= b and not a;
    layer0_outputs(1380) <= b;
    layer0_outputs(1381) <= a or b;
    layer0_outputs(1382) <= 1'b0;
    layer0_outputs(1383) <= 1'b1;
    layer0_outputs(1384) <= not b or a;
    layer0_outputs(1385) <= not b or a;
    layer0_outputs(1386) <= not b;
    layer0_outputs(1387) <= b and not a;
    layer0_outputs(1388) <= 1'b1;
    layer0_outputs(1389) <= a;
    layer0_outputs(1390) <= not (a xor b);
    layer0_outputs(1391) <= not (a or b);
    layer0_outputs(1392) <= not (a or b);
    layer0_outputs(1393) <= 1'b1;
    layer0_outputs(1394) <= a and b;
    layer0_outputs(1395) <= not (a xor b);
    layer0_outputs(1396) <= 1'b1;
    layer0_outputs(1397) <= not b;
    layer0_outputs(1398) <= b and not a;
    layer0_outputs(1399) <= a or b;
    layer0_outputs(1400) <= a xor b;
    layer0_outputs(1401) <= 1'b0;
    layer0_outputs(1402) <= 1'b0;
    layer0_outputs(1403) <= b;
    layer0_outputs(1404) <= not b;
    layer0_outputs(1405) <= not (a xor b);
    layer0_outputs(1406) <= a and not b;
    layer0_outputs(1407) <= not (a and b);
    layer0_outputs(1408) <= a and not b;
    layer0_outputs(1409) <= 1'b1;
    layer0_outputs(1410) <= 1'b1;
    layer0_outputs(1411) <= a or b;
    layer0_outputs(1412) <= 1'b1;
    layer0_outputs(1413) <= b and not a;
    layer0_outputs(1414) <= a xor b;
    layer0_outputs(1415) <= b;
    layer0_outputs(1416) <= not a or b;
    layer0_outputs(1417) <= 1'b1;
    layer0_outputs(1418) <= b and not a;
    layer0_outputs(1419) <= not a or b;
    layer0_outputs(1420) <= a;
    layer0_outputs(1421) <= b and not a;
    layer0_outputs(1422) <= not b;
    layer0_outputs(1423) <= b;
    layer0_outputs(1424) <= not (a or b);
    layer0_outputs(1425) <= not a or b;
    layer0_outputs(1426) <= b and not a;
    layer0_outputs(1427) <= 1'b0;
    layer0_outputs(1428) <= b;
    layer0_outputs(1429) <= not (a and b);
    layer0_outputs(1430) <= not a or b;
    layer0_outputs(1431) <= a or b;
    layer0_outputs(1432) <= b;
    layer0_outputs(1433) <= not (a and b);
    layer0_outputs(1434) <= not a;
    layer0_outputs(1435) <= not (a or b);
    layer0_outputs(1436) <= a and not b;
    layer0_outputs(1437) <= 1'b1;
    layer0_outputs(1438) <= not a or b;
    layer0_outputs(1439) <= not (a or b);
    layer0_outputs(1440) <= a and b;
    layer0_outputs(1441) <= b and not a;
    layer0_outputs(1442) <= not a;
    layer0_outputs(1443) <= b;
    layer0_outputs(1444) <= not a;
    layer0_outputs(1445) <= not (a and b);
    layer0_outputs(1446) <= not (a xor b);
    layer0_outputs(1447) <= a and not b;
    layer0_outputs(1448) <= not a;
    layer0_outputs(1449) <= not b or a;
    layer0_outputs(1450) <= not b;
    layer0_outputs(1451) <= a xor b;
    layer0_outputs(1452) <= a and b;
    layer0_outputs(1453) <= a or b;
    layer0_outputs(1454) <= b;
    layer0_outputs(1455) <= a and b;
    layer0_outputs(1456) <= b;
    layer0_outputs(1457) <= 1'b0;
    layer0_outputs(1458) <= 1'b1;
    layer0_outputs(1459) <= a and not b;
    layer0_outputs(1460) <= a and b;
    layer0_outputs(1461) <= a and b;
    layer0_outputs(1462) <= not (a and b);
    layer0_outputs(1463) <= 1'b1;
    layer0_outputs(1464) <= a;
    layer0_outputs(1465) <= a and b;
    layer0_outputs(1466) <= b and not a;
    layer0_outputs(1467) <= not (a or b);
    layer0_outputs(1468) <= 1'b1;
    layer0_outputs(1469) <= not b;
    layer0_outputs(1470) <= 1'b1;
    layer0_outputs(1471) <= 1'b0;
    layer0_outputs(1472) <= not b or a;
    layer0_outputs(1473) <= b;
    layer0_outputs(1474) <= a;
    layer0_outputs(1475) <= not (a or b);
    layer0_outputs(1476) <= a or b;
    layer0_outputs(1477) <= not (a xor b);
    layer0_outputs(1478) <= 1'b1;
    layer0_outputs(1479) <= not a;
    layer0_outputs(1480) <= not b or a;
    layer0_outputs(1481) <= not b or a;
    layer0_outputs(1482) <= not a or b;
    layer0_outputs(1483) <= not (a xor b);
    layer0_outputs(1484) <= not b;
    layer0_outputs(1485) <= a and b;
    layer0_outputs(1486) <= b;
    layer0_outputs(1487) <= a;
    layer0_outputs(1488) <= a and b;
    layer0_outputs(1489) <= not (a or b);
    layer0_outputs(1490) <= not (a and b);
    layer0_outputs(1491) <= not b;
    layer0_outputs(1492) <= a xor b;
    layer0_outputs(1493) <= not (a and b);
    layer0_outputs(1494) <= a and b;
    layer0_outputs(1495) <= not (a and b);
    layer0_outputs(1496) <= not a or b;
    layer0_outputs(1497) <= a;
    layer0_outputs(1498) <= not (a xor b);
    layer0_outputs(1499) <= not b or a;
    layer0_outputs(1500) <= not b or a;
    layer0_outputs(1501) <= b and not a;
    layer0_outputs(1502) <= b and not a;
    layer0_outputs(1503) <= a xor b;
    layer0_outputs(1504) <= a and b;
    layer0_outputs(1505) <= a xor b;
    layer0_outputs(1506) <= not a or b;
    layer0_outputs(1507) <= not (a or b);
    layer0_outputs(1508) <= not b or a;
    layer0_outputs(1509) <= b;
    layer0_outputs(1510) <= not a;
    layer0_outputs(1511) <= a and b;
    layer0_outputs(1512) <= b and not a;
    layer0_outputs(1513) <= a and b;
    layer0_outputs(1514) <= b and not a;
    layer0_outputs(1515) <= not a;
    layer0_outputs(1516) <= a;
    layer0_outputs(1517) <= not (a and b);
    layer0_outputs(1518) <= not (a or b);
    layer0_outputs(1519) <= b;
    layer0_outputs(1520) <= not (a xor b);
    layer0_outputs(1521) <= a xor b;
    layer0_outputs(1522) <= not a or b;
    layer0_outputs(1523) <= a xor b;
    layer0_outputs(1524) <= b and not a;
    layer0_outputs(1525) <= not (a and b);
    layer0_outputs(1526) <= b;
    layer0_outputs(1527) <= not a or b;
    layer0_outputs(1528) <= not a;
    layer0_outputs(1529) <= a;
    layer0_outputs(1530) <= 1'b1;
    layer0_outputs(1531) <= b and not a;
    layer0_outputs(1532) <= not b or a;
    layer0_outputs(1533) <= not (a or b);
    layer0_outputs(1534) <= a and not b;
    layer0_outputs(1535) <= b;
    layer0_outputs(1536) <= a and b;
    layer0_outputs(1537) <= not a or b;
    layer0_outputs(1538) <= not a or b;
    layer0_outputs(1539) <= a;
    layer0_outputs(1540) <= a and not b;
    layer0_outputs(1541) <= not (a or b);
    layer0_outputs(1542) <= a or b;
    layer0_outputs(1543) <= 1'b1;
    layer0_outputs(1544) <= not b;
    layer0_outputs(1545) <= a and not b;
    layer0_outputs(1546) <= b;
    layer0_outputs(1547) <= not b;
    layer0_outputs(1548) <= b;
    layer0_outputs(1549) <= not b or a;
    layer0_outputs(1550) <= not b or a;
    layer0_outputs(1551) <= not b;
    layer0_outputs(1552) <= 1'b0;
    layer0_outputs(1553) <= 1'b0;
    layer0_outputs(1554) <= 1'b1;
    layer0_outputs(1555) <= a and b;
    layer0_outputs(1556) <= not b;
    layer0_outputs(1557) <= not (a or b);
    layer0_outputs(1558) <= not (a xor b);
    layer0_outputs(1559) <= a and not b;
    layer0_outputs(1560) <= not b or a;
    layer0_outputs(1561) <= not b or a;
    layer0_outputs(1562) <= not a;
    layer0_outputs(1563) <= a and not b;
    layer0_outputs(1564) <= not a or b;
    layer0_outputs(1565) <= b and not a;
    layer0_outputs(1566) <= not (a xor b);
    layer0_outputs(1567) <= b;
    layer0_outputs(1568) <= a or b;
    layer0_outputs(1569) <= 1'b0;
    layer0_outputs(1570) <= not a or b;
    layer0_outputs(1571) <= b;
    layer0_outputs(1572) <= a;
    layer0_outputs(1573) <= not a or b;
    layer0_outputs(1574) <= not b;
    layer0_outputs(1575) <= a and b;
    layer0_outputs(1576) <= not b or a;
    layer0_outputs(1577) <= not a;
    layer0_outputs(1578) <= a;
    layer0_outputs(1579) <= not (a xor b);
    layer0_outputs(1580) <= b;
    layer0_outputs(1581) <= not b;
    layer0_outputs(1582) <= b and not a;
    layer0_outputs(1583) <= not a or b;
    layer0_outputs(1584) <= a and b;
    layer0_outputs(1585) <= b and not a;
    layer0_outputs(1586) <= not (a or b);
    layer0_outputs(1587) <= a;
    layer0_outputs(1588) <= not a or b;
    layer0_outputs(1589) <= not (a xor b);
    layer0_outputs(1590) <= a;
    layer0_outputs(1591) <= a;
    layer0_outputs(1592) <= not (a xor b);
    layer0_outputs(1593) <= not b;
    layer0_outputs(1594) <= b and not a;
    layer0_outputs(1595) <= a or b;
    layer0_outputs(1596) <= 1'b1;
    layer0_outputs(1597) <= b and not a;
    layer0_outputs(1598) <= b and not a;
    layer0_outputs(1599) <= not b;
    layer0_outputs(1600) <= 1'b1;
    layer0_outputs(1601) <= not (a xor b);
    layer0_outputs(1602) <= not a;
    layer0_outputs(1603) <= not b or a;
    layer0_outputs(1604) <= b;
    layer0_outputs(1605) <= a;
    layer0_outputs(1606) <= not a or b;
    layer0_outputs(1607) <= a and not b;
    layer0_outputs(1608) <= not (a and b);
    layer0_outputs(1609) <= a and b;
    layer0_outputs(1610) <= a and b;
    layer0_outputs(1611) <= not b;
    layer0_outputs(1612) <= a and not b;
    layer0_outputs(1613) <= b and not a;
    layer0_outputs(1614) <= 1'b0;
    layer0_outputs(1615) <= not b;
    layer0_outputs(1616) <= not b;
    layer0_outputs(1617) <= a and b;
    layer0_outputs(1618) <= not (a and b);
    layer0_outputs(1619) <= not a or b;
    layer0_outputs(1620) <= not (a or b);
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= b and not a;
    layer0_outputs(1623) <= not a or b;
    layer0_outputs(1624) <= not (a or b);
    layer0_outputs(1625) <= not b;
    layer0_outputs(1626) <= 1'b1;
    layer0_outputs(1627) <= a and b;
    layer0_outputs(1628) <= not b or a;
    layer0_outputs(1629) <= b and not a;
    layer0_outputs(1630) <= not (a or b);
    layer0_outputs(1631) <= b;
    layer0_outputs(1632) <= a and not b;
    layer0_outputs(1633) <= not (a and b);
    layer0_outputs(1634) <= b;
    layer0_outputs(1635) <= 1'b1;
    layer0_outputs(1636) <= 1'b0;
    layer0_outputs(1637) <= a or b;
    layer0_outputs(1638) <= b and not a;
    layer0_outputs(1639) <= not (a or b);
    layer0_outputs(1640) <= not b;
    layer0_outputs(1641) <= a xor b;
    layer0_outputs(1642) <= not (a xor b);
    layer0_outputs(1643) <= a;
    layer0_outputs(1644) <= not (a and b);
    layer0_outputs(1645) <= a and b;
    layer0_outputs(1646) <= not b or a;
    layer0_outputs(1647) <= not b or a;
    layer0_outputs(1648) <= a;
    layer0_outputs(1649) <= a or b;
    layer0_outputs(1650) <= not (a and b);
    layer0_outputs(1651) <= 1'b1;
    layer0_outputs(1652) <= a and b;
    layer0_outputs(1653) <= b;
    layer0_outputs(1654) <= a;
    layer0_outputs(1655) <= not a or b;
    layer0_outputs(1656) <= b and not a;
    layer0_outputs(1657) <= not b;
    layer0_outputs(1658) <= b and not a;
    layer0_outputs(1659) <= not (a and b);
    layer0_outputs(1660) <= not (a xor b);
    layer0_outputs(1661) <= a xor b;
    layer0_outputs(1662) <= not b or a;
    layer0_outputs(1663) <= a;
    layer0_outputs(1664) <= a;
    layer0_outputs(1665) <= a and b;
    layer0_outputs(1666) <= not (a and b);
    layer0_outputs(1667) <= a and b;
    layer0_outputs(1668) <= b and not a;
    layer0_outputs(1669) <= a or b;
    layer0_outputs(1670) <= a;
    layer0_outputs(1671) <= a and b;
    layer0_outputs(1672) <= not b;
    layer0_outputs(1673) <= a;
    layer0_outputs(1674) <= not (a or b);
    layer0_outputs(1675) <= a or b;
    layer0_outputs(1676) <= a and b;
    layer0_outputs(1677) <= not a or b;
    layer0_outputs(1678) <= not b or a;
    layer0_outputs(1679) <= 1'b0;
    layer0_outputs(1680) <= not b;
    layer0_outputs(1681) <= not (a and b);
    layer0_outputs(1682) <= b;
    layer0_outputs(1683) <= b and not a;
    layer0_outputs(1684) <= a and not b;
    layer0_outputs(1685) <= not (a and b);
    layer0_outputs(1686) <= a;
    layer0_outputs(1687) <= not a or b;
    layer0_outputs(1688) <= a xor b;
    layer0_outputs(1689) <= b;
    layer0_outputs(1690) <= 1'b1;
    layer0_outputs(1691) <= 1'b0;
    layer0_outputs(1692) <= 1'b0;
    layer0_outputs(1693) <= a and not b;
    layer0_outputs(1694) <= a xor b;
    layer0_outputs(1695) <= not (a xor b);
    layer0_outputs(1696) <= not (a and b);
    layer0_outputs(1697) <= not (a xor b);
    layer0_outputs(1698) <= b and not a;
    layer0_outputs(1699) <= a or b;
    layer0_outputs(1700) <= a;
    layer0_outputs(1701) <= not a or b;
    layer0_outputs(1702) <= not (a or b);
    layer0_outputs(1703) <= a or b;
    layer0_outputs(1704) <= b;
    layer0_outputs(1705) <= 1'b0;
    layer0_outputs(1706) <= a;
    layer0_outputs(1707) <= not a;
    layer0_outputs(1708) <= 1'b0;
    layer0_outputs(1709) <= a xor b;
    layer0_outputs(1710) <= not a;
    layer0_outputs(1711) <= not b or a;
    layer0_outputs(1712) <= a;
    layer0_outputs(1713) <= a or b;
    layer0_outputs(1714) <= not (a xor b);
    layer0_outputs(1715) <= not a or b;
    layer0_outputs(1716) <= not (a and b);
    layer0_outputs(1717) <= a or b;
    layer0_outputs(1718) <= not a;
    layer0_outputs(1719) <= b and not a;
    layer0_outputs(1720) <= 1'b1;
    layer0_outputs(1721) <= 1'b0;
    layer0_outputs(1722) <= 1'b1;
    layer0_outputs(1723) <= a xor b;
    layer0_outputs(1724) <= a xor b;
    layer0_outputs(1725) <= b and not a;
    layer0_outputs(1726) <= not b;
    layer0_outputs(1727) <= not (a or b);
    layer0_outputs(1728) <= not a or b;
    layer0_outputs(1729) <= a xor b;
    layer0_outputs(1730) <= a and b;
    layer0_outputs(1731) <= a and not b;
    layer0_outputs(1732) <= not (a and b);
    layer0_outputs(1733) <= not a or b;
    layer0_outputs(1734) <= a and not b;
    layer0_outputs(1735) <= 1'b1;
    layer0_outputs(1736) <= a;
    layer0_outputs(1737) <= not a;
    layer0_outputs(1738) <= not (a xor b);
    layer0_outputs(1739) <= b;
    layer0_outputs(1740) <= not a;
    layer0_outputs(1741) <= not (a or b);
    layer0_outputs(1742) <= not (a xor b);
    layer0_outputs(1743) <= not (a and b);
    layer0_outputs(1744) <= b and not a;
    layer0_outputs(1745) <= b;
    layer0_outputs(1746) <= not (a and b);
    layer0_outputs(1747) <= b;
    layer0_outputs(1748) <= not a or b;
    layer0_outputs(1749) <= 1'b0;
    layer0_outputs(1750) <= not (a and b);
    layer0_outputs(1751) <= not (a and b);
    layer0_outputs(1752) <= 1'b0;
    layer0_outputs(1753) <= not a;
    layer0_outputs(1754) <= b;
    layer0_outputs(1755) <= a and b;
    layer0_outputs(1756) <= a;
    layer0_outputs(1757) <= b and not a;
    layer0_outputs(1758) <= b;
    layer0_outputs(1759) <= not a or b;
    layer0_outputs(1760) <= a;
    layer0_outputs(1761) <= not b;
    layer0_outputs(1762) <= not (a xor b);
    layer0_outputs(1763) <= a xor b;
    layer0_outputs(1764) <= not a;
    layer0_outputs(1765) <= a;
    layer0_outputs(1766) <= not a or b;
    layer0_outputs(1767) <= a;
    layer0_outputs(1768) <= b;
    layer0_outputs(1769) <= not a or b;
    layer0_outputs(1770) <= b;
    layer0_outputs(1771) <= 1'b1;
    layer0_outputs(1772) <= a;
    layer0_outputs(1773) <= not a;
    layer0_outputs(1774) <= not (a xor b);
    layer0_outputs(1775) <= not a or b;
    layer0_outputs(1776) <= not a;
    layer0_outputs(1777) <= not (a and b);
    layer0_outputs(1778) <= b;
    layer0_outputs(1779) <= b;
    layer0_outputs(1780) <= b and not a;
    layer0_outputs(1781) <= not (a xor b);
    layer0_outputs(1782) <= a and b;
    layer0_outputs(1783) <= a;
    layer0_outputs(1784) <= not a or b;
    layer0_outputs(1785) <= b and not a;
    layer0_outputs(1786) <= not (a and b);
    layer0_outputs(1787) <= a and b;
    layer0_outputs(1788) <= 1'b1;
    layer0_outputs(1789) <= b and not a;
    layer0_outputs(1790) <= a or b;
    layer0_outputs(1791) <= not a;
    layer0_outputs(1792) <= 1'b0;
    layer0_outputs(1793) <= a;
    layer0_outputs(1794) <= not b;
    layer0_outputs(1795) <= not a;
    layer0_outputs(1796) <= a;
    layer0_outputs(1797) <= 1'b1;
    layer0_outputs(1798) <= not (a or b);
    layer0_outputs(1799) <= a and b;
    layer0_outputs(1800) <= not a;
    layer0_outputs(1801) <= b and not a;
    layer0_outputs(1802) <= a;
    layer0_outputs(1803) <= a xor b;
    layer0_outputs(1804) <= not b;
    layer0_outputs(1805) <= not a;
    layer0_outputs(1806) <= a;
    layer0_outputs(1807) <= a or b;
    layer0_outputs(1808) <= 1'b1;
    layer0_outputs(1809) <= not a or b;
    layer0_outputs(1810) <= not (a xor b);
    layer0_outputs(1811) <= not a;
    layer0_outputs(1812) <= not (a or b);
    layer0_outputs(1813) <= 1'b1;
    layer0_outputs(1814) <= not b or a;
    layer0_outputs(1815) <= a or b;
    layer0_outputs(1816) <= 1'b1;
    layer0_outputs(1817) <= 1'b0;
    layer0_outputs(1818) <= a;
    layer0_outputs(1819) <= not (a xor b);
    layer0_outputs(1820) <= not (a and b);
    layer0_outputs(1821) <= a;
    layer0_outputs(1822) <= not b or a;
    layer0_outputs(1823) <= not (a and b);
    layer0_outputs(1824) <= not b;
    layer0_outputs(1825) <= a and not b;
    layer0_outputs(1826) <= not b;
    layer0_outputs(1827) <= not b;
    layer0_outputs(1828) <= a and not b;
    layer0_outputs(1829) <= not (a xor b);
    layer0_outputs(1830) <= a and not b;
    layer0_outputs(1831) <= 1'b0;
    layer0_outputs(1832) <= not (a xor b);
    layer0_outputs(1833) <= not a or b;
    layer0_outputs(1834) <= a xor b;
    layer0_outputs(1835) <= not (a or b);
    layer0_outputs(1836) <= not b or a;
    layer0_outputs(1837) <= not b or a;
    layer0_outputs(1838) <= b;
    layer0_outputs(1839) <= b;
    layer0_outputs(1840) <= a xor b;
    layer0_outputs(1841) <= not b;
    layer0_outputs(1842) <= not (a xor b);
    layer0_outputs(1843) <= b and not a;
    layer0_outputs(1844) <= not (a and b);
    layer0_outputs(1845) <= b;
    layer0_outputs(1846) <= a or b;
    layer0_outputs(1847) <= 1'b1;
    layer0_outputs(1848) <= not (a and b);
    layer0_outputs(1849) <= a xor b;
    layer0_outputs(1850) <= a and b;
    layer0_outputs(1851) <= b and not a;
    layer0_outputs(1852) <= 1'b0;
    layer0_outputs(1853) <= not b or a;
    layer0_outputs(1854) <= a and b;
    layer0_outputs(1855) <= not b;
    layer0_outputs(1856) <= not (a xor b);
    layer0_outputs(1857) <= a and not b;
    layer0_outputs(1858) <= a and not b;
    layer0_outputs(1859) <= a and b;
    layer0_outputs(1860) <= a and b;
    layer0_outputs(1861) <= not (a or b);
    layer0_outputs(1862) <= a xor b;
    layer0_outputs(1863) <= a or b;
    layer0_outputs(1864) <= not (a and b);
    layer0_outputs(1865) <= not b;
    layer0_outputs(1866) <= a and b;
    layer0_outputs(1867) <= b;
    layer0_outputs(1868) <= 1'b0;
    layer0_outputs(1869) <= not (a xor b);
    layer0_outputs(1870) <= b;
    layer0_outputs(1871) <= a and not b;
    layer0_outputs(1872) <= 1'b0;
    layer0_outputs(1873) <= a xor b;
    layer0_outputs(1874) <= not (a or b);
    layer0_outputs(1875) <= b;
    layer0_outputs(1876) <= b and not a;
    layer0_outputs(1877) <= 1'b0;
    layer0_outputs(1878) <= 1'b0;
    layer0_outputs(1879) <= 1'b1;
    layer0_outputs(1880) <= not (a or b);
    layer0_outputs(1881) <= 1'b1;
    layer0_outputs(1882) <= b;
    layer0_outputs(1883) <= b;
    layer0_outputs(1884) <= not a;
    layer0_outputs(1885) <= a or b;
    layer0_outputs(1886) <= a and not b;
    layer0_outputs(1887) <= not a or b;
    layer0_outputs(1888) <= a;
    layer0_outputs(1889) <= 1'b1;
    layer0_outputs(1890) <= b;
    layer0_outputs(1891) <= not b;
    layer0_outputs(1892) <= not b or a;
    layer0_outputs(1893) <= a or b;
    layer0_outputs(1894) <= not b;
    layer0_outputs(1895) <= a and b;
    layer0_outputs(1896) <= not b;
    layer0_outputs(1897) <= b;
    layer0_outputs(1898) <= not a or b;
    layer0_outputs(1899) <= not b;
    layer0_outputs(1900) <= 1'b1;
    layer0_outputs(1901) <= 1'b0;
    layer0_outputs(1902) <= not b;
    layer0_outputs(1903) <= not b;
    layer0_outputs(1904) <= b and not a;
    layer0_outputs(1905) <= not b or a;
    layer0_outputs(1906) <= a and not b;
    layer0_outputs(1907) <= not b or a;
    layer0_outputs(1908) <= a and not b;
    layer0_outputs(1909) <= not (a and b);
    layer0_outputs(1910) <= not b or a;
    layer0_outputs(1911) <= a;
    layer0_outputs(1912) <= not a or b;
    layer0_outputs(1913) <= a xor b;
    layer0_outputs(1914) <= a and b;
    layer0_outputs(1915) <= a xor b;
    layer0_outputs(1916) <= not (a or b);
    layer0_outputs(1917) <= not a or b;
    layer0_outputs(1918) <= a xor b;
    layer0_outputs(1919) <= not a or b;
    layer0_outputs(1920) <= a and b;
    layer0_outputs(1921) <= not b;
    layer0_outputs(1922) <= not b;
    layer0_outputs(1923) <= not (a and b);
    layer0_outputs(1924) <= a or b;
    layer0_outputs(1925) <= not a;
    layer0_outputs(1926) <= a;
    layer0_outputs(1927) <= 1'b0;
    layer0_outputs(1928) <= 1'b1;
    layer0_outputs(1929) <= a and b;
    layer0_outputs(1930) <= not (a and b);
    layer0_outputs(1931) <= 1'b1;
    layer0_outputs(1932) <= not (a and b);
    layer0_outputs(1933) <= not b;
    layer0_outputs(1934) <= 1'b1;
    layer0_outputs(1935) <= 1'b0;
    layer0_outputs(1936) <= not (a and b);
    layer0_outputs(1937) <= 1'b0;
    layer0_outputs(1938) <= not (a and b);
    layer0_outputs(1939) <= a and not b;
    layer0_outputs(1940) <= 1'b0;
    layer0_outputs(1941) <= b;
    layer0_outputs(1942) <= 1'b1;
    layer0_outputs(1943) <= a xor b;
    layer0_outputs(1944) <= 1'b0;
    layer0_outputs(1945) <= a xor b;
    layer0_outputs(1946) <= not (a or b);
    layer0_outputs(1947) <= not b or a;
    layer0_outputs(1948) <= not (a and b);
    layer0_outputs(1949) <= 1'b0;
    layer0_outputs(1950) <= a and b;
    layer0_outputs(1951) <= 1'b0;
    layer0_outputs(1952) <= a and not b;
    layer0_outputs(1953) <= 1'b1;
    layer0_outputs(1954) <= not b or a;
    layer0_outputs(1955) <= a xor b;
    layer0_outputs(1956) <= 1'b1;
    layer0_outputs(1957) <= 1'b0;
    layer0_outputs(1958) <= 1'b1;
    layer0_outputs(1959) <= 1'b0;
    layer0_outputs(1960) <= b;
    layer0_outputs(1961) <= 1'b0;
    layer0_outputs(1962) <= a or b;
    layer0_outputs(1963) <= 1'b0;
    layer0_outputs(1964) <= not a;
    layer0_outputs(1965) <= b and not a;
    layer0_outputs(1966) <= b and not a;
    layer0_outputs(1967) <= not a or b;
    layer0_outputs(1968) <= b;
    layer0_outputs(1969) <= a;
    layer0_outputs(1970) <= b and not a;
    layer0_outputs(1971) <= 1'b1;
    layer0_outputs(1972) <= not b or a;
    layer0_outputs(1973) <= not (a xor b);
    layer0_outputs(1974) <= a and not b;
    layer0_outputs(1975) <= not (a and b);
    layer0_outputs(1976) <= a or b;
    layer0_outputs(1977) <= 1'b1;
    layer0_outputs(1978) <= not a;
    layer0_outputs(1979) <= not (a and b);
    layer0_outputs(1980) <= a and b;
    layer0_outputs(1981) <= a and b;
    layer0_outputs(1982) <= 1'b1;
    layer0_outputs(1983) <= not b or a;
    layer0_outputs(1984) <= not a;
    layer0_outputs(1985) <= a or b;
    layer0_outputs(1986) <= not (a or b);
    layer0_outputs(1987) <= not (a or b);
    layer0_outputs(1988) <= a or b;
    layer0_outputs(1989) <= not b or a;
    layer0_outputs(1990) <= not b or a;
    layer0_outputs(1991) <= not (a or b);
    layer0_outputs(1992) <= 1'b1;
    layer0_outputs(1993) <= b;
    layer0_outputs(1994) <= a or b;
    layer0_outputs(1995) <= not b;
    layer0_outputs(1996) <= b and not a;
    layer0_outputs(1997) <= a and not b;
    layer0_outputs(1998) <= a or b;
    layer0_outputs(1999) <= not a;
    layer0_outputs(2000) <= a and not b;
    layer0_outputs(2001) <= a and not b;
    layer0_outputs(2002) <= not (a and b);
    layer0_outputs(2003) <= not (a or b);
    layer0_outputs(2004) <= not (a xor b);
    layer0_outputs(2005) <= a;
    layer0_outputs(2006) <= 1'b1;
    layer0_outputs(2007) <= b and not a;
    layer0_outputs(2008) <= not a;
    layer0_outputs(2009) <= a and b;
    layer0_outputs(2010) <= a;
    layer0_outputs(2011) <= a and b;
    layer0_outputs(2012) <= not b;
    layer0_outputs(2013) <= not b or a;
    layer0_outputs(2014) <= 1'b1;
    layer0_outputs(2015) <= a and not b;
    layer0_outputs(2016) <= b and not a;
    layer0_outputs(2017) <= 1'b0;
    layer0_outputs(2018) <= not a;
    layer0_outputs(2019) <= not a or b;
    layer0_outputs(2020) <= b;
    layer0_outputs(2021) <= not (a or b);
    layer0_outputs(2022) <= not (a xor b);
    layer0_outputs(2023) <= b and not a;
    layer0_outputs(2024) <= not (a and b);
    layer0_outputs(2025) <= not b or a;
    layer0_outputs(2026) <= a;
    layer0_outputs(2027) <= not (a and b);
    layer0_outputs(2028) <= a xor b;
    layer0_outputs(2029) <= not b;
    layer0_outputs(2030) <= 1'b0;
    layer0_outputs(2031) <= not a or b;
    layer0_outputs(2032) <= not (a xor b);
    layer0_outputs(2033) <= a;
    layer0_outputs(2034) <= b and not a;
    layer0_outputs(2035) <= a and b;
    layer0_outputs(2036) <= not a;
    layer0_outputs(2037) <= b;
    layer0_outputs(2038) <= 1'b1;
    layer0_outputs(2039) <= a and not b;
    layer0_outputs(2040) <= not (a xor b);
    layer0_outputs(2041) <= not b;
    layer0_outputs(2042) <= a and b;
    layer0_outputs(2043) <= a and not b;
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= b;
    layer0_outputs(2046) <= b and not a;
    layer0_outputs(2047) <= a or b;
    layer0_outputs(2048) <= a;
    layer0_outputs(2049) <= not (a xor b);
    layer0_outputs(2050) <= a xor b;
    layer0_outputs(2051) <= not (a or b);
    layer0_outputs(2052) <= 1'b1;
    layer0_outputs(2053) <= b;
    layer0_outputs(2054) <= 1'b1;
    layer0_outputs(2055) <= not (a or b);
    layer0_outputs(2056) <= b;
    layer0_outputs(2057) <= not (a and b);
    layer0_outputs(2058) <= a;
    layer0_outputs(2059) <= a and b;
    layer0_outputs(2060) <= b;
    layer0_outputs(2061) <= a;
    layer0_outputs(2062) <= a and not b;
    layer0_outputs(2063) <= a;
    layer0_outputs(2064) <= 1'b1;
    layer0_outputs(2065) <= not (a and b);
    layer0_outputs(2066) <= a xor b;
    layer0_outputs(2067) <= 1'b0;
    layer0_outputs(2068) <= not a or b;
    layer0_outputs(2069) <= not a;
    layer0_outputs(2070) <= a and b;
    layer0_outputs(2071) <= a or b;
    layer0_outputs(2072) <= not (a and b);
    layer0_outputs(2073) <= a or b;
    layer0_outputs(2074) <= a and not b;
    layer0_outputs(2075) <= 1'b1;
    layer0_outputs(2076) <= not a or b;
    layer0_outputs(2077) <= not b or a;
    layer0_outputs(2078) <= not a or b;
    layer0_outputs(2079) <= not b or a;
    layer0_outputs(2080) <= 1'b0;
    layer0_outputs(2081) <= not a or b;
    layer0_outputs(2082) <= a and b;
    layer0_outputs(2083) <= b;
    layer0_outputs(2084) <= a;
    layer0_outputs(2085) <= 1'b0;
    layer0_outputs(2086) <= not (a or b);
    layer0_outputs(2087) <= not (a or b);
    layer0_outputs(2088) <= b and not a;
    layer0_outputs(2089) <= b and not a;
    layer0_outputs(2090) <= a or b;
    layer0_outputs(2091) <= a or b;
    layer0_outputs(2092) <= not (a xor b);
    layer0_outputs(2093) <= not (a xor b);
    layer0_outputs(2094) <= a or b;
    layer0_outputs(2095) <= a;
    layer0_outputs(2096) <= a;
    layer0_outputs(2097) <= a xor b;
    layer0_outputs(2098) <= not (a and b);
    layer0_outputs(2099) <= a and not b;
    layer0_outputs(2100) <= not b or a;
    layer0_outputs(2101) <= a and b;
    layer0_outputs(2102) <= a and b;
    layer0_outputs(2103) <= b;
    layer0_outputs(2104) <= not b;
    layer0_outputs(2105) <= b;
    layer0_outputs(2106) <= not (a or b);
    layer0_outputs(2107) <= 1'b0;
    layer0_outputs(2108) <= not a;
    layer0_outputs(2109) <= not (a and b);
    layer0_outputs(2110) <= a xor b;
    layer0_outputs(2111) <= a or b;
    layer0_outputs(2112) <= b;
    layer0_outputs(2113) <= 1'b1;
    layer0_outputs(2114) <= a or b;
    layer0_outputs(2115) <= a xor b;
    layer0_outputs(2116) <= 1'b0;
    layer0_outputs(2117) <= a or b;
    layer0_outputs(2118) <= a xor b;
    layer0_outputs(2119) <= b;
    layer0_outputs(2120) <= b and not a;
    layer0_outputs(2121) <= not (a xor b);
    layer0_outputs(2122) <= b and not a;
    layer0_outputs(2123) <= not b or a;
    layer0_outputs(2124) <= a and not b;
    layer0_outputs(2125) <= b;
    layer0_outputs(2126) <= a and b;
    layer0_outputs(2127) <= 1'b1;
    layer0_outputs(2128) <= not (a xor b);
    layer0_outputs(2129) <= a or b;
    layer0_outputs(2130) <= not a;
    layer0_outputs(2131) <= 1'b1;
    layer0_outputs(2132) <= not (a and b);
    layer0_outputs(2133) <= b and not a;
    layer0_outputs(2134) <= not a;
    layer0_outputs(2135) <= 1'b0;
    layer0_outputs(2136) <= 1'b0;
    layer0_outputs(2137) <= a xor b;
    layer0_outputs(2138) <= b and not a;
    layer0_outputs(2139) <= not b;
    layer0_outputs(2140) <= a and b;
    layer0_outputs(2141) <= not a;
    layer0_outputs(2142) <= not b;
    layer0_outputs(2143) <= b;
    layer0_outputs(2144) <= a;
    layer0_outputs(2145) <= a;
    layer0_outputs(2146) <= not b;
    layer0_outputs(2147) <= not b or a;
    layer0_outputs(2148) <= b;
    layer0_outputs(2149) <= not (a and b);
    layer0_outputs(2150) <= a;
    layer0_outputs(2151) <= b and not a;
    layer0_outputs(2152) <= a and b;
    layer0_outputs(2153) <= b;
    layer0_outputs(2154) <= not (a and b);
    layer0_outputs(2155) <= not a or b;
    layer0_outputs(2156) <= a and not b;
    layer0_outputs(2157) <= 1'b1;
    layer0_outputs(2158) <= a and not b;
    layer0_outputs(2159) <= a and b;
    layer0_outputs(2160) <= a xor b;
    layer0_outputs(2161) <= a xor b;
    layer0_outputs(2162) <= not b or a;
    layer0_outputs(2163) <= a;
    layer0_outputs(2164) <= a xor b;
    layer0_outputs(2165) <= b;
    layer0_outputs(2166) <= 1'b0;
    layer0_outputs(2167) <= not b or a;
    layer0_outputs(2168) <= a xor b;
    layer0_outputs(2169) <= not a;
    layer0_outputs(2170) <= not (a or b);
    layer0_outputs(2171) <= a xor b;
    layer0_outputs(2172) <= not b or a;
    layer0_outputs(2173) <= not b;
    layer0_outputs(2174) <= not b or a;
    layer0_outputs(2175) <= 1'b1;
    layer0_outputs(2176) <= 1'b1;
    layer0_outputs(2177) <= 1'b0;
    layer0_outputs(2178) <= not b or a;
    layer0_outputs(2179) <= b;
    layer0_outputs(2180) <= not (a xor b);
    layer0_outputs(2181) <= 1'b1;
    layer0_outputs(2182) <= a or b;
    layer0_outputs(2183) <= a and not b;
    layer0_outputs(2184) <= not (a xor b);
    layer0_outputs(2185) <= a and b;
    layer0_outputs(2186) <= not (a xor b);
    layer0_outputs(2187) <= a;
    layer0_outputs(2188) <= not (a and b);
    layer0_outputs(2189) <= a;
    layer0_outputs(2190) <= a xor b;
    layer0_outputs(2191) <= not a;
    layer0_outputs(2192) <= a;
    layer0_outputs(2193) <= not a;
    layer0_outputs(2194) <= not b;
    layer0_outputs(2195) <= not (a xor b);
    layer0_outputs(2196) <= not a or b;
    layer0_outputs(2197) <= a or b;
    layer0_outputs(2198) <= not (a xor b);
    layer0_outputs(2199) <= not b;
    layer0_outputs(2200) <= b;
    layer0_outputs(2201) <= a and not b;
    layer0_outputs(2202) <= not a;
    layer0_outputs(2203) <= b and not a;
    layer0_outputs(2204) <= not b;
    layer0_outputs(2205) <= 1'b1;
    layer0_outputs(2206) <= not b or a;
    layer0_outputs(2207) <= a or b;
    layer0_outputs(2208) <= not a or b;
    layer0_outputs(2209) <= not b;
    layer0_outputs(2210) <= b;
    layer0_outputs(2211) <= b;
    layer0_outputs(2212) <= a xor b;
    layer0_outputs(2213) <= not a;
    layer0_outputs(2214) <= not a or b;
    layer0_outputs(2215) <= 1'b1;
    layer0_outputs(2216) <= not (a or b);
    layer0_outputs(2217) <= not (a and b);
    layer0_outputs(2218) <= not b or a;
    layer0_outputs(2219) <= a and b;
    layer0_outputs(2220) <= a;
    layer0_outputs(2221) <= not (a and b);
    layer0_outputs(2222) <= a xor b;
    layer0_outputs(2223) <= b and not a;
    layer0_outputs(2224) <= a or b;
    layer0_outputs(2225) <= not a;
    layer0_outputs(2226) <= not (a or b);
    layer0_outputs(2227) <= not b or a;
    layer0_outputs(2228) <= a or b;
    layer0_outputs(2229) <= a;
    layer0_outputs(2230) <= not b;
    layer0_outputs(2231) <= a or b;
    layer0_outputs(2232) <= not a;
    layer0_outputs(2233) <= b;
    layer0_outputs(2234) <= not (a xor b);
    layer0_outputs(2235) <= not (a xor b);
    layer0_outputs(2236) <= a and not b;
    layer0_outputs(2237) <= not a;
    layer0_outputs(2238) <= not b;
    layer0_outputs(2239) <= not a;
    layer0_outputs(2240) <= a and b;
    layer0_outputs(2241) <= not a or b;
    layer0_outputs(2242) <= not (a or b);
    layer0_outputs(2243) <= not (a xor b);
    layer0_outputs(2244) <= not (a xor b);
    layer0_outputs(2245) <= a and not b;
    layer0_outputs(2246) <= not (a and b);
    layer0_outputs(2247) <= 1'b1;
    layer0_outputs(2248) <= a and not b;
    layer0_outputs(2249) <= a and b;
    layer0_outputs(2250) <= not (a or b);
    layer0_outputs(2251) <= 1'b0;
    layer0_outputs(2252) <= 1'b0;
    layer0_outputs(2253) <= b;
    layer0_outputs(2254) <= not b or a;
    layer0_outputs(2255) <= not a;
    layer0_outputs(2256) <= 1'b1;
    layer0_outputs(2257) <= not a or b;
    layer0_outputs(2258) <= a and not b;
    layer0_outputs(2259) <= a or b;
    layer0_outputs(2260) <= b and not a;
    layer0_outputs(2261) <= not a or b;
    layer0_outputs(2262) <= a and b;
    layer0_outputs(2263) <= not (a or b);
    layer0_outputs(2264) <= b and not a;
    layer0_outputs(2265) <= 1'b0;
    layer0_outputs(2266) <= b;
    layer0_outputs(2267) <= a or b;
    layer0_outputs(2268) <= not b or a;
    layer0_outputs(2269) <= not a or b;
    layer0_outputs(2270) <= not a or b;
    layer0_outputs(2271) <= a;
    layer0_outputs(2272) <= not b or a;
    layer0_outputs(2273) <= 1'b0;
    layer0_outputs(2274) <= a and not b;
    layer0_outputs(2275) <= not a;
    layer0_outputs(2276) <= not (a xor b);
    layer0_outputs(2277) <= not b;
    layer0_outputs(2278) <= 1'b0;
    layer0_outputs(2279) <= not a or b;
    layer0_outputs(2280) <= a;
    layer0_outputs(2281) <= a and not b;
    layer0_outputs(2282) <= 1'b0;
    layer0_outputs(2283) <= not b;
    layer0_outputs(2284) <= 1'b1;
    layer0_outputs(2285) <= 1'b0;
    layer0_outputs(2286) <= not b;
    layer0_outputs(2287) <= not (a or b);
    layer0_outputs(2288) <= 1'b0;
    layer0_outputs(2289) <= a and b;
    layer0_outputs(2290) <= b;
    layer0_outputs(2291) <= a and b;
    layer0_outputs(2292) <= not (a or b);
    layer0_outputs(2293) <= not b;
    layer0_outputs(2294) <= 1'b0;
    layer0_outputs(2295) <= not a;
    layer0_outputs(2296) <= not (a xor b);
    layer0_outputs(2297) <= not b;
    layer0_outputs(2298) <= a;
    layer0_outputs(2299) <= not b;
    layer0_outputs(2300) <= not a;
    layer0_outputs(2301) <= a and not b;
    layer0_outputs(2302) <= not (a and b);
    layer0_outputs(2303) <= not a;
    layer0_outputs(2304) <= not b;
    layer0_outputs(2305) <= not b;
    layer0_outputs(2306) <= a and not b;
    layer0_outputs(2307) <= not (a xor b);
    layer0_outputs(2308) <= b;
    layer0_outputs(2309) <= not (a or b);
    layer0_outputs(2310) <= not a;
    layer0_outputs(2311) <= 1'b1;
    layer0_outputs(2312) <= not b or a;
    layer0_outputs(2313) <= a xor b;
    layer0_outputs(2314) <= a or b;
    layer0_outputs(2315) <= 1'b0;
    layer0_outputs(2316) <= not b;
    layer0_outputs(2317) <= a and b;
    layer0_outputs(2318) <= a;
    layer0_outputs(2319) <= not b;
    layer0_outputs(2320) <= a or b;
    layer0_outputs(2321) <= a;
    layer0_outputs(2322) <= not b;
    layer0_outputs(2323) <= a;
    layer0_outputs(2324) <= not (a and b);
    layer0_outputs(2325) <= b and not a;
    layer0_outputs(2326) <= a and b;
    layer0_outputs(2327) <= b;
    layer0_outputs(2328) <= a and not b;
    layer0_outputs(2329) <= not a or b;
    layer0_outputs(2330) <= b and not a;
    layer0_outputs(2331) <= not (a xor b);
    layer0_outputs(2332) <= not a or b;
    layer0_outputs(2333) <= not b;
    layer0_outputs(2334) <= not b or a;
    layer0_outputs(2335) <= not a;
    layer0_outputs(2336) <= not b or a;
    layer0_outputs(2337) <= 1'b1;
    layer0_outputs(2338) <= 1'b0;
    layer0_outputs(2339) <= not (a or b);
    layer0_outputs(2340) <= not (a and b);
    layer0_outputs(2341) <= not a;
    layer0_outputs(2342) <= not b;
    layer0_outputs(2343) <= a;
    layer0_outputs(2344) <= b and not a;
    layer0_outputs(2345) <= not (a or b);
    layer0_outputs(2346) <= b;
    layer0_outputs(2347) <= not b;
    layer0_outputs(2348) <= a and not b;
    layer0_outputs(2349) <= not a;
    layer0_outputs(2350) <= a;
    layer0_outputs(2351) <= a and not b;
    layer0_outputs(2352) <= b;
    layer0_outputs(2353) <= a and b;
    layer0_outputs(2354) <= b;
    layer0_outputs(2355) <= b and not a;
    layer0_outputs(2356) <= not b;
    layer0_outputs(2357) <= not a;
    layer0_outputs(2358) <= not a or b;
    layer0_outputs(2359) <= not a;
    layer0_outputs(2360) <= a and not b;
    layer0_outputs(2361) <= 1'b1;
    layer0_outputs(2362) <= 1'b0;
    layer0_outputs(2363) <= 1'b0;
    layer0_outputs(2364) <= a and not b;
    layer0_outputs(2365) <= not a;
    layer0_outputs(2366) <= a and not b;
    layer0_outputs(2367) <= not (a or b);
    layer0_outputs(2368) <= not a or b;
    layer0_outputs(2369) <= not b or a;
    layer0_outputs(2370) <= a;
    layer0_outputs(2371) <= a or b;
    layer0_outputs(2372) <= 1'b0;
    layer0_outputs(2373) <= a and b;
    layer0_outputs(2374) <= a;
    layer0_outputs(2375) <= 1'b0;
    layer0_outputs(2376) <= a xor b;
    layer0_outputs(2377) <= 1'b0;
    layer0_outputs(2378) <= not b;
    layer0_outputs(2379) <= a;
    layer0_outputs(2380) <= not (a or b);
    layer0_outputs(2381) <= not (a or b);
    layer0_outputs(2382) <= not a;
    layer0_outputs(2383) <= not b;
    layer0_outputs(2384) <= 1'b0;
    layer0_outputs(2385) <= not (a or b);
    layer0_outputs(2386) <= a or b;
    layer0_outputs(2387) <= 1'b0;
    layer0_outputs(2388) <= not (a or b);
    layer0_outputs(2389) <= 1'b0;
    layer0_outputs(2390) <= a and not b;
    layer0_outputs(2391) <= not (a and b);
    layer0_outputs(2392) <= not (a or b);
    layer0_outputs(2393) <= 1'b0;
    layer0_outputs(2394) <= not a or b;
    layer0_outputs(2395) <= not (a and b);
    layer0_outputs(2396) <= a;
    layer0_outputs(2397) <= a and not b;
    layer0_outputs(2398) <= a xor b;
    layer0_outputs(2399) <= b;
    layer0_outputs(2400) <= b;
    layer0_outputs(2401) <= a or b;
    layer0_outputs(2402) <= 1'b1;
    layer0_outputs(2403) <= b and not a;
    layer0_outputs(2404) <= not (a and b);
    layer0_outputs(2405) <= not a or b;
    layer0_outputs(2406) <= not (a xor b);
    layer0_outputs(2407) <= a;
    layer0_outputs(2408) <= a and not b;
    layer0_outputs(2409) <= b;
    layer0_outputs(2410) <= not b or a;
    layer0_outputs(2411) <= b;
    layer0_outputs(2412) <= 1'b1;
    layer0_outputs(2413) <= 1'b1;
    layer0_outputs(2414) <= not b;
    layer0_outputs(2415) <= not b or a;
    layer0_outputs(2416) <= b and not a;
    layer0_outputs(2417) <= not (a xor b);
    layer0_outputs(2418) <= not (a and b);
    layer0_outputs(2419) <= not b or a;
    layer0_outputs(2420) <= 1'b0;
    layer0_outputs(2421) <= 1'b0;
    layer0_outputs(2422) <= b and not a;
    layer0_outputs(2423) <= not a;
    layer0_outputs(2424) <= not (a or b);
    layer0_outputs(2425) <= b;
    layer0_outputs(2426) <= b;
    layer0_outputs(2427) <= a;
    layer0_outputs(2428) <= a;
    layer0_outputs(2429) <= not (a and b);
    layer0_outputs(2430) <= 1'b0;
    layer0_outputs(2431) <= 1'b0;
    layer0_outputs(2432) <= a;
    layer0_outputs(2433) <= not (a or b);
    layer0_outputs(2434) <= a xor b;
    layer0_outputs(2435) <= a;
    layer0_outputs(2436) <= not (a xor b);
    layer0_outputs(2437) <= 1'b1;
    layer0_outputs(2438) <= a;
    layer0_outputs(2439) <= a and not b;
    layer0_outputs(2440) <= 1'b1;
    layer0_outputs(2441) <= not b;
    layer0_outputs(2442) <= 1'b0;
    layer0_outputs(2443) <= a and not b;
    layer0_outputs(2444) <= a or b;
    layer0_outputs(2445) <= a or b;
    layer0_outputs(2446) <= b and not a;
    layer0_outputs(2447) <= 1'b0;
    layer0_outputs(2448) <= not b or a;
    layer0_outputs(2449) <= b;
    layer0_outputs(2450) <= a;
    layer0_outputs(2451) <= not (a and b);
    layer0_outputs(2452) <= b and not a;
    layer0_outputs(2453) <= not a;
    layer0_outputs(2454) <= b and not a;
    layer0_outputs(2455) <= b;
    layer0_outputs(2456) <= not (a xor b);
    layer0_outputs(2457) <= a or b;
    layer0_outputs(2458) <= not (a xor b);
    layer0_outputs(2459) <= 1'b1;
    layer0_outputs(2460) <= b and not a;
    layer0_outputs(2461) <= not (a or b);
    layer0_outputs(2462) <= b;
    layer0_outputs(2463) <= not a or b;
    layer0_outputs(2464) <= a and not b;
    layer0_outputs(2465) <= not (a and b);
    layer0_outputs(2466) <= b;
    layer0_outputs(2467) <= b and not a;
    layer0_outputs(2468) <= not a or b;
    layer0_outputs(2469) <= 1'b0;
    layer0_outputs(2470) <= b and not a;
    layer0_outputs(2471) <= b and not a;
    layer0_outputs(2472) <= not a;
    layer0_outputs(2473) <= a and not b;
    layer0_outputs(2474) <= a or b;
    layer0_outputs(2475) <= b and not a;
    layer0_outputs(2476) <= b;
    layer0_outputs(2477) <= b;
    layer0_outputs(2478) <= not a;
    layer0_outputs(2479) <= a;
    layer0_outputs(2480) <= a xor b;
    layer0_outputs(2481) <= not a or b;
    layer0_outputs(2482) <= not (a or b);
    layer0_outputs(2483) <= b and not a;
    layer0_outputs(2484) <= a or b;
    layer0_outputs(2485) <= b and not a;
    layer0_outputs(2486) <= a and b;
    layer0_outputs(2487) <= a xor b;
    layer0_outputs(2488) <= not a;
    layer0_outputs(2489) <= not b;
    layer0_outputs(2490) <= not b;
    layer0_outputs(2491) <= not a or b;
    layer0_outputs(2492) <= not (a xor b);
    layer0_outputs(2493) <= not (a and b);
    layer0_outputs(2494) <= 1'b0;
    layer0_outputs(2495) <= b;
    layer0_outputs(2496) <= b;
    layer0_outputs(2497) <= 1'b1;
    layer0_outputs(2498) <= b;
    layer0_outputs(2499) <= a and not b;
    layer0_outputs(2500) <= b;
    layer0_outputs(2501) <= not b;
    layer0_outputs(2502) <= a;
    layer0_outputs(2503) <= not (a xor b);
    layer0_outputs(2504) <= 1'b1;
    layer0_outputs(2505) <= a and not b;
    layer0_outputs(2506) <= not (a xor b);
    layer0_outputs(2507) <= b and not a;
    layer0_outputs(2508) <= a;
    layer0_outputs(2509) <= a or b;
    layer0_outputs(2510) <= not (a xor b);
    layer0_outputs(2511) <= not a;
    layer0_outputs(2512) <= a and not b;
    layer0_outputs(2513) <= a;
    layer0_outputs(2514) <= not a;
    layer0_outputs(2515) <= b;
    layer0_outputs(2516) <= b;
    layer0_outputs(2517) <= not b or a;
    layer0_outputs(2518) <= not (a and b);
    layer0_outputs(2519) <= a and b;
    layer0_outputs(2520) <= 1'b0;
    layer0_outputs(2521) <= a and b;
    layer0_outputs(2522) <= a xor b;
    layer0_outputs(2523) <= b and not a;
    layer0_outputs(2524) <= not a;
    layer0_outputs(2525) <= a and not b;
    layer0_outputs(2526) <= 1'b0;
    layer0_outputs(2527) <= b;
    layer0_outputs(2528) <= not b;
    layer0_outputs(2529) <= 1'b0;
    layer0_outputs(2530) <= 1'b1;
    layer0_outputs(2531) <= not b;
    layer0_outputs(2532) <= not (a and b);
    layer0_outputs(2533) <= a and b;
    layer0_outputs(2534) <= a;
    layer0_outputs(2535) <= a and not b;
    layer0_outputs(2536) <= a or b;
    layer0_outputs(2537) <= a or b;
    layer0_outputs(2538) <= a and not b;
    layer0_outputs(2539) <= a;
    layer0_outputs(2540) <= not (a xor b);
    layer0_outputs(2541) <= a and not b;
    layer0_outputs(2542) <= a and not b;
    layer0_outputs(2543) <= 1'b1;
    layer0_outputs(2544) <= not (a xor b);
    layer0_outputs(2545) <= not b;
    layer0_outputs(2546) <= a xor b;
    layer0_outputs(2547) <= b and not a;
    layer0_outputs(2548) <= 1'b0;
    layer0_outputs(2549) <= 1'b1;
    layer0_outputs(2550) <= 1'b1;
    layer0_outputs(2551) <= not b or a;
    layer0_outputs(2552) <= a and not b;
    layer0_outputs(2553) <= a and b;
    layer0_outputs(2554) <= not b;
    layer0_outputs(2555) <= not b;
    layer0_outputs(2556) <= 1'b0;
    layer0_outputs(2557) <= not (a and b);
    layer0_outputs(2558) <= a;
    layer0_outputs(2559) <= not (a or b);
    layer0_outputs(2560) <= b;
    layer0_outputs(2561) <= b;
    layer0_outputs(2562) <= b and not a;
    layer0_outputs(2563) <= not a;
    layer0_outputs(2564) <= not (a and b);
    layer0_outputs(2565) <= not b or a;
    layer0_outputs(2566) <= a or b;
    layer0_outputs(2567) <= a;
    layer0_outputs(2568) <= b;
    layer0_outputs(2569) <= not b;
    layer0_outputs(2570) <= a or b;
    layer0_outputs(2571) <= 1'b0;
    layer0_outputs(2572) <= not a or b;
    layer0_outputs(2573) <= not a or b;
    layer0_outputs(2574) <= 1'b1;
    layer0_outputs(2575) <= b and not a;
    layer0_outputs(2576) <= 1'b1;
    layer0_outputs(2577) <= 1'b1;
    layer0_outputs(2578) <= not (a or b);
    layer0_outputs(2579) <= a;
    layer0_outputs(2580) <= not (a or b);
    layer0_outputs(2581) <= 1'b0;
    layer0_outputs(2582) <= a;
    layer0_outputs(2583) <= b and not a;
    layer0_outputs(2584) <= 1'b0;
    layer0_outputs(2585) <= a and b;
    layer0_outputs(2586) <= a and b;
    layer0_outputs(2587) <= b and not a;
    layer0_outputs(2588) <= a and b;
    layer0_outputs(2589) <= not (a xor b);
    layer0_outputs(2590) <= not b or a;
    layer0_outputs(2591) <= not b;
    layer0_outputs(2592) <= a and not b;
    layer0_outputs(2593) <= 1'b0;
    layer0_outputs(2594) <= not b;
    layer0_outputs(2595) <= 1'b0;
    layer0_outputs(2596) <= a and not b;
    layer0_outputs(2597) <= not (a and b);
    layer0_outputs(2598) <= 1'b1;
    layer0_outputs(2599) <= 1'b1;
    layer0_outputs(2600) <= not b or a;
    layer0_outputs(2601) <= b;
    layer0_outputs(2602) <= not b or a;
    layer0_outputs(2603) <= 1'b1;
    layer0_outputs(2604) <= a or b;
    layer0_outputs(2605) <= not (a and b);
    layer0_outputs(2606) <= not b or a;
    layer0_outputs(2607) <= 1'b0;
    layer0_outputs(2608) <= a;
    layer0_outputs(2609) <= a;
    layer0_outputs(2610) <= not b or a;
    layer0_outputs(2611) <= 1'b1;
    layer0_outputs(2612) <= a xor b;
    layer0_outputs(2613) <= not (a xor b);
    layer0_outputs(2614) <= not b or a;
    layer0_outputs(2615) <= a and not b;
    layer0_outputs(2616) <= a;
    layer0_outputs(2617) <= a and not b;
    layer0_outputs(2618) <= 1'b0;
    layer0_outputs(2619) <= a and not b;
    layer0_outputs(2620) <= not (a xor b);
    layer0_outputs(2621) <= not b;
    layer0_outputs(2622) <= 1'b0;
    layer0_outputs(2623) <= not a;
    layer0_outputs(2624) <= 1'b0;
    layer0_outputs(2625) <= a;
    layer0_outputs(2626) <= not a;
    layer0_outputs(2627) <= 1'b0;
    layer0_outputs(2628) <= b;
    layer0_outputs(2629) <= not b;
    layer0_outputs(2630) <= a;
    layer0_outputs(2631) <= b;
    layer0_outputs(2632) <= not a or b;
    layer0_outputs(2633) <= not (a or b);
    layer0_outputs(2634) <= 1'b0;
    layer0_outputs(2635) <= not b;
    layer0_outputs(2636) <= not (a and b);
    layer0_outputs(2637) <= not (a xor b);
    layer0_outputs(2638) <= not a;
    layer0_outputs(2639) <= not a or b;
    layer0_outputs(2640) <= a or b;
    layer0_outputs(2641) <= a;
    layer0_outputs(2642) <= b;
    layer0_outputs(2643) <= a and not b;
    layer0_outputs(2644) <= a;
    layer0_outputs(2645) <= not a or b;
    layer0_outputs(2646) <= not b or a;
    layer0_outputs(2647) <= a;
    layer0_outputs(2648) <= 1'b0;
    layer0_outputs(2649) <= not a;
    layer0_outputs(2650) <= not a;
    layer0_outputs(2651) <= not (a xor b);
    layer0_outputs(2652) <= a;
    layer0_outputs(2653) <= not a or b;
    layer0_outputs(2654) <= a or b;
    layer0_outputs(2655) <= not (a and b);
    layer0_outputs(2656) <= not a;
    layer0_outputs(2657) <= a xor b;
    layer0_outputs(2658) <= not b;
    layer0_outputs(2659) <= not (a and b);
    layer0_outputs(2660) <= a xor b;
    layer0_outputs(2661) <= a;
    layer0_outputs(2662) <= not a;
    layer0_outputs(2663) <= not (a and b);
    layer0_outputs(2664) <= not (a or b);
    layer0_outputs(2665) <= not b or a;
    layer0_outputs(2666) <= 1'b1;
    layer0_outputs(2667) <= not a or b;
    layer0_outputs(2668) <= not (a or b);
    layer0_outputs(2669) <= not a;
    layer0_outputs(2670) <= 1'b1;
    layer0_outputs(2671) <= b;
    layer0_outputs(2672) <= b and not a;
    layer0_outputs(2673) <= b and not a;
    layer0_outputs(2674) <= a and b;
    layer0_outputs(2675) <= a;
    layer0_outputs(2676) <= b and not a;
    layer0_outputs(2677) <= not (a and b);
    layer0_outputs(2678) <= not a or b;
    layer0_outputs(2679) <= a and not b;
    layer0_outputs(2680) <= not b or a;
    layer0_outputs(2681) <= 1'b1;
    layer0_outputs(2682) <= b;
    layer0_outputs(2683) <= b;
    layer0_outputs(2684) <= a xor b;
    layer0_outputs(2685) <= a and not b;
    layer0_outputs(2686) <= a and b;
    layer0_outputs(2687) <= a xor b;
    layer0_outputs(2688) <= a or b;
    layer0_outputs(2689) <= a xor b;
    layer0_outputs(2690) <= 1'b1;
    layer0_outputs(2691) <= a;
    layer0_outputs(2692) <= b;
    layer0_outputs(2693) <= 1'b1;
    layer0_outputs(2694) <= not b or a;
    layer0_outputs(2695) <= not (a xor b);
    layer0_outputs(2696) <= not (a and b);
    layer0_outputs(2697) <= a and not b;
    layer0_outputs(2698) <= not b;
    layer0_outputs(2699) <= not b or a;
    layer0_outputs(2700) <= a and not b;
    layer0_outputs(2701) <= not (a xor b);
    layer0_outputs(2702) <= a and not b;
    layer0_outputs(2703) <= not b or a;
    layer0_outputs(2704) <= a xor b;
    layer0_outputs(2705) <= a;
    layer0_outputs(2706) <= not b or a;
    layer0_outputs(2707) <= a;
    layer0_outputs(2708) <= a xor b;
    layer0_outputs(2709) <= not (a or b);
    layer0_outputs(2710) <= not a;
    layer0_outputs(2711) <= a and not b;
    layer0_outputs(2712) <= not b;
    layer0_outputs(2713) <= a;
    layer0_outputs(2714) <= not (a or b);
    layer0_outputs(2715) <= not b or a;
    layer0_outputs(2716) <= a and b;
    layer0_outputs(2717) <= a xor b;
    layer0_outputs(2718) <= a or b;
    layer0_outputs(2719) <= not (a and b);
    layer0_outputs(2720) <= a;
    layer0_outputs(2721) <= b and not a;
    layer0_outputs(2722) <= not a;
    layer0_outputs(2723) <= not a;
    layer0_outputs(2724) <= not b;
    layer0_outputs(2725) <= not a or b;
    layer0_outputs(2726) <= not b;
    layer0_outputs(2727) <= a or b;
    layer0_outputs(2728) <= not (a and b);
    layer0_outputs(2729) <= b;
    layer0_outputs(2730) <= not (a or b);
    layer0_outputs(2731) <= not b;
    layer0_outputs(2732) <= a xor b;
    layer0_outputs(2733) <= not (a and b);
    layer0_outputs(2734) <= a xor b;
    layer0_outputs(2735) <= a and not b;
    layer0_outputs(2736) <= 1'b0;
    layer0_outputs(2737) <= 1'b1;
    layer0_outputs(2738) <= not b or a;
    layer0_outputs(2739) <= b and not a;
    layer0_outputs(2740) <= not a or b;
    layer0_outputs(2741) <= not b;
    layer0_outputs(2742) <= not a;
    layer0_outputs(2743) <= 1'b1;
    layer0_outputs(2744) <= a;
    layer0_outputs(2745) <= b and not a;
    layer0_outputs(2746) <= not b or a;
    layer0_outputs(2747) <= not (a xor b);
    layer0_outputs(2748) <= 1'b0;
    layer0_outputs(2749) <= a and not b;
    layer0_outputs(2750) <= a and not b;
    layer0_outputs(2751) <= b;
    layer0_outputs(2752) <= a and not b;
    layer0_outputs(2753) <= a;
    layer0_outputs(2754) <= a or b;
    layer0_outputs(2755) <= not a or b;
    layer0_outputs(2756) <= b and not a;
    layer0_outputs(2757) <= a;
    layer0_outputs(2758) <= not (a and b);
    layer0_outputs(2759) <= a or b;
    layer0_outputs(2760) <= not b or a;
    layer0_outputs(2761) <= a or b;
    layer0_outputs(2762) <= b;
    layer0_outputs(2763) <= not (a or b);
    layer0_outputs(2764) <= a xor b;
    layer0_outputs(2765) <= 1'b1;
    layer0_outputs(2766) <= not b;
    layer0_outputs(2767) <= not a or b;
    layer0_outputs(2768) <= a or b;
    layer0_outputs(2769) <= not b;
    layer0_outputs(2770) <= not (a or b);
    layer0_outputs(2771) <= b and not a;
    layer0_outputs(2772) <= not (a or b);
    layer0_outputs(2773) <= not b or a;
    layer0_outputs(2774) <= a and not b;
    layer0_outputs(2775) <= a or b;
    layer0_outputs(2776) <= 1'b0;
    layer0_outputs(2777) <= 1'b0;
    layer0_outputs(2778) <= not a;
    layer0_outputs(2779) <= 1'b1;
    layer0_outputs(2780) <= 1'b1;
    layer0_outputs(2781) <= a and not b;
    layer0_outputs(2782) <= not a or b;
    layer0_outputs(2783) <= a and not b;
    layer0_outputs(2784) <= not b;
    layer0_outputs(2785) <= not b;
    layer0_outputs(2786) <= not (a xor b);
    layer0_outputs(2787) <= not a or b;
    layer0_outputs(2788) <= not a or b;
    layer0_outputs(2789) <= a;
    layer0_outputs(2790) <= not b;
    layer0_outputs(2791) <= b;
    layer0_outputs(2792) <= a and not b;
    layer0_outputs(2793) <= not b;
    layer0_outputs(2794) <= 1'b1;
    layer0_outputs(2795) <= not (a xor b);
    layer0_outputs(2796) <= b and not a;
    layer0_outputs(2797) <= b and not a;
    layer0_outputs(2798) <= a and b;
    layer0_outputs(2799) <= b;
    layer0_outputs(2800) <= not (a and b);
    layer0_outputs(2801) <= not (a xor b);
    layer0_outputs(2802) <= not b;
    layer0_outputs(2803) <= b;
    layer0_outputs(2804) <= not a or b;
    layer0_outputs(2805) <= a and not b;
    layer0_outputs(2806) <= not b;
    layer0_outputs(2807) <= not b or a;
    layer0_outputs(2808) <= 1'b1;
    layer0_outputs(2809) <= not a;
    layer0_outputs(2810) <= 1'b1;
    layer0_outputs(2811) <= b;
    layer0_outputs(2812) <= 1'b1;
    layer0_outputs(2813) <= not a or b;
    layer0_outputs(2814) <= not (a or b);
    layer0_outputs(2815) <= not b;
    layer0_outputs(2816) <= not (a and b);
    layer0_outputs(2817) <= not (a xor b);
    layer0_outputs(2818) <= not (a and b);
    layer0_outputs(2819) <= b;
    layer0_outputs(2820) <= not (a or b);
    layer0_outputs(2821) <= a and not b;
    layer0_outputs(2822) <= not (a or b);
    layer0_outputs(2823) <= 1'b1;
    layer0_outputs(2824) <= not a;
    layer0_outputs(2825) <= a or b;
    layer0_outputs(2826) <= b and not a;
    layer0_outputs(2827) <= not (a or b);
    layer0_outputs(2828) <= not (a xor b);
    layer0_outputs(2829) <= not b or a;
    layer0_outputs(2830) <= not a or b;
    layer0_outputs(2831) <= not a or b;
    layer0_outputs(2832) <= a;
    layer0_outputs(2833) <= a and b;
    layer0_outputs(2834) <= a or b;
    layer0_outputs(2835) <= not a or b;
    layer0_outputs(2836) <= not (a or b);
    layer0_outputs(2837) <= not (a xor b);
    layer0_outputs(2838) <= b;
    layer0_outputs(2839) <= 1'b0;
    layer0_outputs(2840) <= a and b;
    layer0_outputs(2841) <= not a;
    layer0_outputs(2842) <= 1'b1;
    layer0_outputs(2843) <= not (a xor b);
    layer0_outputs(2844) <= a and b;
    layer0_outputs(2845) <= not (a or b);
    layer0_outputs(2846) <= not b;
    layer0_outputs(2847) <= not b or a;
    layer0_outputs(2848) <= not (a or b);
    layer0_outputs(2849) <= not b or a;
    layer0_outputs(2850) <= not (a or b);
    layer0_outputs(2851) <= b;
    layer0_outputs(2852) <= not a;
    layer0_outputs(2853) <= not (a or b);
    layer0_outputs(2854) <= a xor b;
    layer0_outputs(2855) <= a and b;
    layer0_outputs(2856) <= a or b;
    layer0_outputs(2857) <= 1'b0;
    layer0_outputs(2858) <= not (a and b);
    layer0_outputs(2859) <= a;
    layer0_outputs(2860) <= not b;
    layer0_outputs(2861) <= a and not b;
    layer0_outputs(2862) <= not (a or b);
    layer0_outputs(2863) <= a xor b;
    layer0_outputs(2864) <= 1'b1;
    layer0_outputs(2865) <= not b or a;
    layer0_outputs(2866) <= a xor b;
    layer0_outputs(2867) <= a;
    layer0_outputs(2868) <= a or b;
    layer0_outputs(2869) <= a or b;
    layer0_outputs(2870) <= b;
    layer0_outputs(2871) <= not a or b;
    layer0_outputs(2872) <= a;
    layer0_outputs(2873) <= a xor b;
    layer0_outputs(2874) <= b;
    layer0_outputs(2875) <= not b;
    layer0_outputs(2876) <= b;
    layer0_outputs(2877) <= 1'b0;
    layer0_outputs(2878) <= not (a xor b);
    layer0_outputs(2879) <= not (a xor b);
    layer0_outputs(2880) <= 1'b0;
    layer0_outputs(2881) <= not a;
    layer0_outputs(2882) <= b;
    layer0_outputs(2883) <= a xor b;
    layer0_outputs(2884) <= a and b;
    layer0_outputs(2885) <= 1'b0;
    layer0_outputs(2886) <= not b;
    layer0_outputs(2887) <= a xor b;
    layer0_outputs(2888) <= not (a or b);
    layer0_outputs(2889) <= not (a xor b);
    layer0_outputs(2890) <= a xor b;
    layer0_outputs(2891) <= a;
    layer0_outputs(2892) <= a and not b;
    layer0_outputs(2893) <= b;
    layer0_outputs(2894) <= a;
    layer0_outputs(2895) <= not a;
    layer0_outputs(2896) <= not (a and b);
    layer0_outputs(2897) <= a or b;
    layer0_outputs(2898) <= a;
    layer0_outputs(2899) <= a and b;
    layer0_outputs(2900) <= 1'b0;
    layer0_outputs(2901) <= not (a or b);
    layer0_outputs(2902) <= not (a xor b);
    layer0_outputs(2903) <= a and b;
    layer0_outputs(2904) <= 1'b1;
    layer0_outputs(2905) <= b;
    layer0_outputs(2906) <= not (a or b);
    layer0_outputs(2907) <= a and not b;
    layer0_outputs(2908) <= b and not a;
    layer0_outputs(2909) <= not b;
    layer0_outputs(2910) <= a or b;
    layer0_outputs(2911) <= b and not a;
    layer0_outputs(2912) <= b and not a;
    layer0_outputs(2913) <= a;
    layer0_outputs(2914) <= not a;
    layer0_outputs(2915) <= a and not b;
    layer0_outputs(2916) <= 1'b0;
    layer0_outputs(2917) <= not a;
    layer0_outputs(2918) <= not a or b;
    layer0_outputs(2919) <= not b;
    layer0_outputs(2920) <= a and not b;
    layer0_outputs(2921) <= a xor b;
    layer0_outputs(2922) <= a and b;
    layer0_outputs(2923) <= 1'b0;
    layer0_outputs(2924) <= not b or a;
    layer0_outputs(2925) <= a and not b;
    layer0_outputs(2926) <= a;
    layer0_outputs(2927) <= a;
    layer0_outputs(2928) <= b and not a;
    layer0_outputs(2929) <= not a;
    layer0_outputs(2930) <= b;
    layer0_outputs(2931) <= not a or b;
    layer0_outputs(2932) <= 1'b0;
    layer0_outputs(2933) <= b;
    layer0_outputs(2934) <= not b;
    layer0_outputs(2935) <= not a or b;
    layer0_outputs(2936) <= 1'b1;
    layer0_outputs(2937) <= not b;
    layer0_outputs(2938) <= b;
    layer0_outputs(2939) <= a;
    layer0_outputs(2940) <= not (a and b);
    layer0_outputs(2941) <= a and b;
    layer0_outputs(2942) <= b;
    layer0_outputs(2943) <= a or b;
    layer0_outputs(2944) <= not b;
    layer0_outputs(2945) <= b and not a;
    layer0_outputs(2946) <= a and not b;
    layer0_outputs(2947) <= not a;
    layer0_outputs(2948) <= 1'b0;
    layer0_outputs(2949) <= not b;
    layer0_outputs(2950) <= not b or a;
    layer0_outputs(2951) <= 1'b1;
    layer0_outputs(2952) <= a;
    layer0_outputs(2953) <= a and b;
    layer0_outputs(2954) <= 1'b0;
    layer0_outputs(2955) <= not (a or b);
    layer0_outputs(2956) <= 1'b1;
    layer0_outputs(2957) <= not a or b;
    layer0_outputs(2958) <= a;
    layer0_outputs(2959) <= not b;
    layer0_outputs(2960) <= not a or b;
    layer0_outputs(2961) <= not a or b;
    layer0_outputs(2962) <= a and not b;
    layer0_outputs(2963) <= not (a and b);
    layer0_outputs(2964) <= a or b;
    layer0_outputs(2965) <= b;
    layer0_outputs(2966) <= not a;
    layer0_outputs(2967) <= a;
    layer0_outputs(2968) <= not b;
    layer0_outputs(2969) <= not (a and b);
    layer0_outputs(2970) <= not (a xor b);
    layer0_outputs(2971) <= b;
    layer0_outputs(2972) <= b;
    layer0_outputs(2973) <= b;
    layer0_outputs(2974) <= not b or a;
    layer0_outputs(2975) <= not (a xor b);
    layer0_outputs(2976) <= not b;
    layer0_outputs(2977) <= not a or b;
    layer0_outputs(2978) <= not a;
    layer0_outputs(2979) <= a and b;
    layer0_outputs(2980) <= a;
    layer0_outputs(2981) <= not (a or b);
    layer0_outputs(2982) <= 1'b0;
    layer0_outputs(2983) <= 1'b0;
    layer0_outputs(2984) <= a;
    layer0_outputs(2985) <= not b;
    layer0_outputs(2986) <= not (a or b);
    layer0_outputs(2987) <= not (a or b);
    layer0_outputs(2988) <= 1'b0;
    layer0_outputs(2989) <= not (a and b);
    layer0_outputs(2990) <= a xor b;
    layer0_outputs(2991) <= 1'b0;
    layer0_outputs(2992) <= a and b;
    layer0_outputs(2993) <= a or b;
    layer0_outputs(2994) <= 1'b1;
    layer0_outputs(2995) <= a;
    layer0_outputs(2996) <= a and b;
    layer0_outputs(2997) <= not (a xor b);
    layer0_outputs(2998) <= not (a and b);
    layer0_outputs(2999) <= not a or b;
    layer0_outputs(3000) <= a and b;
    layer0_outputs(3001) <= b;
    layer0_outputs(3002) <= not b;
    layer0_outputs(3003) <= not (a or b);
    layer0_outputs(3004) <= not a;
    layer0_outputs(3005) <= a and not b;
    layer0_outputs(3006) <= a xor b;
    layer0_outputs(3007) <= not a or b;
    layer0_outputs(3008) <= 1'b1;
    layer0_outputs(3009) <= 1'b1;
    layer0_outputs(3010) <= not (a or b);
    layer0_outputs(3011) <= not a;
    layer0_outputs(3012) <= not b;
    layer0_outputs(3013) <= not a;
    layer0_outputs(3014) <= not a or b;
    layer0_outputs(3015) <= 1'b1;
    layer0_outputs(3016) <= not (a xor b);
    layer0_outputs(3017) <= 1'b1;
    layer0_outputs(3018) <= 1'b1;
    layer0_outputs(3019) <= a and not b;
    layer0_outputs(3020) <= a;
    layer0_outputs(3021) <= 1'b0;
    layer0_outputs(3022) <= a and b;
    layer0_outputs(3023) <= not a or b;
    layer0_outputs(3024) <= not a or b;
    layer0_outputs(3025) <= not (a xor b);
    layer0_outputs(3026) <= a and b;
    layer0_outputs(3027) <= not a or b;
    layer0_outputs(3028) <= a or b;
    layer0_outputs(3029) <= a xor b;
    layer0_outputs(3030) <= b;
    layer0_outputs(3031) <= not b or a;
    layer0_outputs(3032) <= not b or a;
    layer0_outputs(3033) <= b;
    layer0_outputs(3034) <= a and b;
    layer0_outputs(3035) <= not (a and b);
    layer0_outputs(3036) <= not (a and b);
    layer0_outputs(3037) <= not a or b;
    layer0_outputs(3038) <= a;
    layer0_outputs(3039) <= 1'b1;
    layer0_outputs(3040) <= not (a or b);
    layer0_outputs(3041) <= b;
    layer0_outputs(3042) <= not (a and b);
    layer0_outputs(3043) <= not a;
    layer0_outputs(3044) <= a;
    layer0_outputs(3045) <= a and not b;
    layer0_outputs(3046) <= not a;
    layer0_outputs(3047) <= a and not b;
    layer0_outputs(3048) <= not (a xor b);
    layer0_outputs(3049) <= a;
    layer0_outputs(3050) <= a xor b;
    layer0_outputs(3051) <= b and not a;
    layer0_outputs(3052) <= not a;
    layer0_outputs(3053) <= 1'b1;
    layer0_outputs(3054) <= a or b;
    layer0_outputs(3055) <= 1'b0;
    layer0_outputs(3056) <= not (a or b);
    layer0_outputs(3057) <= not a;
    layer0_outputs(3058) <= a and not b;
    layer0_outputs(3059) <= not b;
    layer0_outputs(3060) <= a or b;
    layer0_outputs(3061) <= b and not a;
    layer0_outputs(3062) <= not a;
    layer0_outputs(3063) <= b;
    layer0_outputs(3064) <= a;
    layer0_outputs(3065) <= a xor b;
    layer0_outputs(3066) <= not (a or b);
    layer0_outputs(3067) <= b;
    layer0_outputs(3068) <= not a or b;
    layer0_outputs(3069) <= a xor b;
    layer0_outputs(3070) <= b and not a;
    layer0_outputs(3071) <= not a or b;
    layer0_outputs(3072) <= 1'b1;
    layer0_outputs(3073) <= not a;
    layer0_outputs(3074) <= not a or b;
    layer0_outputs(3075) <= not (a and b);
    layer0_outputs(3076) <= a and not b;
    layer0_outputs(3077) <= not (a and b);
    layer0_outputs(3078) <= not a;
    layer0_outputs(3079) <= a xor b;
    layer0_outputs(3080) <= not a or b;
    layer0_outputs(3081) <= a and not b;
    layer0_outputs(3082) <= a xor b;
    layer0_outputs(3083) <= not (a or b);
    layer0_outputs(3084) <= not b;
    layer0_outputs(3085) <= 1'b0;
    layer0_outputs(3086) <= 1'b1;
    layer0_outputs(3087) <= 1'b0;
    layer0_outputs(3088) <= not (a or b);
    layer0_outputs(3089) <= a and b;
    layer0_outputs(3090) <= 1'b0;
    layer0_outputs(3091) <= a and not b;
    layer0_outputs(3092) <= a and b;
    layer0_outputs(3093) <= not a or b;
    layer0_outputs(3094) <= not b or a;
    layer0_outputs(3095) <= 1'b0;
    layer0_outputs(3096) <= not b;
    layer0_outputs(3097) <= not b or a;
    layer0_outputs(3098) <= a;
    layer0_outputs(3099) <= a;
    layer0_outputs(3100) <= a and b;
    layer0_outputs(3101) <= not (a and b);
    layer0_outputs(3102) <= b and not a;
    layer0_outputs(3103) <= not b or a;
    layer0_outputs(3104) <= a and not b;
    layer0_outputs(3105) <= not b or a;
    layer0_outputs(3106) <= b and not a;
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= a or b;
    layer0_outputs(3109) <= not b or a;
    layer0_outputs(3110) <= 1'b0;
    layer0_outputs(3111) <= a or b;
    layer0_outputs(3112) <= not b;
    layer0_outputs(3113) <= a or b;
    layer0_outputs(3114) <= a;
    layer0_outputs(3115) <= not (a and b);
    layer0_outputs(3116) <= not (a and b);
    layer0_outputs(3117) <= a or b;
    layer0_outputs(3118) <= not b;
    layer0_outputs(3119) <= b;
    layer0_outputs(3120) <= not (a and b);
    layer0_outputs(3121) <= b;
    layer0_outputs(3122) <= 1'b0;
    layer0_outputs(3123) <= a;
    layer0_outputs(3124) <= not a or b;
    layer0_outputs(3125) <= not b or a;
    layer0_outputs(3126) <= 1'b0;
    layer0_outputs(3127) <= a and not b;
    layer0_outputs(3128) <= 1'b0;
    layer0_outputs(3129) <= a xor b;
    layer0_outputs(3130) <= not b or a;
    layer0_outputs(3131) <= 1'b1;
    layer0_outputs(3132) <= not (a or b);
    layer0_outputs(3133) <= not a;
    layer0_outputs(3134) <= a;
    layer0_outputs(3135) <= a;
    layer0_outputs(3136) <= 1'b0;
    layer0_outputs(3137) <= b;
    layer0_outputs(3138) <= not b;
    layer0_outputs(3139) <= a and b;
    layer0_outputs(3140) <= b;
    layer0_outputs(3141) <= b;
    layer0_outputs(3142) <= not a;
    layer0_outputs(3143) <= a or b;
    layer0_outputs(3144) <= a and b;
    layer0_outputs(3145) <= 1'b1;
    layer0_outputs(3146) <= a and b;
    layer0_outputs(3147) <= a and b;
    layer0_outputs(3148) <= 1'b1;
    layer0_outputs(3149) <= a or b;
    layer0_outputs(3150) <= not b;
    layer0_outputs(3151) <= not b or a;
    layer0_outputs(3152) <= not b;
    layer0_outputs(3153) <= a and b;
    layer0_outputs(3154) <= b;
    layer0_outputs(3155) <= not a or b;
    layer0_outputs(3156) <= not b;
    layer0_outputs(3157) <= a and b;
    layer0_outputs(3158) <= not b or a;
    layer0_outputs(3159) <= 1'b1;
    layer0_outputs(3160) <= a and not b;
    layer0_outputs(3161) <= a or b;
    layer0_outputs(3162) <= not b or a;
    layer0_outputs(3163) <= a or b;
    layer0_outputs(3164) <= a and b;
    layer0_outputs(3165) <= not (a xor b);
    layer0_outputs(3166) <= a xor b;
    layer0_outputs(3167) <= not a or b;
    layer0_outputs(3168) <= not a;
    layer0_outputs(3169) <= b;
    layer0_outputs(3170) <= not a;
    layer0_outputs(3171) <= b and not a;
    layer0_outputs(3172) <= b and not a;
    layer0_outputs(3173) <= 1'b0;
    layer0_outputs(3174) <= not b;
    layer0_outputs(3175) <= not b or a;
    layer0_outputs(3176) <= not b or a;
    layer0_outputs(3177) <= a;
    layer0_outputs(3178) <= not a;
    layer0_outputs(3179) <= not b or a;
    layer0_outputs(3180) <= a and not b;
    layer0_outputs(3181) <= 1'b1;
    layer0_outputs(3182) <= a or b;
    layer0_outputs(3183) <= 1'b1;
    layer0_outputs(3184) <= not a;
    layer0_outputs(3185) <= 1'b0;
    layer0_outputs(3186) <= a or b;
    layer0_outputs(3187) <= not b;
    layer0_outputs(3188) <= a xor b;
    layer0_outputs(3189) <= not b;
    layer0_outputs(3190) <= 1'b1;
    layer0_outputs(3191) <= not a;
    layer0_outputs(3192) <= not (a or b);
    layer0_outputs(3193) <= not (a and b);
    layer0_outputs(3194) <= b and not a;
    layer0_outputs(3195) <= a or b;
    layer0_outputs(3196) <= b and not a;
    layer0_outputs(3197) <= a or b;
    layer0_outputs(3198) <= not (a or b);
    layer0_outputs(3199) <= 1'b1;
    layer0_outputs(3200) <= a or b;
    layer0_outputs(3201) <= a xor b;
    layer0_outputs(3202) <= not (a and b);
    layer0_outputs(3203) <= b;
    layer0_outputs(3204) <= 1'b0;
    layer0_outputs(3205) <= not b;
    layer0_outputs(3206) <= not a;
    layer0_outputs(3207) <= a and b;
    layer0_outputs(3208) <= not (a and b);
    layer0_outputs(3209) <= a xor b;
    layer0_outputs(3210) <= 1'b1;
    layer0_outputs(3211) <= not (a xor b);
    layer0_outputs(3212) <= not (a and b);
    layer0_outputs(3213) <= not (a or b);
    layer0_outputs(3214) <= not a;
    layer0_outputs(3215) <= a and not b;
    layer0_outputs(3216) <= b;
    layer0_outputs(3217) <= a xor b;
    layer0_outputs(3218) <= not (a xor b);
    layer0_outputs(3219) <= a xor b;
    layer0_outputs(3220) <= a xor b;
    layer0_outputs(3221) <= a and b;
    layer0_outputs(3222) <= a and not b;
    layer0_outputs(3223) <= a;
    layer0_outputs(3224) <= not (a or b);
    layer0_outputs(3225) <= not a;
    layer0_outputs(3226) <= a and b;
    layer0_outputs(3227) <= 1'b0;
    layer0_outputs(3228) <= not (a and b);
    layer0_outputs(3229) <= b;
    layer0_outputs(3230) <= b;
    layer0_outputs(3231) <= a and b;
    layer0_outputs(3232) <= not a;
    layer0_outputs(3233) <= not b;
    layer0_outputs(3234) <= 1'b0;
    layer0_outputs(3235) <= b and not a;
    layer0_outputs(3236) <= 1'b1;
    layer0_outputs(3237) <= a;
    layer0_outputs(3238) <= 1'b0;
    layer0_outputs(3239) <= 1'b0;
    layer0_outputs(3240) <= 1'b1;
    layer0_outputs(3241) <= 1'b1;
    layer0_outputs(3242) <= not (a xor b);
    layer0_outputs(3243) <= a and not b;
    layer0_outputs(3244) <= not (a and b);
    layer0_outputs(3245) <= a and not b;
    layer0_outputs(3246) <= not b;
    layer0_outputs(3247) <= b;
    layer0_outputs(3248) <= 1'b0;
    layer0_outputs(3249) <= b and not a;
    layer0_outputs(3250) <= not (a and b);
    layer0_outputs(3251) <= b;
    layer0_outputs(3252) <= not (a and b);
    layer0_outputs(3253) <= b and not a;
    layer0_outputs(3254) <= 1'b0;
    layer0_outputs(3255) <= a or b;
    layer0_outputs(3256) <= not b;
    layer0_outputs(3257) <= not a;
    layer0_outputs(3258) <= not (a and b);
    layer0_outputs(3259) <= not b or a;
    layer0_outputs(3260) <= not (a and b);
    layer0_outputs(3261) <= not b or a;
    layer0_outputs(3262) <= not (a and b);
    layer0_outputs(3263) <= a xor b;
    layer0_outputs(3264) <= not (a or b);
    layer0_outputs(3265) <= not b;
    layer0_outputs(3266) <= not a;
    layer0_outputs(3267) <= not a;
    layer0_outputs(3268) <= not a;
    layer0_outputs(3269) <= a;
    layer0_outputs(3270) <= a;
    layer0_outputs(3271) <= not b or a;
    layer0_outputs(3272) <= b;
    layer0_outputs(3273) <= not (a xor b);
    layer0_outputs(3274) <= a and not b;
    layer0_outputs(3275) <= b;
    layer0_outputs(3276) <= a;
    layer0_outputs(3277) <= not a;
    layer0_outputs(3278) <= not (a xor b);
    layer0_outputs(3279) <= 1'b0;
    layer0_outputs(3280) <= not (a xor b);
    layer0_outputs(3281) <= b;
    layer0_outputs(3282) <= a or b;
    layer0_outputs(3283) <= a and b;
    layer0_outputs(3284) <= b and not a;
    layer0_outputs(3285) <= not b;
    layer0_outputs(3286) <= b;
    layer0_outputs(3287) <= a and b;
    layer0_outputs(3288) <= a or b;
    layer0_outputs(3289) <= not (a and b);
    layer0_outputs(3290) <= not b;
    layer0_outputs(3291) <= a or b;
    layer0_outputs(3292) <= 1'b0;
    layer0_outputs(3293) <= a or b;
    layer0_outputs(3294) <= a or b;
    layer0_outputs(3295) <= a and b;
    layer0_outputs(3296) <= b and not a;
    layer0_outputs(3297) <= not a;
    layer0_outputs(3298) <= a or b;
    layer0_outputs(3299) <= 1'b1;
    layer0_outputs(3300) <= a and b;
    layer0_outputs(3301) <= not a;
    layer0_outputs(3302) <= a or b;
    layer0_outputs(3303) <= a or b;
    layer0_outputs(3304) <= 1'b0;
    layer0_outputs(3305) <= b;
    layer0_outputs(3306) <= 1'b0;
    layer0_outputs(3307) <= not a;
    layer0_outputs(3308) <= not a or b;
    layer0_outputs(3309) <= 1'b0;
    layer0_outputs(3310) <= not a;
    layer0_outputs(3311) <= 1'b0;
    layer0_outputs(3312) <= a xor b;
    layer0_outputs(3313) <= not b;
    layer0_outputs(3314) <= not (a or b);
    layer0_outputs(3315) <= not (a or b);
    layer0_outputs(3316) <= a and b;
    layer0_outputs(3317) <= a xor b;
    layer0_outputs(3318) <= b and not a;
    layer0_outputs(3319) <= not (a and b);
    layer0_outputs(3320) <= a and not b;
    layer0_outputs(3321) <= not b;
    layer0_outputs(3322) <= b;
    layer0_outputs(3323) <= not b or a;
    layer0_outputs(3324) <= a and not b;
    layer0_outputs(3325) <= not b or a;
    layer0_outputs(3326) <= not b or a;
    layer0_outputs(3327) <= not a;
    layer0_outputs(3328) <= a and not b;
    layer0_outputs(3329) <= not a or b;
    layer0_outputs(3330) <= a and b;
    layer0_outputs(3331) <= not (a and b);
    layer0_outputs(3332) <= a and not b;
    layer0_outputs(3333) <= a xor b;
    layer0_outputs(3334) <= 1'b1;
    layer0_outputs(3335) <= a;
    layer0_outputs(3336) <= a and not b;
    layer0_outputs(3337) <= not a or b;
    layer0_outputs(3338) <= 1'b1;
    layer0_outputs(3339) <= 1'b0;
    layer0_outputs(3340) <= b and not a;
    layer0_outputs(3341) <= not (a or b);
    layer0_outputs(3342) <= a;
    layer0_outputs(3343) <= b and not a;
    layer0_outputs(3344) <= not a or b;
    layer0_outputs(3345) <= 1'b1;
    layer0_outputs(3346) <= not b;
    layer0_outputs(3347) <= 1'b1;
    layer0_outputs(3348) <= not (a or b);
    layer0_outputs(3349) <= not b or a;
    layer0_outputs(3350) <= not (a xor b);
    layer0_outputs(3351) <= a or b;
    layer0_outputs(3352) <= not (a and b);
    layer0_outputs(3353) <= not b;
    layer0_outputs(3354) <= not b or a;
    layer0_outputs(3355) <= a;
    layer0_outputs(3356) <= not b or a;
    layer0_outputs(3357) <= a xor b;
    layer0_outputs(3358) <= not a;
    layer0_outputs(3359) <= a xor b;
    layer0_outputs(3360) <= not a;
    layer0_outputs(3361) <= 1'b1;
    layer0_outputs(3362) <= b and not a;
    layer0_outputs(3363) <= not (a xor b);
    layer0_outputs(3364) <= a and not b;
    layer0_outputs(3365) <= a and b;
    layer0_outputs(3366) <= 1'b0;
    layer0_outputs(3367) <= not a;
    layer0_outputs(3368) <= not (a or b);
    layer0_outputs(3369) <= b;
    layer0_outputs(3370) <= not (a and b);
    layer0_outputs(3371) <= a xor b;
    layer0_outputs(3372) <= b and not a;
    layer0_outputs(3373) <= b;
    layer0_outputs(3374) <= not (a or b);
    layer0_outputs(3375) <= a and b;
    layer0_outputs(3376) <= not a or b;
    layer0_outputs(3377) <= not b;
    layer0_outputs(3378) <= not (a and b);
    layer0_outputs(3379) <= not a or b;
    layer0_outputs(3380) <= not (a xor b);
    layer0_outputs(3381) <= not (a xor b);
    layer0_outputs(3382) <= a and b;
    layer0_outputs(3383) <= not b;
    layer0_outputs(3384) <= a and not b;
    layer0_outputs(3385) <= a;
    layer0_outputs(3386) <= a;
    layer0_outputs(3387) <= a and b;
    layer0_outputs(3388) <= a and b;
    layer0_outputs(3389) <= not (a or b);
    layer0_outputs(3390) <= not (a xor b);
    layer0_outputs(3391) <= b and not a;
    layer0_outputs(3392) <= not a or b;
    layer0_outputs(3393) <= not a;
    layer0_outputs(3394) <= a and b;
    layer0_outputs(3395) <= not b;
    layer0_outputs(3396) <= a;
    layer0_outputs(3397) <= 1'b1;
    layer0_outputs(3398) <= 1'b1;
    layer0_outputs(3399) <= not (a and b);
    layer0_outputs(3400) <= not (a and b);
    layer0_outputs(3401) <= not a;
    layer0_outputs(3402) <= 1'b1;
    layer0_outputs(3403) <= b;
    layer0_outputs(3404) <= not a or b;
    layer0_outputs(3405) <= a xor b;
    layer0_outputs(3406) <= a or b;
    layer0_outputs(3407) <= a;
    layer0_outputs(3408) <= 1'b1;
    layer0_outputs(3409) <= not b;
    layer0_outputs(3410) <= b;
    layer0_outputs(3411) <= not a;
    layer0_outputs(3412) <= not a or b;
    layer0_outputs(3413) <= a and not b;
    layer0_outputs(3414) <= b;
    layer0_outputs(3415) <= a;
    layer0_outputs(3416) <= not (a and b);
    layer0_outputs(3417) <= a or b;
    layer0_outputs(3418) <= not a or b;
    layer0_outputs(3419) <= 1'b1;
    layer0_outputs(3420) <= a and not b;
    layer0_outputs(3421) <= not a or b;
    layer0_outputs(3422) <= not a;
    layer0_outputs(3423) <= not (a xor b);
    layer0_outputs(3424) <= a;
    layer0_outputs(3425) <= b and not a;
    layer0_outputs(3426) <= 1'b0;
    layer0_outputs(3427) <= a;
    layer0_outputs(3428) <= not a;
    layer0_outputs(3429) <= 1'b1;
    layer0_outputs(3430) <= not (a or b);
    layer0_outputs(3431) <= not b;
    layer0_outputs(3432) <= a;
    layer0_outputs(3433) <= not a;
    layer0_outputs(3434) <= b and not a;
    layer0_outputs(3435) <= a xor b;
    layer0_outputs(3436) <= a and b;
    layer0_outputs(3437) <= not (a xor b);
    layer0_outputs(3438) <= not (a or b);
    layer0_outputs(3439) <= a and b;
    layer0_outputs(3440) <= not (a and b);
    layer0_outputs(3441) <= a or b;
    layer0_outputs(3442) <= not (a or b);
    layer0_outputs(3443) <= not (a xor b);
    layer0_outputs(3444) <= not a;
    layer0_outputs(3445) <= b and not a;
    layer0_outputs(3446) <= 1'b0;
    layer0_outputs(3447) <= not a;
    layer0_outputs(3448) <= not a or b;
    layer0_outputs(3449) <= not a or b;
    layer0_outputs(3450) <= not b or a;
    layer0_outputs(3451) <= not b or a;
    layer0_outputs(3452) <= not b;
    layer0_outputs(3453) <= b and not a;
    layer0_outputs(3454) <= not b or a;
    layer0_outputs(3455) <= not b;
    layer0_outputs(3456) <= not b;
    layer0_outputs(3457) <= a and b;
    layer0_outputs(3458) <= a xor b;
    layer0_outputs(3459) <= a and not b;
    layer0_outputs(3460) <= not a;
    layer0_outputs(3461) <= 1'b0;
    layer0_outputs(3462) <= a or b;
    layer0_outputs(3463) <= not (a or b);
    layer0_outputs(3464) <= not (a or b);
    layer0_outputs(3465) <= a and not b;
    layer0_outputs(3466) <= a and b;
    layer0_outputs(3467) <= not a;
    layer0_outputs(3468) <= b and not a;
    layer0_outputs(3469) <= not b or a;
    layer0_outputs(3470) <= b and not a;
    layer0_outputs(3471) <= not (a or b);
    layer0_outputs(3472) <= not (a or b);
    layer0_outputs(3473) <= b and not a;
    layer0_outputs(3474) <= not a or b;
    layer0_outputs(3475) <= not a or b;
    layer0_outputs(3476) <= a;
    layer0_outputs(3477) <= not b or a;
    layer0_outputs(3478) <= not b;
    layer0_outputs(3479) <= not (a xor b);
    layer0_outputs(3480) <= a xor b;
    layer0_outputs(3481) <= b and not a;
    layer0_outputs(3482) <= b;
    layer0_outputs(3483) <= not b;
    layer0_outputs(3484) <= b and not a;
    layer0_outputs(3485) <= not (a or b);
    layer0_outputs(3486) <= not b;
    layer0_outputs(3487) <= a and b;
    layer0_outputs(3488) <= a and b;
    layer0_outputs(3489) <= a and b;
    layer0_outputs(3490) <= not b;
    layer0_outputs(3491) <= 1'b1;
    layer0_outputs(3492) <= a and b;
    layer0_outputs(3493) <= not (a and b);
    layer0_outputs(3494) <= not b;
    layer0_outputs(3495) <= a xor b;
    layer0_outputs(3496) <= not b or a;
    layer0_outputs(3497) <= b and not a;
    layer0_outputs(3498) <= a and not b;
    layer0_outputs(3499) <= not a;
    layer0_outputs(3500) <= not (a xor b);
    layer0_outputs(3501) <= a xor b;
    layer0_outputs(3502) <= 1'b1;
    layer0_outputs(3503) <= not b or a;
    layer0_outputs(3504) <= not a;
    layer0_outputs(3505) <= a and not b;
    layer0_outputs(3506) <= not b or a;
    layer0_outputs(3507) <= not a;
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= a and not b;
    layer0_outputs(3510) <= a or b;
    layer0_outputs(3511) <= not b or a;
    layer0_outputs(3512) <= b and not a;
    layer0_outputs(3513) <= not a or b;
    layer0_outputs(3514) <= not (a and b);
    layer0_outputs(3515) <= 1'b1;
    layer0_outputs(3516) <= a or b;
    layer0_outputs(3517) <= a xor b;
    layer0_outputs(3518) <= not b;
    layer0_outputs(3519) <= not (a and b);
    layer0_outputs(3520) <= b;
    layer0_outputs(3521) <= 1'b1;
    layer0_outputs(3522) <= 1'b1;
    layer0_outputs(3523) <= a or b;
    layer0_outputs(3524) <= 1'b0;
    layer0_outputs(3525) <= a;
    layer0_outputs(3526) <= a;
    layer0_outputs(3527) <= a;
    layer0_outputs(3528) <= a xor b;
    layer0_outputs(3529) <= not a or b;
    layer0_outputs(3530) <= not a or b;
    layer0_outputs(3531) <= b and not a;
    layer0_outputs(3532) <= a xor b;
    layer0_outputs(3533) <= not a;
    layer0_outputs(3534) <= a;
    layer0_outputs(3535) <= not b;
    layer0_outputs(3536) <= not (a and b);
    layer0_outputs(3537) <= 1'b0;
    layer0_outputs(3538) <= 1'b1;
    layer0_outputs(3539) <= 1'b0;
    layer0_outputs(3540) <= a or b;
    layer0_outputs(3541) <= not a;
    layer0_outputs(3542) <= not a or b;
    layer0_outputs(3543) <= not (a xor b);
    layer0_outputs(3544) <= a and b;
    layer0_outputs(3545) <= a or b;
    layer0_outputs(3546) <= a and not b;
    layer0_outputs(3547) <= a;
    layer0_outputs(3548) <= not b or a;
    layer0_outputs(3549) <= not b;
    layer0_outputs(3550) <= not (a and b);
    layer0_outputs(3551) <= a and b;
    layer0_outputs(3552) <= not (a and b);
    layer0_outputs(3553) <= a and b;
    layer0_outputs(3554) <= 1'b1;
    layer0_outputs(3555) <= b;
    layer0_outputs(3556) <= not a or b;
    layer0_outputs(3557) <= a;
    layer0_outputs(3558) <= not (a or b);
    layer0_outputs(3559) <= not a or b;
    layer0_outputs(3560) <= a or b;
    layer0_outputs(3561) <= not b or a;
    layer0_outputs(3562) <= a and not b;
    layer0_outputs(3563) <= 1'b1;
    layer0_outputs(3564) <= not (a xor b);
    layer0_outputs(3565) <= not b or a;
    layer0_outputs(3566) <= a or b;
    layer0_outputs(3567) <= a and not b;
    layer0_outputs(3568) <= a;
    layer0_outputs(3569) <= a and b;
    layer0_outputs(3570) <= not (a xor b);
    layer0_outputs(3571) <= not (a or b);
    layer0_outputs(3572) <= b;
    layer0_outputs(3573) <= a or b;
    layer0_outputs(3574) <= not b or a;
    layer0_outputs(3575) <= 1'b0;
    layer0_outputs(3576) <= a xor b;
    layer0_outputs(3577) <= not a;
    layer0_outputs(3578) <= not b;
    layer0_outputs(3579) <= a;
    layer0_outputs(3580) <= 1'b1;
    layer0_outputs(3581) <= b;
    layer0_outputs(3582) <= 1'b1;
    layer0_outputs(3583) <= a and not b;
    layer0_outputs(3584) <= not b or a;
    layer0_outputs(3585) <= not b or a;
    layer0_outputs(3586) <= not b;
    layer0_outputs(3587) <= 1'b1;
    layer0_outputs(3588) <= not b;
    layer0_outputs(3589) <= a or b;
    layer0_outputs(3590) <= 1'b1;
    layer0_outputs(3591) <= not a or b;
    layer0_outputs(3592) <= not (a and b);
    layer0_outputs(3593) <= not (a xor b);
    layer0_outputs(3594) <= not (a or b);
    layer0_outputs(3595) <= not a or b;
    layer0_outputs(3596) <= not (a or b);
    layer0_outputs(3597) <= a or b;
    layer0_outputs(3598) <= not a;
    layer0_outputs(3599) <= not (a and b);
    layer0_outputs(3600) <= a xor b;
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= not (a and b);
    layer0_outputs(3603) <= a;
    layer0_outputs(3604) <= a or b;
    layer0_outputs(3605) <= a xor b;
    layer0_outputs(3606) <= a;
    layer0_outputs(3607) <= b;
    layer0_outputs(3608) <= b;
    layer0_outputs(3609) <= b and not a;
    layer0_outputs(3610) <= not (a and b);
    layer0_outputs(3611) <= 1'b0;
    layer0_outputs(3612) <= a and not b;
    layer0_outputs(3613) <= not (a and b);
    layer0_outputs(3614) <= a;
    layer0_outputs(3615) <= not b or a;
    layer0_outputs(3616) <= a and b;
    layer0_outputs(3617) <= not (a or b);
    layer0_outputs(3618) <= a;
    layer0_outputs(3619) <= a xor b;
    layer0_outputs(3620) <= not a;
    layer0_outputs(3621) <= a and b;
    layer0_outputs(3622) <= a;
    layer0_outputs(3623) <= not b;
    layer0_outputs(3624) <= a and not b;
    layer0_outputs(3625) <= a or b;
    layer0_outputs(3626) <= not a;
    layer0_outputs(3627) <= b and not a;
    layer0_outputs(3628) <= not (a and b);
    layer0_outputs(3629) <= 1'b1;
    layer0_outputs(3630) <= 1'b0;
    layer0_outputs(3631) <= b;
    layer0_outputs(3632) <= not (a and b);
    layer0_outputs(3633) <= not b;
    layer0_outputs(3634) <= a or b;
    layer0_outputs(3635) <= not (a xor b);
    layer0_outputs(3636) <= not (a xor b);
    layer0_outputs(3637) <= 1'b1;
    layer0_outputs(3638) <= a;
    layer0_outputs(3639) <= not b;
    layer0_outputs(3640) <= not a or b;
    layer0_outputs(3641) <= a or b;
    layer0_outputs(3642) <= not a or b;
    layer0_outputs(3643) <= not a or b;
    layer0_outputs(3644) <= not (a and b);
    layer0_outputs(3645) <= not b or a;
    layer0_outputs(3646) <= not a or b;
    layer0_outputs(3647) <= not b;
    layer0_outputs(3648) <= not a;
    layer0_outputs(3649) <= not b;
    layer0_outputs(3650) <= 1'b0;
    layer0_outputs(3651) <= 1'b1;
    layer0_outputs(3652) <= not a or b;
    layer0_outputs(3653) <= not (a or b);
    layer0_outputs(3654) <= not a or b;
    layer0_outputs(3655) <= not (a or b);
    layer0_outputs(3656) <= not (a and b);
    layer0_outputs(3657) <= 1'b1;
    layer0_outputs(3658) <= not a or b;
    layer0_outputs(3659) <= not b;
    layer0_outputs(3660) <= a or b;
    layer0_outputs(3661) <= b;
    layer0_outputs(3662) <= not b or a;
    layer0_outputs(3663) <= 1'b1;
    layer0_outputs(3664) <= b and not a;
    layer0_outputs(3665) <= a;
    layer0_outputs(3666) <= a and b;
    layer0_outputs(3667) <= b and not a;
    layer0_outputs(3668) <= b and not a;
    layer0_outputs(3669) <= a;
    layer0_outputs(3670) <= a;
    layer0_outputs(3671) <= not (a and b);
    layer0_outputs(3672) <= 1'b0;
    layer0_outputs(3673) <= b;
    layer0_outputs(3674) <= 1'b0;
    layer0_outputs(3675) <= a and b;
    layer0_outputs(3676) <= 1'b0;
    layer0_outputs(3677) <= 1'b0;
    layer0_outputs(3678) <= 1'b0;
    layer0_outputs(3679) <= not a or b;
    layer0_outputs(3680) <= a xor b;
    layer0_outputs(3681) <= b;
    layer0_outputs(3682) <= not a or b;
    layer0_outputs(3683) <= 1'b1;
    layer0_outputs(3684) <= 1'b0;
    layer0_outputs(3685) <= not (a or b);
    layer0_outputs(3686) <= a or b;
    layer0_outputs(3687) <= a and not b;
    layer0_outputs(3688) <= b;
    layer0_outputs(3689) <= not (a and b);
    layer0_outputs(3690) <= a or b;
    layer0_outputs(3691) <= not b;
    layer0_outputs(3692) <= a and b;
    layer0_outputs(3693) <= not (a or b);
    layer0_outputs(3694) <= a or b;
    layer0_outputs(3695) <= not b;
    layer0_outputs(3696) <= 1'b1;
    layer0_outputs(3697) <= b and not a;
    layer0_outputs(3698) <= a and b;
    layer0_outputs(3699) <= not b or a;
    layer0_outputs(3700) <= 1'b1;
    layer0_outputs(3701) <= not a or b;
    layer0_outputs(3702) <= b;
    layer0_outputs(3703) <= a;
    layer0_outputs(3704) <= not (a and b);
    layer0_outputs(3705) <= b and not a;
    layer0_outputs(3706) <= 1'b0;
    layer0_outputs(3707) <= not b or a;
    layer0_outputs(3708) <= not b;
    layer0_outputs(3709) <= a;
    layer0_outputs(3710) <= a and not b;
    layer0_outputs(3711) <= not b or a;
    layer0_outputs(3712) <= not (a or b);
    layer0_outputs(3713) <= a or b;
    layer0_outputs(3714) <= 1'b0;
    layer0_outputs(3715) <= a xor b;
    layer0_outputs(3716) <= a xor b;
    layer0_outputs(3717) <= a and b;
    layer0_outputs(3718) <= not (a and b);
    layer0_outputs(3719) <= a;
    layer0_outputs(3720) <= not (a or b);
    layer0_outputs(3721) <= a and not b;
    layer0_outputs(3722) <= a or b;
    layer0_outputs(3723) <= b;
    layer0_outputs(3724) <= 1'b1;
    layer0_outputs(3725) <= a;
    layer0_outputs(3726) <= 1'b0;
    layer0_outputs(3727) <= a or b;
    layer0_outputs(3728) <= not (a or b);
    layer0_outputs(3729) <= not (a or b);
    layer0_outputs(3730) <= not b;
    layer0_outputs(3731) <= b and not a;
    layer0_outputs(3732) <= a or b;
    layer0_outputs(3733) <= not a or b;
    layer0_outputs(3734) <= a or b;
    layer0_outputs(3735) <= a and not b;
    layer0_outputs(3736) <= not (a xor b);
    layer0_outputs(3737) <= b and not a;
    layer0_outputs(3738) <= 1'b0;
    layer0_outputs(3739) <= 1'b0;
    layer0_outputs(3740) <= 1'b1;
    layer0_outputs(3741) <= a and not b;
    layer0_outputs(3742) <= a xor b;
    layer0_outputs(3743) <= b and not a;
    layer0_outputs(3744) <= a or b;
    layer0_outputs(3745) <= not a;
    layer0_outputs(3746) <= not (a xor b);
    layer0_outputs(3747) <= b;
    layer0_outputs(3748) <= not a or b;
    layer0_outputs(3749) <= b;
    layer0_outputs(3750) <= a and b;
    layer0_outputs(3751) <= not b or a;
    layer0_outputs(3752) <= a or b;
    layer0_outputs(3753) <= not a;
    layer0_outputs(3754) <= a;
    layer0_outputs(3755) <= not a;
    layer0_outputs(3756) <= not (a or b);
    layer0_outputs(3757) <= b and not a;
    layer0_outputs(3758) <= not a;
    layer0_outputs(3759) <= not (a or b);
    layer0_outputs(3760) <= a;
    layer0_outputs(3761) <= b;
    layer0_outputs(3762) <= a and not b;
    layer0_outputs(3763) <= not b;
    layer0_outputs(3764) <= a or b;
    layer0_outputs(3765) <= not (a and b);
    layer0_outputs(3766) <= b;
    layer0_outputs(3767) <= b and not a;
    layer0_outputs(3768) <= b and not a;
    layer0_outputs(3769) <= 1'b0;
    layer0_outputs(3770) <= a and b;
    layer0_outputs(3771) <= a and b;
    layer0_outputs(3772) <= 1'b1;
    layer0_outputs(3773) <= a;
    layer0_outputs(3774) <= b and not a;
    layer0_outputs(3775) <= not (a and b);
    layer0_outputs(3776) <= a and not b;
    layer0_outputs(3777) <= a or b;
    layer0_outputs(3778) <= b;
    layer0_outputs(3779) <= b;
    layer0_outputs(3780) <= not a;
    layer0_outputs(3781) <= not a or b;
    layer0_outputs(3782) <= not (a xor b);
    layer0_outputs(3783) <= a and not b;
    layer0_outputs(3784) <= not (a xor b);
    layer0_outputs(3785) <= b and not a;
    layer0_outputs(3786) <= a;
    layer0_outputs(3787) <= b;
    layer0_outputs(3788) <= not (a xor b);
    layer0_outputs(3789) <= not (a or b);
    layer0_outputs(3790) <= not a;
    layer0_outputs(3791) <= not (a and b);
    layer0_outputs(3792) <= b;
    layer0_outputs(3793) <= 1'b0;
    layer0_outputs(3794) <= not b;
    layer0_outputs(3795) <= not (a or b);
    layer0_outputs(3796) <= a and not b;
    layer0_outputs(3797) <= a or b;
    layer0_outputs(3798) <= a or b;
    layer0_outputs(3799) <= a and not b;
    layer0_outputs(3800) <= a;
    layer0_outputs(3801) <= a or b;
    layer0_outputs(3802) <= not a or b;
    layer0_outputs(3803) <= not a;
    layer0_outputs(3804) <= 1'b0;
    layer0_outputs(3805) <= 1'b1;
    layer0_outputs(3806) <= not (a and b);
    layer0_outputs(3807) <= not b or a;
    layer0_outputs(3808) <= a and not b;
    layer0_outputs(3809) <= a xor b;
    layer0_outputs(3810) <= b and not a;
    layer0_outputs(3811) <= not (a or b);
    layer0_outputs(3812) <= a;
    layer0_outputs(3813) <= 1'b0;
    layer0_outputs(3814) <= 1'b1;
    layer0_outputs(3815) <= not (a or b);
    layer0_outputs(3816) <= a;
    layer0_outputs(3817) <= not a;
    layer0_outputs(3818) <= not b or a;
    layer0_outputs(3819) <= not a or b;
    layer0_outputs(3820) <= not a;
    layer0_outputs(3821) <= b;
    layer0_outputs(3822) <= 1'b1;
    layer0_outputs(3823) <= not (a or b);
    layer0_outputs(3824) <= not b;
    layer0_outputs(3825) <= not (a or b);
    layer0_outputs(3826) <= not a;
    layer0_outputs(3827) <= 1'b0;
    layer0_outputs(3828) <= not a;
    layer0_outputs(3829) <= not a;
    layer0_outputs(3830) <= 1'b1;
    layer0_outputs(3831) <= b;
    layer0_outputs(3832) <= not (a or b);
    layer0_outputs(3833) <= a xor b;
    layer0_outputs(3834) <= not a or b;
    layer0_outputs(3835) <= not (a or b);
    layer0_outputs(3836) <= a;
    layer0_outputs(3837) <= b;
    layer0_outputs(3838) <= 1'b0;
    layer0_outputs(3839) <= not a;
    layer0_outputs(3840) <= b and not a;
    layer0_outputs(3841) <= not a;
    layer0_outputs(3842) <= a and not b;
    layer0_outputs(3843) <= 1'b1;
    layer0_outputs(3844) <= a xor b;
    layer0_outputs(3845) <= b and not a;
    layer0_outputs(3846) <= not b;
    layer0_outputs(3847) <= 1'b1;
    layer0_outputs(3848) <= b and not a;
    layer0_outputs(3849) <= a;
    layer0_outputs(3850) <= 1'b1;
    layer0_outputs(3851) <= a or b;
    layer0_outputs(3852) <= b;
    layer0_outputs(3853) <= a and not b;
    layer0_outputs(3854) <= a and b;
    layer0_outputs(3855) <= a and not b;
    layer0_outputs(3856) <= b;
    layer0_outputs(3857) <= not b;
    layer0_outputs(3858) <= 1'b0;
    layer0_outputs(3859) <= not a;
    layer0_outputs(3860) <= a or b;
    layer0_outputs(3861) <= not (a and b);
    layer0_outputs(3862) <= 1'b1;
    layer0_outputs(3863) <= 1'b0;
    layer0_outputs(3864) <= 1'b0;
    layer0_outputs(3865) <= not b;
    layer0_outputs(3866) <= not (a or b);
    layer0_outputs(3867) <= b and not a;
    layer0_outputs(3868) <= 1'b0;
    layer0_outputs(3869) <= not b or a;
    layer0_outputs(3870) <= 1'b0;
    layer0_outputs(3871) <= not (a or b);
    layer0_outputs(3872) <= not (a xor b);
    layer0_outputs(3873) <= 1'b0;
    layer0_outputs(3874) <= not (a or b);
    layer0_outputs(3875) <= not (a xor b);
    layer0_outputs(3876) <= a;
    layer0_outputs(3877) <= a and b;
    layer0_outputs(3878) <= 1'b0;
    layer0_outputs(3879) <= not (a xor b);
    layer0_outputs(3880) <= a;
    layer0_outputs(3881) <= a and b;
    layer0_outputs(3882) <= not (a or b);
    layer0_outputs(3883) <= not a;
    layer0_outputs(3884) <= a;
    layer0_outputs(3885) <= not a;
    layer0_outputs(3886) <= 1'b0;
    layer0_outputs(3887) <= a;
    layer0_outputs(3888) <= a and b;
    layer0_outputs(3889) <= a and b;
    layer0_outputs(3890) <= a;
    layer0_outputs(3891) <= not (a or b);
    layer0_outputs(3892) <= not a or b;
    layer0_outputs(3893) <= 1'b0;
    layer0_outputs(3894) <= not (a and b);
    layer0_outputs(3895) <= not b;
    layer0_outputs(3896) <= a and b;
    layer0_outputs(3897) <= 1'b0;
    layer0_outputs(3898) <= not (a or b);
    layer0_outputs(3899) <= 1'b0;
    layer0_outputs(3900) <= a or b;
    layer0_outputs(3901) <= not (a xor b);
    layer0_outputs(3902) <= not b or a;
    layer0_outputs(3903) <= a or b;
    layer0_outputs(3904) <= not a;
    layer0_outputs(3905) <= a and b;
    layer0_outputs(3906) <= a xor b;
    layer0_outputs(3907) <= 1'b1;
    layer0_outputs(3908) <= 1'b0;
    layer0_outputs(3909) <= not (a and b);
    layer0_outputs(3910) <= b;
    layer0_outputs(3911) <= not (a or b);
    layer0_outputs(3912) <= a xor b;
    layer0_outputs(3913) <= a xor b;
    layer0_outputs(3914) <= a;
    layer0_outputs(3915) <= not b;
    layer0_outputs(3916) <= 1'b0;
    layer0_outputs(3917) <= a and not b;
    layer0_outputs(3918) <= a xor b;
    layer0_outputs(3919) <= a or b;
    layer0_outputs(3920) <= b and not a;
    layer0_outputs(3921) <= a xor b;
    layer0_outputs(3922) <= not (a and b);
    layer0_outputs(3923) <= not a;
    layer0_outputs(3924) <= not b or a;
    layer0_outputs(3925) <= not a or b;
    layer0_outputs(3926) <= a and b;
    layer0_outputs(3927) <= a or b;
    layer0_outputs(3928) <= not b or a;
    layer0_outputs(3929) <= not a;
    layer0_outputs(3930) <= b and not a;
    layer0_outputs(3931) <= a and b;
    layer0_outputs(3932) <= 1'b0;
    layer0_outputs(3933) <= not a or b;
    layer0_outputs(3934) <= not (a xor b);
    layer0_outputs(3935) <= not a or b;
    layer0_outputs(3936) <= a;
    layer0_outputs(3937) <= a or b;
    layer0_outputs(3938) <= a;
    layer0_outputs(3939) <= not b or a;
    layer0_outputs(3940) <= 1'b0;
    layer0_outputs(3941) <= not (a or b);
    layer0_outputs(3942) <= not a or b;
    layer0_outputs(3943) <= 1'b0;
    layer0_outputs(3944) <= a or b;
    layer0_outputs(3945) <= not b or a;
    layer0_outputs(3946) <= not a or b;
    layer0_outputs(3947) <= not (a and b);
    layer0_outputs(3948) <= a or b;
    layer0_outputs(3949) <= a and not b;
    layer0_outputs(3950) <= a;
    layer0_outputs(3951) <= not (a and b);
    layer0_outputs(3952) <= a and b;
    layer0_outputs(3953) <= 1'b1;
    layer0_outputs(3954) <= not a or b;
    layer0_outputs(3955) <= a and not b;
    layer0_outputs(3956) <= not b;
    layer0_outputs(3957) <= a;
    layer0_outputs(3958) <= not (a xor b);
    layer0_outputs(3959) <= not b;
    layer0_outputs(3960) <= 1'b1;
    layer0_outputs(3961) <= 1'b0;
    layer0_outputs(3962) <= not (a or b);
    layer0_outputs(3963) <= not a;
    layer0_outputs(3964) <= 1'b0;
    layer0_outputs(3965) <= 1'b1;
    layer0_outputs(3966) <= a or b;
    layer0_outputs(3967) <= a or b;
    layer0_outputs(3968) <= a or b;
    layer0_outputs(3969) <= a or b;
    layer0_outputs(3970) <= a or b;
    layer0_outputs(3971) <= not (a xor b);
    layer0_outputs(3972) <= not b or a;
    layer0_outputs(3973) <= not b or a;
    layer0_outputs(3974) <= a and not b;
    layer0_outputs(3975) <= not b or a;
    layer0_outputs(3976) <= not (a xor b);
    layer0_outputs(3977) <= not a or b;
    layer0_outputs(3978) <= not a or b;
    layer0_outputs(3979) <= not a;
    layer0_outputs(3980) <= a xor b;
    layer0_outputs(3981) <= not a or b;
    layer0_outputs(3982) <= not (a and b);
    layer0_outputs(3983) <= not b or a;
    layer0_outputs(3984) <= 1'b1;
    layer0_outputs(3985) <= not (a or b);
    layer0_outputs(3986) <= 1'b1;
    layer0_outputs(3987) <= not (a xor b);
    layer0_outputs(3988) <= 1'b0;
    layer0_outputs(3989) <= not (a or b);
    layer0_outputs(3990) <= 1'b1;
    layer0_outputs(3991) <= not (a and b);
    layer0_outputs(3992) <= 1'b1;
    layer0_outputs(3993) <= not b or a;
    layer0_outputs(3994) <= not (a xor b);
    layer0_outputs(3995) <= not b;
    layer0_outputs(3996) <= not (a and b);
    layer0_outputs(3997) <= a xor b;
    layer0_outputs(3998) <= not (a and b);
    layer0_outputs(3999) <= b and not a;
    layer0_outputs(4000) <= 1'b1;
    layer0_outputs(4001) <= a or b;
    layer0_outputs(4002) <= not a or b;
    layer0_outputs(4003) <= a or b;
    layer0_outputs(4004) <= a or b;
    layer0_outputs(4005) <= not a or b;
    layer0_outputs(4006) <= not (a and b);
    layer0_outputs(4007) <= a and b;
    layer0_outputs(4008) <= not a;
    layer0_outputs(4009) <= not (a xor b);
    layer0_outputs(4010) <= not b;
    layer0_outputs(4011) <= a;
    layer0_outputs(4012) <= a and b;
    layer0_outputs(4013) <= not a or b;
    layer0_outputs(4014) <= a and not b;
    layer0_outputs(4015) <= a xor b;
    layer0_outputs(4016) <= not b or a;
    layer0_outputs(4017) <= a or b;
    layer0_outputs(4018) <= 1'b0;
    layer0_outputs(4019) <= a;
    layer0_outputs(4020) <= a and b;
    layer0_outputs(4021) <= not (a or b);
    layer0_outputs(4022) <= not (a or b);
    layer0_outputs(4023) <= not b;
    layer0_outputs(4024) <= 1'b1;
    layer0_outputs(4025) <= not (a and b);
    layer0_outputs(4026) <= not b;
    layer0_outputs(4027) <= a or b;
    layer0_outputs(4028) <= not a;
    layer0_outputs(4029) <= a xor b;
    layer0_outputs(4030) <= a xor b;
    layer0_outputs(4031) <= a and b;
    layer0_outputs(4032) <= b;
    layer0_outputs(4033) <= not b or a;
    layer0_outputs(4034) <= a and not b;
    layer0_outputs(4035) <= not (a or b);
    layer0_outputs(4036) <= not (a xor b);
    layer0_outputs(4037) <= not b;
    layer0_outputs(4038) <= not a or b;
    layer0_outputs(4039) <= a or b;
    layer0_outputs(4040) <= not a;
    layer0_outputs(4041) <= not (a and b);
    layer0_outputs(4042) <= 1'b1;
    layer0_outputs(4043) <= not a;
    layer0_outputs(4044) <= not b;
    layer0_outputs(4045) <= not (a xor b);
    layer0_outputs(4046) <= not b;
    layer0_outputs(4047) <= not a or b;
    layer0_outputs(4048) <= a;
    layer0_outputs(4049) <= 1'b0;
    layer0_outputs(4050) <= not (a or b);
    layer0_outputs(4051) <= a xor b;
    layer0_outputs(4052) <= 1'b1;
    layer0_outputs(4053) <= a;
    layer0_outputs(4054) <= 1'b1;
    layer0_outputs(4055) <= not (a and b);
    layer0_outputs(4056) <= not a;
    layer0_outputs(4057) <= a and b;
    layer0_outputs(4058) <= 1'b0;
    layer0_outputs(4059) <= b and not a;
    layer0_outputs(4060) <= not b or a;
    layer0_outputs(4061) <= 1'b1;
    layer0_outputs(4062) <= not a;
    layer0_outputs(4063) <= not b or a;
    layer0_outputs(4064) <= 1'b1;
    layer0_outputs(4065) <= not b or a;
    layer0_outputs(4066) <= a or b;
    layer0_outputs(4067) <= 1'b0;
    layer0_outputs(4068) <= 1'b1;
    layer0_outputs(4069) <= a or b;
    layer0_outputs(4070) <= b and not a;
    layer0_outputs(4071) <= a or b;
    layer0_outputs(4072) <= not b;
    layer0_outputs(4073) <= a or b;
    layer0_outputs(4074) <= not (a xor b);
    layer0_outputs(4075) <= a;
    layer0_outputs(4076) <= not b or a;
    layer0_outputs(4077) <= not (a and b);
    layer0_outputs(4078) <= b and not a;
    layer0_outputs(4079) <= not b;
    layer0_outputs(4080) <= a and b;
    layer0_outputs(4081) <= not (a or b);
    layer0_outputs(4082) <= b;
    layer0_outputs(4083) <= a and not b;
    layer0_outputs(4084) <= a and not b;
    layer0_outputs(4085) <= b and not a;
    layer0_outputs(4086) <= b;
    layer0_outputs(4087) <= not (a and b);
    layer0_outputs(4088) <= b;
    layer0_outputs(4089) <= b;
    layer0_outputs(4090) <= a and not b;
    layer0_outputs(4091) <= not a or b;
    layer0_outputs(4092) <= not a or b;
    layer0_outputs(4093) <= a;
    layer0_outputs(4094) <= not (a or b);
    layer0_outputs(4095) <= not (a xor b);
    layer0_outputs(4096) <= not (a or b);
    layer0_outputs(4097) <= b;
    layer0_outputs(4098) <= not (a xor b);
    layer0_outputs(4099) <= a xor b;
    layer0_outputs(4100) <= a and not b;
    layer0_outputs(4101) <= 1'b1;
    layer0_outputs(4102) <= a xor b;
    layer0_outputs(4103) <= not (a or b);
    layer0_outputs(4104) <= not (a xor b);
    layer0_outputs(4105) <= a and b;
    layer0_outputs(4106) <= not (a or b);
    layer0_outputs(4107) <= 1'b1;
    layer0_outputs(4108) <= a;
    layer0_outputs(4109) <= a;
    layer0_outputs(4110) <= 1'b0;
    layer0_outputs(4111) <= a or b;
    layer0_outputs(4112) <= b;
    layer0_outputs(4113) <= not (a and b);
    layer0_outputs(4114) <= not a or b;
    layer0_outputs(4115) <= not (a or b);
    layer0_outputs(4116) <= not a or b;
    layer0_outputs(4117) <= a and not b;
    layer0_outputs(4118) <= b;
    layer0_outputs(4119) <= not (a or b);
    layer0_outputs(4120) <= not (a and b);
    layer0_outputs(4121) <= 1'b1;
    layer0_outputs(4122) <= a or b;
    layer0_outputs(4123) <= a and b;
    layer0_outputs(4124) <= not (a or b);
    layer0_outputs(4125) <= not (a or b);
    layer0_outputs(4126) <= 1'b1;
    layer0_outputs(4127) <= not (a or b);
    layer0_outputs(4128) <= not b or a;
    layer0_outputs(4129) <= not (a or b);
    layer0_outputs(4130) <= a or b;
    layer0_outputs(4131) <= not (a or b);
    layer0_outputs(4132) <= not b or a;
    layer0_outputs(4133) <= not (a or b);
    layer0_outputs(4134) <= a;
    layer0_outputs(4135) <= not (a and b);
    layer0_outputs(4136) <= a;
    layer0_outputs(4137) <= a;
    layer0_outputs(4138) <= a and b;
    layer0_outputs(4139) <= not a or b;
    layer0_outputs(4140) <= a;
    layer0_outputs(4141) <= a;
    layer0_outputs(4142) <= a and b;
    layer0_outputs(4143) <= b;
    layer0_outputs(4144) <= a and b;
    layer0_outputs(4145) <= 1'b1;
    layer0_outputs(4146) <= not b or a;
    layer0_outputs(4147) <= not a or b;
    layer0_outputs(4148) <= not (a or b);
    layer0_outputs(4149) <= a and b;
    layer0_outputs(4150) <= a and b;
    layer0_outputs(4151) <= not b or a;
    layer0_outputs(4152) <= a;
    layer0_outputs(4153) <= not a;
    layer0_outputs(4154) <= not b or a;
    layer0_outputs(4155) <= a;
    layer0_outputs(4156) <= a or b;
    layer0_outputs(4157) <= not b or a;
    layer0_outputs(4158) <= a xor b;
    layer0_outputs(4159) <= a xor b;
    layer0_outputs(4160) <= 1'b1;
    layer0_outputs(4161) <= a and not b;
    layer0_outputs(4162) <= not (a and b);
    layer0_outputs(4163) <= a xor b;
    layer0_outputs(4164) <= 1'b0;
    layer0_outputs(4165) <= b and not a;
    layer0_outputs(4166) <= b;
    layer0_outputs(4167) <= not (a or b);
    layer0_outputs(4168) <= 1'b0;
    layer0_outputs(4169) <= not a;
    layer0_outputs(4170) <= not b;
    layer0_outputs(4171) <= not a or b;
    layer0_outputs(4172) <= not (a and b);
    layer0_outputs(4173) <= a xor b;
    layer0_outputs(4174) <= b;
    layer0_outputs(4175) <= 1'b1;
    layer0_outputs(4176) <= a and b;
    layer0_outputs(4177) <= b;
    layer0_outputs(4178) <= a xor b;
    layer0_outputs(4179) <= not b or a;
    layer0_outputs(4180) <= a or b;
    layer0_outputs(4181) <= not a or b;
    layer0_outputs(4182) <= 1'b0;
    layer0_outputs(4183) <= a xor b;
    layer0_outputs(4184) <= a or b;
    layer0_outputs(4185) <= a and b;
    layer0_outputs(4186) <= not a or b;
    layer0_outputs(4187) <= a and not b;
    layer0_outputs(4188) <= not (a and b);
    layer0_outputs(4189) <= not (a and b);
    layer0_outputs(4190) <= 1'b0;
    layer0_outputs(4191) <= not (a and b);
    layer0_outputs(4192) <= a and b;
    layer0_outputs(4193) <= a or b;
    layer0_outputs(4194) <= a and not b;
    layer0_outputs(4195) <= not (a xor b);
    layer0_outputs(4196) <= b;
    layer0_outputs(4197) <= not (a and b);
    layer0_outputs(4198) <= 1'b1;
    layer0_outputs(4199) <= a and b;
    layer0_outputs(4200) <= not b;
    layer0_outputs(4201) <= not (a and b);
    layer0_outputs(4202) <= not (a or b);
    layer0_outputs(4203) <= 1'b0;
    layer0_outputs(4204) <= not (a xor b);
    layer0_outputs(4205) <= a xor b;
    layer0_outputs(4206) <= a xor b;
    layer0_outputs(4207) <= 1'b0;
    layer0_outputs(4208) <= a xor b;
    layer0_outputs(4209) <= not a;
    layer0_outputs(4210) <= not (a xor b);
    layer0_outputs(4211) <= not (a and b);
    layer0_outputs(4212) <= not (a xor b);
    layer0_outputs(4213) <= b and not a;
    layer0_outputs(4214) <= not b;
    layer0_outputs(4215) <= 1'b0;
    layer0_outputs(4216) <= a or b;
    layer0_outputs(4217) <= b and not a;
    layer0_outputs(4218) <= a and b;
    layer0_outputs(4219) <= not b;
    layer0_outputs(4220) <= not (a or b);
    layer0_outputs(4221) <= not (a and b);
    layer0_outputs(4222) <= not b or a;
    layer0_outputs(4223) <= b;
    layer0_outputs(4224) <= b;
    layer0_outputs(4225) <= not b or a;
    layer0_outputs(4226) <= b;
    layer0_outputs(4227) <= 1'b0;
    layer0_outputs(4228) <= a or b;
    layer0_outputs(4229) <= not a or b;
    layer0_outputs(4230) <= b and not a;
    layer0_outputs(4231) <= not b;
    layer0_outputs(4232) <= not (a or b);
    layer0_outputs(4233) <= a;
    layer0_outputs(4234) <= not b;
    layer0_outputs(4235) <= not b or a;
    layer0_outputs(4236) <= b;
    layer0_outputs(4237) <= not a or b;
    layer0_outputs(4238) <= a;
    layer0_outputs(4239) <= not a;
    layer0_outputs(4240) <= b and not a;
    layer0_outputs(4241) <= not (a or b);
    layer0_outputs(4242) <= a and not b;
    layer0_outputs(4243) <= a xor b;
    layer0_outputs(4244) <= a xor b;
    layer0_outputs(4245) <= not a or b;
    layer0_outputs(4246) <= a or b;
    layer0_outputs(4247) <= a;
    layer0_outputs(4248) <= 1'b1;
    layer0_outputs(4249) <= b;
    layer0_outputs(4250) <= b;
    layer0_outputs(4251) <= not a;
    layer0_outputs(4252) <= not (a and b);
    layer0_outputs(4253) <= not (a and b);
    layer0_outputs(4254) <= a or b;
    layer0_outputs(4255) <= not b or a;
    layer0_outputs(4256) <= a;
    layer0_outputs(4257) <= not b;
    layer0_outputs(4258) <= not (a or b);
    layer0_outputs(4259) <= not (a xor b);
    layer0_outputs(4260) <= b and not a;
    layer0_outputs(4261) <= not a;
    layer0_outputs(4262) <= not b or a;
    layer0_outputs(4263) <= b;
    layer0_outputs(4264) <= a and not b;
    layer0_outputs(4265) <= 1'b1;
    layer0_outputs(4266) <= not (a and b);
    layer0_outputs(4267) <= 1'b1;
    layer0_outputs(4268) <= a;
    layer0_outputs(4269) <= a xor b;
    layer0_outputs(4270) <= not b or a;
    layer0_outputs(4271) <= a or b;
    layer0_outputs(4272) <= not (a or b);
    layer0_outputs(4273) <= a and not b;
    layer0_outputs(4274) <= b;
    layer0_outputs(4275) <= not (a or b);
    layer0_outputs(4276) <= a xor b;
    layer0_outputs(4277) <= not b;
    layer0_outputs(4278) <= b and not a;
    layer0_outputs(4279) <= not (a or b);
    layer0_outputs(4280) <= not a;
    layer0_outputs(4281) <= a xor b;
    layer0_outputs(4282) <= not b or a;
    layer0_outputs(4283) <= a;
    layer0_outputs(4284) <= not (a xor b);
    layer0_outputs(4285) <= b and not a;
    layer0_outputs(4286) <= 1'b1;
    layer0_outputs(4287) <= not a;
    layer0_outputs(4288) <= not (a or b);
    layer0_outputs(4289) <= not (a or b);
    layer0_outputs(4290) <= a;
    layer0_outputs(4291) <= not (a xor b);
    layer0_outputs(4292) <= 1'b1;
    layer0_outputs(4293) <= a and b;
    layer0_outputs(4294) <= a;
    layer0_outputs(4295) <= b;
    layer0_outputs(4296) <= 1'b1;
    layer0_outputs(4297) <= 1'b1;
    layer0_outputs(4298) <= a;
    layer0_outputs(4299) <= not (a or b);
    layer0_outputs(4300) <= 1'b0;
    layer0_outputs(4301) <= not a;
    layer0_outputs(4302) <= b and not a;
    layer0_outputs(4303) <= 1'b1;
    layer0_outputs(4304) <= a and not b;
    layer0_outputs(4305) <= not a;
    layer0_outputs(4306) <= not a;
    layer0_outputs(4307) <= a or b;
    layer0_outputs(4308) <= a or b;
    layer0_outputs(4309) <= not (a and b);
    layer0_outputs(4310) <= 1'b0;
    layer0_outputs(4311) <= 1'b0;
    layer0_outputs(4312) <= not (a and b);
    layer0_outputs(4313) <= not b or a;
    layer0_outputs(4314) <= b and not a;
    layer0_outputs(4315) <= 1'b0;
    layer0_outputs(4316) <= not a;
    layer0_outputs(4317) <= not (a and b);
    layer0_outputs(4318) <= not b;
    layer0_outputs(4319) <= b and not a;
    layer0_outputs(4320) <= not a;
    layer0_outputs(4321) <= b;
    layer0_outputs(4322) <= not a;
    layer0_outputs(4323) <= 1'b0;
    layer0_outputs(4324) <= not (a and b);
    layer0_outputs(4325) <= b and not a;
    layer0_outputs(4326) <= 1'b0;
    layer0_outputs(4327) <= not b;
    layer0_outputs(4328) <= b and not a;
    layer0_outputs(4329) <= not (a and b);
    layer0_outputs(4330) <= not (a and b);
    layer0_outputs(4331) <= not b or a;
    layer0_outputs(4332) <= not b;
    layer0_outputs(4333) <= a or b;
    layer0_outputs(4334) <= not b;
    layer0_outputs(4335) <= b;
    layer0_outputs(4336) <= not (a xor b);
    layer0_outputs(4337) <= a and not b;
    layer0_outputs(4338) <= a or b;
    layer0_outputs(4339) <= not b or a;
    layer0_outputs(4340) <= not a or b;
    layer0_outputs(4341) <= not a;
    layer0_outputs(4342) <= not a or b;
    layer0_outputs(4343) <= not (a or b);
    layer0_outputs(4344) <= a;
    layer0_outputs(4345) <= b;
    layer0_outputs(4346) <= a or b;
    layer0_outputs(4347) <= 1'b1;
    layer0_outputs(4348) <= not a or b;
    layer0_outputs(4349) <= not (a or b);
    layer0_outputs(4350) <= not b or a;
    layer0_outputs(4351) <= 1'b0;
    layer0_outputs(4352) <= b and not a;
    layer0_outputs(4353) <= not b or a;
    layer0_outputs(4354) <= not a;
    layer0_outputs(4355) <= a xor b;
    layer0_outputs(4356) <= a or b;
    layer0_outputs(4357) <= b and not a;
    layer0_outputs(4358) <= not a;
    layer0_outputs(4359) <= a and b;
    layer0_outputs(4360) <= a or b;
    layer0_outputs(4361) <= not (a and b);
    layer0_outputs(4362) <= not (a xor b);
    layer0_outputs(4363) <= b and not a;
    layer0_outputs(4364) <= a and not b;
    layer0_outputs(4365) <= not (a or b);
    layer0_outputs(4366) <= not (a and b);
    layer0_outputs(4367) <= not b or a;
    layer0_outputs(4368) <= not (a or b);
    layer0_outputs(4369) <= not a or b;
    layer0_outputs(4370) <= a and b;
    layer0_outputs(4371) <= a;
    layer0_outputs(4372) <= b;
    layer0_outputs(4373) <= 1'b1;
    layer0_outputs(4374) <= 1'b1;
    layer0_outputs(4375) <= 1'b1;
    layer0_outputs(4376) <= a;
    layer0_outputs(4377) <= 1'b0;
    layer0_outputs(4378) <= 1'b0;
    layer0_outputs(4379) <= not (a and b);
    layer0_outputs(4380) <= a;
    layer0_outputs(4381) <= b and not a;
    layer0_outputs(4382) <= not a or b;
    layer0_outputs(4383) <= not (a and b);
    layer0_outputs(4384) <= not (a or b);
    layer0_outputs(4385) <= b;
    layer0_outputs(4386) <= not a or b;
    layer0_outputs(4387) <= not a or b;
    layer0_outputs(4388) <= a or b;
    layer0_outputs(4389) <= not a or b;
    layer0_outputs(4390) <= a and not b;
    layer0_outputs(4391) <= b;
    layer0_outputs(4392) <= b;
    layer0_outputs(4393) <= 1'b0;
    layer0_outputs(4394) <= a or b;
    layer0_outputs(4395) <= b and not a;
    layer0_outputs(4396) <= not a;
    layer0_outputs(4397) <= a xor b;
    layer0_outputs(4398) <= not a or b;
    layer0_outputs(4399) <= 1'b1;
    layer0_outputs(4400) <= b;
    layer0_outputs(4401) <= not (a or b);
    layer0_outputs(4402) <= b and not a;
    layer0_outputs(4403) <= b;
    layer0_outputs(4404) <= not (a or b);
    layer0_outputs(4405) <= not a or b;
    layer0_outputs(4406) <= not b;
    layer0_outputs(4407) <= a and not b;
    layer0_outputs(4408) <= a;
    layer0_outputs(4409) <= not (a or b);
    layer0_outputs(4410) <= not b;
    layer0_outputs(4411) <= a and not b;
    layer0_outputs(4412) <= a or b;
    layer0_outputs(4413) <= 1'b1;
    layer0_outputs(4414) <= a xor b;
    layer0_outputs(4415) <= a or b;
    layer0_outputs(4416) <= not a;
    layer0_outputs(4417) <= 1'b0;
    layer0_outputs(4418) <= a or b;
    layer0_outputs(4419) <= not (a and b);
    layer0_outputs(4420) <= a or b;
    layer0_outputs(4421) <= not b;
    layer0_outputs(4422) <= a xor b;
    layer0_outputs(4423) <= not b or a;
    layer0_outputs(4424) <= a;
    layer0_outputs(4425) <= not b;
    layer0_outputs(4426) <= a and b;
    layer0_outputs(4427) <= not a;
    layer0_outputs(4428) <= not a or b;
    layer0_outputs(4429) <= not b;
    layer0_outputs(4430) <= 1'b0;
    layer0_outputs(4431) <= not (a or b);
    layer0_outputs(4432) <= a and b;
    layer0_outputs(4433) <= 1'b1;
    layer0_outputs(4434) <= b;
    layer0_outputs(4435) <= a;
    layer0_outputs(4436) <= not (a xor b);
    layer0_outputs(4437) <= not b;
    layer0_outputs(4438) <= a xor b;
    layer0_outputs(4439) <= not a;
    layer0_outputs(4440) <= not (a xor b);
    layer0_outputs(4441) <= not b;
    layer0_outputs(4442) <= a;
    layer0_outputs(4443) <= not (a or b);
    layer0_outputs(4444) <= not (a xor b);
    layer0_outputs(4445) <= not (a or b);
    layer0_outputs(4446) <= not b or a;
    layer0_outputs(4447) <= not a;
    layer0_outputs(4448) <= not (a or b);
    layer0_outputs(4449) <= a or b;
    layer0_outputs(4450) <= a and not b;
    layer0_outputs(4451) <= 1'b1;
    layer0_outputs(4452) <= not b;
    layer0_outputs(4453) <= not b;
    layer0_outputs(4454) <= not (a or b);
    layer0_outputs(4455) <= a xor b;
    layer0_outputs(4456) <= not (a or b);
    layer0_outputs(4457) <= a and not b;
    layer0_outputs(4458) <= a xor b;
    layer0_outputs(4459) <= not a;
    layer0_outputs(4460) <= not (a xor b);
    layer0_outputs(4461) <= not (a or b);
    layer0_outputs(4462) <= not (a or b);
    layer0_outputs(4463) <= not (a or b);
    layer0_outputs(4464) <= a and b;
    layer0_outputs(4465) <= a and not b;
    layer0_outputs(4466) <= a and not b;
    layer0_outputs(4467) <= 1'b1;
    layer0_outputs(4468) <= not (a or b);
    layer0_outputs(4469) <= b;
    layer0_outputs(4470) <= a xor b;
    layer0_outputs(4471) <= a and b;
    layer0_outputs(4472) <= b and not a;
    layer0_outputs(4473) <= not b or a;
    layer0_outputs(4474) <= not a;
    layer0_outputs(4475) <= not b;
    layer0_outputs(4476) <= b;
    layer0_outputs(4477) <= not a;
    layer0_outputs(4478) <= b and not a;
    layer0_outputs(4479) <= 1'b1;
    layer0_outputs(4480) <= not a or b;
    layer0_outputs(4481) <= not a;
    layer0_outputs(4482) <= not (a xor b);
    layer0_outputs(4483) <= a and b;
    layer0_outputs(4484) <= not b;
    layer0_outputs(4485) <= a xor b;
    layer0_outputs(4486) <= b;
    layer0_outputs(4487) <= b and not a;
    layer0_outputs(4488) <= not a;
    layer0_outputs(4489) <= b;
    layer0_outputs(4490) <= 1'b1;
    layer0_outputs(4491) <= 1'b1;
    layer0_outputs(4492) <= a and b;
    layer0_outputs(4493) <= a and not b;
    layer0_outputs(4494) <= b;
    layer0_outputs(4495) <= a;
    layer0_outputs(4496) <= a and not b;
    layer0_outputs(4497) <= not (a xor b);
    layer0_outputs(4498) <= not b or a;
    layer0_outputs(4499) <= not (a and b);
    layer0_outputs(4500) <= a or b;
    layer0_outputs(4501) <= 1'b0;
    layer0_outputs(4502) <= not a;
    layer0_outputs(4503) <= a;
    layer0_outputs(4504) <= a and b;
    layer0_outputs(4505) <= a xor b;
    layer0_outputs(4506) <= not (a or b);
    layer0_outputs(4507) <= a xor b;
    layer0_outputs(4508) <= not (a xor b);
    layer0_outputs(4509) <= not (a and b);
    layer0_outputs(4510) <= not b;
    layer0_outputs(4511) <= not a or b;
    layer0_outputs(4512) <= a or b;
    layer0_outputs(4513) <= not a or b;
    layer0_outputs(4514) <= a and b;
    layer0_outputs(4515) <= a xor b;
    layer0_outputs(4516) <= not a;
    layer0_outputs(4517) <= a and b;
    layer0_outputs(4518) <= a or b;
    layer0_outputs(4519) <= a xor b;
    layer0_outputs(4520) <= b;
    layer0_outputs(4521) <= b and not a;
    layer0_outputs(4522) <= not b;
    layer0_outputs(4523) <= 1'b1;
    layer0_outputs(4524) <= 1'b1;
    layer0_outputs(4525) <= not a or b;
    layer0_outputs(4526) <= not a;
    layer0_outputs(4527) <= not b;
    layer0_outputs(4528) <= not b;
    layer0_outputs(4529) <= not (a and b);
    layer0_outputs(4530) <= a;
    layer0_outputs(4531) <= 1'b0;
    layer0_outputs(4532) <= not b;
    layer0_outputs(4533) <= not b or a;
    layer0_outputs(4534) <= a and b;
    layer0_outputs(4535) <= not a or b;
    layer0_outputs(4536) <= not b;
    layer0_outputs(4537) <= a or b;
    layer0_outputs(4538) <= b;
    layer0_outputs(4539) <= not a;
    layer0_outputs(4540) <= 1'b1;
    layer0_outputs(4541) <= b;
    layer0_outputs(4542) <= not (a xor b);
    layer0_outputs(4543) <= not b or a;
    layer0_outputs(4544) <= a or b;
    layer0_outputs(4545) <= a or b;
    layer0_outputs(4546) <= not a;
    layer0_outputs(4547) <= not a or b;
    layer0_outputs(4548) <= a or b;
    layer0_outputs(4549) <= a;
    layer0_outputs(4550) <= not a or b;
    layer0_outputs(4551) <= a and b;
    layer0_outputs(4552) <= not (a or b);
    layer0_outputs(4553) <= a and b;
    layer0_outputs(4554) <= b;
    layer0_outputs(4555) <= 1'b0;
    layer0_outputs(4556) <= b;
    layer0_outputs(4557) <= not a or b;
    layer0_outputs(4558) <= b;
    layer0_outputs(4559) <= a xor b;
    layer0_outputs(4560) <= not b or a;
    layer0_outputs(4561) <= a;
    layer0_outputs(4562) <= b and not a;
    layer0_outputs(4563) <= 1'b0;
    layer0_outputs(4564) <= 1'b0;
    layer0_outputs(4565) <= a;
    layer0_outputs(4566) <= a or b;
    layer0_outputs(4567) <= b;
    layer0_outputs(4568) <= not b or a;
    layer0_outputs(4569) <= not a or b;
    layer0_outputs(4570) <= not (a and b);
    layer0_outputs(4571) <= b;
    layer0_outputs(4572) <= 1'b1;
    layer0_outputs(4573) <= a xor b;
    layer0_outputs(4574) <= a or b;
    layer0_outputs(4575) <= 1'b0;
    layer0_outputs(4576) <= 1'b0;
    layer0_outputs(4577) <= b;
    layer0_outputs(4578) <= not b or a;
    layer0_outputs(4579) <= not a or b;
    layer0_outputs(4580) <= not a;
    layer0_outputs(4581) <= not b or a;
    layer0_outputs(4582) <= a and not b;
    layer0_outputs(4583) <= not (a or b);
    layer0_outputs(4584) <= a;
    layer0_outputs(4585) <= not b or a;
    layer0_outputs(4586) <= a and not b;
    layer0_outputs(4587) <= not (a or b);
    layer0_outputs(4588) <= 1'b1;
    layer0_outputs(4589) <= a and b;
    layer0_outputs(4590) <= b;
    layer0_outputs(4591) <= not a;
    layer0_outputs(4592) <= not b or a;
    layer0_outputs(4593) <= a;
    layer0_outputs(4594) <= not b;
    layer0_outputs(4595) <= a xor b;
    layer0_outputs(4596) <= a and b;
    layer0_outputs(4597) <= a or b;
    layer0_outputs(4598) <= a;
    layer0_outputs(4599) <= a;
    layer0_outputs(4600) <= a xor b;
    layer0_outputs(4601) <= a and b;
    layer0_outputs(4602) <= not (a or b);
    layer0_outputs(4603) <= b;
    layer0_outputs(4604) <= not b or a;
    layer0_outputs(4605) <= b and not a;
    layer0_outputs(4606) <= a and b;
    layer0_outputs(4607) <= not b;
    layer0_outputs(4608) <= 1'b0;
    layer0_outputs(4609) <= not b or a;
    layer0_outputs(4610) <= a or b;
    layer0_outputs(4611) <= not (a xor b);
    layer0_outputs(4612) <= a and not b;
    layer0_outputs(4613) <= a and b;
    layer0_outputs(4614) <= 1'b1;
    layer0_outputs(4615) <= b and not a;
    layer0_outputs(4616) <= b and not a;
    layer0_outputs(4617) <= not (a or b);
    layer0_outputs(4618) <= a xor b;
    layer0_outputs(4619) <= not (a and b);
    layer0_outputs(4620) <= not a or b;
    layer0_outputs(4621) <= a and b;
    layer0_outputs(4622) <= b;
    layer0_outputs(4623) <= a or b;
    layer0_outputs(4624) <= b;
    layer0_outputs(4625) <= a and b;
    layer0_outputs(4626) <= a;
    layer0_outputs(4627) <= 1'b1;
    layer0_outputs(4628) <= 1'b1;
    layer0_outputs(4629) <= a;
    layer0_outputs(4630) <= not a;
    layer0_outputs(4631) <= not (a or b);
    layer0_outputs(4632) <= not (a xor b);
    layer0_outputs(4633) <= a or b;
    layer0_outputs(4634) <= not (a xor b);
    layer0_outputs(4635) <= not a or b;
    layer0_outputs(4636) <= not (a xor b);
    layer0_outputs(4637) <= a and b;
    layer0_outputs(4638) <= 1'b1;
    layer0_outputs(4639) <= a or b;
    layer0_outputs(4640) <= not (a and b);
    layer0_outputs(4641) <= 1'b0;
    layer0_outputs(4642) <= a xor b;
    layer0_outputs(4643) <= not (a and b);
    layer0_outputs(4644) <= 1'b0;
    layer0_outputs(4645) <= 1'b0;
    layer0_outputs(4646) <= a or b;
    layer0_outputs(4647) <= not b or a;
    layer0_outputs(4648) <= a xor b;
    layer0_outputs(4649) <= not b;
    layer0_outputs(4650) <= not b;
    layer0_outputs(4651) <= b and not a;
    layer0_outputs(4652) <= b;
    layer0_outputs(4653) <= not (a or b);
    layer0_outputs(4654) <= b;
    layer0_outputs(4655) <= b and not a;
    layer0_outputs(4656) <= a;
    layer0_outputs(4657) <= not b;
    layer0_outputs(4658) <= 1'b1;
    layer0_outputs(4659) <= b and not a;
    layer0_outputs(4660) <= a;
    layer0_outputs(4661) <= not a;
    layer0_outputs(4662) <= b and not a;
    layer0_outputs(4663) <= a and b;
    layer0_outputs(4664) <= 1'b1;
    layer0_outputs(4665) <= b and not a;
    layer0_outputs(4666) <= 1'b0;
    layer0_outputs(4667) <= not (a or b);
    layer0_outputs(4668) <= b and not a;
    layer0_outputs(4669) <= a xor b;
    layer0_outputs(4670) <= not (a xor b);
    layer0_outputs(4671) <= not (a or b);
    layer0_outputs(4672) <= 1'b0;
    layer0_outputs(4673) <= a;
    layer0_outputs(4674) <= not a;
    layer0_outputs(4675) <= b;
    layer0_outputs(4676) <= not a;
    layer0_outputs(4677) <= a xor b;
    layer0_outputs(4678) <= not a;
    layer0_outputs(4679) <= a and not b;
    layer0_outputs(4680) <= not (a and b);
    layer0_outputs(4681) <= a and not b;
    layer0_outputs(4682) <= b;
    layer0_outputs(4683) <= b;
    layer0_outputs(4684) <= not a or b;
    layer0_outputs(4685) <= b;
    layer0_outputs(4686) <= 1'b0;
    layer0_outputs(4687) <= not (a and b);
    layer0_outputs(4688) <= not b;
    layer0_outputs(4689) <= 1'b1;
    layer0_outputs(4690) <= 1'b0;
    layer0_outputs(4691) <= not (a xor b);
    layer0_outputs(4692) <= not (a and b);
    layer0_outputs(4693) <= a and not b;
    layer0_outputs(4694) <= 1'b0;
    layer0_outputs(4695) <= 1'b1;
    layer0_outputs(4696) <= b;
    layer0_outputs(4697) <= b;
    layer0_outputs(4698) <= not a or b;
    layer0_outputs(4699) <= 1'b1;
    layer0_outputs(4700) <= a;
    layer0_outputs(4701) <= a;
    layer0_outputs(4702) <= not a or b;
    layer0_outputs(4703) <= not a;
    layer0_outputs(4704) <= not a or b;
    layer0_outputs(4705) <= not (a and b);
    layer0_outputs(4706) <= not b;
    layer0_outputs(4707) <= not a or b;
    layer0_outputs(4708) <= a;
    layer0_outputs(4709) <= b and not a;
    layer0_outputs(4710) <= not (a xor b);
    layer0_outputs(4711) <= not (a and b);
    layer0_outputs(4712) <= not a;
    layer0_outputs(4713) <= a and b;
    layer0_outputs(4714) <= not a or b;
    layer0_outputs(4715) <= a and b;
    layer0_outputs(4716) <= not a or b;
    layer0_outputs(4717) <= not (a or b);
    layer0_outputs(4718) <= not b;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= a and b;
    layer0_outputs(4721) <= not a;
    layer0_outputs(4722) <= 1'b1;
    layer0_outputs(4723) <= not b or a;
    layer0_outputs(4724) <= not (a xor b);
    layer0_outputs(4725) <= b and not a;
    layer0_outputs(4726) <= a or b;
    layer0_outputs(4727) <= b;
    layer0_outputs(4728) <= a and b;
    layer0_outputs(4729) <= a and b;
    layer0_outputs(4730) <= not (a xor b);
    layer0_outputs(4731) <= not a or b;
    layer0_outputs(4732) <= not b or a;
    layer0_outputs(4733) <= not a or b;
    layer0_outputs(4734) <= 1'b0;
    layer0_outputs(4735) <= 1'b0;
    layer0_outputs(4736) <= not b or a;
    layer0_outputs(4737) <= a and b;
    layer0_outputs(4738) <= b;
    layer0_outputs(4739) <= a xor b;
    layer0_outputs(4740) <= 1'b0;
    layer0_outputs(4741) <= not a or b;
    layer0_outputs(4742) <= a or b;
    layer0_outputs(4743) <= not (a and b);
    layer0_outputs(4744) <= a and not b;
    layer0_outputs(4745) <= b;
    layer0_outputs(4746) <= 1'b1;
    layer0_outputs(4747) <= a and not b;
    layer0_outputs(4748) <= b;
    layer0_outputs(4749) <= a;
    layer0_outputs(4750) <= a or b;
    layer0_outputs(4751) <= a xor b;
    layer0_outputs(4752) <= a;
    layer0_outputs(4753) <= a or b;
    layer0_outputs(4754) <= a and b;
    layer0_outputs(4755) <= b and not a;
    layer0_outputs(4756) <= a;
    layer0_outputs(4757) <= not (a xor b);
    layer0_outputs(4758) <= a;
    layer0_outputs(4759) <= 1'b0;
    layer0_outputs(4760) <= not a or b;
    layer0_outputs(4761) <= a xor b;
    layer0_outputs(4762) <= not (a xor b);
    layer0_outputs(4763) <= not b;
    layer0_outputs(4764) <= not (a and b);
    layer0_outputs(4765) <= a or b;
    layer0_outputs(4766) <= not b;
    layer0_outputs(4767) <= a;
    layer0_outputs(4768) <= not a or b;
    layer0_outputs(4769) <= a xor b;
    layer0_outputs(4770) <= a xor b;
    layer0_outputs(4771) <= a or b;
    layer0_outputs(4772) <= a;
    layer0_outputs(4773) <= a and b;
    layer0_outputs(4774) <= 1'b0;
    layer0_outputs(4775) <= a;
    layer0_outputs(4776) <= not (a xor b);
    layer0_outputs(4777) <= a and b;
    layer0_outputs(4778) <= not a;
    layer0_outputs(4779) <= 1'b1;
    layer0_outputs(4780) <= 1'b1;
    layer0_outputs(4781) <= not (a and b);
    layer0_outputs(4782) <= not b or a;
    layer0_outputs(4783) <= a and not b;
    layer0_outputs(4784) <= not b or a;
    layer0_outputs(4785) <= b;
    layer0_outputs(4786) <= not b;
    layer0_outputs(4787) <= 1'b0;
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= b;
    layer0_outputs(4790) <= 1'b0;
    layer0_outputs(4791) <= a and not b;
    layer0_outputs(4792) <= a or b;
    layer0_outputs(4793) <= 1'b1;
    layer0_outputs(4794) <= not b or a;
    layer0_outputs(4795) <= b;
    layer0_outputs(4796) <= b;
    layer0_outputs(4797) <= not (a and b);
    layer0_outputs(4798) <= not (a and b);
    layer0_outputs(4799) <= 1'b1;
    layer0_outputs(4800) <= a and b;
    layer0_outputs(4801) <= not a;
    layer0_outputs(4802) <= not (a or b);
    layer0_outputs(4803) <= b;
    layer0_outputs(4804) <= a and not b;
    layer0_outputs(4805) <= not (a xor b);
    layer0_outputs(4806) <= b and not a;
    layer0_outputs(4807) <= not a;
    layer0_outputs(4808) <= 1'b0;
    layer0_outputs(4809) <= b;
    layer0_outputs(4810) <= not (a xor b);
    layer0_outputs(4811) <= b;
    layer0_outputs(4812) <= a and not b;
    layer0_outputs(4813) <= b;
    layer0_outputs(4814) <= 1'b0;
    layer0_outputs(4815) <= 1'b0;
    layer0_outputs(4816) <= not (a or b);
    layer0_outputs(4817) <= a and b;
    layer0_outputs(4818) <= b and not a;
    layer0_outputs(4819) <= not (a and b);
    layer0_outputs(4820) <= not (a and b);
    layer0_outputs(4821) <= a and b;
    layer0_outputs(4822) <= not b or a;
    layer0_outputs(4823) <= not (a or b);
    layer0_outputs(4824) <= 1'b0;
    layer0_outputs(4825) <= not a;
    layer0_outputs(4826) <= a and b;
    layer0_outputs(4827) <= b and not a;
    layer0_outputs(4828) <= 1'b0;
    layer0_outputs(4829) <= b and not a;
    layer0_outputs(4830) <= a and not b;
    layer0_outputs(4831) <= 1'b1;
    layer0_outputs(4832) <= not b;
    layer0_outputs(4833) <= not b;
    layer0_outputs(4834) <= not (a xor b);
    layer0_outputs(4835) <= not (a and b);
    layer0_outputs(4836) <= not (a xor b);
    layer0_outputs(4837) <= 1'b1;
    layer0_outputs(4838) <= a or b;
    layer0_outputs(4839) <= a xor b;
    layer0_outputs(4840) <= 1'b1;
    layer0_outputs(4841) <= a xor b;
    layer0_outputs(4842) <= not a;
    layer0_outputs(4843) <= b and not a;
    layer0_outputs(4844) <= not b or a;
    layer0_outputs(4845) <= a;
    layer0_outputs(4846) <= not (a xor b);
    layer0_outputs(4847) <= 1'b0;
    layer0_outputs(4848) <= a and not b;
    layer0_outputs(4849) <= not b;
    layer0_outputs(4850) <= a;
    layer0_outputs(4851) <= not b;
    layer0_outputs(4852) <= b;
    layer0_outputs(4853) <= not b;
    layer0_outputs(4854) <= not (a and b);
    layer0_outputs(4855) <= a and b;
    layer0_outputs(4856) <= a;
    layer0_outputs(4857) <= not a;
    layer0_outputs(4858) <= not (a and b);
    layer0_outputs(4859) <= not b;
    layer0_outputs(4860) <= a and not b;
    layer0_outputs(4861) <= b and not a;
    layer0_outputs(4862) <= not a;
    layer0_outputs(4863) <= a and not b;
    layer0_outputs(4864) <= not (a xor b);
    layer0_outputs(4865) <= not (a and b);
    layer0_outputs(4866) <= 1'b1;
    layer0_outputs(4867) <= a xor b;
    layer0_outputs(4868) <= 1'b0;
    layer0_outputs(4869) <= 1'b1;
    layer0_outputs(4870) <= 1'b1;
    layer0_outputs(4871) <= not b;
    layer0_outputs(4872) <= b;
    layer0_outputs(4873) <= 1'b0;
    layer0_outputs(4874) <= not a;
    layer0_outputs(4875) <= not (a and b);
    layer0_outputs(4876) <= 1'b0;
    layer0_outputs(4877) <= a;
    layer0_outputs(4878) <= not a;
    layer0_outputs(4879) <= a xor b;
    layer0_outputs(4880) <= a and b;
    layer0_outputs(4881) <= not b or a;
    layer0_outputs(4882) <= not a or b;
    layer0_outputs(4883) <= not (a xor b);
    layer0_outputs(4884) <= not a;
    layer0_outputs(4885) <= a and not b;
    layer0_outputs(4886) <= not (a or b);
    layer0_outputs(4887) <= 1'b1;
    layer0_outputs(4888) <= b;
    layer0_outputs(4889) <= 1'b1;
    layer0_outputs(4890) <= a or b;
    layer0_outputs(4891) <= 1'b0;
    layer0_outputs(4892) <= b and not a;
    layer0_outputs(4893) <= b and not a;
    layer0_outputs(4894) <= not a;
    layer0_outputs(4895) <= 1'b0;
    layer0_outputs(4896) <= not a;
    layer0_outputs(4897) <= not a;
    layer0_outputs(4898) <= not b or a;
    layer0_outputs(4899) <= not b;
    layer0_outputs(4900) <= a;
    layer0_outputs(4901) <= a and b;
    layer0_outputs(4902) <= a xor b;
    layer0_outputs(4903) <= not (a xor b);
    layer0_outputs(4904) <= 1'b1;
    layer0_outputs(4905) <= not b or a;
    layer0_outputs(4906) <= b;
    layer0_outputs(4907) <= not (a and b);
    layer0_outputs(4908) <= not b or a;
    layer0_outputs(4909) <= a and not b;
    layer0_outputs(4910) <= 1'b1;
    layer0_outputs(4911) <= a or b;
    layer0_outputs(4912) <= not a or b;
    layer0_outputs(4913) <= not a or b;
    layer0_outputs(4914) <= b and not a;
    layer0_outputs(4915) <= b and not a;
    layer0_outputs(4916) <= not (a or b);
    layer0_outputs(4917) <= a xor b;
    layer0_outputs(4918) <= not a;
    layer0_outputs(4919) <= a or b;
    layer0_outputs(4920) <= 1'b1;
    layer0_outputs(4921) <= not (a or b);
    layer0_outputs(4922) <= not b or a;
    layer0_outputs(4923) <= not a;
    layer0_outputs(4924) <= not (a xor b);
    layer0_outputs(4925) <= 1'b0;
    layer0_outputs(4926) <= a and b;
    layer0_outputs(4927) <= a and not b;
    layer0_outputs(4928) <= a or b;
    layer0_outputs(4929) <= 1'b0;
    layer0_outputs(4930) <= a or b;
    layer0_outputs(4931) <= 1'b0;
    layer0_outputs(4932) <= not (a xor b);
    layer0_outputs(4933) <= not b or a;
    layer0_outputs(4934) <= 1'b0;
    layer0_outputs(4935) <= not (a or b);
    layer0_outputs(4936) <= 1'b1;
    layer0_outputs(4937) <= 1'b0;
    layer0_outputs(4938) <= a or b;
    layer0_outputs(4939) <= a or b;
    layer0_outputs(4940) <= a;
    layer0_outputs(4941) <= not a;
    layer0_outputs(4942) <= a or b;
    layer0_outputs(4943) <= not b;
    layer0_outputs(4944) <= 1'b1;
    layer0_outputs(4945) <= 1'b1;
    layer0_outputs(4946) <= not b or a;
    layer0_outputs(4947) <= b;
    layer0_outputs(4948) <= not b;
    layer0_outputs(4949) <= not b or a;
    layer0_outputs(4950) <= not (a and b);
    layer0_outputs(4951) <= b and not a;
    layer0_outputs(4952) <= 1'b1;
    layer0_outputs(4953) <= a;
    layer0_outputs(4954) <= not b or a;
    layer0_outputs(4955) <= 1'b1;
    layer0_outputs(4956) <= a xor b;
    layer0_outputs(4957) <= a;
    layer0_outputs(4958) <= a;
    layer0_outputs(4959) <= not a;
    layer0_outputs(4960) <= not a;
    layer0_outputs(4961) <= a and not b;
    layer0_outputs(4962) <= not (a and b);
    layer0_outputs(4963) <= b;
    layer0_outputs(4964) <= not a or b;
    layer0_outputs(4965) <= b;
    layer0_outputs(4966) <= a and b;
    layer0_outputs(4967) <= not (a or b);
    layer0_outputs(4968) <= a and not b;
    layer0_outputs(4969) <= not (a xor b);
    layer0_outputs(4970) <= b and not a;
    layer0_outputs(4971) <= a and not b;
    layer0_outputs(4972) <= a and b;
    layer0_outputs(4973) <= a;
    layer0_outputs(4974) <= a or b;
    layer0_outputs(4975) <= b;
    layer0_outputs(4976) <= not (a xor b);
    layer0_outputs(4977) <= a or b;
    layer0_outputs(4978) <= a and b;
    layer0_outputs(4979) <= not a;
    layer0_outputs(4980) <= b;
    layer0_outputs(4981) <= a or b;
    layer0_outputs(4982) <= not (a or b);
    layer0_outputs(4983) <= 1'b1;
    layer0_outputs(4984) <= 1'b0;
    layer0_outputs(4985) <= b;
    layer0_outputs(4986) <= b and not a;
    layer0_outputs(4987) <= a xor b;
    layer0_outputs(4988) <= 1'b0;
    layer0_outputs(4989) <= b;
    layer0_outputs(4990) <= a;
    layer0_outputs(4991) <= a;
    layer0_outputs(4992) <= not a or b;
    layer0_outputs(4993) <= not b;
    layer0_outputs(4994) <= a and not b;
    layer0_outputs(4995) <= not b or a;
    layer0_outputs(4996) <= a;
    layer0_outputs(4997) <= a and not b;
    layer0_outputs(4998) <= not b or a;
    layer0_outputs(4999) <= not b or a;
    layer0_outputs(5000) <= not b;
    layer0_outputs(5001) <= 1'b0;
    layer0_outputs(5002) <= b;
    layer0_outputs(5003) <= not b or a;
    layer0_outputs(5004) <= a and not b;
    layer0_outputs(5005) <= not (a and b);
    layer0_outputs(5006) <= 1'b1;
    layer0_outputs(5007) <= b;
    layer0_outputs(5008) <= b;
    layer0_outputs(5009) <= not (a and b);
    layer0_outputs(5010) <= not b or a;
    layer0_outputs(5011) <= a and b;
    layer0_outputs(5012) <= not b or a;
    layer0_outputs(5013) <= a and b;
    layer0_outputs(5014) <= not (a and b);
    layer0_outputs(5015) <= a xor b;
    layer0_outputs(5016) <= not b;
    layer0_outputs(5017) <= 1'b1;
    layer0_outputs(5018) <= not b;
    layer0_outputs(5019) <= not b;
    layer0_outputs(5020) <= 1'b1;
    layer0_outputs(5021) <= b;
    layer0_outputs(5022) <= not (a xor b);
    layer0_outputs(5023) <= 1'b0;
    layer0_outputs(5024) <= not b;
    layer0_outputs(5025) <= 1'b0;
    layer0_outputs(5026) <= not (a and b);
    layer0_outputs(5027) <= not (a or b);
    layer0_outputs(5028) <= not a or b;
    layer0_outputs(5029) <= 1'b1;
    layer0_outputs(5030) <= b and not a;
    layer0_outputs(5031) <= not (a and b);
    layer0_outputs(5032) <= a or b;
    layer0_outputs(5033) <= 1'b1;
    layer0_outputs(5034) <= 1'b1;
    layer0_outputs(5035) <= not (a and b);
    layer0_outputs(5036) <= not (a or b);
    layer0_outputs(5037) <= 1'b1;
    layer0_outputs(5038) <= not b;
    layer0_outputs(5039) <= 1'b0;
    layer0_outputs(5040) <= not (a or b);
    layer0_outputs(5041) <= a or b;
    layer0_outputs(5042) <= not b;
    layer0_outputs(5043) <= not (a xor b);
    layer0_outputs(5044) <= 1'b1;
    layer0_outputs(5045) <= not b;
    layer0_outputs(5046) <= 1'b0;
    layer0_outputs(5047) <= a;
    layer0_outputs(5048) <= b;
    layer0_outputs(5049) <= not (a or b);
    layer0_outputs(5050) <= a;
    layer0_outputs(5051) <= 1'b1;
    layer0_outputs(5052) <= a and not b;
    layer0_outputs(5053) <= a xor b;
    layer0_outputs(5054) <= not b;
    layer0_outputs(5055) <= a and not b;
    layer0_outputs(5056) <= b and not a;
    layer0_outputs(5057) <= not (a and b);
    layer0_outputs(5058) <= a or b;
    layer0_outputs(5059) <= not a;
    layer0_outputs(5060) <= 1'b1;
    layer0_outputs(5061) <= not a or b;
    layer0_outputs(5062) <= 1'b0;
    layer0_outputs(5063) <= a;
    layer0_outputs(5064) <= a or b;
    layer0_outputs(5065) <= not b or a;
    layer0_outputs(5066) <= 1'b0;
    layer0_outputs(5067) <= not a;
    layer0_outputs(5068) <= not b or a;
    layer0_outputs(5069) <= not (a and b);
    layer0_outputs(5070) <= not (a or b);
    layer0_outputs(5071) <= a;
    layer0_outputs(5072) <= not (a or b);
    layer0_outputs(5073) <= not b;
    layer0_outputs(5074) <= b;
    layer0_outputs(5075) <= a and not b;
    layer0_outputs(5076) <= not (a xor b);
    layer0_outputs(5077) <= b and not a;
    layer0_outputs(5078) <= not a or b;
    layer0_outputs(5079) <= b;
    layer0_outputs(5080) <= b and not a;
    layer0_outputs(5081) <= b and not a;
    layer0_outputs(5082) <= 1'b1;
    layer0_outputs(5083) <= not (a xor b);
    layer0_outputs(5084) <= a and b;
    layer0_outputs(5085) <= 1'b1;
    layer0_outputs(5086) <= not a;
    layer0_outputs(5087) <= a and not b;
    layer0_outputs(5088) <= a xor b;
    layer0_outputs(5089) <= not (a xor b);
    layer0_outputs(5090) <= b and not a;
    layer0_outputs(5091) <= not b;
    layer0_outputs(5092) <= a and b;
    layer0_outputs(5093) <= a and not b;
    layer0_outputs(5094) <= a or b;
    layer0_outputs(5095) <= b;
    layer0_outputs(5096) <= 1'b0;
    layer0_outputs(5097) <= a and not b;
    layer0_outputs(5098) <= 1'b0;
    layer0_outputs(5099) <= not (a and b);
    layer0_outputs(5100) <= not b;
    layer0_outputs(5101) <= 1'b0;
    layer0_outputs(5102) <= not (a and b);
    layer0_outputs(5103) <= not (a or b);
    layer0_outputs(5104) <= b;
    layer0_outputs(5105) <= not (a or b);
    layer0_outputs(5106) <= not a;
    layer0_outputs(5107) <= not (a or b);
    layer0_outputs(5108) <= a or b;
    layer0_outputs(5109) <= not b or a;
    layer0_outputs(5110) <= a and not b;
    layer0_outputs(5111) <= a;
    layer0_outputs(5112) <= a and b;
    layer0_outputs(5113) <= 1'b0;
    layer0_outputs(5114) <= a and not b;
    layer0_outputs(5115) <= a and not b;
    layer0_outputs(5116) <= not (a or b);
    layer0_outputs(5117) <= b and not a;
    layer0_outputs(5118) <= 1'b1;
    layer0_outputs(5119) <= not a or b;
    layer0_outputs(5120) <= not a;
    layer0_outputs(5121) <= a;
    layer0_outputs(5122) <= not a or b;
    layer0_outputs(5123) <= 1'b0;
    layer0_outputs(5124) <= not (a xor b);
    layer0_outputs(5125) <= not b or a;
    layer0_outputs(5126) <= not (a xor b);
    layer0_outputs(5127) <= a and b;
    layer0_outputs(5128) <= 1'b0;
    layer0_outputs(5129) <= a xor b;
    layer0_outputs(5130) <= a or b;
    layer0_outputs(5131) <= b and not a;
    layer0_outputs(5132) <= not b;
    layer0_outputs(5133) <= not b or a;
    layer0_outputs(5134) <= a;
    layer0_outputs(5135) <= b and not a;
    layer0_outputs(5136) <= a or b;
    layer0_outputs(5137) <= a and not b;
    layer0_outputs(5138) <= 1'b0;
    layer0_outputs(5139) <= 1'b1;
    layer0_outputs(5140) <= a and b;
    layer0_outputs(5141) <= not b;
    layer0_outputs(5142) <= not (a or b);
    layer0_outputs(5143) <= not (a or b);
    layer0_outputs(5144) <= not b or a;
    layer0_outputs(5145) <= 1'b0;
    layer0_outputs(5146) <= not (a and b);
    layer0_outputs(5147) <= a or b;
    layer0_outputs(5148) <= a or b;
    layer0_outputs(5149) <= not b or a;
    layer0_outputs(5150) <= 1'b1;
    layer0_outputs(5151) <= not b or a;
    layer0_outputs(5152) <= b;
    layer0_outputs(5153) <= not a or b;
    layer0_outputs(5154) <= not a or b;
    layer0_outputs(5155) <= b;
    layer0_outputs(5156) <= a;
    layer0_outputs(5157) <= not b or a;
    layer0_outputs(5158) <= not a;
    layer0_outputs(5159) <= not b or a;
    layer0_outputs(5160) <= not a or b;
    layer0_outputs(5161) <= not b or a;
    layer0_outputs(5162) <= not b;
    layer0_outputs(5163) <= b;
    layer0_outputs(5164) <= 1'b1;
    layer0_outputs(5165) <= b and not a;
    layer0_outputs(5166) <= a xor b;
    layer0_outputs(5167) <= not b;
    layer0_outputs(5168) <= not b or a;
    layer0_outputs(5169) <= a xor b;
    layer0_outputs(5170) <= a or b;
    layer0_outputs(5171) <= 1'b1;
    layer0_outputs(5172) <= not a or b;
    layer0_outputs(5173) <= b;
    layer0_outputs(5174) <= b;
    layer0_outputs(5175) <= b and not a;
    layer0_outputs(5176) <= not a;
    layer0_outputs(5177) <= not a or b;
    layer0_outputs(5178) <= b and not a;
    layer0_outputs(5179) <= a and b;
    layer0_outputs(5180) <= b;
    layer0_outputs(5181) <= not a or b;
    layer0_outputs(5182) <= not a;
    layer0_outputs(5183) <= not a or b;
    layer0_outputs(5184) <= b;
    layer0_outputs(5185) <= a and not b;
    layer0_outputs(5186) <= a xor b;
    layer0_outputs(5187) <= b and not a;
    layer0_outputs(5188) <= a;
    layer0_outputs(5189) <= a xor b;
    layer0_outputs(5190) <= b;
    layer0_outputs(5191) <= not b or a;
    layer0_outputs(5192) <= not (a or b);
    layer0_outputs(5193) <= a xor b;
    layer0_outputs(5194) <= 1'b0;
    layer0_outputs(5195) <= b and not a;
    layer0_outputs(5196) <= 1'b1;
    layer0_outputs(5197) <= not a;
    layer0_outputs(5198) <= 1'b1;
    layer0_outputs(5199) <= a or b;
    layer0_outputs(5200) <= a and b;
    layer0_outputs(5201) <= a or b;
    layer0_outputs(5202) <= a and not b;
    layer0_outputs(5203) <= not b;
    layer0_outputs(5204) <= 1'b0;
    layer0_outputs(5205) <= not (a xor b);
    layer0_outputs(5206) <= not b;
    layer0_outputs(5207) <= 1'b0;
    layer0_outputs(5208) <= not (a and b);
    layer0_outputs(5209) <= 1'b1;
    layer0_outputs(5210) <= not a or b;
    layer0_outputs(5211) <= a and not b;
    layer0_outputs(5212) <= b;
    layer0_outputs(5213) <= not a;
    layer0_outputs(5214) <= b and not a;
    layer0_outputs(5215) <= a or b;
    layer0_outputs(5216) <= a xor b;
    layer0_outputs(5217) <= 1'b1;
    layer0_outputs(5218) <= not a or b;
    layer0_outputs(5219) <= b and not a;
    layer0_outputs(5220) <= 1'b1;
    layer0_outputs(5221) <= b;
    layer0_outputs(5222) <= a xor b;
    layer0_outputs(5223) <= not b or a;
    layer0_outputs(5224) <= not (a or b);
    layer0_outputs(5225) <= a and not b;
    layer0_outputs(5226) <= a and not b;
    layer0_outputs(5227) <= b and not a;
    layer0_outputs(5228) <= a and not b;
    layer0_outputs(5229) <= not b or a;
    layer0_outputs(5230) <= not (a xor b);
    layer0_outputs(5231) <= a xor b;
    layer0_outputs(5232) <= b and not a;
    layer0_outputs(5233) <= a xor b;
    layer0_outputs(5234) <= 1'b1;
    layer0_outputs(5235) <= not (a xor b);
    layer0_outputs(5236) <= a or b;
    layer0_outputs(5237) <= a xor b;
    layer0_outputs(5238) <= 1'b0;
    layer0_outputs(5239) <= a or b;
    layer0_outputs(5240) <= not b or a;
    layer0_outputs(5241) <= not a;
    layer0_outputs(5242) <= not b or a;
    layer0_outputs(5243) <= not (a or b);
    layer0_outputs(5244) <= not (a and b);
    layer0_outputs(5245) <= a or b;
    layer0_outputs(5246) <= 1'b1;
    layer0_outputs(5247) <= 1'b1;
    layer0_outputs(5248) <= b and not a;
    layer0_outputs(5249) <= a and not b;
    layer0_outputs(5250) <= 1'b0;
    layer0_outputs(5251) <= not (a xor b);
    layer0_outputs(5252) <= a and b;
    layer0_outputs(5253) <= not (a xor b);
    layer0_outputs(5254) <= 1'b1;
    layer0_outputs(5255) <= not b or a;
    layer0_outputs(5256) <= not a or b;
    layer0_outputs(5257) <= not b;
    layer0_outputs(5258) <= 1'b0;
    layer0_outputs(5259) <= not b;
    layer0_outputs(5260) <= a xor b;
    layer0_outputs(5261) <= 1'b1;
    layer0_outputs(5262) <= 1'b0;
    layer0_outputs(5263) <= not b or a;
    layer0_outputs(5264) <= not (a xor b);
    layer0_outputs(5265) <= 1'b1;
    layer0_outputs(5266) <= not a or b;
    layer0_outputs(5267) <= not b;
    layer0_outputs(5268) <= not b or a;
    layer0_outputs(5269) <= 1'b0;
    layer0_outputs(5270) <= 1'b0;
    layer0_outputs(5271) <= not b or a;
    layer0_outputs(5272) <= b;
    layer0_outputs(5273) <= a;
    layer0_outputs(5274) <= 1'b0;
    layer0_outputs(5275) <= 1'b1;
    layer0_outputs(5276) <= not a or b;
    layer0_outputs(5277) <= not (a xor b);
    layer0_outputs(5278) <= not (a xor b);
    layer0_outputs(5279) <= not a or b;
    layer0_outputs(5280) <= a;
    layer0_outputs(5281) <= a and not b;
    layer0_outputs(5282) <= a xor b;
    layer0_outputs(5283) <= a;
    layer0_outputs(5284) <= 1'b0;
    layer0_outputs(5285) <= a;
    layer0_outputs(5286) <= b;
    layer0_outputs(5287) <= not (a or b);
    layer0_outputs(5288) <= 1'b0;
    layer0_outputs(5289) <= not a or b;
    layer0_outputs(5290) <= a and not b;
    layer0_outputs(5291) <= a;
    layer0_outputs(5292) <= a xor b;
    layer0_outputs(5293) <= not a;
    layer0_outputs(5294) <= a or b;
    layer0_outputs(5295) <= 1'b0;
    layer0_outputs(5296) <= a xor b;
    layer0_outputs(5297) <= 1'b1;
    layer0_outputs(5298) <= not (a or b);
    layer0_outputs(5299) <= a xor b;
    layer0_outputs(5300) <= a or b;
    layer0_outputs(5301) <= b and not a;
    layer0_outputs(5302) <= not (a xor b);
    layer0_outputs(5303) <= a or b;
    layer0_outputs(5304) <= 1'b1;
    layer0_outputs(5305) <= a;
    layer0_outputs(5306) <= not (a xor b);
    layer0_outputs(5307) <= not a;
    layer0_outputs(5308) <= 1'b1;
    layer0_outputs(5309) <= not (a or b);
    layer0_outputs(5310) <= 1'b0;
    layer0_outputs(5311) <= a and b;
    layer0_outputs(5312) <= b;
    layer0_outputs(5313) <= not (a xor b);
    layer0_outputs(5314) <= not b or a;
    layer0_outputs(5315) <= b;
    layer0_outputs(5316) <= not a or b;
    layer0_outputs(5317) <= 1'b1;
    layer0_outputs(5318) <= not (a or b);
    layer0_outputs(5319) <= not a or b;
    layer0_outputs(5320) <= a or b;
    layer0_outputs(5321) <= not b;
    layer0_outputs(5322) <= not (a or b);
    layer0_outputs(5323) <= not (a or b);
    layer0_outputs(5324) <= not b or a;
    layer0_outputs(5325) <= b;
    layer0_outputs(5326) <= not a or b;
    layer0_outputs(5327) <= a or b;
    layer0_outputs(5328) <= not b;
    layer0_outputs(5329) <= not b or a;
    layer0_outputs(5330) <= a and not b;
    layer0_outputs(5331) <= not (a xor b);
    layer0_outputs(5332) <= not (a and b);
    layer0_outputs(5333) <= a;
    layer0_outputs(5334) <= 1'b1;
    layer0_outputs(5335) <= not a;
    layer0_outputs(5336) <= 1'b0;
    layer0_outputs(5337) <= a or b;
    layer0_outputs(5338) <= not b or a;
    layer0_outputs(5339) <= 1'b0;
    layer0_outputs(5340) <= not (a xor b);
    layer0_outputs(5341) <= a or b;
    layer0_outputs(5342) <= not a or b;
    layer0_outputs(5343) <= a and b;
    layer0_outputs(5344) <= b;
    layer0_outputs(5345) <= a and b;
    layer0_outputs(5346) <= a and not b;
    layer0_outputs(5347) <= 1'b0;
    layer0_outputs(5348) <= not (a or b);
    layer0_outputs(5349) <= a and not b;
    layer0_outputs(5350) <= not a;
    layer0_outputs(5351) <= a or b;
    layer0_outputs(5352) <= b and not a;
    layer0_outputs(5353) <= not (a and b);
    layer0_outputs(5354) <= a and b;
    layer0_outputs(5355) <= not a;
    layer0_outputs(5356) <= a xor b;
    layer0_outputs(5357) <= b and not a;
    layer0_outputs(5358) <= not (a or b);
    layer0_outputs(5359) <= not (a xor b);
    layer0_outputs(5360) <= not a;
    layer0_outputs(5361) <= not (a or b);
    layer0_outputs(5362) <= b;
    layer0_outputs(5363) <= not b;
    layer0_outputs(5364) <= 1'b1;
    layer0_outputs(5365) <= a;
    layer0_outputs(5366) <= not (a or b);
    layer0_outputs(5367) <= not a or b;
    layer0_outputs(5368) <= not (a or b);
    layer0_outputs(5369) <= a and b;
    layer0_outputs(5370) <= a and b;
    layer0_outputs(5371) <= a or b;
    layer0_outputs(5372) <= 1'b1;
    layer0_outputs(5373) <= a or b;
    layer0_outputs(5374) <= not b or a;
    layer0_outputs(5375) <= not (a xor b);
    layer0_outputs(5376) <= 1'b1;
    layer0_outputs(5377) <= 1'b0;
    layer0_outputs(5378) <= 1'b1;
    layer0_outputs(5379) <= not a or b;
    layer0_outputs(5380) <= not b or a;
    layer0_outputs(5381) <= not b;
    layer0_outputs(5382) <= a and not b;
    layer0_outputs(5383) <= 1'b0;
    layer0_outputs(5384) <= not a;
    layer0_outputs(5385) <= a xor b;
    layer0_outputs(5386) <= not b or a;
    layer0_outputs(5387) <= a;
    layer0_outputs(5388) <= a and b;
    layer0_outputs(5389) <= 1'b0;
    layer0_outputs(5390) <= not b or a;
    layer0_outputs(5391) <= b;
    layer0_outputs(5392) <= not a;
    layer0_outputs(5393) <= not (a or b);
    layer0_outputs(5394) <= 1'b1;
    layer0_outputs(5395) <= not b;
    layer0_outputs(5396) <= not a or b;
    layer0_outputs(5397) <= a;
    layer0_outputs(5398) <= 1'b1;
    layer0_outputs(5399) <= a and not b;
    layer0_outputs(5400) <= not b;
    layer0_outputs(5401) <= not a;
    layer0_outputs(5402) <= not a;
    layer0_outputs(5403) <= b and not a;
    layer0_outputs(5404) <= not (a and b);
    layer0_outputs(5405) <= a;
    layer0_outputs(5406) <= not a or b;
    layer0_outputs(5407) <= not a;
    layer0_outputs(5408) <= 1'b0;
    layer0_outputs(5409) <= not b or a;
    layer0_outputs(5410) <= not (a or b);
    layer0_outputs(5411) <= not (a and b);
    layer0_outputs(5412) <= a;
    layer0_outputs(5413) <= b;
    layer0_outputs(5414) <= a or b;
    layer0_outputs(5415) <= a xor b;
    layer0_outputs(5416) <= a;
    layer0_outputs(5417) <= a and not b;
    layer0_outputs(5418) <= not (a xor b);
    layer0_outputs(5419) <= a and b;
    layer0_outputs(5420) <= a and b;
    layer0_outputs(5421) <= a and b;
    layer0_outputs(5422) <= not a;
    layer0_outputs(5423) <= b;
    layer0_outputs(5424) <= 1'b1;
    layer0_outputs(5425) <= not a;
    layer0_outputs(5426) <= a and b;
    layer0_outputs(5427) <= not b;
    layer0_outputs(5428) <= a xor b;
    layer0_outputs(5429) <= not a;
    layer0_outputs(5430) <= not b;
    layer0_outputs(5431) <= not b;
    layer0_outputs(5432) <= b;
    layer0_outputs(5433) <= a xor b;
    layer0_outputs(5434) <= b and not a;
    layer0_outputs(5435) <= not a or b;
    layer0_outputs(5436) <= a;
    layer0_outputs(5437) <= a xor b;
    layer0_outputs(5438) <= a and not b;
    layer0_outputs(5439) <= 1'b0;
    layer0_outputs(5440) <= not b;
    layer0_outputs(5441) <= 1'b0;
    layer0_outputs(5442) <= not a or b;
    layer0_outputs(5443) <= not (a xor b);
    layer0_outputs(5444) <= not b;
    layer0_outputs(5445) <= a xor b;
    layer0_outputs(5446) <= a or b;
    layer0_outputs(5447) <= a and not b;
    layer0_outputs(5448) <= a or b;
    layer0_outputs(5449) <= a and not b;
    layer0_outputs(5450) <= not (a and b);
    layer0_outputs(5451) <= 1'b0;
    layer0_outputs(5452) <= not a or b;
    layer0_outputs(5453) <= a xor b;
    layer0_outputs(5454) <= a xor b;
    layer0_outputs(5455) <= not (a xor b);
    layer0_outputs(5456) <= a and not b;
    layer0_outputs(5457) <= not (a and b);
    layer0_outputs(5458) <= not a or b;
    layer0_outputs(5459) <= a and b;
    layer0_outputs(5460) <= 1'b1;
    layer0_outputs(5461) <= not a or b;
    layer0_outputs(5462) <= 1'b1;
    layer0_outputs(5463) <= b and not a;
    layer0_outputs(5464) <= a;
    layer0_outputs(5465) <= a xor b;
    layer0_outputs(5466) <= 1'b1;
    layer0_outputs(5467) <= 1'b1;
    layer0_outputs(5468) <= a or b;
    layer0_outputs(5469) <= 1'b0;
    layer0_outputs(5470) <= a or b;
    layer0_outputs(5471) <= not a;
    layer0_outputs(5472) <= a and not b;
    layer0_outputs(5473) <= a and b;
    layer0_outputs(5474) <= a or b;
    layer0_outputs(5475) <= not (a and b);
    layer0_outputs(5476) <= b and not a;
    layer0_outputs(5477) <= a or b;
    layer0_outputs(5478) <= not a;
    layer0_outputs(5479) <= 1'b0;
    layer0_outputs(5480) <= not (a or b);
    layer0_outputs(5481) <= 1'b0;
    layer0_outputs(5482) <= b and not a;
    layer0_outputs(5483) <= not a or b;
    layer0_outputs(5484) <= b;
    layer0_outputs(5485) <= 1'b1;
    layer0_outputs(5486) <= b and not a;
    layer0_outputs(5487) <= b;
    layer0_outputs(5488) <= 1'b1;
    layer0_outputs(5489) <= not (a and b);
    layer0_outputs(5490) <= b and not a;
    layer0_outputs(5491) <= a and not b;
    layer0_outputs(5492) <= a xor b;
    layer0_outputs(5493) <= b;
    layer0_outputs(5494) <= a xor b;
    layer0_outputs(5495) <= a and b;
    layer0_outputs(5496) <= not (a xor b);
    layer0_outputs(5497) <= not a or b;
    layer0_outputs(5498) <= not b;
    layer0_outputs(5499) <= 1'b1;
    layer0_outputs(5500) <= not (a or b);
    layer0_outputs(5501) <= a xor b;
    layer0_outputs(5502) <= b and not a;
    layer0_outputs(5503) <= not (a or b);
    layer0_outputs(5504) <= not (a or b);
    layer0_outputs(5505) <= a and not b;
    layer0_outputs(5506) <= a or b;
    layer0_outputs(5507) <= a and b;
    layer0_outputs(5508) <= 1'b0;
    layer0_outputs(5509) <= b and not a;
    layer0_outputs(5510) <= not a or b;
    layer0_outputs(5511) <= 1'b1;
    layer0_outputs(5512) <= not a or b;
    layer0_outputs(5513) <= not b;
    layer0_outputs(5514) <= not b or a;
    layer0_outputs(5515) <= a or b;
    layer0_outputs(5516) <= a;
    layer0_outputs(5517) <= not a or b;
    layer0_outputs(5518) <= a xor b;
    layer0_outputs(5519) <= b and not a;
    layer0_outputs(5520) <= 1'b1;
    layer0_outputs(5521) <= not (a or b);
    layer0_outputs(5522) <= a or b;
    layer0_outputs(5523) <= not (a xor b);
    layer0_outputs(5524) <= a and not b;
    layer0_outputs(5525) <= not b;
    layer0_outputs(5526) <= not b or a;
    layer0_outputs(5527) <= a and not b;
    layer0_outputs(5528) <= not a;
    layer0_outputs(5529) <= not b or a;
    layer0_outputs(5530) <= 1'b0;
    layer0_outputs(5531) <= not a or b;
    layer0_outputs(5532) <= b;
    layer0_outputs(5533) <= not a;
    layer0_outputs(5534) <= 1'b1;
    layer0_outputs(5535) <= a or b;
    layer0_outputs(5536) <= not b;
    layer0_outputs(5537) <= not a;
    layer0_outputs(5538) <= not b;
    layer0_outputs(5539) <= a or b;
    layer0_outputs(5540) <= a xor b;
    layer0_outputs(5541) <= not b;
    layer0_outputs(5542) <= a or b;
    layer0_outputs(5543) <= a or b;
    layer0_outputs(5544) <= not (a and b);
    layer0_outputs(5545) <= 1'b0;
    layer0_outputs(5546) <= 1'b1;
    layer0_outputs(5547) <= not (a or b);
    layer0_outputs(5548) <= a and not b;
    layer0_outputs(5549) <= not b;
    layer0_outputs(5550) <= 1'b0;
    layer0_outputs(5551) <= a and not b;
    layer0_outputs(5552) <= not a or b;
    layer0_outputs(5553) <= not (a and b);
    layer0_outputs(5554) <= a xor b;
    layer0_outputs(5555) <= 1'b1;
    layer0_outputs(5556) <= b;
    layer0_outputs(5557) <= b;
    layer0_outputs(5558) <= a;
    layer0_outputs(5559) <= not b or a;
    layer0_outputs(5560) <= a or b;
    layer0_outputs(5561) <= 1'b0;
    layer0_outputs(5562) <= a and not b;
    layer0_outputs(5563) <= not (a xor b);
    layer0_outputs(5564) <= a;
    layer0_outputs(5565) <= not a;
    layer0_outputs(5566) <= 1'b1;
    layer0_outputs(5567) <= a and not b;
    layer0_outputs(5568) <= not b;
    layer0_outputs(5569) <= not b;
    layer0_outputs(5570) <= 1'b1;
    layer0_outputs(5571) <= a xor b;
    layer0_outputs(5572) <= not (a or b);
    layer0_outputs(5573) <= not b or a;
    layer0_outputs(5574) <= a or b;
    layer0_outputs(5575) <= b;
    layer0_outputs(5576) <= a;
    layer0_outputs(5577) <= not (a or b);
    layer0_outputs(5578) <= a xor b;
    layer0_outputs(5579) <= b;
    layer0_outputs(5580) <= not (a xor b);
    layer0_outputs(5581) <= 1'b0;
    layer0_outputs(5582) <= not (a or b);
    layer0_outputs(5583) <= a and b;
    layer0_outputs(5584) <= 1'b1;
    layer0_outputs(5585) <= not b or a;
    layer0_outputs(5586) <= a;
    layer0_outputs(5587) <= not a;
    layer0_outputs(5588) <= not b;
    layer0_outputs(5589) <= not (a and b);
    layer0_outputs(5590) <= not (a xor b);
    layer0_outputs(5591) <= not (a or b);
    layer0_outputs(5592) <= not a or b;
    layer0_outputs(5593) <= a xor b;
    layer0_outputs(5594) <= not b or a;
    layer0_outputs(5595) <= not (a or b);
    layer0_outputs(5596) <= not (a or b);
    layer0_outputs(5597) <= a and b;
    layer0_outputs(5598) <= a;
    layer0_outputs(5599) <= not (a or b);
    layer0_outputs(5600) <= 1'b0;
    layer0_outputs(5601) <= a and not b;
    layer0_outputs(5602) <= not (a xor b);
    layer0_outputs(5603) <= a and b;
    layer0_outputs(5604) <= not (a or b);
    layer0_outputs(5605) <= b and not a;
    layer0_outputs(5606) <= not b;
    layer0_outputs(5607) <= not (a and b);
    layer0_outputs(5608) <= a xor b;
    layer0_outputs(5609) <= not (a and b);
    layer0_outputs(5610) <= a;
    layer0_outputs(5611) <= 1'b0;
    layer0_outputs(5612) <= 1'b0;
    layer0_outputs(5613) <= b;
    layer0_outputs(5614) <= not (a xor b);
    layer0_outputs(5615) <= a and b;
    layer0_outputs(5616) <= a or b;
    layer0_outputs(5617) <= not a or b;
    layer0_outputs(5618) <= not a or b;
    layer0_outputs(5619) <= a or b;
    layer0_outputs(5620) <= not (a and b);
    layer0_outputs(5621) <= not a;
    layer0_outputs(5622) <= a and b;
    layer0_outputs(5623) <= b and not a;
    layer0_outputs(5624) <= not b;
    layer0_outputs(5625) <= not (a and b);
    layer0_outputs(5626) <= not (a or b);
    layer0_outputs(5627) <= b;
    layer0_outputs(5628) <= a and b;
    layer0_outputs(5629) <= not (a or b);
    layer0_outputs(5630) <= not a;
    layer0_outputs(5631) <= a;
    layer0_outputs(5632) <= a and b;
    layer0_outputs(5633) <= a;
    layer0_outputs(5634) <= not (a or b);
    layer0_outputs(5635) <= 1'b1;
    layer0_outputs(5636) <= not (a or b);
    layer0_outputs(5637) <= 1'b0;
    layer0_outputs(5638) <= not b or a;
    layer0_outputs(5639) <= 1'b0;
    layer0_outputs(5640) <= a and not b;
    layer0_outputs(5641) <= a and not b;
    layer0_outputs(5642) <= not a or b;
    layer0_outputs(5643) <= 1'b0;
    layer0_outputs(5644) <= not a;
    layer0_outputs(5645) <= 1'b0;
    layer0_outputs(5646) <= not a or b;
    layer0_outputs(5647) <= 1'b1;
    layer0_outputs(5648) <= not a or b;
    layer0_outputs(5649) <= a xor b;
    layer0_outputs(5650) <= not (a or b);
    layer0_outputs(5651) <= 1'b1;
    layer0_outputs(5652) <= 1'b0;
    layer0_outputs(5653) <= a or b;
    layer0_outputs(5654) <= not a or b;
    layer0_outputs(5655) <= not a or b;
    layer0_outputs(5656) <= a or b;
    layer0_outputs(5657) <= not b;
    layer0_outputs(5658) <= a xor b;
    layer0_outputs(5659) <= not (a and b);
    layer0_outputs(5660) <= b;
    layer0_outputs(5661) <= 1'b0;
    layer0_outputs(5662) <= a xor b;
    layer0_outputs(5663) <= not a;
    layer0_outputs(5664) <= not b;
    layer0_outputs(5665) <= not (a and b);
    layer0_outputs(5666) <= a;
    layer0_outputs(5667) <= 1'b0;
    layer0_outputs(5668) <= not (a or b);
    layer0_outputs(5669) <= not b or a;
    layer0_outputs(5670) <= not a or b;
    layer0_outputs(5671) <= not b or a;
    layer0_outputs(5672) <= 1'b0;
    layer0_outputs(5673) <= a or b;
    layer0_outputs(5674) <= a and b;
    layer0_outputs(5675) <= 1'b0;
    layer0_outputs(5676) <= a or b;
    layer0_outputs(5677) <= b;
    layer0_outputs(5678) <= 1'b0;
    layer0_outputs(5679) <= b;
    layer0_outputs(5680) <= a and not b;
    layer0_outputs(5681) <= 1'b0;
    layer0_outputs(5682) <= not a;
    layer0_outputs(5683) <= not a or b;
    layer0_outputs(5684) <= a or b;
    layer0_outputs(5685) <= not a;
    layer0_outputs(5686) <= 1'b0;
    layer0_outputs(5687) <= not b;
    layer0_outputs(5688) <= a xor b;
    layer0_outputs(5689) <= a;
    layer0_outputs(5690) <= not a or b;
    layer0_outputs(5691) <= not (a or b);
    layer0_outputs(5692) <= a or b;
    layer0_outputs(5693) <= a and b;
    layer0_outputs(5694) <= a;
    layer0_outputs(5695) <= not (a xor b);
    layer0_outputs(5696) <= not (a or b);
    layer0_outputs(5697) <= not b or a;
    layer0_outputs(5698) <= not (a xor b);
    layer0_outputs(5699) <= not b or a;
    layer0_outputs(5700) <= a and not b;
    layer0_outputs(5701) <= 1'b0;
    layer0_outputs(5702) <= a xor b;
    layer0_outputs(5703) <= not (a xor b);
    layer0_outputs(5704) <= not a or b;
    layer0_outputs(5705) <= 1'b1;
    layer0_outputs(5706) <= 1'b1;
    layer0_outputs(5707) <= not (a and b);
    layer0_outputs(5708) <= a and not b;
    layer0_outputs(5709) <= not (a or b);
    layer0_outputs(5710) <= 1'b1;
    layer0_outputs(5711) <= not (a or b);
    layer0_outputs(5712) <= b;
    layer0_outputs(5713) <= b;
    layer0_outputs(5714) <= a xor b;
    layer0_outputs(5715) <= 1'b0;
    layer0_outputs(5716) <= not a or b;
    layer0_outputs(5717) <= b and not a;
    layer0_outputs(5718) <= b;
    layer0_outputs(5719) <= 1'b1;
    layer0_outputs(5720) <= not a;
    layer0_outputs(5721) <= not a;
    layer0_outputs(5722) <= not a;
    layer0_outputs(5723) <= b;
    layer0_outputs(5724) <= 1'b0;
    layer0_outputs(5725) <= not (a or b);
    layer0_outputs(5726) <= not (a xor b);
    layer0_outputs(5727) <= a;
    layer0_outputs(5728) <= not a or b;
    layer0_outputs(5729) <= not a or b;
    layer0_outputs(5730) <= a;
    layer0_outputs(5731) <= 1'b1;
    layer0_outputs(5732) <= a and not b;
    layer0_outputs(5733) <= a xor b;
    layer0_outputs(5734) <= not (a or b);
    layer0_outputs(5735) <= not a;
    layer0_outputs(5736) <= b;
    layer0_outputs(5737) <= 1'b0;
    layer0_outputs(5738) <= not b or a;
    layer0_outputs(5739) <= b and not a;
    layer0_outputs(5740) <= not b;
    layer0_outputs(5741) <= 1'b0;
    layer0_outputs(5742) <= a;
    layer0_outputs(5743) <= not b or a;
    layer0_outputs(5744) <= not a;
    layer0_outputs(5745) <= not a or b;
    layer0_outputs(5746) <= 1'b1;
    layer0_outputs(5747) <= not b or a;
    layer0_outputs(5748) <= not b;
    layer0_outputs(5749) <= not b;
    layer0_outputs(5750) <= a xor b;
    layer0_outputs(5751) <= not (a or b);
    layer0_outputs(5752) <= not a;
    layer0_outputs(5753) <= not (a xor b);
    layer0_outputs(5754) <= 1'b1;
    layer0_outputs(5755) <= b;
    layer0_outputs(5756) <= not b;
    layer0_outputs(5757) <= a xor b;
    layer0_outputs(5758) <= not b;
    layer0_outputs(5759) <= a or b;
    layer0_outputs(5760) <= 1'b0;
    layer0_outputs(5761) <= b;
    layer0_outputs(5762) <= a and not b;
    layer0_outputs(5763) <= not (a and b);
    layer0_outputs(5764) <= b and not a;
    layer0_outputs(5765) <= a and not b;
    layer0_outputs(5766) <= not a or b;
    layer0_outputs(5767) <= a and b;
    layer0_outputs(5768) <= b;
    layer0_outputs(5769) <= not (a and b);
    layer0_outputs(5770) <= not (a and b);
    layer0_outputs(5771) <= not (a or b);
    layer0_outputs(5772) <= not b or a;
    layer0_outputs(5773) <= a and b;
    layer0_outputs(5774) <= not a;
    layer0_outputs(5775) <= a or b;
    layer0_outputs(5776) <= a or b;
    layer0_outputs(5777) <= not (a and b);
    layer0_outputs(5778) <= b;
    layer0_outputs(5779) <= a and b;
    layer0_outputs(5780) <= not (a and b);
    layer0_outputs(5781) <= not a or b;
    layer0_outputs(5782) <= a;
    layer0_outputs(5783) <= not a or b;
    layer0_outputs(5784) <= not a or b;
    layer0_outputs(5785) <= not a or b;
    layer0_outputs(5786) <= 1'b0;
    layer0_outputs(5787) <= not (a xor b);
    layer0_outputs(5788) <= not (a or b);
    layer0_outputs(5789) <= b;
    layer0_outputs(5790) <= not a;
    layer0_outputs(5791) <= not a;
    layer0_outputs(5792) <= a and not b;
    layer0_outputs(5793) <= a and not b;
    layer0_outputs(5794) <= not b or a;
    layer0_outputs(5795) <= not a or b;
    layer0_outputs(5796) <= a;
    layer0_outputs(5797) <= a xor b;
    layer0_outputs(5798) <= a;
    layer0_outputs(5799) <= not b or a;
    layer0_outputs(5800) <= a xor b;
    layer0_outputs(5801) <= b;
    layer0_outputs(5802) <= 1'b1;
    layer0_outputs(5803) <= not (a or b);
    layer0_outputs(5804) <= 1'b0;
    layer0_outputs(5805) <= 1'b1;
    layer0_outputs(5806) <= not (a xor b);
    layer0_outputs(5807) <= 1'b1;
    layer0_outputs(5808) <= not a or b;
    layer0_outputs(5809) <= not (a and b);
    layer0_outputs(5810) <= a or b;
    layer0_outputs(5811) <= a and b;
    layer0_outputs(5812) <= 1'b1;
    layer0_outputs(5813) <= not a or b;
    layer0_outputs(5814) <= not a or b;
    layer0_outputs(5815) <= not a;
    layer0_outputs(5816) <= b;
    layer0_outputs(5817) <= 1'b0;
    layer0_outputs(5818) <= not (a and b);
    layer0_outputs(5819) <= 1'b1;
    layer0_outputs(5820) <= not (a xor b);
    layer0_outputs(5821) <= not a or b;
    layer0_outputs(5822) <= b;
    layer0_outputs(5823) <= a;
    layer0_outputs(5824) <= not a;
    layer0_outputs(5825) <= a and not b;
    layer0_outputs(5826) <= a or b;
    layer0_outputs(5827) <= a or b;
    layer0_outputs(5828) <= a;
    layer0_outputs(5829) <= a xor b;
    layer0_outputs(5830) <= b;
    layer0_outputs(5831) <= a;
    layer0_outputs(5832) <= 1'b0;
    layer0_outputs(5833) <= 1'b1;
    layer0_outputs(5834) <= not (a xor b);
    layer0_outputs(5835) <= not (a or b);
    layer0_outputs(5836) <= not b;
    layer0_outputs(5837) <= a and b;
    layer0_outputs(5838) <= 1'b1;
    layer0_outputs(5839) <= not (a xor b);
    layer0_outputs(5840) <= not (a and b);
    layer0_outputs(5841) <= not b;
    layer0_outputs(5842) <= a;
    layer0_outputs(5843) <= b and not a;
    layer0_outputs(5844) <= a or b;
    layer0_outputs(5845) <= not a or b;
    layer0_outputs(5846) <= not a or b;
    layer0_outputs(5847) <= not a;
    layer0_outputs(5848) <= b and not a;
    layer0_outputs(5849) <= not (a or b);
    layer0_outputs(5850) <= b;
    layer0_outputs(5851) <= a xor b;
    layer0_outputs(5852) <= 1'b0;
    layer0_outputs(5853) <= not a or b;
    layer0_outputs(5854) <= a xor b;
    layer0_outputs(5855) <= a and b;
    layer0_outputs(5856) <= not b;
    layer0_outputs(5857) <= not (a and b);
    layer0_outputs(5858) <= a xor b;
    layer0_outputs(5859) <= a;
    layer0_outputs(5860) <= b;
    layer0_outputs(5861) <= 1'b1;
    layer0_outputs(5862) <= b;
    layer0_outputs(5863) <= not (a or b);
    layer0_outputs(5864) <= not (a and b);
    layer0_outputs(5865) <= a and not b;
    layer0_outputs(5866) <= a;
    layer0_outputs(5867) <= a and not b;
    layer0_outputs(5868) <= a and b;
    layer0_outputs(5869) <= not (a or b);
    layer0_outputs(5870) <= 1'b0;
    layer0_outputs(5871) <= not b;
    layer0_outputs(5872) <= not (a xor b);
    layer0_outputs(5873) <= not a or b;
    layer0_outputs(5874) <= 1'b0;
    layer0_outputs(5875) <= a;
    layer0_outputs(5876) <= not (a or b);
    layer0_outputs(5877) <= b and not a;
    layer0_outputs(5878) <= a and b;
    layer0_outputs(5879) <= not a;
    layer0_outputs(5880) <= a xor b;
    layer0_outputs(5881) <= 1'b1;
    layer0_outputs(5882) <= a xor b;
    layer0_outputs(5883) <= not b or a;
    layer0_outputs(5884) <= a or b;
    layer0_outputs(5885) <= a or b;
    layer0_outputs(5886) <= not a or b;
    layer0_outputs(5887) <= not a;
    layer0_outputs(5888) <= a;
    layer0_outputs(5889) <= a and not b;
    layer0_outputs(5890) <= not (a and b);
    layer0_outputs(5891) <= not (a and b);
    layer0_outputs(5892) <= a xor b;
    layer0_outputs(5893) <= not (a xor b);
    layer0_outputs(5894) <= a and b;
    layer0_outputs(5895) <= b;
    layer0_outputs(5896) <= a or b;
    layer0_outputs(5897) <= a;
    layer0_outputs(5898) <= b;
    layer0_outputs(5899) <= a or b;
    layer0_outputs(5900) <= a xor b;
    layer0_outputs(5901) <= not b;
    layer0_outputs(5902) <= not (a xor b);
    layer0_outputs(5903) <= not (a and b);
    layer0_outputs(5904) <= not a or b;
    layer0_outputs(5905) <= a;
    layer0_outputs(5906) <= b and not a;
    layer0_outputs(5907) <= not a;
    layer0_outputs(5908) <= not b or a;
    layer0_outputs(5909) <= not (a and b);
    layer0_outputs(5910) <= 1'b0;
    layer0_outputs(5911) <= not (a or b);
    layer0_outputs(5912) <= 1'b0;
    layer0_outputs(5913) <= a and b;
    layer0_outputs(5914) <= not b or a;
    layer0_outputs(5915) <= a xor b;
    layer0_outputs(5916) <= a xor b;
    layer0_outputs(5917) <= a or b;
    layer0_outputs(5918) <= b;
    layer0_outputs(5919) <= a and b;
    layer0_outputs(5920) <= not b;
    layer0_outputs(5921) <= not a;
    layer0_outputs(5922) <= not a;
    layer0_outputs(5923) <= a;
    layer0_outputs(5924) <= b;
    layer0_outputs(5925) <= not (a and b);
    layer0_outputs(5926) <= not b;
    layer0_outputs(5927) <= a;
    layer0_outputs(5928) <= not a;
    layer0_outputs(5929) <= not a;
    layer0_outputs(5930) <= a xor b;
    layer0_outputs(5931) <= a or b;
    layer0_outputs(5932) <= a or b;
    layer0_outputs(5933) <= not a or b;
    layer0_outputs(5934) <= b;
    layer0_outputs(5935) <= b and not a;
    layer0_outputs(5936) <= not (a or b);
    layer0_outputs(5937) <= a or b;
    layer0_outputs(5938) <= 1'b0;
    layer0_outputs(5939) <= b;
    layer0_outputs(5940) <= not b or a;
    layer0_outputs(5941) <= not a or b;
    layer0_outputs(5942) <= not (a xor b);
    layer0_outputs(5943) <= a and not b;
    layer0_outputs(5944) <= a;
    layer0_outputs(5945) <= b;
    layer0_outputs(5946) <= b;
    layer0_outputs(5947) <= a xor b;
    layer0_outputs(5948) <= not (a and b);
    layer0_outputs(5949) <= b and not a;
    layer0_outputs(5950) <= b;
    layer0_outputs(5951) <= b and not a;
    layer0_outputs(5952) <= not a;
    layer0_outputs(5953) <= a and not b;
    layer0_outputs(5954) <= a and b;
    layer0_outputs(5955) <= not (a xor b);
    layer0_outputs(5956) <= a and b;
    layer0_outputs(5957) <= 1'b1;
    layer0_outputs(5958) <= not b;
    layer0_outputs(5959) <= a or b;
    layer0_outputs(5960) <= a and b;
    layer0_outputs(5961) <= not a;
    layer0_outputs(5962) <= not (a or b);
    layer0_outputs(5963) <= a;
    layer0_outputs(5964) <= a and b;
    layer0_outputs(5965) <= 1'b0;
    layer0_outputs(5966) <= not a;
    layer0_outputs(5967) <= not a;
    layer0_outputs(5968) <= a xor b;
    layer0_outputs(5969) <= 1'b0;
    layer0_outputs(5970) <= a and b;
    layer0_outputs(5971) <= a;
    layer0_outputs(5972) <= not a or b;
    layer0_outputs(5973) <= a xor b;
    layer0_outputs(5974) <= not (a and b);
    layer0_outputs(5975) <= not a;
    layer0_outputs(5976) <= not b or a;
    layer0_outputs(5977) <= not b;
    layer0_outputs(5978) <= not a or b;
    layer0_outputs(5979) <= a;
    layer0_outputs(5980) <= not a;
    layer0_outputs(5981) <= a or b;
    layer0_outputs(5982) <= not (a or b);
    layer0_outputs(5983) <= b and not a;
    layer0_outputs(5984) <= not a;
    layer0_outputs(5985) <= not (a or b);
    layer0_outputs(5986) <= b;
    layer0_outputs(5987) <= not b;
    layer0_outputs(5988) <= 1'b0;
    layer0_outputs(5989) <= 1'b1;
    layer0_outputs(5990) <= a;
    layer0_outputs(5991) <= a or b;
    layer0_outputs(5992) <= not a or b;
    layer0_outputs(5993) <= not a;
    layer0_outputs(5994) <= a or b;
    layer0_outputs(5995) <= a and b;
    layer0_outputs(5996) <= not (a and b);
    layer0_outputs(5997) <= not (a or b);
    layer0_outputs(5998) <= not b or a;
    layer0_outputs(5999) <= 1'b1;
    layer0_outputs(6000) <= 1'b0;
    layer0_outputs(6001) <= not b;
    layer0_outputs(6002) <= not a;
    layer0_outputs(6003) <= not a;
    layer0_outputs(6004) <= not a or b;
    layer0_outputs(6005) <= b;
    layer0_outputs(6006) <= not (a or b);
    layer0_outputs(6007) <= not b;
    layer0_outputs(6008) <= not b;
    layer0_outputs(6009) <= not (a and b);
    layer0_outputs(6010) <= a and b;
    layer0_outputs(6011) <= 1'b1;
    layer0_outputs(6012) <= b and not a;
    layer0_outputs(6013) <= b and not a;
    layer0_outputs(6014) <= a;
    layer0_outputs(6015) <= a or b;
    layer0_outputs(6016) <= a or b;
    layer0_outputs(6017) <= b;
    layer0_outputs(6018) <= not b or a;
    layer0_outputs(6019) <= a or b;
    layer0_outputs(6020) <= not (a and b);
    layer0_outputs(6021) <= not a or b;
    layer0_outputs(6022) <= 1'b1;
    layer0_outputs(6023) <= 1'b1;
    layer0_outputs(6024) <= not a;
    layer0_outputs(6025) <= 1'b0;
    layer0_outputs(6026) <= not b;
    layer0_outputs(6027) <= a and not b;
    layer0_outputs(6028) <= 1'b0;
    layer0_outputs(6029) <= not b or a;
    layer0_outputs(6030) <= not a or b;
    layer0_outputs(6031) <= not a or b;
    layer0_outputs(6032) <= not b or a;
    layer0_outputs(6033) <= not (a or b);
    layer0_outputs(6034) <= not b or a;
    layer0_outputs(6035) <= not (a or b);
    layer0_outputs(6036) <= b and not a;
    layer0_outputs(6037) <= not (a or b);
    layer0_outputs(6038) <= not a;
    layer0_outputs(6039) <= not b or a;
    layer0_outputs(6040) <= b;
    layer0_outputs(6041) <= a xor b;
    layer0_outputs(6042) <= b and not a;
    layer0_outputs(6043) <= not b;
    layer0_outputs(6044) <= a and not b;
    layer0_outputs(6045) <= a or b;
    layer0_outputs(6046) <= b and not a;
    layer0_outputs(6047) <= not a or b;
    layer0_outputs(6048) <= not (a or b);
    layer0_outputs(6049) <= 1'b0;
    layer0_outputs(6050) <= not a or b;
    layer0_outputs(6051) <= a or b;
    layer0_outputs(6052) <= not b or a;
    layer0_outputs(6053) <= a and b;
    layer0_outputs(6054) <= not a;
    layer0_outputs(6055) <= not b;
    layer0_outputs(6056) <= a or b;
    layer0_outputs(6057) <= not b;
    layer0_outputs(6058) <= b;
    layer0_outputs(6059) <= a and not b;
    layer0_outputs(6060) <= 1'b1;
    layer0_outputs(6061) <= 1'b0;
    layer0_outputs(6062) <= not a or b;
    layer0_outputs(6063) <= a xor b;
    layer0_outputs(6064) <= not b;
    layer0_outputs(6065) <= not (a or b);
    layer0_outputs(6066) <= not b or a;
    layer0_outputs(6067) <= a and b;
    layer0_outputs(6068) <= a or b;
    layer0_outputs(6069) <= not b;
    layer0_outputs(6070) <= not (a or b);
    layer0_outputs(6071) <= not (a xor b);
    layer0_outputs(6072) <= not a or b;
    layer0_outputs(6073) <= a and not b;
    layer0_outputs(6074) <= not (a or b);
    layer0_outputs(6075) <= a or b;
    layer0_outputs(6076) <= a and not b;
    layer0_outputs(6077) <= b and not a;
    layer0_outputs(6078) <= not (a or b);
    layer0_outputs(6079) <= a and b;
    layer0_outputs(6080) <= 1'b1;
    layer0_outputs(6081) <= a and not b;
    layer0_outputs(6082) <= b and not a;
    layer0_outputs(6083) <= not b;
    layer0_outputs(6084) <= 1'b0;
    layer0_outputs(6085) <= not a;
    layer0_outputs(6086) <= 1'b0;
    layer0_outputs(6087) <= 1'b0;
    layer0_outputs(6088) <= 1'b1;
    layer0_outputs(6089) <= 1'b1;
    layer0_outputs(6090) <= not a;
    layer0_outputs(6091) <= a and not b;
    layer0_outputs(6092) <= not (a xor b);
    layer0_outputs(6093) <= b and not a;
    layer0_outputs(6094) <= not (a and b);
    layer0_outputs(6095) <= 1'b0;
    layer0_outputs(6096) <= not b;
    layer0_outputs(6097) <= not (a or b);
    layer0_outputs(6098) <= 1'b0;
    layer0_outputs(6099) <= a and not b;
    layer0_outputs(6100) <= a or b;
    layer0_outputs(6101) <= a and not b;
    layer0_outputs(6102) <= a or b;
    layer0_outputs(6103) <= b;
    layer0_outputs(6104) <= b and not a;
    layer0_outputs(6105) <= a and b;
    layer0_outputs(6106) <= 1'b1;
    layer0_outputs(6107) <= not (a or b);
    layer0_outputs(6108) <= not (a and b);
    layer0_outputs(6109) <= not a;
    layer0_outputs(6110) <= not (a and b);
    layer0_outputs(6111) <= not a;
    layer0_outputs(6112) <= not (a or b);
    layer0_outputs(6113) <= b;
    layer0_outputs(6114) <= not b;
    layer0_outputs(6115) <= not b or a;
    layer0_outputs(6116) <= a and not b;
    layer0_outputs(6117) <= b and not a;
    layer0_outputs(6118) <= not (a and b);
    layer0_outputs(6119) <= a;
    layer0_outputs(6120) <= a or b;
    layer0_outputs(6121) <= b and not a;
    layer0_outputs(6122) <= not (a and b);
    layer0_outputs(6123) <= not (a xor b);
    layer0_outputs(6124) <= a xor b;
    layer0_outputs(6125) <= 1'b0;
    layer0_outputs(6126) <= 1'b0;
    layer0_outputs(6127) <= a or b;
    layer0_outputs(6128) <= 1'b0;
    layer0_outputs(6129) <= 1'b0;
    layer0_outputs(6130) <= not a or b;
    layer0_outputs(6131) <= a;
    layer0_outputs(6132) <= not b;
    layer0_outputs(6133) <= not (a or b);
    layer0_outputs(6134) <= a or b;
    layer0_outputs(6135) <= not (a xor b);
    layer0_outputs(6136) <= a or b;
    layer0_outputs(6137) <= not (a or b);
    layer0_outputs(6138) <= not (a or b);
    layer0_outputs(6139) <= a or b;
    layer0_outputs(6140) <= not a;
    layer0_outputs(6141) <= not a;
    layer0_outputs(6142) <= not b;
    layer0_outputs(6143) <= 1'b1;
    layer0_outputs(6144) <= not (a or b);
    layer0_outputs(6145) <= not b;
    layer0_outputs(6146) <= not b;
    layer0_outputs(6147) <= a xor b;
    layer0_outputs(6148) <= 1'b1;
    layer0_outputs(6149) <= a;
    layer0_outputs(6150) <= a or b;
    layer0_outputs(6151) <= not b;
    layer0_outputs(6152) <= a or b;
    layer0_outputs(6153) <= b and not a;
    layer0_outputs(6154) <= 1'b0;
    layer0_outputs(6155) <= b;
    layer0_outputs(6156) <= 1'b1;
    layer0_outputs(6157) <= a and not b;
    layer0_outputs(6158) <= not (a or b);
    layer0_outputs(6159) <= not b;
    layer0_outputs(6160) <= a and not b;
    layer0_outputs(6161) <= not a or b;
    layer0_outputs(6162) <= a xor b;
    layer0_outputs(6163) <= 1'b0;
    layer0_outputs(6164) <= not (a and b);
    layer0_outputs(6165) <= a;
    layer0_outputs(6166) <= not (a or b);
    layer0_outputs(6167) <= a and b;
    layer0_outputs(6168) <= a xor b;
    layer0_outputs(6169) <= a xor b;
    layer0_outputs(6170) <= 1'b1;
    layer0_outputs(6171) <= not (a and b);
    layer0_outputs(6172) <= 1'b1;
    layer0_outputs(6173) <= not (a or b);
    layer0_outputs(6174) <= b and not a;
    layer0_outputs(6175) <= b and not a;
    layer0_outputs(6176) <= not b or a;
    layer0_outputs(6177) <= not (a and b);
    layer0_outputs(6178) <= 1'b1;
    layer0_outputs(6179) <= a;
    layer0_outputs(6180) <= not (a or b);
    layer0_outputs(6181) <= not b or a;
    layer0_outputs(6182) <= not (a and b);
    layer0_outputs(6183) <= not b or a;
    layer0_outputs(6184) <= b;
    layer0_outputs(6185) <= not a;
    layer0_outputs(6186) <= not a;
    layer0_outputs(6187) <= b and not a;
    layer0_outputs(6188) <= not a or b;
    layer0_outputs(6189) <= not (a xor b);
    layer0_outputs(6190) <= a and b;
    layer0_outputs(6191) <= not a or b;
    layer0_outputs(6192) <= a;
    layer0_outputs(6193) <= not (a or b);
    layer0_outputs(6194) <= not (a and b);
    layer0_outputs(6195) <= a;
    layer0_outputs(6196) <= a and b;
    layer0_outputs(6197) <= not (a and b);
    layer0_outputs(6198) <= a xor b;
    layer0_outputs(6199) <= not (a xor b);
    layer0_outputs(6200) <= not b or a;
    layer0_outputs(6201) <= 1'b1;
    layer0_outputs(6202) <= not b or a;
    layer0_outputs(6203) <= 1'b1;
    layer0_outputs(6204) <= not b;
    layer0_outputs(6205) <= 1'b0;
    layer0_outputs(6206) <= a and b;
    layer0_outputs(6207) <= not b;
    layer0_outputs(6208) <= not b;
    layer0_outputs(6209) <= not b or a;
    layer0_outputs(6210) <= not b;
    layer0_outputs(6211) <= a or b;
    layer0_outputs(6212) <= a and not b;
    layer0_outputs(6213) <= a or b;
    layer0_outputs(6214) <= a;
    layer0_outputs(6215) <= not a;
    layer0_outputs(6216) <= not a;
    layer0_outputs(6217) <= a;
    layer0_outputs(6218) <= b and not a;
    layer0_outputs(6219) <= not (a xor b);
    layer0_outputs(6220) <= b;
    layer0_outputs(6221) <= not (a and b);
    layer0_outputs(6222) <= not b or a;
    layer0_outputs(6223) <= not b;
    layer0_outputs(6224) <= not b or a;
    layer0_outputs(6225) <= not a;
    layer0_outputs(6226) <= 1'b1;
    layer0_outputs(6227) <= 1'b1;
    layer0_outputs(6228) <= a and not b;
    layer0_outputs(6229) <= a and b;
    layer0_outputs(6230) <= a;
    layer0_outputs(6231) <= a or b;
    layer0_outputs(6232) <= not b or a;
    layer0_outputs(6233) <= not (a xor b);
    layer0_outputs(6234) <= a and not b;
    layer0_outputs(6235) <= a;
    layer0_outputs(6236) <= not a;
    layer0_outputs(6237) <= not (a xor b);
    layer0_outputs(6238) <= a xor b;
    layer0_outputs(6239) <= 1'b0;
    layer0_outputs(6240) <= b;
    layer0_outputs(6241) <= not b;
    layer0_outputs(6242) <= 1'b0;
    layer0_outputs(6243) <= a and b;
    layer0_outputs(6244) <= a;
    layer0_outputs(6245) <= not (a xor b);
    layer0_outputs(6246) <= b and not a;
    layer0_outputs(6247) <= b and not a;
    layer0_outputs(6248) <= 1'b0;
    layer0_outputs(6249) <= not b;
    layer0_outputs(6250) <= b;
    layer0_outputs(6251) <= a and b;
    layer0_outputs(6252) <= not (a and b);
    layer0_outputs(6253) <= 1'b0;
    layer0_outputs(6254) <= 1'b0;
    layer0_outputs(6255) <= not (a xor b);
    layer0_outputs(6256) <= not b;
    layer0_outputs(6257) <= 1'b1;
    layer0_outputs(6258) <= not b or a;
    layer0_outputs(6259) <= not (a or b);
    layer0_outputs(6260) <= not (a or b);
    layer0_outputs(6261) <= not b or a;
    layer0_outputs(6262) <= not (a or b);
    layer0_outputs(6263) <= a and not b;
    layer0_outputs(6264) <= a and b;
    layer0_outputs(6265) <= not (a and b);
    layer0_outputs(6266) <= a;
    layer0_outputs(6267) <= 1'b1;
    layer0_outputs(6268) <= a and b;
    layer0_outputs(6269) <= not (a or b);
    layer0_outputs(6270) <= a xor b;
    layer0_outputs(6271) <= a and b;
    layer0_outputs(6272) <= a and b;
    layer0_outputs(6273) <= 1'b1;
    layer0_outputs(6274) <= a;
    layer0_outputs(6275) <= b and not a;
    layer0_outputs(6276) <= not b or a;
    layer0_outputs(6277) <= b;
    layer0_outputs(6278) <= 1'b1;
    layer0_outputs(6279) <= a;
    layer0_outputs(6280) <= not b;
    layer0_outputs(6281) <= not a or b;
    layer0_outputs(6282) <= not (a or b);
    layer0_outputs(6283) <= not a or b;
    layer0_outputs(6284) <= a;
    layer0_outputs(6285) <= 1'b0;
    layer0_outputs(6286) <= not (a xor b);
    layer0_outputs(6287) <= not b;
    layer0_outputs(6288) <= b and not a;
    layer0_outputs(6289) <= 1'b0;
    layer0_outputs(6290) <= not b or a;
    layer0_outputs(6291) <= not a or b;
    layer0_outputs(6292) <= 1'b1;
    layer0_outputs(6293) <= b;
    layer0_outputs(6294) <= a and b;
    layer0_outputs(6295) <= not (a xor b);
    layer0_outputs(6296) <= 1'b0;
    layer0_outputs(6297) <= a or b;
    layer0_outputs(6298) <= 1'b1;
    layer0_outputs(6299) <= not b;
    layer0_outputs(6300) <= not (a xor b);
    layer0_outputs(6301) <= not (a xor b);
    layer0_outputs(6302) <= b and not a;
    layer0_outputs(6303) <= not b;
    layer0_outputs(6304) <= 1'b1;
    layer0_outputs(6305) <= b and not a;
    layer0_outputs(6306) <= a xor b;
    layer0_outputs(6307) <= not a or b;
    layer0_outputs(6308) <= not (a and b);
    layer0_outputs(6309) <= not a or b;
    layer0_outputs(6310) <= b;
    layer0_outputs(6311) <= not (a or b);
    layer0_outputs(6312) <= not b or a;
    layer0_outputs(6313) <= not b or a;
    layer0_outputs(6314) <= not b or a;
    layer0_outputs(6315) <= not b or a;
    layer0_outputs(6316) <= not b or a;
    layer0_outputs(6317) <= a or b;
    layer0_outputs(6318) <= not (a or b);
    layer0_outputs(6319) <= b;
    layer0_outputs(6320) <= 1'b0;
    layer0_outputs(6321) <= 1'b1;
    layer0_outputs(6322) <= a and not b;
    layer0_outputs(6323) <= a and not b;
    layer0_outputs(6324) <= a xor b;
    layer0_outputs(6325) <= a or b;
    layer0_outputs(6326) <= not (a xor b);
    layer0_outputs(6327) <= a and b;
    layer0_outputs(6328) <= not a or b;
    layer0_outputs(6329) <= a xor b;
    layer0_outputs(6330) <= not (a and b);
    layer0_outputs(6331) <= b;
    layer0_outputs(6332) <= 1'b1;
    layer0_outputs(6333) <= b and not a;
    layer0_outputs(6334) <= b;
    layer0_outputs(6335) <= b and not a;
    layer0_outputs(6336) <= not a;
    layer0_outputs(6337) <= 1'b1;
    layer0_outputs(6338) <= a;
    layer0_outputs(6339) <= not b;
    layer0_outputs(6340) <= b and not a;
    layer0_outputs(6341) <= not a;
    layer0_outputs(6342) <= 1'b0;
    layer0_outputs(6343) <= a;
    layer0_outputs(6344) <= a;
    layer0_outputs(6345) <= not a;
    layer0_outputs(6346) <= not (a xor b);
    layer0_outputs(6347) <= not b;
    layer0_outputs(6348) <= not a;
    layer0_outputs(6349) <= a and not b;
    layer0_outputs(6350) <= not b or a;
    layer0_outputs(6351) <= not (a and b);
    layer0_outputs(6352) <= a and not b;
    layer0_outputs(6353) <= 1'b0;
    layer0_outputs(6354) <= a and not b;
    layer0_outputs(6355) <= 1'b1;
    layer0_outputs(6356) <= 1'b0;
    layer0_outputs(6357) <= not a or b;
    layer0_outputs(6358) <= not a or b;
    layer0_outputs(6359) <= not b or a;
    layer0_outputs(6360) <= a or b;
    layer0_outputs(6361) <= not a or b;
    layer0_outputs(6362) <= not a;
    layer0_outputs(6363) <= 1'b1;
    layer0_outputs(6364) <= a or b;
    layer0_outputs(6365) <= 1'b0;
    layer0_outputs(6366) <= a and not b;
    layer0_outputs(6367) <= not a;
    layer0_outputs(6368) <= not (a or b);
    layer0_outputs(6369) <= b and not a;
    layer0_outputs(6370) <= 1'b0;
    layer0_outputs(6371) <= a;
    layer0_outputs(6372) <= not b;
    layer0_outputs(6373) <= 1'b0;
    layer0_outputs(6374) <= a and b;
    layer0_outputs(6375) <= not (a xor b);
    layer0_outputs(6376) <= not a or b;
    layer0_outputs(6377) <= 1'b1;
    layer0_outputs(6378) <= 1'b1;
    layer0_outputs(6379) <= not a;
    layer0_outputs(6380) <= 1'b1;
    layer0_outputs(6381) <= 1'b1;
    layer0_outputs(6382) <= a and not b;
    layer0_outputs(6383) <= a;
    layer0_outputs(6384) <= 1'b0;
    layer0_outputs(6385) <= b and not a;
    layer0_outputs(6386) <= 1'b0;
    layer0_outputs(6387) <= b and not a;
    layer0_outputs(6388) <= a and not b;
    layer0_outputs(6389) <= not b;
    layer0_outputs(6390) <= a;
    layer0_outputs(6391) <= b and not a;
    layer0_outputs(6392) <= a or b;
    layer0_outputs(6393) <= b;
    layer0_outputs(6394) <= a or b;
    layer0_outputs(6395) <= not a;
    layer0_outputs(6396) <= not b;
    layer0_outputs(6397) <= b;
    layer0_outputs(6398) <= b;
    layer0_outputs(6399) <= 1'b1;
    layer0_outputs(6400) <= a and not b;
    layer0_outputs(6401) <= 1'b1;
    layer0_outputs(6402) <= not a or b;
    layer0_outputs(6403) <= a;
    layer0_outputs(6404) <= not (a or b);
    layer0_outputs(6405) <= not (a and b);
    layer0_outputs(6406) <= a or b;
    layer0_outputs(6407) <= a or b;
    layer0_outputs(6408) <= a and b;
    layer0_outputs(6409) <= a and not b;
    layer0_outputs(6410) <= not b or a;
    layer0_outputs(6411) <= a and not b;
    layer0_outputs(6412) <= 1'b1;
    layer0_outputs(6413) <= not a or b;
    layer0_outputs(6414) <= 1'b1;
    layer0_outputs(6415) <= not (a or b);
    layer0_outputs(6416) <= not (a and b);
    layer0_outputs(6417) <= a and b;
    layer0_outputs(6418) <= a or b;
    layer0_outputs(6419) <= 1'b0;
    layer0_outputs(6420) <= b;
    layer0_outputs(6421) <= not a or b;
    layer0_outputs(6422) <= a and b;
    layer0_outputs(6423) <= a and b;
    layer0_outputs(6424) <= b and not a;
    layer0_outputs(6425) <= not b or a;
    layer0_outputs(6426) <= not (a xor b);
    layer0_outputs(6427) <= a or b;
    layer0_outputs(6428) <= a xor b;
    layer0_outputs(6429) <= not b;
    layer0_outputs(6430) <= a and not b;
    layer0_outputs(6431) <= not b or a;
    layer0_outputs(6432) <= a and b;
    layer0_outputs(6433) <= not b or a;
    layer0_outputs(6434) <= not (a and b);
    layer0_outputs(6435) <= b and not a;
    layer0_outputs(6436) <= not b or a;
    layer0_outputs(6437) <= not b;
    layer0_outputs(6438) <= a xor b;
    layer0_outputs(6439) <= b;
    layer0_outputs(6440) <= a or b;
    layer0_outputs(6441) <= not (a and b);
    layer0_outputs(6442) <= 1'b0;
    layer0_outputs(6443) <= not (a and b);
    layer0_outputs(6444) <= not a or b;
    layer0_outputs(6445) <= b;
    layer0_outputs(6446) <= not (a or b);
    layer0_outputs(6447) <= a;
    layer0_outputs(6448) <= 1'b1;
    layer0_outputs(6449) <= b and not a;
    layer0_outputs(6450) <= a and b;
    layer0_outputs(6451) <= b and not a;
    layer0_outputs(6452) <= a and not b;
    layer0_outputs(6453) <= a and not b;
    layer0_outputs(6454) <= not a or b;
    layer0_outputs(6455) <= not a or b;
    layer0_outputs(6456) <= not b;
    layer0_outputs(6457) <= not a or b;
    layer0_outputs(6458) <= not a;
    layer0_outputs(6459) <= b;
    layer0_outputs(6460) <= not (a or b);
    layer0_outputs(6461) <= b and not a;
    layer0_outputs(6462) <= not (a xor b);
    layer0_outputs(6463) <= a and b;
    layer0_outputs(6464) <= b;
    layer0_outputs(6465) <= a;
    layer0_outputs(6466) <= not b or a;
    layer0_outputs(6467) <= not a or b;
    layer0_outputs(6468) <= a xor b;
    layer0_outputs(6469) <= a xor b;
    layer0_outputs(6470) <= a and not b;
    layer0_outputs(6471) <= 1'b0;
    layer0_outputs(6472) <= a or b;
    layer0_outputs(6473) <= not (a and b);
    layer0_outputs(6474) <= not (a and b);
    layer0_outputs(6475) <= 1'b0;
    layer0_outputs(6476) <= a and not b;
    layer0_outputs(6477) <= a xor b;
    layer0_outputs(6478) <= a;
    layer0_outputs(6479) <= a and not b;
    layer0_outputs(6480) <= a and not b;
    layer0_outputs(6481) <= a and b;
    layer0_outputs(6482) <= not b;
    layer0_outputs(6483) <= b;
    layer0_outputs(6484) <= not a;
    layer0_outputs(6485) <= a or b;
    layer0_outputs(6486) <= a and not b;
    layer0_outputs(6487) <= b;
    layer0_outputs(6488) <= not a;
    layer0_outputs(6489) <= a xor b;
    layer0_outputs(6490) <= a xor b;
    layer0_outputs(6491) <= a xor b;
    layer0_outputs(6492) <= not b;
    layer0_outputs(6493) <= not b;
    layer0_outputs(6494) <= 1'b0;
    layer0_outputs(6495) <= not (a or b);
    layer0_outputs(6496) <= not (a and b);
    layer0_outputs(6497) <= not a;
    layer0_outputs(6498) <= a xor b;
    layer0_outputs(6499) <= not b or a;
    layer0_outputs(6500) <= b;
    layer0_outputs(6501) <= not b or a;
    layer0_outputs(6502) <= a xor b;
    layer0_outputs(6503) <= a and not b;
    layer0_outputs(6504) <= b and not a;
    layer0_outputs(6505) <= a or b;
    layer0_outputs(6506) <= b;
    layer0_outputs(6507) <= a xor b;
    layer0_outputs(6508) <= 1'b0;
    layer0_outputs(6509) <= 1'b0;
    layer0_outputs(6510) <= 1'b0;
    layer0_outputs(6511) <= not b;
    layer0_outputs(6512) <= not b;
    layer0_outputs(6513) <= a;
    layer0_outputs(6514) <= a;
    layer0_outputs(6515) <= not b;
    layer0_outputs(6516) <= 1'b1;
    layer0_outputs(6517) <= 1'b1;
    layer0_outputs(6518) <= not (a xor b);
    layer0_outputs(6519) <= not b;
    layer0_outputs(6520) <= not (a or b);
    layer0_outputs(6521) <= not (a xor b);
    layer0_outputs(6522) <= a xor b;
    layer0_outputs(6523) <= b;
    layer0_outputs(6524) <= a and b;
    layer0_outputs(6525) <= not a;
    layer0_outputs(6526) <= 1'b1;
    layer0_outputs(6527) <= not (a and b);
    layer0_outputs(6528) <= 1'b0;
    layer0_outputs(6529) <= 1'b0;
    layer0_outputs(6530) <= a and not b;
    layer0_outputs(6531) <= not a or b;
    layer0_outputs(6532) <= not (a and b);
    layer0_outputs(6533) <= a and b;
    layer0_outputs(6534) <= not b or a;
    layer0_outputs(6535) <= a or b;
    layer0_outputs(6536) <= not a or b;
    layer0_outputs(6537) <= a xor b;
    layer0_outputs(6538) <= not a;
    layer0_outputs(6539) <= b;
    layer0_outputs(6540) <= 1'b0;
    layer0_outputs(6541) <= not a or b;
    layer0_outputs(6542) <= a xor b;
    layer0_outputs(6543) <= a;
    layer0_outputs(6544) <= b;
    layer0_outputs(6545) <= not (a and b);
    layer0_outputs(6546) <= a and not b;
    layer0_outputs(6547) <= not b;
    layer0_outputs(6548) <= not b or a;
    layer0_outputs(6549) <= not (a xor b);
    layer0_outputs(6550) <= b and not a;
    layer0_outputs(6551) <= a;
    layer0_outputs(6552) <= a xor b;
    layer0_outputs(6553) <= b and not a;
    layer0_outputs(6554) <= not b;
    layer0_outputs(6555) <= a or b;
    layer0_outputs(6556) <= not (a and b);
    layer0_outputs(6557) <= not b or a;
    layer0_outputs(6558) <= not (a and b);
    layer0_outputs(6559) <= a;
    layer0_outputs(6560) <= a and not b;
    layer0_outputs(6561) <= not b or a;
    layer0_outputs(6562) <= not a;
    layer0_outputs(6563) <= a;
    layer0_outputs(6564) <= a or b;
    layer0_outputs(6565) <= not a;
    layer0_outputs(6566) <= a and b;
    layer0_outputs(6567) <= not b or a;
    layer0_outputs(6568) <= not b;
    layer0_outputs(6569) <= 1'b1;
    layer0_outputs(6570) <= not b or a;
    layer0_outputs(6571) <= not b;
    layer0_outputs(6572) <= b;
    layer0_outputs(6573) <= a and not b;
    layer0_outputs(6574) <= not b;
    layer0_outputs(6575) <= 1'b0;
    layer0_outputs(6576) <= not (a and b);
    layer0_outputs(6577) <= not (a and b);
    layer0_outputs(6578) <= a or b;
    layer0_outputs(6579) <= not b or a;
    layer0_outputs(6580) <= b;
    layer0_outputs(6581) <= a or b;
    layer0_outputs(6582) <= not b;
    layer0_outputs(6583) <= 1'b1;
    layer0_outputs(6584) <= not (a xor b);
    layer0_outputs(6585) <= not (a or b);
    layer0_outputs(6586) <= b and not a;
    layer0_outputs(6587) <= 1'b1;
    layer0_outputs(6588) <= not a or b;
    layer0_outputs(6589) <= not a;
    layer0_outputs(6590) <= not (a xor b);
    layer0_outputs(6591) <= not b;
    layer0_outputs(6592) <= not a;
    layer0_outputs(6593) <= not b or a;
    layer0_outputs(6594) <= a and b;
    layer0_outputs(6595) <= a xor b;
    layer0_outputs(6596) <= b;
    layer0_outputs(6597) <= b and not a;
    layer0_outputs(6598) <= 1'b0;
    layer0_outputs(6599) <= a;
    layer0_outputs(6600) <= not (a or b);
    layer0_outputs(6601) <= not (a and b);
    layer0_outputs(6602) <= not a;
    layer0_outputs(6603) <= not a;
    layer0_outputs(6604) <= not b or a;
    layer0_outputs(6605) <= a and not b;
    layer0_outputs(6606) <= not a;
    layer0_outputs(6607) <= a or b;
    layer0_outputs(6608) <= not b or a;
    layer0_outputs(6609) <= a;
    layer0_outputs(6610) <= not (a or b);
    layer0_outputs(6611) <= not (a and b);
    layer0_outputs(6612) <= not (a or b);
    layer0_outputs(6613) <= a and b;
    layer0_outputs(6614) <= 1'b0;
    layer0_outputs(6615) <= a;
    layer0_outputs(6616) <= not a;
    layer0_outputs(6617) <= a;
    layer0_outputs(6618) <= not a;
    layer0_outputs(6619) <= a and b;
    layer0_outputs(6620) <= b;
    layer0_outputs(6621) <= not (a xor b);
    layer0_outputs(6622) <= a and b;
    layer0_outputs(6623) <= not a;
    layer0_outputs(6624) <= a or b;
    layer0_outputs(6625) <= b;
    layer0_outputs(6626) <= b and not a;
    layer0_outputs(6627) <= not (a and b);
    layer0_outputs(6628) <= not (a or b);
    layer0_outputs(6629) <= 1'b1;
    layer0_outputs(6630) <= not (a and b);
    layer0_outputs(6631) <= a;
    layer0_outputs(6632) <= not b or a;
    layer0_outputs(6633) <= a and not b;
    layer0_outputs(6634) <= not (a or b);
    layer0_outputs(6635) <= not b or a;
    layer0_outputs(6636) <= not (a or b);
    layer0_outputs(6637) <= a and b;
    layer0_outputs(6638) <= not a or b;
    layer0_outputs(6639) <= a;
    layer0_outputs(6640) <= 1'b1;
    layer0_outputs(6641) <= b and not a;
    layer0_outputs(6642) <= b and not a;
    layer0_outputs(6643) <= not (a or b);
    layer0_outputs(6644) <= a or b;
    layer0_outputs(6645) <= not b or a;
    layer0_outputs(6646) <= not a or b;
    layer0_outputs(6647) <= 1'b1;
    layer0_outputs(6648) <= a and not b;
    layer0_outputs(6649) <= not b or a;
    layer0_outputs(6650) <= not a or b;
    layer0_outputs(6651) <= 1'b1;
    layer0_outputs(6652) <= not a;
    layer0_outputs(6653) <= a and b;
    layer0_outputs(6654) <= a or b;
    layer0_outputs(6655) <= 1'b1;
    layer0_outputs(6656) <= not a;
    layer0_outputs(6657) <= 1'b0;
    layer0_outputs(6658) <= not b or a;
    layer0_outputs(6659) <= a or b;
    layer0_outputs(6660) <= not (a xor b);
    layer0_outputs(6661) <= not (a or b);
    layer0_outputs(6662) <= b and not a;
    layer0_outputs(6663) <= a and b;
    layer0_outputs(6664) <= not b;
    layer0_outputs(6665) <= not (a and b);
    layer0_outputs(6666) <= 1'b1;
    layer0_outputs(6667) <= a and not b;
    layer0_outputs(6668) <= a or b;
    layer0_outputs(6669) <= 1'b0;
    layer0_outputs(6670) <= a;
    layer0_outputs(6671) <= b;
    layer0_outputs(6672) <= a;
    layer0_outputs(6673) <= a and b;
    layer0_outputs(6674) <= b;
    layer0_outputs(6675) <= a and not b;
    layer0_outputs(6676) <= not b or a;
    layer0_outputs(6677) <= a;
    layer0_outputs(6678) <= a or b;
    layer0_outputs(6679) <= not b or a;
    layer0_outputs(6680) <= not (a or b);
    layer0_outputs(6681) <= not (a xor b);
    layer0_outputs(6682) <= not a;
    layer0_outputs(6683) <= not a;
    layer0_outputs(6684) <= not a or b;
    layer0_outputs(6685) <= not b;
    layer0_outputs(6686) <= not (a and b);
    layer0_outputs(6687) <= not b or a;
    layer0_outputs(6688) <= not b;
    layer0_outputs(6689) <= b and not a;
    layer0_outputs(6690) <= not a;
    layer0_outputs(6691) <= a and b;
    layer0_outputs(6692) <= not b or a;
    layer0_outputs(6693) <= b and not a;
    layer0_outputs(6694) <= not a;
    layer0_outputs(6695) <= not a or b;
    layer0_outputs(6696) <= b;
    layer0_outputs(6697) <= b;
    layer0_outputs(6698) <= not b;
    layer0_outputs(6699) <= not b or a;
    layer0_outputs(6700) <= not b or a;
    layer0_outputs(6701) <= a and not b;
    layer0_outputs(6702) <= not b;
    layer0_outputs(6703) <= a and b;
    layer0_outputs(6704) <= not a or b;
    layer0_outputs(6705) <= 1'b1;
    layer0_outputs(6706) <= 1'b0;
    layer0_outputs(6707) <= a;
    layer0_outputs(6708) <= a;
    layer0_outputs(6709) <= b;
    layer0_outputs(6710) <= a and b;
    layer0_outputs(6711) <= 1'b0;
    layer0_outputs(6712) <= 1'b0;
    layer0_outputs(6713) <= not (a xor b);
    layer0_outputs(6714) <= not (a xor b);
    layer0_outputs(6715) <= 1'b1;
    layer0_outputs(6716) <= a and not b;
    layer0_outputs(6717) <= not (a and b);
    layer0_outputs(6718) <= 1'b0;
    layer0_outputs(6719) <= not (a or b);
    layer0_outputs(6720) <= b and not a;
    layer0_outputs(6721) <= not (a xor b);
    layer0_outputs(6722) <= not (a and b);
    layer0_outputs(6723) <= a or b;
    layer0_outputs(6724) <= 1'b1;
    layer0_outputs(6725) <= not b;
    layer0_outputs(6726) <= a and b;
    layer0_outputs(6727) <= 1'b1;
    layer0_outputs(6728) <= a;
    layer0_outputs(6729) <= a and not b;
    layer0_outputs(6730) <= not (a xor b);
    layer0_outputs(6731) <= not a or b;
    layer0_outputs(6732) <= a;
    layer0_outputs(6733) <= not (a or b);
    layer0_outputs(6734) <= not (a or b);
    layer0_outputs(6735) <= a;
    layer0_outputs(6736) <= not (a xor b);
    layer0_outputs(6737) <= not (a or b);
    layer0_outputs(6738) <= 1'b1;
    layer0_outputs(6739) <= not b;
    layer0_outputs(6740) <= not b;
    layer0_outputs(6741) <= not (a and b);
    layer0_outputs(6742) <= 1'b1;
    layer0_outputs(6743) <= not a;
    layer0_outputs(6744) <= not b;
    layer0_outputs(6745) <= a;
    layer0_outputs(6746) <= b;
    layer0_outputs(6747) <= 1'b1;
    layer0_outputs(6748) <= a and not b;
    layer0_outputs(6749) <= a;
    layer0_outputs(6750) <= a and not b;
    layer0_outputs(6751) <= not (a xor b);
    layer0_outputs(6752) <= not b;
    layer0_outputs(6753) <= not (a xor b);
    layer0_outputs(6754) <= a;
    layer0_outputs(6755) <= b and not a;
    layer0_outputs(6756) <= a and b;
    layer0_outputs(6757) <= 1'b0;
    layer0_outputs(6758) <= b and not a;
    layer0_outputs(6759) <= a xor b;
    layer0_outputs(6760) <= a;
    layer0_outputs(6761) <= not b or a;
    layer0_outputs(6762) <= not (a xor b);
    layer0_outputs(6763) <= not a or b;
    layer0_outputs(6764) <= a;
    layer0_outputs(6765) <= not (a and b);
    layer0_outputs(6766) <= not (a xor b);
    layer0_outputs(6767) <= a;
    layer0_outputs(6768) <= a or b;
    layer0_outputs(6769) <= 1'b0;
    layer0_outputs(6770) <= a xor b;
    layer0_outputs(6771) <= a and b;
    layer0_outputs(6772) <= b;
    layer0_outputs(6773) <= not b or a;
    layer0_outputs(6774) <= not a;
    layer0_outputs(6775) <= not (a or b);
    layer0_outputs(6776) <= a or b;
    layer0_outputs(6777) <= not a;
    layer0_outputs(6778) <= not b or a;
    layer0_outputs(6779) <= 1'b1;
    layer0_outputs(6780) <= not (a and b);
    layer0_outputs(6781) <= a xor b;
    layer0_outputs(6782) <= not b;
    layer0_outputs(6783) <= not (a or b);
    layer0_outputs(6784) <= a;
    layer0_outputs(6785) <= 1'b1;
    layer0_outputs(6786) <= 1'b0;
    layer0_outputs(6787) <= a and not b;
    layer0_outputs(6788) <= a and b;
    layer0_outputs(6789) <= not (a xor b);
    layer0_outputs(6790) <= b and not a;
    layer0_outputs(6791) <= not (a or b);
    layer0_outputs(6792) <= b;
    layer0_outputs(6793) <= not (a and b);
    layer0_outputs(6794) <= b;
    layer0_outputs(6795) <= not b or a;
    layer0_outputs(6796) <= a and b;
    layer0_outputs(6797) <= not b or a;
    layer0_outputs(6798) <= a and b;
    layer0_outputs(6799) <= a xor b;
    layer0_outputs(6800) <= a xor b;
    layer0_outputs(6801) <= not (a xor b);
    layer0_outputs(6802) <= 1'b1;
    layer0_outputs(6803) <= not a or b;
    layer0_outputs(6804) <= not a or b;
    layer0_outputs(6805) <= 1'b1;
    layer0_outputs(6806) <= b;
    layer0_outputs(6807) <= a;
    layer0_outputs(6808) <= not (a or b);
    layer0_outputs(6809) <= not (a or b);
    layer0_outputs(6810) <= a or b;
    layer0_outputs(6811) <= a;
    layer0_outputs(6812) <= not a or b;
    layer0_outputs(6813) <= a and not b;
    layer0_outputs(6814) <= a or b;
    layer0_outputs(6815) <= a;
    layer0_outputs(6816) <= b and not a;
    layer0_outputs(6817) <= b and not a;
    layer0_outputs(6818) <= not b or a;
    layer0_outputs(6819) <= not a or b;
    layer0_outputs(6820) <= a xor b;
    layer0_outputs(6821) <= 1'b0;
    layer0_outputs(6822) <= 1'b0;
    layer0_outputs(6823) <= not b;
    layer0_outputs(6824) <= not b or a;
    layer0_outputs(6825) <= not (a and b);
    layer0_outputs(6826) <= a and b;
    layer0_outputs(6827) <= not b;
    layer0_outputs(6828) <= a and not b;
    layer0_outputs(6829) <= not a;
    layer0_outputs(6830) <= not b or a;
    layer0_outputs(6831) <= not (a and b);
    layer0_outputs(6832) <= 1'b0;
    layer0_outputs(6833) <= a and b;
    layer0_outputs(6834) <= a xor b;
    layer0_outputs(6835) <= not (a or b);
    layer0_outputs(6836) <= a and b;
    layer0_outputs(6837) <= not b;
    layer0_outputs(6838) <= not (a or b);
    layer0_outputs(6839) <= not a or b;
    layer0_outputs(6840) <= not a or b;
    layer0_outputs(6841) <= not (a and b);
    layer0_outputs(6842) <= a;
    layer0_outputs(6843) <= a;
    layer0_outputs(6844) <= not b;
    layer0_outputs(6845) <= not (a xor b);
    layer0_outputs(6846) <= a;
    layer0_outputs(6847) <= 1'b1;
    layer0_outputs(6848) <= not a;
    layer0_outputs(6849) <= a or b;
    layer0_outputs(6850) <= a and b;
    layer0_outputs(6851) <= a and not b;
    layer0_outputs(6852) <= 1'b1;
    layer0_outputs(6853) <= not (a and b);
    layer0_outputs(6854) <= not (a and b);
    layer0_outputs(6855) <= a or b;
    layer0_outputs(6856) <= b and not a;
    layer0_outputs(6857) <= not b;
    layer0_outputs(6858) <= b and not a;
    layer0_outputs(6859) <= not (a and b);
    layer0_outputs(6860) <= b;
    layer0_outputs(6861) <= b and not a;
    layer0_outputs(6862) <= not b or a;
    layer0_outputs(6863) <= not a;
    layer0_outputs(6864) <= not (a xor b);
    layer0_outputs(6865) <= a;
    layer0_outputs(6866) <= not b;
    layer0_outputs(6867) <= a and b;
    layer0_outputs(6868) <= not (a and b);
    layer0_outputs(6869) <= not a;
    layer0_outputs(6870) <= a or b;
    layer0_outputs(6871) <= not (a or b);
    layer0_outputs(6872) <= not (a or b);
    layer0_outputs(6873) <= a;
    layer0_outputs(6874) <= not a or b;
    layer0_outputs(6875) <= not a or b;
    layer0_outputs(6876) <= b and not a;
    layer0_outputs(6877) <= not (a and b);
    layer0_outputs(6878) <= not b or a;
    layer0_outputs(6879) <= not (a xor b);
    layer0_outputs(6880) <= a;
    layer0_outputs(6881) <= 1'b0;
    layer0_outputs(6882) <= not a;
    layer0_outputs(6883) <= 1'b0;
    layer0_outputs(6884) <= 1'b1;
    layer0_outputs(6885) <= a and not b;
    layer0_outputs(6886) <= a or b;
    layer0_outputs(6887) <= not a;
    layer0_outputs(6888) <= not (a or b);
    layer0_outputs(6889) <= a;
    layer0_outputs(6890) <= not b;
    layer0_outputs(6891) <= a xor b;
    layer0_outputs(6892) <= a and not b;
    layer0_outputs(6893) <= a and b;
    layer0_outputs(6894) <= 1'b0;
    layer0_outputs(6895) <= a and b;
    layer0_outputs(6896) <= not a;
    layer0_outputs(6897) <= a or b;
    layer0_outputs(6898) <= b and not a;
    layer0_outputs(6899) <= 1'b1;
    layer0_outputs(6900) <= not (a xor b);
    layer0_outputs(6901) <= not (a xor b);
    layer0_outputs(6902) <= 1'b0;
    layer0_outputs(6903) <= not (a or b);
    layer0_outputs(6904) <= not (a xor b);
    layer0_outputs(6905) <= not b or a;
    layer0_outputs(6906) <= not a;
    layer0_outputs(6907) <= a and not b;
    layer0_outputs(6908) <= not b or a;
    layer0_outputs(6909) <= not (a and b);
    layer0_outputs(6910) <= a or b;
    layer0_outputs(6911) <= not (a and b);
    layer0_outputs(6912) <= b and not a;
    layer0_outputs(6913) <= a and b;
    layer0_outputs(6914) <= 1'b0;
    layer0_outputs(6915) <= a;
    layer0_outputs(6916) <= 1'b1;
    layer0_outputs(6917) <= a xor b;
    layer0_outputs(6918) <= not (a and b);
    layer0_outputs(6919) <= not b or a;
    layer0_outputs(6920) <= b and not a;
    layer0_outputs(6921) <= not (a and b);
    layer0_outputs(6922) <= not b or a;
    layer0_outputs(6923) <= b and not a;
    layer0_outputs(6924) <= 1'b0;
    layer0_outputs(6925) <= 1'b0;
    layer0_outputs(6926) <= a xor b;
    layer0_outputs(6927) <= not a;
    layer0_outputs(6928) <= not b or a;
    layer0_outputs(6929) <= not a or b;
    layer0_outputs(6930) <= not b or a;
    layer0_outputs(6931) <= a or b;
    layer0_outputs(6932) <= 1'b1;
    layer0_outputs(6933) <= not a or b;
    layer0_outputs(6934) <= not a or b;
    layer0_outputs(6935) <= not (a xor b);
    layer0_outputs(6936) <= b and not a;
    layer0_outputs(6937) <= a and b;
    layer0_outputs(6938) <= 1'b1;
    layer0_outputs(6939) <= b and not a;
    layer0_outputs(6940) <= 1'b0;
    layer0_outputs(6941) <= not b;
    layer0_outputs(6942) <= b and not a;
    layer0_outputs(6943) <= 1'b0;
    layer0_outputs(6944) <= a;
    layer0_outputs(6945) <= not (a and b);
    layer0_outputs(6946) <= not b or a;
    layer0_outputs(6947) <= not (a and b);
    layer0_outputs(6948) <= a;
    layer0_outputs(6949) <= not (a xor b);
    layer0_outputs(6950) <= b and not a;
    layer0_outputs(6951) <= a or b;
    layer0_outputs(6952) <= 1'b0;
    layer0_outputs(6953) <= a and b;
    layer0_outputs(6954) <= b and not a;
    layer0_outputs(6955) <= not (a and b);
    layer0_outputs(6956) <= a or b;
    layer0_outputs(6957) <= not b;
    layer0_outputs(6958) <= 1'b1;
    layer0_outputs(6959) <= not b or a;
    layer0_outputs(6960) <= not b or a;
    layer0_outputs(6961) <= not b or a;
    layer0_outputs(6962) <= b;
    layer0_outputs(6963) <= not (a or b);
    layer0_outputs(6964) <= a and b;
    layer0_outputs(6965) <= not a;
    layer0_outputs(6966) <= a xor b;
    layer0_outputs(6967) <= a and b;
    layer0_outputs(6968) <= a or b;
    layer0_outputs(6969) <= b;
    layer0_outputs(6970) <= not a or b;
    layer0_outputs(6971) <= a;
    layer0_outputs(6972) <= not (a xor b);
    layer0_outputs(6973) <= a xor b;
    layer0_outputs(6974) <= b;
    layer0_outputs(6975) <= a and b;
    layer0_outputs(6976) <= a or b;
    layer0_outputs(6977) <= b and not a;
    layer0_outputs(6978) <= a;
    layer0_outputs(6979) <= not b;
    layer0_outputs(6980) <= 1'b0;
    layer0_outputs(6981) <= a and b;
    layer0_outputs(6982) <= a and not b;
    layer0_outputs(6983) <= a and not b;
    layer0_outputs(6984) <= not a or b;
    layer0_outputs(6985) <= not (a or b);
    layer0_outputs(6986) <= a and b;
    layer0_outputs(6987) <= a and not b;
    layer0_outputs(6988) <= not b;
    layer0_outputs(6989) <= not b;
    layer0_outputs(6990) <= a xor b;
    layer0_outputs(6991) <= a or b;
    layer0_outputs(6992) <= not (a or b);
    layer0_outputs(6993) <= not (a and b);
    layer0_outputs(6994) <= 1'b0;
    layer0_outputs(6995) <= not b or a;
    layer0_outputs(6996) <= not b or a;
    layer0_outputs(6997) <= not b;
    layer0_outputs(6998) <= b;
    layer0_outputs(6999) <= 1'b0;
    layer0_outputs(7000) <= b;
    layer0_outputs(7001) <= b and not a;
    layer0_outputs(7002) <= not a;
    layer0_outputs(7003) <= b and not a;
    layer0_outputs(7004) <= a or b;
    layer0_outputs(7005) <= a and not b;
    layer0_outputs(7006) <= 1'b1;
    layer0_outputs(7007) <= not b;
    layer0_outputs(7008) <= not (a xor b);
    layer0_outputs(7009) <= a or b;
    layer0_outputs(7010) <= 1'b0;
    layer0_outputs(7011) <= a or b;
    layer0_outputs(7012) <= b and not a;
    layer0_outputs(7013) <= a or b;
    layer0_outputs(7014) <= not (a xor b);
    layer0_outputs(7015) <= not b;
    layer0_outputs(7016) <= a xor b;
    layer0_outputs(7017) <= 1'b0;
    layer0_outputs(7018) <= not a;
    layer0_outputs(7019) <= a xor b;
    layer0_outputs(7020) <= a or b;
    layer0_outputs(7021) <= not a or b;
    layer0_outputs(7022) <= 1'b0;
    layer0_outputs(7023) <= not b or a;
    layer0_outputs(7024) <= a or b;
    layer0_outputs(7025) <= not b or a;
    layer0_outputs(7026) <= not a;
    layer0_outputs(7027) <= not b or a;
    layer0_outputs(7028) <= a and not b;
    layer0_outputs(7029) <= a xor b;
    layer0_outputs(7030) <= b and not a;
    layer0_outputs(7031) <= 1'b0;
    layer0_outputs(7032) <= not b;
    layer0_outputs(7033) <= not (a xor b);
    layer0_outputs(7034) <= 1'b0;
    layer0_outputs(7035) <= not (a or b);
    layer0_outputs(7036) <= a or b;
    layer0_outputs(7037) <= not (a or b);
    layer0_outputs(7038) <= not a;
    layer0_outputs(7039) <= not (a xor b);
    layer0_outputs(7040) <= not (a and b);
    layer0_outputs(7041) <= not (a xor b);
    layer0_outputs(7042) <= not a;
    layer0_outputs(7043) <= not a or b;
    layer0_outputs(7044) <= a and b;
    layer0_outputs(7045) <= not (a or b);
    layer0_outputs(7046) <= not (a or b);
    layer0_outputs(7047) <= not (a xor b);
    layer0_outputs(7048) <= not a or b;
    layer0_outputs(7049) <= not b or a;
    layer0_outputs(7050) <= not b or a;
    layer0_outputs(7051) <= b;
    layer0_outputs(7052) <= not a;
    layer0_outputs(7053) <= a;
    layer0_outputs(7054) <= not a;
    layer0_outputs(7055) <= a or b;
    layer0_outputs(7056) <= a;
    layer0_outputs(7057) <= b;
    layer0_outputs(7058) <= a;
    layer0_outputs(7059) <= not a;
    layer0_outputs(7060) <= not (a and b);
    layer0_outputs(7061) <= not b;
    layer0_outputs(7062) <= not a;
    layer0_outputs(7063) <= not a;
    layer0_outputs(7064) <= a and not b;
    layer0_outputs(7065) <= a and b;
    layer0_outputs(7066) <= not a;
    layer0_outputs(7067) <= not b or a;
    layer0_outputs(7068) <= b and not a;
    layer0_outputs(7069) <= a and not b;
    layer0_outputs(7070) <= a xor b;
    layer0_outputs(7071) <= 1'b0;
    layer0_outputs(7072) <= a;
    layer0_outputs(7073) <= a or b;
    layer0_outputs(7074) <= b and not a;
    layer0_outputs(7075) <= b and not a;
    layer0_outputs(7076) <= b and not a;
    layer0_outputs(7077) <= a and not b;
    layer0_outputs(7078) <= a or b;
    layer0_outputs(7079) <= not a or b;
    layer0_outputs(7080) <= a and not b;
    layer0_outputs(7081) <= 1'b1;
    layer0_outputs(7082) <= 1'b0;
    layer0_outputs(7083) <= b and not a;
    layer0_outputs(7084) <= b and not a;
    layer0_outputs(7085) <= a and b;
    layer0_outputs(7086) <= 1'b1;
    layer0_outputs(7087) <= not b;
    layer0_outputs(7088) <= b and not a;
    layer0_outputs(7089) <= a and not b;
    layer0_outputs(7090) <= a and not b;
    layer0_outputs(7091) <= a and not b;
    layer0_outputs(7092) <= a or b;
    layer0_outputs(7093) <= not (a or b);
    layer0_outputs(7094) <= a;
    layer0_outputs(7095) <= not b or a;
    layer0_outputs(7096) <= b and not a;
    layer0_outputs(7097) <= a and not b;
    layer0_outputs(7098) <= not a;
    layer0_outputs(7099) <= not a or b;
    layer0_outputs(7100) <= not (a and b);
    layer0_outputs(7101) <= not a;
    layer0_outputs(7102) <= a;
    layer0_outputs(7103) <= a;
    layer0_outputs(7104) <= a and b;
    layer0_outputs(7105) <= not (a xor b);
    layer0_outputs(7106) <= b;
    layer0_outputs(7107) <= a and b;
    layer0_outputs(7108) <= b and not a;
    layer0_outputs(7109) <= b;
    layer0_outputs(7110) <= 1'b0;
    layer0_outputs(7111) <= not a or b;
    layer0_outputs(7112) <= not (a and b);
    layer0_outputs(7113) <= not a or b;
    layer0_outputs(7114) <= not (a or b);
    layer0_outputs(7115) <= not (a or b);
    layer0_outputs(7116) <= a and not b;
    layer0_outputs(7117) <= not (a and b);
    layer0_outputs(7118) <= b;
    layer0_outputs(7119) <= a or b;
    layer0_outputs(7120) <= b;
    layer0_outputs(7121) <= not (a or b);
    layer0_outputs(7122) <= b;
    layer0_outputs(7123) <= not (a or b);
    layer0_outputs(7124) <= not (a or b);
    layer0_outputs(7125) <= not a or b;
    layer0_outputs(7126) <= not a or b;
    layer0_outputs(7127) <= not b;
    layer0_outputs(7128) <= not a;
    layer0_outputs(7129) <= a;
    layer0_outputs(7130) <= 1'b0;
    layer0_outputs(7131) <= a;
    layer0_outputs(7132) <= not (a or b);
    layer0_outputs(7133) <= not a or b;
    layer0_outputs(7134) <= not (a or b);
    layer0_outputs(7135) <= not b or a;
    layer0_outputs(7136) <= not (a xor b);
    layer0_outputs(7137) <= a and b;
    layer0_outputs(7138) <= not a;
    layer0_outputs(7139) <= a and b;
    layer0_outputs(7140) <= b;
    layer0_outputs(7141) <= b;
    layer0_outputs(7142) <= a or b;
    layer0_outputs(7143) <= a and not b;
    layer0_outputs(7144) <= 1'b1;
    layer0_outputs(7145) <= not (a and b);
    layer0_outputs(7146) <= not b;
    layer0_outputs(7147) <= 1'b1;
    layer0_outputs(7148) <= 1'b1;
    layer0_outputs(7149) <= 1'b0;
    layer0_outputs(7150) <= 1'b1;
    layer0_outputs(7151) <= a or b;
    layer0_outputs(7152) <= not (a xor b);
    layer0_outputs(7153) <= not a or b;
    layer0_outputs(7154) <= a;
    layer0_outputs(7155) <= a;
    layer0_outputs(7156) <= b;
    layer0_outputs(7157) <= not (a and b);
    layer0_outputs(7158) <= not a;
    layer0_outputs(7159) <= b;
    layer0_outputs(7160) <= b;
    layer0_outputs(7161) <= not (a xor b);
    layer0_outputs(7162) <= not a or b;
    layer0_outputs(7163) <= a and not b;
    layer0_outputs(7164) <= 1'b0;
    layer0_outputs(7165) <= not a;
    layer0_outputs(7166) <= not (a or b);
    layer0_outputs(7167) <= not (a xor b);
    layer0_outputs(7168) <= not (a and b);
    layer0_outputs(7169) <= a and b;
    layer0_outputs(7170) <= a or b;
    layer0_outputs(7171) <= b and not a;
    layer0_outputs(7172) <= not (a and b);
    layer0_outputs(7173) <= b and not a;
    layer0_outputs(7174) <= not a or b;
    layer0_outputs(7175) <= a and not b;
    layer0_outputs(7176) <= a and b;
    layer0_outputs(7177) <= a xor b;
    layer0_outputs(7178) <= a or b;
    layer0_outputs(7179) <= b and not a;
    layer0_outputs(7180) <= a and b;
    layer0_outputs(7181) <= a or b;
    layer0_outputs(7182) <= not a or b;
    layer0_outputs(7183) <= not a or b;
    layer0_outputs(7184) <= a and not b;
    layer0_outputs(7185) <= a;
    layer0_outputs(7186) <= 1'b1;
    layer0_outputs(7187) <= not (a and b);
    layer0_outputs(7188) <= not (a or b);
    layer0_outputs(7189) <= not a;
    layer0_outputs(7190) <= not (a and b);
    layer0_outputs(7191) <= not b;
    layer0_outputs(7192) <= b;
    layer0_outputs(7193) <= 1'b0;
    layer0_outputs(7194) <= not (a or b);
    layer0_outputs(7195) <= 1'b0;
    layer0_outputs(7196) <= 1'b0;
    layer0_outputs(7197) <= a or b;
    layer0_outputs(7198) <= b and not a;
    layer0_outputs(7199) <= not (a or b);
    layer0_outputs(7200) <= a or b;
    layer0_outputs(7201) <= a;
    layer0_outputs(7202) <= a or b;
    layer0_outputs(7203) <= 1'b0;
    layer0_outputs(7204) <= 1'b1;
    layer0_outputs(7205) <= 1'b0;
    layer0_outputs(7206) <= not b or a;
    layer0_outputs(7207) <= 1'b0;
    layer0_outputs(7208) <= not b or a;
    layer0_outputs(7209) <= not (a or b);
    layer0_outputs(7210) <= not (a xor b);
    layer0_outputs(7211) <= a;
    layer0_outputs(7212) <= not (a xor b);
    layer0_outputs(7213) <= not a or b;
    layer0_outputs(7214) <= a or b;
    layer0_outputs(7215) <= a or b;
    layer0_outputs(7216) <= a;
    layer0_outputs(7217) <= not b;
    layer0_outputs(7218) <= a xor b;
    layer0_outputs(7219) <= not (a and b);
    layer0_outputs(7220) <= b;
    layer0_outputs(7221) <= a or b;
    layer0_outputs(7222) <= not (a and b);
    layer0_outputs(7223) <= a and not b;
    layer0_outputs(7224) <= a xor b;
    layer0_outputs(7225) <= b and not a;
    layer0_outputs(7226) <= not b;
    layer0_outputs(7227) <= b and not a;
    layer0_outputs(7228) <= a xor b;
    layer0_outputs(7229) <= a and not b;
    layer0_outputs(7230) <= not a;
    layer0_outputs(7231) <= a and not b;
    layer0_outputs(7232) <= b and not a;
    layer0_outputs(7233) <= not (a or b);
    layer0_outputs(7234) <= not b or a;
    layer0_outputs(7235) <= not b or a;
    layer0_outputs(7236) <= not b or a;
    layer0_outputs(7237) <= 1'b1;
    layer0_outputs(7238) <= a;
    layer0_outputs(7239) <= not (a and b);
    layer0_outputs(7240) <= not b or a;
    layer0_outputs(7241) <= not b or a;
    layer0_outputs(7242) <= 1'b1;
    layer0_outputs(7243) <= not b;
    layer0_outputs(7244) <= not (a xor b);
    layer0_outputs(7245) <= b;
    layer0_outputs(7246) <= a and b;
    layer0_outputs(7247) <= b;
    layer0_outputs(7248) <= not b or a;
    layer0_outputs(7249) <= not (a or b);
    layer0_outputs(7250) <= a and not b;
    layer0_outputs(7251) <= a or b;
    layer0_outputs(7252) <= a or b;
    layer0_outputs(7253) <= not a;
    layer0_outputs(7254) <= a or b;
    layer0_outputs(7255) <= 1'b1;
    layer0_outputs(7256) <= not b;
    layer0_outputs(7257) <= a;
    layer0_outputs(7258) <= a and b;
    layer0_outputs(7259) <= not (a or b);
    layer0_outputs(7260) <= not a or b;
    layer0_outputs(7261) <= a;
    layer0_outputs(7262) <= 1'b1;
    layer0_outputs(7263) <= 1'b1;
    layer0_outputs(7264) <= 1'b1;
    layer0_outputs(7265) <= not (a and b);
    layer0_outputs(7266) <= a or b;
    layer0_outputs(7267) <= not b;
    layer0_outputs(7268) <= a xor b;
    layer0_outputs(7269) <= 1'b1;
    layer0_outputs(7270) <= not a or b;
    layer0_outputs(7271) <= b;
    layer0_outputs(7272) <= not b or a;
    layer0_outputs(7273) <= not (a and b);
    layer0_outputs(7274) <= a;
    layer0_outputs(7275) <= not (a xor b);
    layer0_outputs(7276) <= not a or b;
    layer0_outputs(7277) <= b and not a;
    layer0_outputs(7278) <= 1'b1;
    layer0_outputs(7279) <= not (a xor b);
    layer0_outputs(7280) <= not (a xor b);
    layer0_outputs(7281) <= b;
    layer0_outputs(7282) <= a xor b;
    layer0_outputs(7283) <= a xor b;
    layer0_outputs(7284) <= not a or b;
    layer0_outputs(7285) <= a xor b;
    layer0_outputs(7286) <= not a;
    layer0_outputs(7287) <= a;
    layer0_outputs(7288) <= a;
    layer0_outputs(7289) <= 1'b1;
    layer0_outputs(7290) <= a xor b;
    layer0_outputs(7291) <= a xor b;
    layer0_outputs(7292) <= not a;
    layer0_outputs(7293) <= not a;
    layer0_outputs(7294) <= not b;
    layer0_outputs(7295) <= b;
    layer0_outputs(7296) <= not b or a;
    layer0_outputs(7297) <= 1'b1;
    layer0_outputs(7298) <= a;
    layer0_outputs(7299) <= b and not a;
    layer0_outputs(7300) <= b;
    layer0_outputs(7301) <= a;
    layer0_outputs(7302) <= not a or b;
    layer0_outputs(7303) <= not (a or b);
    layer0_outputs(7304) <= not (a and b);
    layer0_outputs(7305) <= 1'b0;
    layer0_outputs(7306) <= not (a xor b);
    layer0_outputs(7307) <= not b or a;
    layer0_outputs(7308) <= b;
    layer0_outputs(7309) <= not (a and b);
    layer0_outputs(7310) <= not b;
    layer0_outputs(7311) <= a or b;
    layer0_outputs(7312) <= a xor b;
    layer0_outputs(7313) <= not (a and b);
    layer0_outputs(7314) <= 1'b1;
    layer0_outputs(7315) <= not a;
    layer0_outputs(7316) <= not a;
    layer0_outputs(7317) <= 1'b0;
    layer0_outputs(7318) <= not (a or b);
    layer0_outputs(7319) <= b and not a;
    layer0_outputs(7320) <= 1'b0;
    layer0_outputs(7321) <= not b;
    layer0_outputs(7322) <= not b or a;
    layer0_outputs(7323) <= a and not b;
    layer0_outputs(7324) <= a;
    layer0_outputs(7325) <= not b;
    layer0_outputs(7326) <= a and not b;
    layer0_outputs(7327) <= not (a or b);
    layer0_outputs(7328) <= 1'b0;
    layer0_outputs(7329) <= a xor b;
    layer0_outputs(7330) <= a xor b;
    layer0_outputs(7331) <= a;
    layer0_outputs(7332) <= a and b;
    layer0_outputs(7333) <= not b or a;
    layer0_outputs(7334) <= not a or b;
    layer0_outputs(7335) <= not a;
    layer0_outputs(7336) <= not a or b;
    layer0_outputs(7337) <= b;
    layer0_outputs(7338) <= not (a xor b);
    layer0_outputs(7339) <= a and b;
    layer0_outputs(7340) <= 1'b0;
    layer0_outputs(7341) <= not b or a;
    layer0_outputs(7342) <= 1'b1;
    layer0_outputs(7343) <= not b;
    layer0_outputs(7344) <= b and not a;
    layer0_outputs(7345) <= 1'b1;
    layer0_outputs(7346) <= a or b;
    layer0_outputs(7347) <= not a or b;
    layer0_outputs(7348) <= a and b;
    layer0_outputs(7349) <= not b;
    layer0_outputs(7350) <= b;
    layer0_outputs(7351) <= a xor b;
    layer0_outputs(7352) <= not b or a;
    layer0_outputs(7353) <= not (a and b);
    layer0_outputs(7354) <= not (a xor b);
    layer0_outputs(7355) <= a and not b;
    layer0_outputs(7356) <= 1'b1;
    layer0_outputs(7357) <= not b or a;
    layer0_outputs(7358) <= b;
    layer0_outputs(7359) <= b;
    layer0_outputs(7360) <= a xor b;
    layer0_outputs(7361) <= not b or a;
    layer0_outputs(7362) <= a;
    layer0_outputs(7363) <= not a;
    layer0_outputs(7364) <= a and b;
    layer0_outputs(7365) <= a or b;
    layer0_outputs(7366) <= a or b;
    layer0_outputs(7367) <= not b;
    layer0_outputs(7368) <= 1'b1;
    layer0_outputs(7369) <= not a;
    layer0_outputs(7370) <= 1'b1;
    layer0_outputs(7371) <= not (a and b);
    layer0_outputs(7372) <= a or b;
    layer0_outputs(7373) <= 1'b1;
    layer0_outputs(7374) <= a xor b;
    layer0_outputs(7375) <= not b or a;
    layer0_outputs(7376) <= b;
    layer0_outputs(7377) <= not a;
    layer0_outputs(7378) <= not a;
    layer0_outputs(7379) <= a xor b;
    layer0_outputs(7380) <= b and not a;
    layer0_outputs(7381) <= not (a xor b);
    layer0_outputs(7382) <= a and not b;
    layer0_outputs(7383) <= a;
    layer0_outputs(7384) <= 1'b1;
    layer0_outputs(7385) <= b;
    layer0_outputs(7386) <= a and not b;
    layer0_outputs(7387) <= 1'b0;
    layer0_outputs(7388) <= not b;
    layer0_outputs(7389) <= b;
    layer0_outputs(7390) <= 1'b0;
    layer0_outputs(7391) <= not (a xor b);
    layer0_outputs(7392) <= not b or a;
    layer0_outputs(7393) <= not (a and b);
    layer0_outputs(7394) <= not a;
    layer0_outputs(7395) <= not (a and b);
    layer0_outputs(7396) <= a and b;
    layer0_outputs(7397) <= not a;
    layer0_outputs(7398) <= a and b;
    layer0_outputs(7399) <= 1'b0;
    layer0_outputs(7400) <= not b;
    layer0_outputs(7401) <= 1'b0;
    layer0_outputs(7402) <= not (a or b);
    layer0_outputs(7403) <= b and not a;
    layer0_outputs(7404) <= a and not b;
    layer0_outputs(7405) <= a or b;
    layer0_outputs(7406) <= a and not b;
    layer0_outputs(7407) <= not b;
    layer0_outputs(7408) <= not (a and b);
    layer0_outputs(7409) <= a xor b;
    layer0_outputs(7410) <= a and not b;
    layer0_outputs(7411) <= a xor b;
    layer0_outputs(7412) <= b;
    layer0_outputs(7413) <= not a or b;
    layer0_outputs(7414) <= a and b;
    layer0_outputs(7415) <= 1'b0;
    layer0_outputs(7416) <= 1'b0;
    layer0_outputs(7417) <= b;
    layer0_outputs(7418) <= not a or b;
    layer0_outputs(7419) <= not (a xor b);
    layer0_outputs(7420) <= a and not b;
    layer0_outputs(7421) <= not (a and b);
    layer0_outputs(7422) <= a or b;
    layer0_outputs(7423) <= a;
    layer0_outputs(7424) <= a;
    layer0_outputs(7425) <= 1'b1;
    layer0_outputs(7426) <= not a;
    layer0_outputs(7427) <= not (a and b);
    layer0_outputs(7428) <= a or b;
    layer0_outputs(7429) <= not a;
    layer0_outputs(7430) <= a and b;
    layer0_outputs(7431) <= not a or b;
    layer0_outputs(7432) <= a;
    layer0_outputs(7433) <= 1'b0;
    layer0_outputs(7434) <= b;
    layer0_outputs(7435) <= a xor b;
    layer0_outputs(7436) <= not a or b;
    layer0_outputs(7437) <= not (a and b);
    layer0_outputs(7438) <= a and b;
    layer0_outputs(7439) <= not b;
    layer0_outputs(7440) <= 1'b1;
    layer0_outputs(7441) <= b;
    layer0_outputs(7442) <= b;
    layer0_outputs(7443) <= b and not a;
    layer0_outputs(7444) <= 1'b1;
    layer0_outputs(7445) <= a and not b;
    layer0_outputs(7446) <= not (a and b);
    layer0_outputs(7447) <= a or b;
    layer0_outputs(7448) <= not a;
    layer0_outputs(7449) <= b;
    layer0_outputs(7450) <= 1'b1;
    layer0_outputs(7451) <= not a or b;
    layer0_outputs(7452) <= not (a or b);
    layer0_outputs(7453) <= a;
    layer0_outputs(7454) <= 1'b1;
    layer0_outputs(7455) <= not b or a;
    layer0_outputs(7456) <= a or b;
    layer0_outputs(7457) <= not (a or b);
    layer0_outputs(7458) <= not (a and b);
    layer0_outputs(7459) <= 1'b1;
    layer0_outputs(7460) <= b;
    layer0_outputs(7461) <= a xor b;
    layer0_outputs(7462) <= not b or a;
    layer0_outputs(7463) <= not a or b;
    layer0_outputs(7464) <= not b or a;
    layer0_outputs(7465) <= 1'b0;
    layer0_outputs(7466) <= b and not a;
    layer0_outputs(7467) <= a and b;
    layer0_outputs(7468) <= b;
    layer0_outputs(7469) <= not a;
    layer0_outputs(7470) <= not (a and b);
    layer0_outputs(7471) <= a or b;
    layer0_outputs(7472) <= a xor b;
    layer0_outputs(7473) <= a and not b;
    layer0_outputs(7474) <= not b or a;
    layer0_outputs(7475) <= not (a xor b);
    layer0_outputs(7476) <= b and not a;
    layer0_outputs(7477) <= 1'b0;
    layer0_outputs(7478) <= not (a or b);
    layer0_outputs(7479) <= b;
    layer0_outputs(7480) <= a or b;
    layer0_outputs(7481) <= not b;
    layer0_outputs(7482) <= b and not a;
    layer0_outputs(7483) <= 1'b0;
    layer0_outputs(7484) <= b;
    layer0_outputs(7485) <= not b or a;
    layer0_outputs(7486) <= not b or a;
    layer0_outputs(7487) <= not a;
    layer0_outputs(7488) <= 1'b1;
    layer0_outputs(7489) <= not a or b;
    layer0_outputs(7490) <= not (a or b);
    layer0_outputs(7491) <= b and not a;
    layer0_outputs(7492) <= not a;
    layer0_outputs(7493) <= a xor b;
    layer0_outputs(7494) <= a;
    layer0_outputs(7495) <= not (a and b);
    layer0_outputs(7496) <= not (a xor b);
    layer0_outputs(7497) <= a xor b;
    layer0_outputs(7498) <= not a or b;
    layer0_outputs(7499) <= not b;
    layer0_outputs(7500) <= a and not b;
    layer0_outputs(7501) <= not a or b;
    layer0_outputs(7502) <= b;
    layer0_outputs(7503) <= not (a and b);
    layer0_outputs(7504) <= 1'b1;
    layer0_outputs(7505) <= not a or b;
    layer0_outputs(7506) <= not (a and b);
    layer0_outputs(7507) <= not (a or b);
    layer0_outputs(7508) <= not (a or b);
    layer0_outputs(7509) <= 1'b0;
    layer0_outputs(7510) <= 1'b1;
    layer0_outputs(7511) <= a and not b;
    layer0_outputs(7512) <= not b;
    layer0_outputs(7513) <= not a or b;
    layer0_outputs(7514) <= a and b;
    layer0_outputs(7515) <= not a or b;
    layer0_outputs(7516) <= not b or a;
    layer0_outputs(7517) <= not b or a;
    layer0_outputs(7518) <= not b;
    layer0_outputs(7519) <= a and not b;
    layer0_outputs(7520) <= not (a or b);
    layer0_outputs(7521) <= not (a xor b);
    layer0_outputs(7522) <= a and not b;
    layer0_outputs(7523) <= a;
    layer0_outputs(7524) <= 1'b1;
    layer0_outputs(7525) <= 1'b0;
    layer0_outputs(7526) <= 1'b1;
    layer0_outputs(7527) <= 1'b1;
    layer0_outputs(7528) <= not (a or b);
    layer0_outputs(7529) <= a and b;
    layer0_outputs(7530) <= not (a and b);
    layer0_outputs(7531) <= a xor b;
    layer0_outputs(7532) <= not b;
    layer0_outputs(7533) <= not (a xor b);
    layer0_outputs(7534) <= 1'b1;
    layer0_outputs(7535) <= a;
    layer0_outputs(7536) <= b;
    layer0_outputs(7537) <= a and not b;
    layer0_outputs(7538) <= 1'b0;
    layer0_outputs(7539) <= not a;
    layer0_outputs(7540) <= a or b;
    layer0_outputs(7541) <= not a;
    layer0_outputs(7542) <= not a or b;
    layer0_outputs(7543) <= 1'b1;
    layer0_outputs(7544) <= 1'b1;
    layer0_outputs(7545) <= 1'b0;
    layer0_outputs(7546) <= not (a or b);
    layer0_outputs(7547) <= not a or b;
    layer0_outputs(7548) <= not b or a;
    layer0_outputs(7549) <= 1'b0;
    layer0_outputs(7550) <= not b;
    layer0_outputs(7551) <= not (a and b);
    layer0_outputs(7552) <= not a or b;
    layer0_outputs(7553) <= a xor b;
    layer0_outputs(7554) <= not b;
    layer0_outputs(7555) <= not (a and b);
    layer0_outputs(7556) <= not (a or b);
    layer0_outputs(7557) <= not b;
    layer0_outputs(7558) <= not b or a;
    layer0_outputs(7559) <= a and not b;
    layer0_outputs(7560) <= not b;
    layer0_outputs(7561) <= not (a or b);
    layer0_outputs(7562) <= a or b;
    layer0_outputs(7563) <= not b or a;
    layer0_outputs(7564) <= not a or b;
    layer0_outputs(7565) <= a xor b;
    layer0_outputs(7566) <= not (a or b);
    layer0_outputs(7567) <= not a;
    layer0_outputs(7568) <= a xor b;
    layer0_outputs(7569) <= b and not a;
    layer0_outputs(7570) <= not b or a;
    layer0_outputs(7571) <= not b or a;
    layer0_outputs(7572) <= a;
    layer0_outputs(7573) <= a xor b;
    layer0_outputs(7574) <= not a or b;
    layer0_outputs(7575) <= not b or a;
    layer0_outputs(7576) <= not b;
    layer0_outputs(7577) <= a or b;
    layer0_outputs(7578) <= 1'b1;
    layer0_outputs(7579) <= a xor b;
    layer0_outputs(7580) <= 1'b0;
    layer0_outputs(7581) <= not b or a;
    layer0_outputs(7582) <= not b;
    layer0_outputs(7583) <= not a;
    layer0_outputs(7584) <= not (a or b);
    layer0_outputs(7585) <= not a;
    layer0_outputs(7586) <= not b or a;
    layer0_outputs(7587) <= not b;
    layer0_outputs(7588) <= 1'b1;
    layer0_outputs(7589) <= not (a xor b);
    layer0_outputs(7590) <= b;
    layer0_outputs(7591) <= a xor b;
    layer0_outputs(7592) <= a xor b;
    layer0_outputs(7593) <= not a;
    layer0_outputs(7594) <= a or b;
    layer0_outputs(7595) <= a xor b;
    layer0_outputs(7596) <= not a;
    layer0_outputs(7597) <= not (a or b);
    layer0_outputs(7598) <= not (a and b);
    layer0_outputs(7599) <= a or b;
    layer0_outputs(7600) <= not a;
    layer0_outputs(7601) <= not b or a;
    layer0_outputs(7602) <= not a;
    layer0_outputs(7603) <= not b or a;
    layer0_outputs(7604) <= not b;
    layer0_outputs(7605) <= b and not a;
    layer0_outputs(7606) <= 1'b1;
    layer0_outputs(7607) <= not (a and b);
    layer0_outputs(7608) <= b;
    layer0_outputs(7609) <= not (a or b);
    layer0_outputs(7610) <= b;
    layer0_outputs(7611) <= b and not a;
    layer0_outputs(7612) <= 1'b1;
    layer0_outputs(7613) <= a and not b;
    layer0_outputs(7614) <= a;
    layer0_outputs(7615) <= b;
    layer0_outputs(7616) <= not (a or b);
    layer0_outputs(7617) <= a;
    layer0_outputs(7618) <= not (a or b);
    layer0_outputs(7619) <= not b;
    layer0_outputs(7620) <= not (a or b);
    layer0_outputs(7621) <= a and not b;
    layer0_outputs(7622) <= a and not b;
    layer0_outputs(7623) <= not (a xor b);
    layer0_outputs(7624) <= 1'b1;
    layer0_outputs(7625) <= 1'b0;
    layer0_outputs(7626) <= not a;
    layer0_outputs(7627) <= not b or a;
    layer0_outputs(7628) <= a and b;
    layer0_outputs(7629) <= 1'b0;
    layer0_outputs(7630) <= not (a and b);
    layer0_outputs(7631) <= not (a and b);
    layer0_outputs(7632) <= a xor b;
    layer0_outputs(7633) <= not (a and b);
    layer0_outputs(7634) <= a xor b;
    layer0_outputs(7635) <= not a or b;
    layer0_outputs(7636) <= not a;
    layer0_outputs(7637) <= a xor b;
    layer0_outputs(7638) <= b and not a;
    layer0_outputs(7639) <= not (a or b);
    layer0_outputs(7640) <= a or b;
    layer0_outputs(7641) <= not b or a;
    layer0_outputs(7642) <= not b or a;
    layer0_outputs(7643) <= a and not b;
    layer0_outputs(7644) <= not (a and b);
    layer0_outputs(7645) <= b;
    layer0_outputs(7646) <= a and not b;
    layer0_outputs(7647) <= not a;
    layer0_outputs(7648) <= 1'b0;
    layer0_outputs(7649) <= a;
    layer0_outputs(7650) <= not b or a;
    layer0_outputs(7651) <= not a;
    layer0_outputs(7652) <= not (a or b);
    layer0_outputs(7653) <= not b or a;
    layer0_outputs(7654) <= b;
    layer0_outputs(7655) <= 1'b1;
    layer0_outputs(7656) <= not b;
    layer0_outputs(7657) <= not (a or b);
    layer0_outputs(7658) <= 1'b1;
    layer0_outputs(7659) <= not a;
    layer0_outputs(7660) <= not b or a;
    layer0_outputs(7661) <= 1'b1;
    layer0_outputs(7662) <= b;
    layer0_outputs(7663) <= a and b;
    layer0_outputs(7664) <= a or b;
    layer0_outputs(7665) <= a and b;
    layer0_outputs(7666) <= not b;
    layer0_outputs(7667) <= a xor b;
    layer0_outputs(7668) <= not (a and b);
    layer0_outputs(7669) <= a and not b;
    layer0_outputs(7670) <= a;
    layer0_outputs(7671) <= 1'b0;
    layer0_outputs(7672) <= a;
    layer0_outputs(7673) <= not a;
    layer0_outputs(7674) <= a and not b;
    layer0_outputs(7675) <= not (a xor b);
    layer0_outputs(7676) <= not (a and b);
    layer0_outputs(7677) <= not b;
    layer0_outputs(7678) <= not a;
    layer0_outputs(7679) <= b;
    layer0_outputs(7680) <= b and not a;
    layer0_outputs(7681) <= a;
    layer0_outputs(7682) <= 1'b1;
    layer0_outputs(7683) <= not b;
    layer0_outputs(7684) <= 1'b0;
    layer0_outputs(7685) <= not a or b;
    layer0_outputs(7686) <= a xor b;
    layer0_outputs(7687) <= b;
    layer0_outputs(7688) <= 1'b1;
    layer0_outputs(7689) <= not (a or b);
    layer0_outputs(7690) <= 1'b0;
    layer0_outputs(7691) <= not a;
    layer0_outputs(7692) <= not (a or b);
    layer0_outputs(7693) <= not a or b;
    layer0_outputs(7694) <= b and not a;
    layer0_outputs(7695) <= not a or b;
    layer0_outputs(7696) <= a;
    layer0_outputs(7697) <= a and not b;
    layer0_outputs(7698) <= not a;
    layer0_outputs(7699) <= not a or b;
    layer0_outputs(7700) <= b;
    layer0_outputs(7701) <= not b;
    layer0_outputs(7702) <= 1'b1;
    layer0_outputs(7703) <= a or b;
    layer0_outputs(7704) <= a;
    layer0_outputs(7705) <= a and not b;
    layer0_outputs(7706) <= not b;
    layer0_outputs(7707) <= b;
    layer0_outputs(7708) <= b;
    layer0_outputs(7709) <= 1'b0;
    layer0_outputs(7710) <= not a;
    layer0_outputs(7711) <= not b or a;
    layer0_outputs(7712) <= b;
    layer0_outputs(7713) <= a and b;
    layer0_outputs(7714) <= not b;
    layer0_outputs(7715) <= not a;
    layer0_outputs(7716) <= b and not a;
    layer0_outputs(7717) <= a and not b;
    layer0_outputs(7718) <= b and not a;
    layer0_outputs(7719) <= 1'b0;
    layer0_outputs(7720) <= not a;
    layer0_outputs(7721) <= not (a and b);
    layer0_outputs(7722) <= a xor b;
    layer0_outputs(7723) <= not b;
    layer0_outputs(7724) <= not (a or b);
    layer0_outputs(7725) <= a and b;
    layer0_outputs(7726) <= not b or a;
    layer0_outputs(7727) <= a;
    layer0_outputs(7728) <= 1'b0;
    layer0_outputs(7729) <= b;
    layer0_outputs(7730) <= b and not a;
    layer0_outputs(7731) <= not (a and b);
    layer0_outputs(7732) <= 1'b1;
    layer0_outputs(7733) <= 1'b0;
    layer0_outputs(7734) <= a and not b;
    layer0_outputs(7735) <= a and b;
    layer0_outputs(7736) <= not a or b;
    layer0_outputs(7737) <= 1'b0;
    layer0_outputs(7738) <= 1'b1;
    layer0_outputs(7739) <= not a or b;
    layer0_outputs(7740) <= not (a and b);
    layer0_outputs(7741) <= not b or a;
    layer0_outputs(7742) <= 1'b1;
    layer0_outputs(7743) <= not b;
    layer0_outputs(7744) <= not b;
    layer0_outputs(7745) <= not a;
    layer0_outputs(7746) <= a or b;
    layer0_outputs(7747) <= b and not a;
    layer0_outputs(7748) <= a;
    layer0_outputs(7749) <= b and not a;
    layer0_outputs(7750) <= b;
    layer0_outputs(7751) <= a xor b;
    layer0_outputs(7752) <= a;
    layer0_outputs(7753) <= b;
    layer0_outputs(7754) <= not (a or b);
    layer0_outputs(7755) <= not a or b;
    layer0_outputs(7756) <= not a;
    layer0_outputs(7757) <= 1'b1;
    layer0_outputs(7758) <= b;
    layer0_outputs(7759) <= not a or b;
    layer0_outputs(7760) <= a xor b;
    layer0_outputs(7761) <= not (a xor b);
    layer0_outputs(7762) <= b;
    layer0_outputs(7763) <= a or b;
    layer0_outputs(7764) <= 1'b0;
    layer0_outputs(7765) <= b;
    layer0_outputs(7766) <= a;
    layer0_outputs(7767) <= 1'b0;
    layer0_outputs(7768) <= not b or a;
    layer0_outputs(7769) <= a or b;
    layer0_outputs(7770) <= a xor b;
    layer0_outputs(7771) <= b;
    layer0_outputs(7772) <= 1'b1;
    layer0_outputs(7773) <= 1'b0;
    layer0_outputs(7774) <= not (a or b);
    layer0_outputs(7775) <= a and not b;
    layer0_outputs(7776) <= not (a or b);
    layer0_outputs(7777) <= a and not b;
    layer0_outputs(7778) <= not (a and b);
    layer0_outputs(7779) <= a xor b;
    layer0_outputs(7780) <= not a;
    layer0_outputs(7781) <= a or b;
    layer0_outputs(7782) <= a xor b;
    layer0_outputs(7783) <= a xor b;
    layer0_outputs(7784) <= 1'b0;
    layer0_outputs(7785) <= a or b;
    layer0_outputs(7786) <= a or b;
    layer0_outputs(7787) <= b and not a;
    layer0_outputs(7788) <= b;
    layer0_outputs(7789) <= a;
    layer0_outputs(7790) <= a and not b;
    layer0_outputs(7791) <= not a or b;
    layer0_outputs(7792) <= not (a or b);
    layer0_outputs(7793) <= a or b;
    layer0_outputs(7794) <= 1'b1;
    layer0_outputs(7795) <= b;
    layer0_outputs(7796) <= not b;
    layer0_outputs(7797) <= not b;
    layer0_outputs(7798) <= not (a xor b);
    layer0_outputs(7799) <= not a or b;
    layer0_outputs(7800) <= b;
    layer0_outputs(7801) <= not b;
    layer0_outputs(7802) <= a or b;
    layer0_outputs(7803) <= not b;
    layer0_outputs(7804) <= b;
    layer0_outputs(7805) <= a and b;
    layer0_outputs(7806) <= not b;
    layer0_outputs(7807) <= not (a xor b);
    layer0_outputs(7808) <= not (a xor b);
    layer0_outputs(7809) <= 1'b1;
    layer0_outputs(7810) <= not (a and b);
    layer0_outputs(7811) <= not (a and b);
    layer0_outputs(7812) <= not (a or b);
    layer0_outputs(7813) <= not (a and b);
    layer0_outputs(7814) <= 1'b0;
    layer0_outputs(7815) <= a and not b;
    layer0_outputs(7816) <= a and b;
    layer0_outputs(7817) <= not (a and b);
    layer0_outputs(7818) <= 1'b0;
    layer0_outputs(7819) <= b and not a;
    layer0_outputs(7820) <= 1'b1;
    layer0_outputs(7821) <= a and b;
    layer0_outputs(7822) <= a and b;
    layer0_outputs(7823) <= not b or a;
    layer0_outputs(7824) <= not (a or b);
    layer0_outputs(7825) <= b;
    layer0_outputs(7826) <= not (a xor b);
    layer0_outputs(7827) <= not (a xor b);
    layer0_outputs(7828) <= 1'b1;
    layer0_outputs(7829) <= b and not a;
    layer0_outputs(7830) <= 1'b1;
    layer0_outputs(7831) <= not a or b;
    layer0_outputs(7832) <= b and not a;
    layer0_outputs(7833) <= 1'b0;
    layer0_outputs(7834) <= not (a and b);
    layer0_outputs(7835) <= b;
    layer0_outputs(7836) <= not a or b;
    layer0_outputs(7837) <= a and b;
    layer0_outputs(7838) <= a and not b;
    layer0_outputs(7839) <= 1'b1;
    layer0_outputs(7840) <= b and not a;
    layer0_outputs(7841) <= not (a and b);
    layer0_outputs(7842) <= not (a or b);
    layer0_outputs(7843) <= not b;
    layer0_outputs(7844) <= a xor b;
    layer0_outputs(7845) <= 1'b0;
    layer0_outputs(7846) <= a;
    layer0_outputs(7847) <= not b or a;
    layer0_outputs(7848) <= not b;
    layer0_outputs(7849) <= not (a and b);
    layer0_outputs(7850) <= not b;
    layer0_outputs(7851) <= not b or a;
    layer0_outputs(7852) <= a or b;
    layer0_outputs(7853) <= not b;
    layer0_outputs(7854) <= b and not a;
    layer0_outputs(7855) <= a xor b;
    layer0_outputs(7856) <= a or b;
    layer0_outputs(7857) <= 1'b0;
    layer0_outputs(7858) <= not (a or b);
    layer0_outputs(7859) <= a and b;
    layer0_outputs(7860) <= a and not b;
    layer0_outputs(7861) <= a;
    layer0_outputs(7862) <= a xor b;
    layer0_outputs(7863) <= not (a or b);
    layer0_outputs(7864) <= not (a or b);
    layer0_outputs(7865) <= 1'b1;
    layer0_outputs(7866) <= a or b;
    layer0_outputs(7867) <= b;
    layer0_outputs(7868) <= a;
    layer0_outputs(7869) <= a and b;
    layer0_outputs(7870) <= a and not b;
    layer0_outputs(7871) <= a xor b;
    layer0_outputs(7872) <= not a or b;
    layer0_outputs(7873) <= b and not a;
    layer0_outputs(7874) <= b;
    layer0_outputs(7875) <= a and b;
    layer0_outputs(7876) <= a and not b;
    layer0_outputs(7877) <= not b or a;
    layer0_outputs(7878) <= not b or a;
    layer0_outputs(7879) <= a and b;
    layer0_outputs(7880) <= b and not a;
    layer0_outputs(7881) <= not b;
    layer0_outputs(7882) <= b;
    layer0_outputs(7883) <= not a or b;
    layer0_outputs(7884) <= not (a or b);
    layer0_outputs(7885) <= not (a and b);
    layer0_outputs(7886) <= not b or a;
    layer0_outputs(7887) <= not (a xor b);
    layer0_outputs(7888) <= not (a and b);
    layer0_outputs(7889) <= 1'b0;
    layer0_outputs(7890) <= 1'b0;
    layer0_outputs(7891) <= a or b;
    layer0_outputs(7892) <= a and not b;
    layer0_outputs(7893) <= a or b;
    layer0_outputs(7894) <= a and not b;
    layer0_outputs(7895) <= a;
    layer0_outputs(7896) <= a and b;
    layer0_outputs(7897) <= a or b;
    layer0_outputs(7898) <= not a;
    layer0_outputs(7899) <= 1'b0;
    layer0_outputs(7900) <= a or b;
    layer0_outputs(7901) <= a and not b;
    layer0_outputs(7902) <= not a or b;
    layer0_outputs(7903) <= not a;
    layer0_outputs(7904) <= 1'b0;
    layer0_outputs(7905) <= not (a xor b);
    layer0_outputs(7906) <= not (a and b);
    layer0_outputs(7907) <= not (a and b);
    layer0_outputs(7908) <= 1'b0;
    layer0_outputs(7909) <= b;
    layer0_outputs(7910) <= a or b;
    layer0_outputs(7911) <= not a or b;
    layer0_outputs(7912) <= a or b;
    layer0_outputs(7913) <= not (a and b);
    layer0_outputs(7914) <= a xor b;
    layer0_outputs(7915) <= 1'b0;
    layer0_outputs(7916) <= not a;
    layer0_outputs(7917) <= a or b;
    layer0_outputs(7918) <= 1'b0;
    layer0_outputs(7919) <= 1'b1;
    layer0_outputs(7920) <= not (a and b);
    layer0_outputs(7921) <= a or b;
    layer0_outputs(7922) <= not (a or b);
    layer0_outputs(7923) <= not b or a;
    layer0_outputs(7924) <= not b;
    layer0_outputs(7925) <= 1'b0;
    layer0_outputs(7926) <= b;
    layer0_outputs(7927) <= not a;
    layer0_outputs(7928) <= a and b;
    layer0_outputs(7929) <= not (a xor b);
    layer0_outputs(7930) <= a and b;
    layer0_outputs(7931) <= a and b;
    layer0_outputs(7932) <= a xor b;
    layer0_outputs(7933) <= 1'b0;
    layer0_outputs(7934) <= a;
    layer0_outputs(7935) <= not (a xor b);
    layer0_outputs(7936) <= not (a or b);
    layer0_outputs(7937) <= not a;
    layer0_outputs(7938) <= not a;
    layer0_outputs(7939) <= 1'b1;
    layer0_outputs(7940) <= not b or a;
    layer0_outputs(7941) <= a;
    layer0_outputs(7942) <= a and b;
    layer0_outputs(7943) <= a;
    layer0_outputs(7944) <= not b;
    layer0_outputs(7945) <= b and not a;
    layer0_outputs(7946) <= not b or a;
    layer0_outputs(7947) <= b and not a;
    layer0_outputs(7948) <= a and b;
    layer0_outputs(7949) <= not (a xor b);
    layer0_outputs(7950) <= b and not a;
    layer0_outputs(7951) <= a and b;
    layer0_outputs(7952) <= not b or a;
    layer0_outputs(7953) <= 1'b1;
    layer0_outputs(7954) <= 1'b0;
    layer0_outputs(7955) <= not a;
    layer0_outputs(7956) <= 1'b0;
    layer0_outputs(7957) <= not b;
    layer0_outputs(7958) <= a and b;
    layer0_outputs(7959) <= a or b;
    layer0_outputs(7960) <= a and not b;
    layer0_outputs(7961) <= b and not a;
    layer0_outputs(7962) <= 1'b1;
    layer0_outputs(7963) <= not a or b;
    layer0_outputs(7964) <= not b;
    layer0_outputs(7965) <= not b;
    layer0_outputs(7966) <= b;
    layer0_outputs(7967) <= a xor b;
    layer0_outputs(7968) <= a;
    layer0_outputs(7969) <= 1'b0;
    layer0_outputs(7970) <= a;
    layer0_outputs(7971) <= not (a and b);
    layer0_outputs(7972) <= not (a and b);
    layer0_outputs(7973) <= not b;
    layer0_outputs(7974) <= b and not a;
    layer0_outputs(7975) <= not (a xor b);
    layer0_outputs(7976) <= not (a and b);
    layer0_outputs(7977) <= b and not a;
    layer0_outputs(7978) <= a;
    layer0_outputs(7979) <= not a or b;
    layer0_outputs(7980) <= not b;
    layer0_outputs(7981) <= 1'b1;
    layer0_outputs(7982) <= a xor b;
    layer0_outputs(7983) <= 1'b1;
    layer0_outputs(7984) <= b;
    layer0_outputs(7985) <= not a;
    layer0_outputs(7986) <= 1'b0;
    layer0_outputs(7987) <= b;
    layer0_outputs(7988) <= a or b;
    layer0_outputs(7989) <= not (a and b);
    layer0_outputs(7990) <= a;
    layer0_outputs(7991) <= not (a and b);
    layer0_outputs(7992) <= a xor b;
    layer0_outputs(7993) <= b;
    layer0_outputs(7994) <= not (a or b);
    layer0_outputs(7995) <= not (a or b);
    layer0_outputs(7996) <= not (a or b);
    layer0_outputs(7997) <= a and not b;
    layer0_outputs(7998) <= not a or b;
    layer0_outputs(7999) <= not b or a;
    layer0_outputs(8000) <= not (a or b);
    layer0_outputs(8001) <= a and not b;
    layer0_outputs(8002) <= not a;
    layer0_outputs(8003) <= not (a xor b);
    layer0_outputs(8004) <= 1'b1;
    layer0_outputs(8005) <= 1'b0;
    layer0_outputs(8006) <= not (a and b);
    layer0_outputs(8007) <= not (a or b);
    layer0_outputs(8008) <= 1'b1;
    layer0_outputs(8009) <= not a;
    layer0_outputs(8010) <= not (a xor b);
    layer0_outputs(8011) <= 1'b1;
    layer0_outputs(8012) <= a or b;
    layer0_outputs(8013) <= a or b;
    layer0_outputs(8014) <= b;
    layer0_outputs(8015) <= a;
    layer0_outputs(8016) <= not b or a;
    layer0_outputs(8017) <= not (a or b);
    layer0_outputs(8018) <= 1'b0;
    layer0_outputs(8019) <= not (a and b);
    layer0_outputs(8020) <= a or b;
    layer0_outputs(8021) <= a or b;
    layer0_outputs(8022) <= not b or a;
    layer0_outputs(8023) <= not b;
    layer0_outputs(8024) <= 1'b0;
    layer0_outputs(8025) <= not b or a;
    layer0_outputs(8026) <= b;
    layer0_outputs(8027) <= not a or b;
    layer0_outputs(8028) <= b and not a;
    layer0_outputs(8029) <= not a or b;
    layer0_outputs(8030) <= a or b;
    layer0_outputs(8031) <= a or b;
    layer0_outputs(8032) <= a and b;
    layer0_outputs(8033) <= 1'b0;
    layer0_outputs(8034) <= not (a or b);
    layer0_outputs(8035) <= not (a xor b);
    layer0_outputs(8036) <= 1'b1;
    layer0_outputs(8037) <= a;
    layer0_outputs(8038) <= not (a or b);
    layer0_outputs(8039) <= not a;
    layer0_outputs(8040) <= not (a and b);
    layer0_outputs(8041) <= not a;
    layer0_outputs(8042) <= not a or b;
    layer0_outputs(8043) <= b;
    layer0_outputs(8044) <= not (a xor b);
    layer0_outputs(8045) <= not b or a;
    layer0_outputs(8046) <= not a;
    layer0_outputs(8047) <= 1'b0;
    layer0_outputs(8048) <= not b or a;
    layer0_outputs(8049) <= 1'b0;
    layer0_outputs(8050) <= a or b;
    layer0_outputs(8051) <= a and b;
    layer0_outputs(8052) <= a and b;
    layer0_outputs(8053) <= 1'b0;
    layer0_outputs(8054) <= a;
    layer0_outputs(8055) <= not b or a;
    layer0_outputs(8056) <= not (a or b);
    layer0_outputs(8057) <= b;
    layer0_outputs(8058) <= not b;
    layer0_outputs(8059) <= a or b;
    layer0_outputs(8060) <= not (a and b);
    layer0_outputs(8061) <= 1'b0;
    layer0_outputs(8062) <= a;
    layer0_outputs(8063) <= b;
    layer0_outputs(8064) <= not (a xor b);
    layer0_outputs(8065) <= not b or a;
    layer0_outputs(8066) <= not (a and b);
    layer0_outputs(8067) <= not b or a;
    layer0_outputs(8068) <= not a;
    layer0_outputs(8069) <= a;
    layer0_outputs(8070) <= 1'b0;
    layer0_outputs(8071) <= a or b;
    layer0_outputs(8072) <= not a or b;
    layer0_outputs(8073) <= not b;
    layer0_outputs(8074) <= 1'b1;
    layer0_outputs(8075) <= a xor b;
    layer0_outputs(8076) <= not (a or b);
    layer0_outputs(8077) <= b and not a;
    layer0_outputs(8078) <= not b or a;
    layer0_outputs(8079) <= a xor b;
    layer0_outputs(8080) <= a or b;
    layer0_outputs(8081) <= not a or b;
    layer0_outputs(8082) <= a;
    layer0_outputs(8083) <= 1'b0;
    layer0_outputs(8084) <= a xor b;
    layer0_outputs(8085) <= b and not a;
    layer0_outputs(8086) <= not a;
    layer0_outputs(8087) <= not b;
    layer0_outputs(8088) <= 1'b1;
    layer0_outputs(8089) <= a and not b;
    layer0_outputs(8090) <= b;
    layer0_outputs(8091) <= a and b;
    layer0_outputs(8092) <= a xor b;
    layer0_outputs(8093) <= a;
    layer0_outputs(8094) <= not b;
    layer0_outputs(8095) <= b;
    layer0_outputs(8096) <= not (a xor b);
    layer0_outputs(8097) <= 1'b0;
    layer0_outputs(8098) <= not b;
    layer0_outputs(8099) <= a or b;
    layer0_outputs(8100) <= a and b;
    layer0_outputs(8101) <= b;
    layer0_outputs(8102) <= 1'b0;
    layer0_outputs(8103) <= not (a or b);
    layer0_outputs(8104) <= not b or a;
    layer0_outputs(8105) <= not a;
    layer0_outputs(8106) <= 1'b1;
    layer0_outputs(8107) <= a and not b;
    layer0_outputs(8108) <= a;
    layer0_outputs(8109) <= 1'b0;
    layer0_outputs(8110) <= not b or a;
    layer0_outputs(8111) <= a;
    layer0_outputs(8112) <= a;
    layer0_outputs(8113) <= not (a xor b);
    layer0_outputs(8114) <= a and not b;
    layer0_outputs(8115) <= not b;
    layer0_outputs(8116) <= not (a and b);
    layer0_outputs(8117) <= not (a or b);
    layer0_outputs(8118) <= b and not a;
    layer0_outputs(8119) <= not (a and b);
    layer0_outputs(8120) <= 1'b0;
    layer0_outputs(8121) <= a xor b;
    layer0_outputs(8122) <= not a;
    layer0_outputs(8123) <= b;
    layer0_outputs(8124) <= not b;
    layer0_outputs(8125) <= not (a or b);
    layer0_outputs(8126) <= a or b;
    layer0_outputs(8127) <= b;
    layer0_outputs(8128) <= a;
    layer0_outputs(8129) <= a and not b;
    layer0_outputs(8130) <= not (a and b);
    layer0_outputs(8131) <= not b;
    layer0_outputs(8132) <= b;
    layer0_outputs(8133) <= not a;
    layer0_outputs(8134) <= b;
    layer0_outputs(8135) <= a and not b;
    layer0_outputs(8136) <= 1'b1;
    layer0_outputs(8137) <= not b;
    layer0_outputs(8138) <= not (a or b);
    layer0_outputs(8139) <= not a;
    layer0_outputs(8140) <= 1'b1;
    layer0_outputs(8141) <= not (a xor b);
    layer0_outputs(8142) <= 1'b1;
    layer0_outputs(8143) <= 1'b1;
    layer0_outputs(8144) <= not (a or b);
    layer0_outputs(8145) <= a and b;
    layer0_outputs(8146) <= b and not a;
    layer0_outputs(8147) <= a and not b;
    layer0_outputs(8148) <= not a;
    layer0_outputs(8149) <= a;
    layer0_outputs(8150) <= a and not b;
    layer0_outputs(8151) <= 1'b0;
    layer0_outputs(8152) <= not (a xor b);
    layer0_outputs(8153) <= 1'b1;
    layer0_outputs(8154) <= b and not a;
    layer0_outputs(8155) <= 1'b0;
    layer0_outputs(8156) <= 1'b1;
    layer0_outputs(8157) <= b;
    layer0_outputs(8158) <= not b;
    layer0_outputs(8159) <= b;
    layer0_outputs(8160) <= b and not a;
    layer0_outputs(8161) <= a and not b;
    layer0_outputs(8162) <= not a;
    layer0_outputs(8163) <= 1'b1;
    layer0_outputs(8164) <= b;
    layer0_outputs(8165) <= not b;
    layer0_outputs(8166) <= b and not a;
    layer0_outputs(8167) <= a;
    layer0_outputs(8168) <= 1'b1;
    layer0_outputs(8169) <= not a or b;
    layer0_outputs(8170) <= a;
    layer0_outputs(8171) <= b;
    layer0_outputs(8172) <= a;
    layer0_outputs(8173) <= a or b;
    layer0_outputs(8174) <= 1'b0;
    layer0_outputs(8175) <= a and not b;
    layer0_outputs(8176) <= a and not b;
    layer0_outputs(8177) <= not b or a;
    layer0_outputs(8178) <= not b or a;
    layer0_outputs(8179) <= not (a or b);
    layer0_outputs(8180) <= not a or b;
    layer0_outputs(8181) <= not a;
    layer0_outputs(8182) <= 1'b1;
    layer0_outputs(8183) <= a or b;
    layer0_outputs(8184) <= 1'b1;
    layer0_outputs(8185) <= not a;
    layer0_outputs(8186) <= not b or a;
    layer0_outputs(8187) <= not (a xor b);
    layer0_outputs(8188) <= a xor b;
    layer0_outputs(8189) <= 1'b0;
    layer0_outputs(8190) <= 1'b0;
    layer0_outputs(8191) <= b;
    layer0_outputs(8192) <= a and b;
    layer0_outputs(8193) <= a;
    layer0_outputs(8194) <= not (a and b);
    layer0_outputs(8195) <= a;
    layer0_outputs(8196) <= a xor b;
    layer0_outputs(8197) <= not (a or b);
    layer0_outputs(8198) <= not (a and b);
    layer0_outputs(8199) <= 1'b0;
    layer0_outputs(8200) <= not (a and b);
    layer0_outputs(8201) <= 1'b1;
    layer0_outputs(8202) <= a and b;
    layer0_outputs(8203) <= a or b;
    layer0_outputs(8204) <= not (a or b);
    layer0_outputs(8205) <= 1'b0;
    layer0_outputs(8206) <= not (a or b);
    layer0_outputs(8207) <= a;
    layer0_outputs(8208) <= a xor b;
    layer0_outputs(8209) <= a xor b;
    layer0_outputs(8210) <= not a or b;
    layer0_outputs(8211) <= not b or a;
    layer0_outputs(8212) <= a xor b;
    layer0_outputs(8213) <= a and not b;
    layer0_outputs(8214) <= 1'b1;
    layer0_outputs(8215) <= a and not b;
    layer0_outputs(8216) <= not b;
    layer0_outputs(8217) <= not b or a;
    layer0_outputs(8218) <= not b;
    layer0_outputs(8219) <= not (a or b);
    layer0_outputs(8220) <= not (a and b);
    layer0_outputs(8221) <= not a;
    layer0_outputs(8222) <= a xor b;
    layer0_outputs(8223) <= a and not b;
    layer0_outputs(8224) <= a xor b;
    layer0_outputs(8225) <= not (a and b);
    layer0_outputs(8226) <= not a;
    layer0_outputs(8227) <= not b;
    layer0_outputs(8228) <= b;
    layer0_outputs(8229) <= not a or b;
    layer0_outputs(8230) <= not (a and b);
    layer0_outputs(8231) <= a or b;
    layer0_outputs(8232) <= not (a and b);
    layer0_outputs(8233) <= b and not a;
    layer0_outputs(8234) <= a and b;
    layer0_outputs(8235) <= not b or a;
    layer0_outputs(8236) <= not (a and b);
    layer0_outputs(8237) <= 1'b1;
    layer0_outputs(8238) <= a and b;
    layer0_outputs(8239) <= not a or b;
    layer0_outputs(8240) <= not a or b;
    layer0_outputs(8241) <= not (a and b);
    layer0_outputs(8242) <= not (a or b);
    layer0_outputs(8243) <= not a or b;
    layer0_outputs(8244) <= not (a xor b);
    layer0_outputs(8245) <= not (a and b);
    layer0_outputs(8246) <= a or b;
    layer0_outputs(8247) <= a;
    layer0_outputs(8248) <= 1'b1;
    layer0_outputs(8249) <= a and not b;
    layer0_outputs(8250) <= not a;
    layer0_outputs(8251) <= not a or b;
    layer0_outputs(8252) <= a or b;
    layer0_outputs(8253) <= not a;
    layer0_outputs(8254) <= not (a or b);
    layer0_outputs(8255) <= a or b;
    layer0_outputs(8256) <= not a;
    layer0_outputs(8257) <= not (a xor b);
    layer0_outputs(8258) <= not b;
    layer0_outputs(8259) <= a and not b;
    layer0_outputs(8260) <= a xor b;
    layer0_outputs(8261) <= not (a or b);
    layer0_outputs(8262) <= a;
    layer0_outputs(8263) <= b;
    layer0_outputs(8264) <= 1'b1;
    layer0_outputs(8265) <= not a;
    layer0_outputs(8266) <= a or b;
    layer0_outputs(8267) <= not a or b;
    layer0_outputs(8268) <= not (a and b);
    layer0_outputs(8269) <= a;
    layer0_outputs(8270) <= 1'b0;
    layer0_outputs(8271) <= not b or a;
    layer0_outputs(8272) <= not (a or b);
    layer0_outputs(8273) <= 1'b1;
    layer0_outputs(8274) <= b and not a;
    layer0_outputs(8275) <= 1'b0;
    layer0_outputs(8276) <= b;
    layer0_outputs(8277) <= not a;
    layer0_outputs(8278) <= a;
    layer0_outputs(8279) <= not (a xor b);
    layer0_outputs(8280) <= a and b;
    layer0_outputs(8281) <= a;
    layer0_outputs(8282) <= not a;
    layer0_outputs(8283) <= not b or a;
    layer0_outputs(8284) <= not b;
    layer0_outputs(8285) <= a xor b;
    layer0_outputs(8286) <= 1'b1;
    layer0_outputs(8287) <= a or b;
    layer0_outputs(8288) <= b and not a;
    layer0_outputs(8289) <= not (a and b);
    layer0_outputs(8290) <= not (a or b);
    layer0_outputs(8291) <= a;
    layer0_outputs(8292) <= not b or a;
    layer0_outputs(8293) <= 1'b1;
    layer0_outputs(8294) <= not a;
    layer0_outputs(8295) <= 1'b1;
    layer0_outputs(8296) <= not a or b;
    layer0_outputs(8297) <= b;
    layer0_outputs(8298) <= 1'b0;
    layer0_outputs(8299) <= not (a xor b);
    layer0_outputs(8300) <= b;
    layer0_outputs(8301) <= a or b;
    layer0_outputs(8302) <= a or b;
    layer0_outputs(8303) <= 1'b0;
    layer0_outputs(8304) <= not (a and b);
    layer0_outputs(8305) <= not (a and b);
    layer0_outputs(8306) <= not a or b;
    layer0_outputs(8307) <= b and not a;
    layer0_outputs(8308) <= a or b;
    layer0_outputs(8309) <= a and not b;
    layer0_outputs(8310) <= not (a or b);
    layer0_outputs(8311) <= not b;
    layer0_outputs(8312) <= not (a and b);
    layer0_outputs(8313) <= not b;
    layer0_outputs(8314) <= not (a and b);
    layer0_outputs(8315) <= not (a or b);
    layer0_outputs(8316) <= a and not b;
    layer0_outputs(8317) <= a and b;
    layer0_outputs(8318) <= not a;
    layer0_outputs(8319) <= a xor b;
    layer0_outputs(8320) <= 1'b0;
    layer0_outputs(8321) <= 1'b0;
    layer0_outputs(8322) <= 1'b0;
    layer0_outputs(8323) <= not b or a;
    layer0_outputs(8324) <= a;
    layer0_outputs(8325) <= a and not b;
    layer0_outputs(8326) <= a and b;
    layer0_outputs(8327) <= not (a xor b);
    layer0_outputs(8328) <= not (a and b);
    layer0_outputs(8329) <= a;
    layer0_outputs(8330) <= a and not b;
    layer0_outputs(8331) <= b;
    layer0_outputs(8332) <= not a or b;
    layer0_outputs(8333) <= not b;
    layer0_outputs(8334) <= 1'b0;
    layer0_outputs(8335) <= a;
    layer0_outputs(8336) <= not a;
    layer0_outputs(8337) <= b;
    layer0_outputs(8338) <= not a or b;
    layer0_outputs(8339) <= not a or b;
    layer0_outputs(8340) <= not (a xor b);
    layer0_outputs(8341) <= not b;
    layer0_outputs(8342) <= not (a xor b);
    layer0_outputs(8343) <= not (a and b);
    layer0_outputs(8344) <= a or b;
    layer0_outputs(8345) <= a and b;
    layer0_outputs(8346) <= b and not a;
    layer0_outputs(8347) <= 1'b1;
    layer0_outputs(8348) <= not b;
    layer0_outputs(8349) <= not a;
    layer0_outputs(8350) <= b and not a;
    layer0_outputs(8351) <= not b;
    layer0_outputs(8352) <= not (a and b);
    layer0_outputs(8353) <= a or b;
    layer0_outputs(8354) <= 1'b1;
    layer0_outputs(8355) <= 1'b0;
    layer0_outputs(8356) <= not b;
    layer0_outputs(8357) <= a and not b;
    layer0_outputs(8358) <= not a or b;
    layer0_outputs(8359) <= a and not b;
    layer0_outputs(8360) <= b and not a;
    layer0_outputs(8361) <= a and b;
    layer0_outputs(8362) <= a and not b;
    layer0_outputs(8363) <= not (a and b);
    layer0_outputs(8364) <= not (a and b);
    layer0_outputs(8365) <= not b;
    layer0_outputs(8366) <= b and not a;
    layer0_outputs(8367) <= a and not b;
    layer0_outputs(8368) <= not b or a;
    layer0_outputs(8369) <= a or b;
    layer0_outputs(8370) <= not a or b;
    layer0_outputs(8371) <= not b or a;
    layer0_outputs(8372) <= a or b;
    layer0_outputs(8373) <= not (a or b);
    layer0_outputs(8374) <= 1'b1;
    layer0_outputs(8375) <= not (a or b);
    layer0_outputs(8376) <= not b;
    layer0_outputs(8377) <= a xor b;
    layer0_outputs(8378) <= not a;
    layer0_outputs(8379) <= 1'b1;
    layer0_outputs(8380) <= 1'b1;
    layer0_outputs(8381) <= 1'b0;
    layer0_outputs(8382) <= 1'b0;
    layer0_outputs(8383) <= not (a and b);
    layer0_outputs(8384) <= a;
    layer0_outputs(8385) <= a and b;
    layer0_outputs(8386) <= not b;
    layer0_outputs(8387) <= a and b;
    layer0_outputs(8388) <= b;
    layer0_outputs(8389) <= not b;
    layer0_outputs(8390) <= a;
    layer0_outputs(8391) <= a xor b;
    layer0_outputs(8392) <= not (a xor b);
    layer0_outputs(8393) <= not a or b;
    layer0_outputs(8394) <= b;
    layer0_outputs(8395) <= a xor b;
    layer0_outputs(8396) <= not (a and b);
    layer0_outputs(8397) <= a or b;
    layer0_outputs(8398) <= a;
    layer0_outputs(8399) <= a and not b;
    layer0_outputs(8400) <= not (a xor b);
    layer0_outputs(8401) <= not (a xor b);
    layer0_outputs(8402) <= b and not a;
    layer0_outputs(8403) <= a and b;
    layer0_outputs(8404) <= not a or b;
    layer0_outputs(8405) <= 1'b0;
    layer0_outputs(8406) <= b and not a;
    layer0_outputs(8407) <= not (a xor b);
    layer0_outputs(8408) <= not a or b;
    layer0_outputs(8409) <= a and not b;
    layer0_outputs(8410) <= b;
    layer0_outputs(8411) <= 1'b1;
    layer0_outputs(8412) <= not (a and b);
    layer0_outputs(8413) <= b and not a;
    layer0_outputs(8414) <= not b or a;
    layer0_outputs(8415) <= not b;
    layer0_outputs(8416) <= not (a xor b);
    layer0_outputs(8417) <= 1'b1;
    layer0_outputs(8418) <= not (a and b);
    layer0_outputs(8419) <= a;
    layer0_outputs(8420) <= b and not a;
    layer0_outputs(8421) <= not (a or b);
    layer0_outputs(8422) <= not a or b;
    layer0_outputs(8423) <= 1'b0;
    layer0_outputs(8424) <= a xor b;
    layer0_outputs(8425) <= b and not a;
    layer0_outputs(8426) <= a;
    layer0_outputs(8427) <= b and not a;
    layer0_outputs(8428) <= a xor b;
    layer0_outputs(8429) <= not b or a;
    layer0_outputs(8430) <= a xor b;
    layer0_outputs(8431) <= a;
    layer0_outputs(8432) <= a;
    layer0_outputs(8433) <= b and not a;
    layer0_outputs(8434) <= not (a xor b);
    layer0_outputs(8435) <= not a;
    layer0_outputs(8436) <= 1'b1;
    layer0_outputs(8437) <= b and not a;
    layer0_outputs(8438) <= not b;
    layer0_outputs(8439) <= 1'b1;
    layer0_outputs(8440) <= not (a xor b);
    layer0_outputs(8441) <= a or b;
    layer0_outputs(8442) <= 1'b1;
    layer0_outputs(8443) <= a or b;
    layer0_outputs(8444) <= a and not b;
    layer0_outputs(8445) <= not (a and b);
    layer0_outputs(8446) <= 1'b1;
    layer0_outputs(8447) <= b;
    layer0_outputs(8448) <= 1'b0;
    layer0_outputs(8449) <= 1'b1;
    layer0_outputs(8450) <= b;
    layer0_outputs(8451) <= b and not a;
    layer0_outputs(8452) <= b;
    layer0_outputs(8453) <= b and not a;
    layer0_outputs(8454) <= not b or a;
    layer0_outputs(8455) <= not (a and b);
    layer0_outputs(8456) <= not b or a;
    layer0_outputs(8457) <= a and b;
    layer0_outputs(8458) <= b;
    layer0_outputs(8459) <= a and b;
    layer0_outputs(8460) <= not (a or b);
    layer0_outputs(8461) <= not a;
    layer0_outputs(8462) <= not (a and b);
    layer0_outputs(8463) <= not (a and b);
    layer0_outputs(8464) <= a or b;
    layer0_outputs(8465) <= b;
    layer0_outputs(8466) <= b;
    layer0_outputs(8467) <= a and b;
    layer0_outputs(8468) <= not a;
    layer0_outputs(8469) <= not a;
    layer0_outputs(8470) <= not (a and b);
    layer0_outputs(8471) <= not a or b;
    layer0_outputs(8472) <= a and b;
    layer0_outputs(8473) <= a or b;
    layer0_outputs(8474) <= a and b;
    layer0_outputs(8475) <= not (a and b);
    layer0_outputs(8476) <= a xor b;
    layer0_outputs(8477) <= b;
    layer0_outputs(8478) <= not (a or b);
    layer0_outputs(8479) <= not b or a;
    layer0_outputs(8480) <= 1'b0;
    layer0_outputs(8481) <= not (a xor b);
    layer0_outputs(8482) <= a and not b;
    layer0_outputs(8483) <= b;
    layer0_outputs(8484) <= not b;
    layer0_outputs(8485) <= a or b;
    layer0_outputs(8486) <= not a;
    layer0_outputs(8487) <= not (a or b);
    layer0_outputs(8488) <= not (a and b);
    layer0_outputs(8489) <= not (a and b);
    layer0_outputs(8490) <= not (a xor b);
    layer0_outputs(8491) <= a xor b;
    layer0_outputs(8492) <= 1'b0;
    layer0_outputs(8493) <= 1'b0;
    layer0_outputs(8494) <= b;
    layer0_outputs(8495) <= a;
    layer0_outputs(8496) <= not (a and b);
    layer0_outputs(8497) <= not a;
    layer0_outputs(8498) <= not b;
    layer0_outputs(8499) <= a and b;
    layer0_outputs(8500) <= not (a or b);
    layer0_outputs(8501) <= not b;
    layer0_outputs(8502) <= 1'b1;
    layer0_outputs(8503) <= a xor b;
    layer0_outputs(8504) <= b;
    layer0_outputs(8505) <= not (a xor b);
    layer0_outputs(8506) <= a and not b;
    layer0_outputs(8507) <= a xor b;
    layer0_outputs(8508) <= a;
    layer0_outputs(8509) <= not b;
    layer0_outputs(8510) <= a xor b;
    layer0_outputs(8511) <= not b;
    layer0_outputs(8512) <= a;
    layer0_outputs(8513) <= not (a or b);
    layer0_outputs(8514) <= not (a xor b);
    layer0_outputs(8515) <= 1'b1;
    layer0_outputs(8516) <= not a;
    layer0_outputs(8517) <= not (a or b);
    layer0_outputs(8518) <= 1'b0;
    layer0_outputs(8519) <= not (a and b);
    layer0_outputs(8520) <= not a or b;
    layer0_outputs(8521) <= not b;
    layer0_outputs(8522) <= a or b;
    layer0_outputs(8523) <= not b;
    layer0_outputs(8524) <= not b;
    layer0_outputs(8525) <= b;
    layer0_outputs(8526) <= a and b;
    layer0_outputs(8527) <= b and not a;
    layer0_outputs(8528) <= not (a and b);
    layer0_outputs(8529) <= a xor b;
    layer0_outputs(8530) <= not (a and b);
    layer0_outputs(8531) <= not (a xor b);
    layer0_outputs(8532) <= a;
    layer0_outputs(8533) <= not (a and b);
    layer0_outputs(8534) <= not b or a;
    layer0_outputs(8535) <= 1'b1;
    layer0_outputs(8536) <= a or b;
    layer0_outputs(8537) <= not b or a;
    layer0_outputs(8538) <= 1'b1;
    layer0_outputs(8539) <= not a;
    layer0_outputs(8540) <= a and not b;
    layer0_outputs(8541) <= not (a and b);
    layer0_outputs(8542) <= b;
    layer0_outputs(8543) <= a xor b;
    layer0_outputs(8544) <= not (a or b);
    layer0_outputs(8545) <= not (a or b);
    layer0_outputs(8546) <= a;
    layer0_outputs(8547) <= b and not a;
    layer0_outputs(8548) <= a;
    layer0_outputs(8549) <= not a;
    layer0_outputs(8550) <= not a;
    layer0_outputs(8551) <= a xor b;
    layer0_outputs(8552) <= not (a xor b);
    layer0_outputs(8553) <= b and not a;
    layer0_outputs(8554) <= not b;
    layer0_outputs(8555) <= not a;
    layer0_outputs(8556) <= 1'b1;
    layer0_outputs(8557) <= not a;
    layer0_outputs(8558) <= b and not a;
    layer0_outputs(8559) <= not b;
    layer0_outputs(8560) <= not (a or b);
    layer0_outputs(8561) <= 1'b1;
    layer0_outputs(8562) <= not (a or b);
    layer0_outputs(8563) <= a or b;
    layer0_outputs(8564) <= not (a and b);
    layer0_outputs(8565) <= not a or b;
    layer0_outputs(8566) <= not (a or b);
    layer0_outputs(8567) <= a;
    layer0_outputs(8568) <= not (a xor b);
    layer0_outputs(8569) <= not (a or b);
    layer0_outputs(8570) <= a or b;
    layer0_outputs(8571) <= a or b;
    layer0_outputs(8572) <= 1'b1;
    layer0_outputs(8573) <= b and not a;
    layer0_outputs(8574) <= not a;
    layer0_outputs(8575) <= not (a or b);
    layer0_outputs(8576) <= a;
    layer0_outputs(8577) <= not b;
    layer0_outputs(8578) <= a xor b;
    layer0_outputs(8579) <= 1'b0;
    layer0_outputs(8580) <= 1'b1;
    layer0_outputs(8581) <= not (a xor b);
    layer0_outputs(8582) <= a xor b;
    layer0_outputs(8583) <= a and b;
    layer0_outputs(8584) <= a and b;
    layer0_outputs(8585) <= a;
    layer0_outputs(8586) <= b and not a;
    layer0_outputs(8587) <= b;
    layer0_outputs(8588) <= a and b;
    layer0_outputs(8589) <= a and b;
    layer0_outputs(8590) <= a;
    layer0_outputs(8591) <= b and not a;
    layer0_outputs(8592) <= not a or b;
    layer0_outputs(8593) <= a or b;
    layer0_outputs(8594) <= a xor b;
    layer0_outputs(8595) <= 1'b0;
    layer0_outputs(8596) <= not a;
    layer0_outputs(8597) <= 1'b1;
    layer0_outputs(8598) <= a;
    layer0_outputs(8599) <= not b;
    layer0_outputs(8600) <= not (a xor b);
    layer0_outputs(8601) <= not b;
    layer0_outputs(8602) <= not b;
    layer0_outputs(8603) <= a and b;
    layer0_outputs(8604) <= 1'b1;
    layer0_outputs(8605) <= not (a and b);
    layer0_outputs(8606) <= not (a or b);
    layer0_outputs(8607) <= not (a and b);
    layer0_outputs(8608) <= not (a xor b);
    layer0_outputs(8609) <= not b;
    layer0_outputs(8610) <= b and not a;
    layer0_outputs(8611) <= a and b;
    layer0_outputs(8612) <= 1'b1;
    layer0_outputs(8613) <= not b or a;
    layer0_outputs(8614) <= not b or a;
    layer0_outputs(8615) <= a or b;
    layer0_outputs(8616) <= not a or b;
    layer0_outputs(8617) <= 1'b0;
    layer0_outputs(8618) <= not b;
    layer0_outputs(8619) <= not (a xor b);
    layer0_outputs(8620) <= a xor b;
    layer0_outputs(8621) <= 1'b0;
    layer0_outputs(8622) <= 1'b1;
    layer0_outputs(8623) <= 1'b1;
    layer0_outputs(8624) <= a;
    layer0_outputs(8625) <= b and not a;
    layer0_outputs(8626) <= b;
    layer0_outputs(8627) <= a and b;
    layer0_outputs(8628) <= a and b;
    layer0_outputs(8629) <= 1'b0;
    layer0_outputs(8630) <= a and b;
    layer0_outputs(8631) <= a and not b;
    layer0_outputs(8632) <= 1'b1;
    layer0_outputs(8633) <= not a or b;
    layer0_outputs(8634) <= not a;
    layer0_outputs(8635) <= 1'b1;
    layer0_outputs(8636) <= a or b;
    layer0_outputs(8637) <= not b;
    layer0_outputs(8638) <= b and not a;
    layer0_outputs(8639) <= b;
    layer0_outputs(8640) <= not a;
    layer0_outputs(8641) <= a or b;
    layer0_outputs(8642) <= 1'b0;
    layer0_outputs(8643) <= a or b;
    layer0_outputs(8644) <= not b;
    layer0_outputs(8645) <= not a;
    layer0_outputs(8646) <= not a;
    layer0_outputs(8647) <= a xor b;
    layer0_outputs(8648) <= a or b;
    layer0_outputs(8649) <= not (a or b);
    layer0_outputs(8650) <= not b;
    layer0_outputs(8651) <= 1'b1;
    layer0_outputs(8652) <= not (a or b);
    layer0_outputs(8653) <= not b;
    layer0_outputs(8654) <= 1'b0;
    layer0_outputs(8655) <= b;
    layer0_outputs(8656) <= not a or b;
    layer0_outputs(8657) <= a xor b;
    layer0_outputs(8658) <= not a or b;
    layer0_outputs(8659) <= 1'b1;
    layer0_outputs(8660) <= 1'b0;
    layer0_outputs(8661) <= not b;
    layer0_outputs(8662) <= a and not b;
    layer0_outputs(8663) <= a;
    layer0_outputs(8664) <= b and not a;
    layer0_outputs(8665) <= a or b;
    layer0_outputs(8666) <= a and b;
    layer0_outputs(8667) <= b;
    layer0_outputs(8668) <= b;
    layer0_outputs(8669) <= not (a and b);
    layer0_outputs(8670) <= not (a and b);
    layer0_outputs(8671) <= 1'b0;
    layer0_outputs(8672) <= a or b;
    layer0_outputs(8673) <= a or b;
    layer0_outputs(8674) <= 1'b1;
    layer0_outputs(8675) <= not a or b;
    layer0_outputs(8676) <= not b;
    layer0_outputs(8677) <= a and b;
    layer0_outputs(8678) <= not a or b;
    layer0_outputs(8679) <= not b;
    layer0_outputs(8680) <= a or b;
    layer0_outputs(8681) <= a and b;
    layer0_outputs(8682) <= a xor b;
    layer0_outputs(8683) <= not a or b;
    layer0_outputs(8684) <= not a or b;
    layer0_outputs(8685) <= a and b;
    layer0_outputs(8686) <= not a;
    layer0_outputs(8687) <= a or b;
    layer0_outputs(8688) <= not b or a;
    layer0_outputs(8689) <= not (a and b);
    layer0_outputs(8690) <= a and not b;
    layer0_outputs(8691) <= not (a or b);
    layer0_outputs(8692) <= 1'b1;
    layer0_outputs(8693) <= not (a and b);
    layer0_outputs(8694) <= 1'b0;
    layer0_outputs(8695) <= b;
    layer0_outputs(8696) <= not a or b;
    layer0_outputs(8697) <= a or b;
    layer0_outputs(8698) <= not a;
    layer0_outputs(8699) <= a and not b;
    layer0_outputs(8700) <= 1'b1;
    layer0_outputs(8701) <= not a;
    layer0_outputs(8702) <= not b;
    layer0_outputs(8703) <= not a;
    layer0_outputs(8704) <= not b;
    layer0_outputs(8705) <= not (a or b);
    layer0_outputs(8706) <= a and b;
    layer0_outputs(8707) <= a or b;
    layer0_outputs(8708) <= a and b;
    layer0_outputs(8709) <= b and not a;
    layer0_outputs(8710) <= not (a and b);
    layer0_outputs(8711) <= 1'b1;
    layer0_outputs(8712) <= b and not a;
    layer0_outputs(8713) <= 1'b1;
    layer0_outputs(8714) <= a;
    layer0_outputs(8715) <= not b;
    layer0_outputs(8716) <= b;
    layer0_outputs(8717) <= b;
    layer0_outputs(8718) <= not a;
    layer0_outputs(8719) <= a and b;
    layer0_outputs(8720) <= not b or a;
    layer0_outputs(8721) <= 1'b1;
    layer0_outputs(8722) <= 1'b0;
    layer0_outputs(8723) <= 1'b1;
    layer0_outputs(8724) <= not (a or b);
    layer0_outputs(8725) <= not a;
    layer0_outputs(8726) <= b;
    layer0_outputs(8727) <= a and b;
    layer0_outputs(8728) <= 1'b0;
    layer0_outputs(8729) <= a xor b;
    layer0_outputs(8730) <= not (a and b);
    layer0_outputs(8731) <= a;
    layer0_outputs(8732) <= a and not b;
    layer0_outputs(8733) <= not b;
    layer0_outputs(8734) <= not b;
    layer0_outputs(8735) <= not (a or b);
    layer0_outputs(8736) <= 1'b1;
    layer0_outputs(8737) <= not a;
    layer0_outputs(8738) <= not a or b;
    layer0_outputs(8739) <= not b;
    layer0_outputs(8740) <= a and b;
    layer0_outputs(8741) <= a and b;
    layer0_outputs(8742) <= not (a or b);
    layer0_outputs(8743) <= not (a xor b);
    layer0_outputs(8744) <= not b;
    layer0_outputs(8745) <= b and not a;
    layer0_outputs(8746) <= 1'b0;
    layer0_outputs(8747) <= a xor b;
    layer0_outputs(8748) <= not a;
    layer0_outputs(8749) <= not b;
    layer0_outputs(8750) <= not (a and b);
    layer0_outputs(8751) <= not b;
    layer0_outputs(8752) <= a xor b;
    layer0_outputs(8753) <= not (a or b);
    layer0_outputs(8754) <= a or b;
    layer0_outputs(8755) <= not (a and b);
    layer0_outputs(8756) <= a or b;
    layer0_outputs(8757) <= not (a xor b);
    layer0_outputs(8758) <= a and b;
    layer0_outputs(8759) <= not (a and b);
    layer0_outputs(8760) <= b;
    layer0_outputs(8761) <= not (a or b);
    layer0_outputs(8762) <= not (a and b);
    layer0_outputs(8763) <= a or b;
    layer0_outputs(8764) <= not (a or b);
    layer0_outputs(8765) <= 1'b1;
    layer0_outputs(8766) <= 1'b0;
    layer0_outputs(8767) <= a and b;
    layer0_outputs(8768) <= a and b;
    layer0_outputs(8769) <= b;
    layer0_outputs(8770) <= not a or b;
    layer0_outputs(8771) <= 1'b1;
    layer0_outputs(8772) <= not a or b;
    layer0_outputs(8773) <= a and not b;
    layer0_outputs(8774) <= not a;
    layer0_outputs(8775) <= not a or b;
    layer0_outputs(8776) <= a;
    layer0_outputs(8777) <= not a or b;
    layer0_outputs(8778) <= a or b;
    layer0_outputs(8779) <= a and not b;
    layer0_outputs(8780) <= not (a xor b);
    layer0_outputs(8781) <= not (a and b);
    layer0_outputs(8782) <= 1'b0;
    layer0_outputs(8783) <= not (a or b);
    layer0_outputs(8784) <= not b;
    layer0_outputs(8785) <= b;
    layer0_outputs(8786) <= a;
    layer0_outputs(8787) <= a xor b;
    layer0_outputs(8788) <= 1'b0;
    layer0_outputs(8789) <= a and not b;
    layer0_outputs(8790) <= 1'b0;
    layer0_outputs(8791) <= not (a and b);
    layer0_outputs(8792) <= a or b;
    layer0_outputs(8793) <= 1'b0;
    layer0_outputs(8794) <= not b;
    layer0_outputs(8795) <= not (a xor b);
    layer0_outputs(8796) <= 1'b1;
    layer0_outputs(8797) <= a and b;
    layer0_outputs(8798) <= b;
    layer0_outputs(8799) <= a;
    layer0_outputs(8800) <= b and not a;
    layer0_outputs(8801) <= a or b;
    layer0_outputs(8802) <= not a or b;
    layer0_outputs(8803) <= a or b;
    layer0_outputs(8804) <= b;
    layer0_outputs(8805) <= a and b;
    layer0_outputs(8806) <= b and not a;
    layer0_outputs(8807) <= a or b;
    layer0_outputs(8808) <= b and not a;
    layer0_outputs(8809) <= a and not b;
    layer0_outputs(8810) <= a;
    layer0_outputs(8811) <= not (a or b);
    layer0_outputs(8812) <= not (a xor b);
    layer0_outputs(8813) <= not a;
    layer0_outputs(8814) <= a xor b;
    layer0_outputs(8815) <= not (a or b);
    layer0_outputs(8816) <= a xor b;
    layer0_outputs(8817) <= 1'b0;
    layer0_outputs(8818) <= not (a and b);
    layer0_outputs(8819) <= not b;
    layer0_outputs(8820) <= not a;
    layer0_outputs(8821) <= a or b;
    layer0_outputs(8822) <= b and not a;
    layer0_outputs(8823) <= not b or a;
    layer0_outputs(8824) <= not b;
    layer0_outputs(8825) <= not (a xor b);
    layer0_outputs(8826) <= a;
    layer0_outputs(8827) <= b and not a;
    layer0_outputs(8828) <= a and not b;
    layer0_outputs(8829) <= not (a and b);
    layer0_outputs(8830) <= a and b;
    layer0_outputs(8831) <= b and not a;
    layer0_outputs(8832) <= a and not b;
    layer0_outputs(8833) <= b and not a;
    layer0_outputs(8834) <= not b or a;
    layer0_outputs(8835) <= not b;
    layer0_outputs(8836) <= not a;
    layer0_outputs(8837) <= not a or b;
    layer0_outputs(8838) <= not a or b;
    layer0_outputs(8839) <= a;
    layer0_outputs(8840) <= not a or b;
    layer0_outputs(8841) <= not a;
    layer0_outputs(8842) <= not a or b;
    layer0_outputs(8843) <= a and not b;
    layer0_outputs(8844) <= not a;
    layer0_outputs(8845) <= a xor b;
    layer0_outputs(8846) <= b and not a;
    layer0_outputs(8847) <= not a or b;
    layer0_outputs(8848) <= not b;
    layer0_outputs(8849) <= not a or b;
    layer0_outputs(8850) <= a xor b;
    layer0_outputs(8851) <= not a;
    layer0_outputs(8852) <= not b;
    layer0_outputs(8853) <= a;
    layer0_outputs(8854) <= not (a or b);
    layer0_outputs(8855) <= a;
    layer0_outputs(8856) <= b;
    layer0_outputs(8857) <= not a or b;
    layer0_outputs(8858) <= not (a and b);
    layer0_outputs(8859) <= not a;
    layer0_outputs(8860) <= not (a and b);
    layer0_outputs(8861) <= a xor b;
    layer0_outputs(8862) <= 1'b1;
    layer0_outputs(8863) <= b and not a;
    layer0_outputs(8864) <= not b or a;
    layer0_outputs(8865) <= a and b;
    layer0_outputs(8866) <= 1'b1;
    layer0_outputs(8867) <= b and not a;
    layer0_outputs(8868) <= not b or a;
    layer0_outputs(8869) <= not (a and b);
    layer0_outputs(8870) <= not b or a;
    layer0_outputs(8871) <= not b;
    layer0_outputs(8872) <= not (a or b);
    layer0_outputs(8873) <= a and not b;
    layer0_outputs(8874) <= not b;
    layer0_outputs(8875) <= b;
    layer0_outputs(8876) <= not a or b;
    layer0_outputs(8877) <= not (a xor b);
    layer0_outputs(8878) <= not a or b;
    layer0_outputs(8879) <= 1'b0;
    layer0_outputs(8880) <= not b or a;
    layer0_outputs(8881) <= not a or b;
    layer0_outputs(8882) <= not b;
    layer0_outputs(8883) <= a and not b;
    layer0_outputs(8884) <= not (a or b);
    layer0_outputs(8885) <= not a or b;
    layer0_outputs(8886) <= b and not a;
    layer0_outputs(8887) <= not a;
    layer0_outputs(8888) <= a and not b;
    layer0_outputs(8889) <= b and not a;
    layer0_outputs(8890) <= 1'b0;
    layer0_outputs(8891) <= b;
    layer0_outputs(8892) <= not (a or b);
    layer0_outputs(8893) <= b and not a;
    layer0_outputs(8894) <= not (a and b);
    layer0_outputs(8895) <= a and not b;
    layer0_outputs(8896) <= not b or a;
    layer0_outputs(8897) <= not (a or b);
    layer0_outputs(8898) <= not b;
    layer0_outputs(8899) <= 1'b1;
    layer0_outputs(8900) <= a;
    layer0_outputs(8901) <= not (a and b);
    layer0_outputs(8902) <= b;
    layer0_outputs(8903) <= a and not b;
    layer0_outputs(8904) <= not (a or b);
    layer0_outputs(8905) <= 1'b0;
    layer0_outputs(8906) <= not b;
    layer0_outputs(8907) <= b and not a;
    layer0_outputs(8908) <= a or b;
    layer0_outputs(8909) <= b;
    layer0_outputs(8910) <= not a;
    layer0_outputs(8911) <= not (a and b);
    layer0_outputs(8912) <= a or b;
    layer0_outputs(8913) <= a or b;
    layer0_outputs(8914) <= not a;
    layer0_outputs(8915) <= a;
    layer0_outputs(8916) <= a or b;
    layer0_outputs(8917) <= not (a xor b);
    layer0_outputs(8918) <= a or b;
    layer0_outputs(8919) <= a xor b;
    layer0_outputs(8920) <= 1'b1;
    layer0_outputs(8921) <= a and b;
    layer0_outputs(8922) <= b;
    layer0_outputs(8923) <= not (a xor b);
    layer0_outputs(8924) <= a and not b;
    layer0_outputs(8925) <= b and not a;
    layer0_outputs(8926) <= a and not b;
    layer0_outputs(8927) <= not (a xor b);
    layer0_outputs(8928) <= not a;
    layer0_outputs(8929) <= not (a and b);
    layer0_outputs(8930) <= 1'b0;
    layer0_outputs(8931) <= not b or a;
    layer0_outputs(8932) <= not a;
    layer0_outputs(8933) <= 1'b0;
    layer0_outputs(8934) <= a and b;
    layer0_outputs(8935) <= not (a or b);
    layer0_outputs(8936) <= 1'b0;
    layer0_outputs(8937) <= a or b;
    layer0_outputs(8938) <= not (a or b);
    layer0_outputs(8939) <= not a or b;
    layer0_outputs(8940) <= a xor b;
    layer0_outputs(8941) <= 1'b0;
    layer0_outputs(8942) <= not a or b;
    layer0_outputs(8943) <= a;
    layer0_outputs(8944) <= not a;
    layer0_outputs(8945) <= a;
    layer0_outputs(8946) <= a and not b;
    layer0_outputs(8947) <= a or b;
    layer0_outputs(8948) <= a or b;
    layer0_outputs(8949) <= not b or a;
    layer0_outputs(8950) <= b and not a;
    layer0_outputs(8951) <= b;
    layer0_outputs(8952) <= not b;
    layer0_outputs(8953) <= a or b;
    layer0_outputs(8954) <= not b;
    layer0_outputs(8955) <= not (a xor b);
    layer0_outputs(8956) <= not (a and b);
    layer0_outputs(8957) <= a and not b;
    layer0_outputs(8958) <= a;
    layer0_outputs(8959) <= not (a xor b);
    layer0_outputs(8960) <= a xor b;
    layer0_outputs(8961) <= 1'b1;
    layer0_outputs(8962) <= a and not b;
    layer0_outputs(8963) <= a xor b;
    layer0_outputs(8964) <= 1'b0;
    layer0_outputs(8965) <= b and not a;
    layer0_outputs(8966) <= a and not b;
    layer0_outputs(8967) <= not b;
    layer0_outputs(8968) <= a;
    layer0_outputs(8969) <= b;
    layer0_outputs(8970) <= a xor b;
    layer0_outputs(8971) <= a xor b;
    layer0_outputs(8972) <= b;
    layer0_outputs(8973) <= not (a or b);
    layer0_outputs(8974) <= 1'b1;
    layer0_outputs(8975) <= not b;
    layer0_outputs(8976) <= not b;
    layer0_outputs(8977) <= not b or a;
    layer0_outputs(8978) <= a and not b;
    layer0_outputs(8979) <= 1'b1;
    layer0_outputs(8980) <= a or b;
    layer0_outputs(8981) <= a and not b;
    layer0_outputs(8982) <= not (a and b);
    layer0_outputs(8983) <= not (a xor b);
    layer0_outputs(8984) <= not a;
    layer0_outputs(8985) <= a xor b;
    layer0_outputs(8986) <= a or b;
    layer0_outputs(8987) <= 1'b0;
    layer0_outputs(8988) <= 1'b1;
    layer0_outputs(8989) <= not (a and b);
    layer0_outputs(8990) <= a and b;
    layer0_outputs(8991) <= 1'b0;
    layer0_outputs(8992) <= b;
    layer0_outputs(8993) <= not (a xor b);
    layer0_outputs(8994) <= a;
    layer0_outputs(8995) <= 1'b1;
    layer0_outputs(8996) <= not a;
    layer0_outputs(8997) <= a;
    layer0_outputs(8998) <= 1'b1;
    layer0_outputs(8999) <= not a;
    layer0_outputs(9000) <= a and not b;
    layer0_outputs(9001) <= b and not a;
    layer0_outputs(9002) <= not (a xor b);
    layer0_outputs(9003) <= b;
    layer0_outputs(9004) <= 1'b0;
    layer0_outputs(9005) <= not a;
    layer0_outputs(9006) <= not b or a;
    layer0_outputs(9007) <= not (a xor b);
    layer0_outputs(9008) <= a and b;
    layer0_outputs(9009) <= a;
    layer0_outputs(9010) <= 1'b1;
    layer0_outputs(9011) <= not (a or b);
    layer0_outputs(9012) <= not b;
    layer0_outputs(9013) <= a;
    layer0_outputs(9014) <= not (a and b);
    layer0_outputs(9015) <= a or b;
    layer0_outputs(9016) <= not a or b;
    layer0_outputs(9017) <= 1'b0;
    layer0_outputs(9018) <= not a or b;
    layer0_outputs(9019) <= a or b;
    layer0_outputs(9020) <= not (a and b);
    layer0_outputs(9021) <= not a;
    layer0_outputs(9022) <= not (a and b);
    layer0_outputs(9023) <= not (a xor b);
    layer0_outputs(9024) <= not (a xor b);
    layer0_outputs(9025) <= not b or a;
    layer0_outputs(9026) <= a and b;
    layer0_outputs(9027) <= a;
    layer0_outputs(9028) <= a and b;
    layer0_outputs(9029) <= a or b;
    layer0_outputs(9030) <= b and not a;
    layer0_outputs(9031) <= a xor b;
    layer0_outputs(9032) <= b;
    layer0_outputs(9033) <= not (a or b);
    layer0_outputs(9034) <= a and b;
    layer0_outputs(9035) <= a;
    layer0_outputs(9036) <= a xor b;
    layer0_outputs(9037) <= b;
    layer0_outputs(9038) <= a or b;
    layer0_outputs(9039) <= not b;
    layer0_outputs(9040) <= 1'b0;
    layer0_outputs(9041) <= not b or a;
    layer0_outputs(9042) <= not a or b;
    layer0_outputs(9043) <= a and not b;
    layer0_outputs(9044) <= 1'b0;
    layer0_outputs(9045) <= not a;
    layer0_outputs(9046) <= not (a and b);
    layer0_outputs(9047) <= not b;
    layer0_outputs(9048) <= b;
    layer0_outputs(9049) <= a;
    layer0_outputs(9050) <= 1'b0;
    layer0_outputs(9051) <= not a;
    layer0_outputs(9052) <= not a or b;
    layer0_outputs(9053) <= not (a xor b);
    layer0_outputs(9054) <= a and not b;
    layer0_outputs(9055) <= 1'b0;
    layer0_outputs(9056) <= 1'b0;
    layer0_outputs(9057) <= 1'b1;
    layer0_outputs(9058) <= not a;
    layer0_outputs(9059) <= a xor b;
    layer0_outputs(9060) <= a or b;
    layer0_outputs(9061) <= not (a or b);
    layer0_outputs(9062) <= 1'b0;
    layer0_outputs(9063) <= 1'b0;
    layer0_outputs(9064) <= b;
    layer0_outputs(9065) <= a xor b;
    layer0_outputs(9066) <= a;
    layer0_outputs(9067) <= b and not a;
    layer0_outputs(9068) <= a and not b;
    layer0_outputs(9069) <= a;
    layer0_outputs(9070) <= not (a xor b);
    layer0_outputs(9071) <= a xor b;
    layer0_outputs(9072) <= not (a or b);
    layer0_outputs(9073) <= b and not a;
    layer0_outputs(9074) <= not a or b;
    layer0_outputs(9075) <= not (a and b);
    layer0_outputs(9076) <= a and not b;
    layer0_outputs(9077) <= not a;
    layer0_outputs(9078) <= not (a xor b);
    layer0_outputs(9079) <= not (a or b);
    layer0_outputs(9080) <= a and b;
    layer0_outputs(9081) <= a;
    layer0_outputs(9082) <= not a;
    layer0_outputs(9083) <= not a or b;
    layer0_outputs(9084) <= a and b;
    layer0_outputs(9085) <= b;
    layer0_outputs(9086) <= not b;
    layer0_outputs(9087) <= 1'b1;
    layer0_outputs(9088) <= not (a xor b);
    layer0_outputs(9089) <= not a or b;
    layer0_outputs(9090) <= not b;
    layer0_outputs(9091) <= not a;
    layer0_outputs(9092) <= a or b;
    layer0_outputs(9093) <= not a;
    layer0_outputs(9094) <= a;
    layer0_outputs(9095) <= a;
    layer0_outputs(9096) <= a or b;
    layer0_outputs(9097) <= not (a and b);
    layer0_outputs(9098) <= not b;
    layer0_outputs(9099) <= a and not b;
    layer0_outputs(9100) <= a and not b;
    layer0_outputs(9101) <= a and not b;
    layer0_outputs(9102) <= not b;
    layer0_outputs(9103) <= not a;
    layer0_outputs(9104) <= a and not b;
    layer0_outputs(9105) <= not (a or b);
    layer0_outputs(9106) <= not a;
    layer0_outputs(9107) <= 1'b0;
    layer0_outputs(9108) <= b;
    layer0_outputs(9109) <= a;
    layer0_outputs(9110) <= a xor b;
    layer0_outputs(9111) <= not (a or b);
    layer0_outputs(9112) <= 1'b0;
    layer0_outputs(9113) <= not b;
    layer0_outputs(9114) <= not a;
    layer0_outputs(9115) <= 1'b0;
    layer0_outputs(9116) <= a or b;
    layer0_outputs(9117) <= a xor b;
    layer0_outputs(9118) <= 1'b1;
    layer0_outputs(9119) <= 1'b0;
    layer0_outputs(9120) <= a and b;
    layer0_outputs(9121) <= not a or b;
    layer0_outputs(9122) <= 1'b0;
    layer0_outputs(9123) <= not b;
    layer0_outputs(9124) <= not b;
    layer0_outputs(9125) <= not (a or b);
    layer0_outputs(9126) <= a;
    layer0_outputs(9127) <= 1'b1;
    layer0_outputs(9128) <= a xor b;
    layer0_outputs(9129) <= a or b;
    layer0_outputs(9130) <= not a;
    layer0_outputs(9131) <= not (a or b);
    layer0_outputs(9132) <= a;
    layer0_outputs(9133) <= a and not b;
    layer0_outputs(9134) <= not (a and b);
    layer0_outputs(9135) <= not b or a;
    layer0_outputs(9136) <= not b or a;
    layer0_outputs(9137) <= a xor b;
    layer0_outputs(9138) <= not (a or b);
    layer0_outputs(9139) <= 1'b1;
    layer0_outputs(9140) <= a and b;
    layer0_outputs(9141) <= b;
    layer0_outputs(9142) <= not a;
    layer0_outputs(9143) <= a xor b;
    layer0_outputs(9144) <= 1'b0;
    layer0_outputs(9145) <= not (a and b);
    layer0_outputs(9146) <= a or b;
    layer0_outputs(9147) <= a;
    layer0_outputs(9148) <= 1'b0;
    layer0_outputs(9149) <= not b;
    layer0_outputs(9150) <= a xor b;
    layer0_outputs(9151) <= a or b;
    layer0_outputs(9152) <= not b or a;
    layer0_outputs(9153) <= b;
    layer0_outputs(9154) <= not (a and b);
    layer0_outputs(9155) <= a and not b;
    layer0_outputs(9156) <= 1'b0;
    layer0_outputs(9157) <= b;
    layer0_outputs(9158) <= not (a or b);
    layer0_outputs(9159) <= not (a xor b);
    layer0_outputs(9160) <= not b;
    layer0_outputs(9161) <= a or b;
    layer0_outputs(9162) <= not b;
    layer0_outputs(9163) <= a or b;
    layer0_outputs(9164) <= a and not b;
    layer0_outputs(9165) <= b;
    layer0_outputs(9166) <= 1'b1;
    layer0_outputs(9167) <= 1'b0;
    layer0_outputs(9168) <= not b or a;
    layer0_outputs(9169) <= not a or b;
    layer0_outputs(9170) <= a and b;
    layer0_outputs(9171) <= 1'b0;
    layer0_outputs(9172) <= not b;
    layer0_outputs(9173) <= b and not a;
    layer0_outputs(9174) <= not b;
    layer0_outputs(9175) <= 1'b0;
    layer0_outputs(9176) <= a and not b;
    layer0_outputs(9177) <= not b;
    layer0_outputs(9178) <= a;
    layer0_outputs(9179) <= not b or a;
    layer0_outputs(9180) <= a and not b;
    layer0_outputs(9181) <= a;
    layer0_outputs(9182) <= a;
    layer0_outputs(9183) <= not a or b;
    layer0_outputs(9184) <= not a or b;
    layer0_outputs(9185) <= b and not a;
    layer0_outputs(9186) <= a;
    layer0_outputs(9187) <= a;
    layer0_outputs(9188) <= 1'b1;
    layer0_outputs(9189) <= not b or a;
    layer0_outputs(9190) <= b;
    layer0_outputs(9191) <= 1'b0;
    layer0_outputs(9192) <= a and b;
    layer0_outputs(9193) <= a;
    layer0_outputs(9194) <= a and not b;
    layer0_outputs(9195) <= not a or b;
    layer0_outputs(9196) <= a and b;
    layer0_outputs(9197) <= not (a xor b);
    layer0_outputs(9198) <= not a;
    layer0_outputs(9199) <= b;
    layer0_outputs(9200) <= a and not b;
    layer0_outputs(9201) <= not a or b;
    layer0_outputs(9202) <= a xor b;
    layer0_outputs(9203) <= 1'b1;
    layer0_outputs(9204) <= b;
    layer0_outputs(9205) <= 1'b1;
    layer0_outputs(9206) <= not b or a;
    layer0_outputs(9207) <= a and not b;
    layer0_outputs(9208) <= not b;
    layer0_outputs(9209) <= not (a and b);
    layer0_outputs(9210) <= not b or a;
    layer0_outputs(9211) <= b and not a;
    layer0_outputs(9212) <= a and not b;
    layer0_outputs(9213) <= not a or b;
    layer0_outputs(9214) <= b;
    layer0_outputs(9215) <= b and not a;
    layer0_outputs(9216) <= a xor b;
    layer0_outputs(9217) <= not a;
    layer0_outputs(9218) <= not (a or b);
    layer0_outputs(9219) <= a and b;
    layer0_outputs(9220) <= not a or b;
    layer0_outputs(9221) <= a or b;
    layer0_outputs(9222) <= a;
    layer0_outputs(9223) <= a;
    layer0_outputs(9224) <= not b or a;
    layer0_outputs(9225) <= not (a xor b);
    layer0_outputs(9226) <= not (a xor b);
    layer0_outputs(9227) <= b;
    layer0_outputs(9228) <= 1'b0;
    layer0_outputs(9229) <= not b or a;
    layer0_outputs(9230) <= not (a and b);
    layer0_outputs(9231) <= 1'b1;
    layer0_outputs(9232) <= not (a and b);
    layer0_outputs(9233) <= b;
    layer0_outputs(9234) <= a;
    layer0_outputs(9235) <= b;
    layer0_outputs(9236) <= not b;
    layer0_outputs(9237) <= 1'b1;
    layer0_outputs(9238) <= a;
    layer0_outputs(9239) <= not a or b;
    layer0_outputs(9240) <= b;
    layer0_outputs(9241) <= a or b;
    layer0_outputs(9242) <= a or b;
    layer0_outputs(9243) <= a or b;
    layer0_outputs(9244) <= not (a and b);
    layer0_outputs(9245) <= not (a or b);
    layer0_outputs(9246) <= b and not a;
    layer0_outputs(9247) <= not (a and b);
    layer0_outputs(9248) <= a xor b;
    layer0_outputs(9249) <= 1'b0;
    layer0_outputs(9250) <= b and not a;
    layer0_outputs(9251) <= 1'b1;
    layer0_outputs(9252) <= a and b;
    layer0_outputs(9253) <= a and b;
    layer0_outputs(9254) <= not (a xor b);
    layer0_outputs(9255) <= not (a and b);
    layer0_outputs(9256) <= not (a or b);
    layer0_outputs(9257) <= 1'b1;
    layer0_outputs(9258) <= a or b;
    layer0_outputs(9259) <= b;
    layer0_outputs(9260) <= not (a and b);
    layer0_outputs(9261) <= b and not a;
    layer0_outputs(9262) <= not (a or b);
    layer0_outputs(9263) <= not a;
    layer0_outputs(9264) <= 1'b0;
    layer0_outputs(9265) <= a xor b;
    layer0_outputs(9266) <= not b or a;
    layer0_outputs(9267) <= b;
    layer0_outputs(9268) <= not a;
    layer0_outputs(9269) <= b and not a;
    layer0_outputs(9270) <= not (a or b);
    layer0_outputs(9271) <= not a;
    layer0_outputs(9272) <= 1'b0;
    layer0_outputs(9273) <= a or b;
    layer0_outputs(9274) <= a xor b;
    layer0_outputs(9275) <= not b;
    layer0_outputs(9276) <= not a;
    layer0_outputs(9277) <= not (a and b);
    layer0_outputs(9278) <= a and not b;
    layer0_outputs(9279) <= b;
    layer0_outputs(9280) <= b;
    layer0_outputs(9281) <= not (a or b);
    layer0_outputs(9282) <= 1'b1;
    layer0_outputs(9283) <= a;
    layer0_outputs(9284) <= not a;
    layer0_outputs(9285) <= a;
    layer0_outputs(9286) <= 1'b0;
    layer0_outputs(9287) <= not a or b;
    layer0_outputs(9288) <= a xor b;
    layer0_outputs(9289) <= not b or a;
    layer0_outputs(9290) <= 1'b1;
    layer0_outputs(9291) <= a and b;
    layer0_outputs(9292) <= 1'b0;
    layer0_outputs(9293) <= not (a xor b);
    layer0_outputs(9294) <= a or b;
    layer0_outputs(9295) <= a and not b;
    layer0_outputs(9296) <= 1'b1;
    layer0_outputs(9297) <= a and not b;
    layer0_outputs(9298) <= not (a or b);
    layer0_outputs(9299) <= b and not a;
    layer0_outputs(9300) <= not a;
    layer0_outputs(9301) <= not (a or b);
    layer0_outputs(9302) <= a and b;
    layer0_outputs(9303) <= not a or b;
    layer0_outputs(9304) <= a or b;
    layer0_outputs(9305) <= 1'b0;
    layer0_outputs(9306) <= not (a xor b);
    layer0_outputs(9307) <= a and b;
    layer0_outputs(9308) <= not a or b;
    layer0_outputs(9309) <= a and not b;
    layer0_outputs(9310) <= not (a xor b);
    layer0_outputs(9311) <= b and not a;
    layer0_outputs(9312) <= b and not a;
    layer0_outputs(9313) <= b;
    layer0_outputs(9314) <= a;
    layer0_outputs(9315) <= not (a and b);
    layer0_outputs(9316) <= not b or a;
    layer0_outputs(9317) <= b and not a;
    layer0_outputs(9318) <= a and not b;
    layer0_outputs(9319) <= a;
    layer0_outputs(9320) <= a and not b;
    layer0_outputs(9321) <= a;
    layer0_outputs(9322) <= a xor b;
    layer0_outputs(9323) <= a and not b;
    layer0_outputs(9324) <= 1'b0;
    layer0_outputs(9325) <= not b;
    layer0_outputs(9326) <= not (a xor b);
    layer0_outputs(9327) <= not b or a;
    layer0_outputs(9328) <= not b or a;
    layer0_outputs(9329) <= b;
    layer0_outputs(9330) <= a or b;
    layer0_outputs(9331) <= a and not b;
    layer0_outputs(9332) <= not b;
    layer0_outputs(9333) <= 1'b1;
    layer0_outputs(9334) <= a or b;
    layer0_outputs(9335) <= a or b;
    layer0_outputs(9336) <= a;
    layer0_outputs(9337) <= a and not b;
    layer0_outputs(9338) <= a and b;
    layer0_outputs(9339) <= not (a and b);
    layer0_outputs(9340) <= not a;
    layer0_outputs(9341) <= not (a and b);
    layer0_outputs(9342) <= a;
    layer0_outputs(9343) <= not b;
    layer0_outputs(9344) <= not b or a;
    layer0_outputs(9345) <= b;
    layer0_outputs(9346) <= not (a or b);
    layer0_outputs(9347) <= a;
    layer0_outputs(9348) <= not (a xor b);
    layer0_outputs(9349) <= not (a and b);
    layer0_outputs(9350) <= not b;
    layer0_outputs(9351) <= a or b;
    layer0_outputs(9352) <= not (a or b);
    layer0_outputs(9353) <= not b or a;
    layer0_outputs(9354) <= b;
    layer0_outputs(9355) <= not a;
    layer0_outputs(9356) <= 1'b0;
    layer0_outputs(9357) <= a and b;
    layer0_outputs(9358) <= 1'b1;
    layer0_outputs(9359) <= not b or a;
    layer0_outputs(9360) <= a or b;
    layer0_outputs(9361) <= b and not a;
    layer0_outputs(9362) <= not b or a;
    layer0_outputs(9363) <= a and b;
    layer0_outputs(9364) <= not a or b;
    layer0_outputs(9365) <= 1'b1;
    layer0_outputs(9366) <= not a or b;
    layer0_outputs(9367) <= not a;
    layer0_outputs(9368) <= not (a and b);
    layer0_outputs(9369) <= not a or b;
    layer0_outputs(9370) <= a and b;
    layer0_outputs(9371) <= a xor b;
    layer0_outputs(9372) <= b;
    layer0_outputs(9373) <= not (a or b);
    layer0_outputs(9374) <= b and not a;
    layer0_outputs(9375) <= a or b;
    layer0_outputs(9376) <= not a;
    layer0_outputs(9377) <= not (a and b);
    layer0_outputs(9378) <= not (a and b);
    layer0_outputs(9379) <= a xor b;
    layer0_outputs(9380) <= not (a or b);
    layer0_outputs(9381) <= 1'b0;
    layer0_outputs(9382) <= not b;
    layer0_outputs(9383) <= a;
    layer0_outputs(9384) <= not (a and b);
    layer0_outputs(9385) <= not (a or b);
    layer0_outputs(9386) <= a and not b;
    layer0_outputs(9387) <= not a;
    layer0_outputs(9388) <= not a;
    layer0_outputs(9389) <= a;
    layer0_outputs(9390) <= not (a xor b);
    layer0_outputs(9391) <= b;
    layer0_outputs(9392) <= a or b;
    layer0_outputs(9393) <= not a or b;
    layer0_outputs(9394) <= not (a and b);
    layer0_outputs(9395) <= a xor b;
    layer0_outputs(9396) <= b and not a;
    layer0_outputs(9397) <= not b or a;
    layer0_outputs(9398) <= a or b;
    layer0_outputs(9399) <= a and not b;
    layer0_outputs(9400) <= 1'b1;
    layer0_outputs(9401) <= not (a xor b);
    layer0_outputs(9402) <= a or b;
    layer0_outputs(9403) <= not (a xor b);
    layer0_outputs(9404) <= a;
    layer0_outputs(9405) <= b and not a;
    layer0_outputs(9406) <= b;
    layer0_outputs(9407) <= not a;
    layer0_outputs(9408) <= b;
    layer0_outputs(9409) <= b and not a;
    layer0_outputs(9410) <= not b;
    layer0_outputs(9411) <= a and b;
    layer0_outputs(9412) <= a and b;
    layer0_outputs(9413) <= b;
    layer0_outputs(9414) <= b;
    layer0_outputs(9415) <= not a;
    layer0_outputs(9416) <= a xor b;
    layer0_outputs(9417) <= b;
    layer0_outputs(9418) <= not a or b;
    layer0_outputs(9419) <= a and not b;
    layer0_outputs(9420) <= b;
    layer0_outputs(9421) <= not (a or b);
    layer0_outputs(9422) <= not b;
    layer0_outputs(9423) <= b and not a;
    layer0_outputs(9424) <= not b;
    layer0_outputs(9425) <= not a or b;
    layer0_outputs(9426) <= a and not b;
    layer0_outputs(9427) <= not (a and b);
    layer0_outputs(9428) <= not b;
    layer0_outputs(9429) <= not b;
    layer0_outputs(9430) <= a;
    layer0_outputs(9431) <= a and not b;
    layer0_outputs(9432) <= 1'b1;
    layer0_outputs(9433) <= not (a xor b);
    layer0_outputs(9434) <= 1'b1;
    layer0_outputs(9435) <= not b;
    layer0_outputs(9436) <= 1'b1;
    layer0_outputs(9437) <= b and not a;
    layer0_outputs(9438) <= a and not b;
    layer0_outputs(9439) <= not (a xor b);
    layer0_outputs(9440) <= b;
    layer0_outputs(9441) <= not a;
    layer0_outputs(9442) <= a and b;
    layer0_outputs(9443) <= not (a xor b);
    layer0_outputs(9444) <= not a;
    layer0_outputs(9445) <= not (a xor b);
    layer0_outputs(9446) <= not a;
    layer0_outputs(9447) <= not b or a;
    layer0_outputs(9448) <= a xor b;
    layer0_outputs(9449) <= not a or b;
    layer0_outputs(9450) <= a and b;
    layer0_outputs(9451) <= 1'b1;
    layer0_outputs(9452) <= not a or b;
    layer0_outputs(9453) <= 1'b1;
    layer0_outputs(9454) <= a or b;
    layer0_outputs(9455) <= a;
    layer0_outputs(9456) <= b;
    layer0_outputs(9457) <= a and b;
    layer0_outputs(9458) <= a and b;
    layer0_outputs(9459) <= a and b;
    layer0_outputs(9460) <= a xor b;
    layer0_outputs(9461) <= not (a and b);
    layer0_outputs(9462) <= not (a and b);
    layer0_outputs(9463) <= not a;
    layer0_outputs(9464) <= a;
    layer0_outputs(9465) <= not (a and b);
    layer0_outputs(9466) <= not a;
    layer0_outputs(9467) <= not a;
    layer0_outputs(9468) <= a;
    layer0_outputs(9469) <= 1'b0;
    layer0_outputs(9470) <= not (a or b);
    layer0_outputs(9471) <= 1'b0;
    layer0_outputs(9472) <= a and not b;
    layer0_outputs(9473) <= not a;
    layer0_outputs(9474) <= b;
    layer0_outputs(9475) <= b and not a;
    layer0_outputs(9476) <= not (a or b);
    layer0_outputs(9477) <= not (a and b);
    layer0_outputs(9478) <= b and not a;
    layer0_outputs(9479) <= 1'b0;
    layer0_outputs(9480) <= b and not a;
    layer0_outputs(9481) <= a and not b;
    layer0_outputs(9482) <= b;
    layer0_outputs(9483) <= a and not b;
    layer0_outputs(9484) <= b and not a;
    layer0_outputs(9485) <= not (a and b);
    layer0_outputs(9486) <= a and b;
    layer0_outputs(9487) <= not (a xor b);
    layer0_outputs(9488) <= a;
    layer0_outputs(9489) <= a and not b;
    layer0_outputs(9490) <= a and b;
    layer0_outputs(9491) <= 1'b0;
    layer0_outputs(9492) <= a xor b;
    layer0_outputs(9493) <= b;
    layer0_outputs(9494) <= a xor b;
    layer0_outputs(9495) <= b and not a;
    layer0_outputs(9496) <= a or b;
    layer0_outputs(9497) <= b and not a;
    layer0_outputs(9498) <= not (a and b);
    layer0_outputs(9499) <= b;
    layer0_outputs(9500) <= 1'b1;
    layer0_outputs(9501) <= 1'b0;
    layer0_outputs(9502) <= not (a or b);
    layer0_outputs(9503) <= a and b;
    layer0_outputs(9504) <= 1'b1;
    layer0_outputs(9505) <= not (a or b);
    layer0_outputs(9506) <= not b or a;
    layer0_outputs(9507) <= not b;
    layer0_outputs(9508) <= a and b;
    layer0_outputs(9509) <= a and b;
    layer0_outputs(9510) <= not (a xor b);
    layer0_outputs(9511) <= a and not b;
    layer0_outputs(9512) <= a and not b;
    layer0_outputs(9513) <= not (a or b);
    layer0_outputs(9514) <= not (a and b);
    layer0_outputs(9515) <= not b;
    layer0_outputs(9516) <= a xor b;
    layer0_outputs(9517) <= not b;
    layer0_outputs(9518) <= not a or b;
    layer0_outputs(9519) <= b;
    layer0_outputs(9520) <= 1'b1;
    layer0_outputs(9521) <= not b or a;
    layer0_outputs(9522) <= not a;
    layer0_outputs(9523) <= a or b;
    layer0_outputs(9524) <= b and not a;
    layer0_outputs(9525) <= not b;
    layer0_outputs(9526) <= 1'b0;
    layer0_outputs(9527) <= not b or a;
    layer0_outputs(9528) <= 1'b0;
    layer0_outputs(9529) <= b;
    layer0_outputs(9530) <= b;
    layer0_outputs(9531) <= not (a and b);
    layer0_outputs(9532) <= not (a or b);
    layer0_outputs(9533) <= a;
    layer0_outputs(9534) <= not a;
    layer0_outputs(9535) <= a xor b;
    layer0_outputs(9536) <= a and b;
    layer0_outputs(9537) <= a and not b;
    layer0_outputs(9538) <= 1'b1;
    layer0_outputs(9539) <= b;
    layer0_outputs(9540) <= a and not b;
    layer0_outputs(9541) <= not (a xor b);
    layer0_outputs(9542) <= not a or b;
    layer0_outputs(9543) <= not a or b;
    layer0_outputs(9544) <= a and not b;
    layer0_outputs(9545) <= 1'b1;
    layer0_outputs(9546) <= b;
    layer0_outputs(9547) <= b;
    layer0_outputs(9548) <= not b;
    layer0_outputs(9549) <= not (a or b);
    layer0_outputs(9550) <= a and b;
    layer0_outputs(9551) <= 1'b0;
    layer0_outputs(9552) <= 1'b1;
    layer0_outputs(9553) <= not b;
    layer0_outputs(9554) <= not (a xor b);
    layer0_outputs(9555) <= 1'b0;
    layer0_outputs(9556) <= not b;
    layer0_outputs(9557) <= not (a or b);
    layer0_outputs(9558) <= a and not b;
    layer0_outputs(9559) <= a xor b;
    layer0_outputs(9560) <= 1'b1;
    layer0_outputs(9561) <= not a;
    layer0_outputs(9562) <= a xor b;
    layer0_outputs(9563) <= 1'b1;
    layer0_outputs(9564) <= b;
    layer0_outputs(9565) <= a xor b;
    layer0_outputs(9566) <= a xor b;
    layer0_outputs(9567) <= b and not a;
    layer0_outputs(9568) <= a and b;
    layer0_outputs(9569) <= not a;
    layer0_outputs(9570) <= a;
    layer0_outputs(9571) <= not (a and b);
    layer0_outputs(9572) <= not (a or b);
    layer0_outputs(9573) <= a or b;
    layer0_outputs(9574) <= not a;
    layer0_outputs(9575) <= a and b;
    layer0_outputs(9576) <= not (a or b);
    layer0_outputs(9577) <= not b;
    layer0_outputs(9578) <= not b;
    layer0_outputs(9579) <= not (a xor b);
    layer0_outputs(9580) <= not a or b;
    layer0_outputs(9581) <= b;
    layer0_outputs(9582) <= b and not a;
    layer0_outputs(9583) <= not (a and b);
    layer0_outputs(9584) <= b;
    layer0_outputs(9585) <= not a or b;
    layer0_outputs(9586) <= not (a xor b);
    layer0_outputs(9587) <= not (a xor b);
    layer0_outputs(9588) <= b and not a;
    layer0_outputs(9589) <= 1'b1;
    layer0_outputs(9590) <= a and b;
    layer0_outputs(9591) <= not a or b;
    layer0_outputs(9592) <= b and not a;
    layer0_outputs(9593) <= not (a and b);
    layer0_outputs(9594) <= not a;
    layer0_outputs(9595) <= a;
    layer0_outputs(9596) <= not (a or b);
    layer0_outputs(9597) <= not (a and b);
    layer0_outputs(9598) <= a and b;
    layer0_outputs(9599) <= not b;
    layer0_outputs(9600) <= not (a and b);
    layer0_outputs(9601) <= a or b;
    layer0_outputs(9602) <= not b or a;
    layer0_outputs(9603) <= not a;
    layer0_outputs(9604) <= not (a xor b);
    layer0_outputs(9605) <= not a;
    layer0_outputs(9606) <= not (a or b);
    layer0_outputs(9607) <= a and b;
    layer0_outputs(9608) <= not (a or b);
    layer0_outputs(9609) <= 1'b0;
    layer0_outputs(9610) <= a xor b;
    layer0_outputs(9611) <= 1'b1;
    layer0_outputs(9612) <= not a;
    layer0_outputs(9613) <= 1'b1;
    layer0_outputs(9614) <= a or b;
    layer0_outputs(9615) <= not (a xor b);
    layer0_outputs(9616) <= a or b;
    layer0_outputs(9617) <= not a or b;
    layer0_outputs(9618) <= not b or a;
    layer0_outputs(9619) <= a;
    layer0_outputs(9620) <= not a;
    layer0_outputs(9621) <= not b or a;
    layer0_outputs(9622) <= a and not b;
    layer0_outputs(9623) <= b and not a;
    layer0_outputs(9624) <= a xor b;
    layer0_outputs(9625) <= not (a or b);
    layer0_outputs(9626) <= not b;
    layer0_outputs(9627) <= 1'b1;
    layer0_outputs(9628) <= 1'b1;
    layer0_outputs(9629) <= b and not a;
    layer0_outputs(9630) <= a or b;
    layer0_outputs(9631) <= 1'b0;
    layer0_outputs(9632) <= a xor b;
    layer0_outputs(9633) <= not (a and b);
    layer0_outputs(9634) <= a or b;
    layer0_outputs(9635) <= a xor b;
    layer0_outputs(9636) <= a;
    layer0_outputs(9637) <= not b;
    layer0_outputs(9638) <= 1'b0;
    layer0_outputs(9639) <= not (a or b);
    layer0_outputs(9640) <= a and b;
    layer0_outputs(9641) <= a or b;
    layer0_outputs(9642) <= not b or a;
    layer0_outputs(9643) <= not (a or b);
    layer0_outputs(9644) <= 1'b0;
    layer0_outputs(9645) <= 1'b1;
    layer0_outputs(9646) <= not b or a;
    layer0_outputs(9647) <= b and not a;
    layer0_outputs(9648) <= 1'b1;
    layer0_outputs(9649) <= b;
    layer0_outputs(9650) <= not (a and b);
    layer0_outputs(9651) <= b;
    layer0_outputs(9652) <= not (a xor b);
    layer0_outputs(9653) <= a and b;
    layer0_outputs(9654) <= not (a and b);
    layer0_outputs(9655) <= 1'b1;
    layer0_outputs(9656) <= a or b;
    layer0_outputs(9657) <= not (a and b);
    layer0_outputs(9658) <= b;
    layer0_outputs(9659) <= not a;
    layer0_outputs(9660) <= a xor b;
    layer0_outputs(9661) <= not (a or b);
    layer0_outputs(9662) <= 1'b1;
    layer0_outputs(9663) <= not b;
    layer0_outputs(9664) <= not (a and b);
    layer0_outputs(9665) <= 1'b1;
    layer0_outputs(9666) <= 1'b0;
    layer0_outputs(9667) <= a;
    layer0_outputs(9668) <= b and not a;
    layer0_outputs(9669) <= not b;
    layer0_outputs(9670) <= not (a xor b);
    layer0_outputs(9671) <= not a;
    layer0_outputs(9672) <= not (a xor b);
    layer0_outputs(9673) <= not b;
    layer0_outputs(9674) <= b;
    layer0_outputs(9675) <= not (a or b);
    layer0_outputs(9676) <= not (a and b);
    layer0_outputs(9677) <= not a;
    layer0_outputs(9678) <= a and b;
    layer0_outputs(9679) <= not (a and b);
    layer0_outputs(9680) <= not b;
    layer0_outputs(9681) <= not (a xor b);
    layer0_outputs(9682) <= not b or a;
    layer0_outputs(9683) <= b;
    layer0_outputs(9684) <= 1'b1;
    layer0_outputs(9685) <= a or b;
    layer0_outputs(9686) <= not a;
    layer0_outputs(9687) <= not a;
    layer0_outputs(9688) <= b;
    layer0_outputs(9689) <= a and not b;
    layer0_outputs(9690) <= not b;
    layer0_outputs(9691) <= not a;
    layer0_outputs(9692) <= not (a and b);
    layer0_outputs(9693) <= not b;
    layer0_outputs(9694) <= not (a xor b);
    layer0_outputs(9695) <= not (a or b);
    layer0_outputs(9696) <= not b;
    layer0_outputs(9697) <= a and b;
    layer0_outputs(9698) <= not a or b;
    layer0_outputs(9699) <= not (a or b);
    layer0_outputs(9700) <= not (a xor b);
    layer0_outputs(9701) <= b;
    layer0_outputs(9702) <= 1'b0;
    layer0_outputs(9703) <= 1'b0;
    layer0_outputs(9704) <= not (a and b);
    layer0_outputs(9705) <= not (a or b);
    layer0_outputs(9706) <= not (a or b);
    layer0_outputs(9707) <= a and not b;
    layer0_outputs(9708) <= not (a and b);
    layer0_outputs(9709) <= not (a xor b);
    layer0_outputs(9710) <= a and not b;
    layer0_outputs(9711) <= not (a xor b);
    layer0_outputs(9712) <= not (a xor b);
    layer0_outputs(9713) <= b;
    layer0_outputs(9714) <= not (a or b);
    layer0_outputs(9715) <= a or b;
    layer0_outputs(9716) <= b and not a;
    layer0_outputs(9717) <= a or b;
    layer0_outputs(9718) <= not b or a;
    layer0_outputs(9719) <= b;
    layer0_outputs(9720) <= 1'b1;
    layer0_outputs(9721) <= a or b;
    layer0_outputs(9722) <= 1'b0;
    layer0_outputs(9723) <= not a;
    layer0_outputs(9724) <= not b;
    layer0_outputs(9725) <= not b;
    layer0_outputs(9726) <= a xor b;
    layer0_outputs(9727) <= a and b;
    layer0_outputs(9728) <= a xor b;
    layer0_outputs(9729) <= not a or b;
    layer0_outputs(9730) <= not a or b;
    layer0_outputs(9731) <= a xor b;
    layer0_outputs(9732) <= not a or b;
    layer0_outputs(9733) <= b and not a;
    layer0_outputs(9734) <= 1'b0;
    layer0_outputs(9735) <= not (a xor b);
    layer0_outputs(9736) <= b;
    layer0_outputs(9737) <= a or b;
    layer0_outputs(9738) <= 1'b0;
    layer0_outputs(9739) <= not (a and b);
    layer0_outputs(9740) <= not a or b;
    layer0_outputs(9741) <= not (a or b);
    layer0_outputs(9742) <= not b;
    layer0_outputs(9743) <= b and not a;
    layer0_outputs(9744) <= not a or b;
    layer0_outputs(9745) <= a and b;
    layer0_outputs(9746) <= a or b;
    layer0_outputs(9747) <= a and b;
    layer0_outputs(9748) <= not a or b;
    layer0_outputs(9749) <= not (a and b);
    layer0_outputs(9750) <= not (a or b);
    layer0_outputs(9751) <= not a or b;
    layer0_outputs(9752) <= 1'b1;
    layer0_outputs(9753) <= a or b;
    layer0_outputs(9754) <= 1'b0;
    layer0_outputs(9755) <= not a or b;
    layer0_outputs(9756) <= b and not a;
    layer0_outputs(9757) <= not a;
    layer0_outputs(9758) <= not a or b;
    layer0_outputs(9759) <= b;
    layer0_outputs(9760) <= a and not b;
    layer0_outputs(9761) <= not b;
    layer0_outputs(9762) <= 1'b0;
    layer0_outputs(9763) <= b and not a;
    layer0_outputs(9764) <= b;
    layer0_outputs(9765) <= a and not b;
    layer0_outputs(9766) <= 1'b1;
    layer0_outputs(9767) <= not a;
    layer0_outputs(9768) <= a and not b;
    layer0_outputs(9769) <= 1'b1;
    layer0_outputs(9770) <= not b;
    layer0_outputs(9771) <= a xor b;
    layer0_outputs(9772) <= a and b;
    layer0_outputs(9773) <= not (a or b);
    layer0_outputs(9774) <= not (a xor b);
    layer0_outputs(9775) <= b and not a;
    layer0_outputs(9776) <= 1'b1;
    layer0_outputs(9777) <= not a;
    layer0_outputs(9778) <= a and b;
    layer0_outputs(9779) <= 1'b0;
    layer0_outputs(9780) <= not b or a;
    layer0_outputs(9781) <= not b;
    layer0_outputs(9782) <= not (a and b);
    layer0_outputs(9783) <= not a;
    layer0_outputs(9784) <= b and not a;
    layer0_outputs(9785) <= not (a xor b);
    layer0_outputs(9786) <= not a;
    layer0_outputs(9787) <= not a;
    layer0_outputs(9788) <= a;
    layer0_outputs(9789) <= not (a and b);
    layer0_outputs(9790) <= a or b;
    layer0_outputs(9791) <= a and not b;
    layer0_outputs(9792) <= b;
    layer0_outputs(9793) <= a or b;
    layer0_outputs(9794) <= not (a and b);
    layer0_outputs(9795) <= not b or a;
    layer0_outputs(9796) <= not b or a;
    layer0_outputs(9797) <= a and not b;
    layer0_outputs(9798) <= not (a xor b);
    layer0_outputs(9799) <= not (a xor b);
    layer0_outputs(9800) <= b;
    layer0_outputs(9801) <= not a;
    layer0_outputs(9802) <= not b or a;
    layer0_outputs(9803) <= not a;
    layer0_outputs(9804) <= not a or b;
    layer0_outputs(9805) <= b and not a;
    layer0_outputs(9806) <= 1'b1;
    layer0_outputs(9807) <= 1'b1;
    layer0_outputs(9808) <= not b or a;
    layer0_outputs(9809) <= not (a or b);
    layer0_outputs(9810) <= not a;
    layer0_outputs(9811) <= not (a or b);
    layer0_outputs(9812) <= not b;
    layer0_outputs(9813) <= b;
    layer0_outputs(9814) <= a;
    layer0_outputs(9815) <= not b;
    layer0_outputs(9816) <= a and not b;
    layer0_outputs(9817) <= not (a and b);
    layer0_outputs(9818) <= not b;
    layer0_outputs(9819) <= b;
    layer0_outputs(9820) <= 1'b0;
    layer0_outputs(9821) <= a;
    layer0_outputs(9822) <= not a;
    layer0_outputs(9823) <= a xor b;
    layer0_outputs(9824) <= a;
    layer0_outputs(9825) <= b;
    layer0_outputs(9826) <= a;
    layer0_outputs(9827) <= b and not a;
    layer0_outputs(9828) <= 1'b1;
    layer0_outputs(9829) <= a;
    layer0_outputs(9830) <= a or b;
    layer0_outputs(9831) <= not a or b;
    layer0_outputs(9832) <= b;
    layer0_outputs(9833) <= not (a or b);
    layer0_outputs(9834) <= not (a and b);
    layer0_outputs(9835) <= a;
    layer0_outputs(9836) <= a xor b;
    layer0_outputs(9837) <= 1'b0;
    layer0_outputs(9838) <= b and not a;
    layer0_outputs(9839) <= b;
    layer0_outputs(9840) <= not (a or b);
    layer0_outputs(9841) <= 1'b0;
    layer0_outputs(9842) <= not b;
    layer0_outputs(9843) <= b;
    layer0_outputs(9844) <= not (a xor b);
    layer0_outputs(9845) <= a or b;
    layer0_outputs(9846) <= a or b;
    layer0_outputs(9847) <= a and b;
    layer0_outputs(9848) <= not a;
    layer0_outputs(9849) <= not (a and b);
    layer0_outputs(9850) <= b;
    layer0_outputs(9851) <= not b or a;
    layer0_outputs(9852) <= a xor b;
    layer0_outputs(9853) <= not (a xor b);
    layer0_outputs(9854) <= a xor b;
    layer0_outputs(9855) <= a and not b;
    layer0_outputs(9856) <= b and not a;
    layer0_outputs(9857) <= 1'b1;
    layer0_outputs(9858) <= not a;
    layer0_outputs(9859) <= a xor b;
    layer0_outputs(9860) <= a and not b;
    layer0_outputs(9861) <= not a or b;
    layer0_outputs(9862) <= not b;
    layer0_outputs(9863) <= 1'b0;
    layer0_outputs(9864) <= not (a or b);
    layer0_outputs(9865) <= 1'b0;
    layer0_outputs(9866) <= a and not b;
    layer0_outputs(9867) <= not (a or b);
    layer0_outputs(9868) <= b;
    layer0_outputs(9869) <= not b;
    layer0_outputs(9870) <= not a;
    layer0_outputs(9871) <= 1'b0;
    layer0_outputs(9872) <= not (a and b);
    layer0_outputs(9873) <= a and b;
    layer0_outputs(9874) <= b and not a;
    layer0_outputs(9875) <= not (a and b);
    layer0_outputs(9876) <= not a or b;
    layer0_outputs(9877) <= 1'b1;
    layer0_outputs(9878) <= not a;
    layer0_outputs(9879) <= 1'b0;
    layer0_outputs(9880) <= a or b;
    layer0_outputs(9881) <= not a or b;
    layer0_outputs(9882) <= b;
    layer0_outputs(9883) <= not a or b;
    layer0_outputs(9884) <= not (a or b);
    layer0_outputs(9885) <= 1'b0;
    layer0_outputs(9886) <= not b or a;
    layer0_outputs(9887) <= 1'b1;
    layer0_outputs(9888) <= 1'b0;
    layer0_outputs(9889) <= not (a or b);
    layer0_outputs(9890) <= not (a or b);
    layer0_outputs(9891) <= a and b;
    layer0_outputs(9892) <= not b or a;
    layer0_outputs(9893) <= not a or b;
    layer0_outputs(9894) <= not b or a;
    layer0_outputs(9895) <= a and b;
    layer0_outputs(9896) <= not (a or b);
    layer0_outputs(9897) <= a and b;
    layer0_outputs(9898) <= a or b;
    layer0_outputs(9899) <= not (a and b);
    layer0_outputs(9900) <= not b or a;
    layer0_outputs(9901) <= not a or b;
    layer0_outputs(9902) <= a and b;
    layer0_outputs(9903) <= a or b;
    layer0_outputs(9904) <= 1'b1;
    layer0_outputs(9905) <= 1'b0;
    layer0_outputs(9906) <= 1'b1;
    layer0_outputs(9907) <= a and b;
    layer0_outputs(9908) <= b;
    layer0_outputs(9909) <= a or b;
    layer0_outputs(9910) <= a and b;
    layer0_outputs(9911) <= not (a or b);
    layer0_outputs(9912) <= not b or a;
    layer0_outputs(9913) <= not b;
    layer0_outputs(9914) <= a;
    layer0_outputs(9915) <= a xor b;
    layer0_outputs(9916) <= not (a xor b);
    layer0_outputs(9917) <= not (a or b);
    layer0_outputs(9918) <= not (a or b);
    layer0_outputs(9919) <= not a;
    layer0_outputs(9920) <= not (a xor b);
    layer0_outputs(9921) <= b;
    layer0_outputs(9922) <= not b or a;
    layer0_outputs(9923) <= a or b;
    layer0_outputs(9924) <= not a;
    layer0_outputs(9925) <= a and not b;
    layer0_outputs(9926) <= a and b;
    layer0_outputs(9927) <= b;
    layer0_outputs(9928) <= not (a or b);
    layer0_outputs(9929) <= a and not b;
    layer0_outputs(9930) <= 1'b1;
    layer0_outputs(9931) <= not b or a;
    layer0_outputs(9932) <= not (a or b);
    layer0_outputs(9933) <= a or b;
    layer0_outputs(9934) <= b;
    layer0_outputs(9935) <= not b;
    layer0_outputs(9936) <= a;
    layer0_outputs(9937) <= b;
    layer0_outputs(9938) <= a or b;
    layer0_outputs(9939) <= not a;
    layer0_outputs(9940) <= not (a or b);
    layer0_outputs(9941) <= 1'b0;
    layer0_outputs(9942) <= a;
    layer0_outputs(9943) <= b;
    layer0_outputs(9944) <= b and not a;
    layer0_outputs(9945) <= b;
    layer0_outputs(9946) <= not a;
    layer0_outputs(9947) <= not a or b;
    layer0_outputs(9948) <= 1'b1;
    layer0_outputs(9949) <= not b or a;
    layer0_outputs(9950) <= not a or b;
    layer0_outputs(9951) <= not (a or b);
    layer0_outputs(9952) <= not (a and b);
    layer0_outputs(9953) <= not b or a;
    layer0_outputs(9954) <= not b;
    layer0_outputs(9955) <= 1'b0;
    layer0_outputs(9956) <= not b;
    layer0_outputs(9957) <= a;
    layer0_outputs(9958) <= a or b;
    layer0_outputs(9959) <= a and b;
    layer0_outputs(9960) <= not a or b;
    layer0_outputs(9961) <= not a;
    layer0_outputs(9962) <= a and b;
    layer0_outputs(9963) <= not (a and b);
    layer0_outputs(9964) <= a or b;
    layer0_outputs(9965) <= a or b;
    layer0_outputs(9966) <= not b;
    layer0_outputs(9967) <= not b;
    layer0_outputs(9968) <= 1'b1;
    layer0_outputs(9969) <= a and b;
    layer0_outputs(9970) <= not b;
    layer0_outputs(9971) <= b;
    layer0_outputs(9972) <= not b or a;
    layer0_outputs(9973) <= not (a and b);
    layer0_outputs(9974) <= 1'b1;
    layer0_outputs(9975) <= a and b;
    layer0_outputs(9976) <= 1'b1;
    layer0_outputs(9977) <= not a;
    layer0_outputs(9978) <= 1'b1;
    layer0_outputs(9979) <= 1'b1;
    layer0_outputs(9980) <= not (a and b);
    layer0_outputs(9981) <= not b;
    layer0_outputs(9982) <= a or b;
    layer0_outputs(9983) <= not a;
    layer0_outputs(9984) <= b;
    layer0_outputs(9985) <= not a;
    layer0_outputs(9986) <= a xor b;
    layer0_outputs(9987) <= not b;
    layer0_outputs(9988) <= b;
    layer0_outputs(9989) <= not (a xor b);
    layer0_outputs(9990) <= not a or b;
    layer0_outputs(9991) <= not (a or b);
    layer0_outputs(9992) <= not a;
    layer0_outputs(9993) <= not (a or b);
    layer0_outputs(9994) <= not (a and b);
    layer0_outputs(9995) <= a and not b;
    layer0_outputs(9996) <= 1'b1;
    layer0_outputs(9997) <= b;
    layer0_outputs(9998) <= b;
    layer0_outputs(9999) <= not b or a;
    layer0_outputs(10000) <= a and not b;
    layer0_outputs(10001) <= a and not b;
    layer0_outputs(10002) <= b;
    layer0_outputs(10003) <= not (a xor b);
    layer0_outputs(10004) <= a;
    layer0_outputs(10005) <= 1'b0;
    layer0_outputs(10006) <= a;
    layer0_outputs(10007) <= not b;
    layer0_outputs(10008) <= a and not b;
    layer0_outputs(10009) <= not a or b;
    layer0_outputs(10010) <= 1'b0;
    layer0_outputs(10011) <= a and b;
    layer0_outputs(10012) <= 1'b0;
    layer0_outputs(10013) <= not b or a;
    layer0_outputs(10014) <= not a;
    layer0_outputs(10015) <= a;
    layer0_outputs(10016) <= not a or b;
    layer0_outputs(10017) <= 1'b0;
    layer0_outputs(10018) <= not b or a;
    layer0_outputs(10019) <= not (a xor b);
    layer0_outputs(10020) <= not a;
    layer0_outputs(10021) <= a;
    layer0_outputs(10022) <= a or b;
    layer0_outputs(10023) <= 1'b1;
    layer0_outputs(10024) <= not b or a;
    layer0_outputs(10025) <= a;
    layer0_outputs(10026) <= a;
    layer0_outputs(10027) <= not (a and b);
    layer0_outputs(10028) <= not a;
    layer0_outputs(10029) <= not a;
    layer0_outputs(10030) <= b and not a;
    layer0_outputs(10031) <= a and b;
    layer0_outputs(10032) <= not a;
    layer0_outputs(10033) <= not b;
    layer0_outputs(10034) <= b and not a;
    layer0_outputs(10035) <= not a;
    layer0_outputs(10036) <= not (a or b);
    layer0_outputs(10037) <= 1'b1;
    layer0_outputs(10038) <= not a;
    layer0_outputs(10039) <= not (a xor b);
    layer0_outputs(10040) <= not (a or b);
    layer0_outputs(10041) <= b and not a;
    layer0_outputs(10042) <= 1'b1;
    layer0_outputs(10043) <= a xor b;
    layer0_outputs(10044) <= b and not a;
    layer0_outputs(10045) <= not b;
    layer0_outputs(10046) <= 1'b1;
    layer0_outputs(10047) <= not b or a;
    layer0_outputs(10048) <= a or b;
    layer0_outputs(10049) <= not b;
    layer0_outputs(10050) <= a;
    layer0_outputs(10051) <= not a;
    layer0_outputs(10052) <= not b or a;
    layer0_outputs(10053) <= 1'b0;
    layer0_outputs(10054) <= not (a xor b);
    layer0_outputs(10055) <= a xor b;
    layer0_outputs(10056) <= not a;
    layer0_outputs(10057) <= a or b;
    layer0_outputs(10058) <= not (a and b);
    layer0_outputs(10059) <= not a;
    layer0_outputs(10060) <= a or b;
    layer0_outputs(10061) <= not (a and b);
    layer0_outputs(10062) <= not (a and b);
    layer0_outputs(10063) <= a xor b;
    layer0_outputs(10064) <= a and not b;
    layer0_outputs(10065) <= 1'b1;
    layer0_outputs(10066) <= 1'b1;
    layer0_outputs(10067) <= a or b;
    layer0_outputs(10068) <= not a or b;
    layer0_outputs(10069) <= not (a or b);
    layer0_outputs(10070) <= a and not b;
    layer0_outputs(10071) <= 1'b0;
    layer0_outputs(10072) <= not a;
    layer0_outputs(10073) <= not a or b;
    layer0_outputs(10074) <= not b;
    layer0_outputs(10075) <= not b;
    layer0_outputs(10076) <= not b or a;
    layer0_outputs(10077) <= b and not a;
    layer0_outputs(10078) <= not (a and b);
    layer0_outputs(10079) <= 1'b0;
    layer0_outputs(10080) <= a xor b;
    layer0_outputs(10081) <= b and not a;
    layer0_outputs(10082) <= 1'b1;
    layer0_outputs(10083) <= a and b;
    layer0_outputs(10084) <= a xor b;
    layer0_outputs(10085) <= a xor b;
    layer0_outputs(10086) <= 1'b0;
    layer0_outputs(10087) <= 1'b0;
    layer0_outputs(10088) <= not (a or b);
    layer0_outputs(10089) <= not b or a;
    layer0_outputs(10090) <= a or b;
    layer0_outputs(10091) <= not b or a;
    layer0_outputs(10092) <= not (a or b);
    layer0_outputs(10093) <= 1'b1;
    layer0_outputs(10094) <= not (a and b);
    layer0_outputs(10095) <= not (a and b);
    layer0_outputs(10096) <= b;
    layer0_outputs(10097) <= not b;
    layer0_outputs(10098) <= not b;
    layer0_outputs(10099) <= not (a or b);
    layer0_outputs(10100) <= not b;
    layer0_outputs(10101) <= not (a or b);
    layer0_outputs(10102) <= a xor b;
    layer0_outputs(10103) <= 1'b1;
    layer0_outputs(10104) <= not b;
    layer0_outputs(10105) <= a;
    layer0_outputs(10106) <= a or b;
    layer0_outputs(10107) <= b and not a;
    layer0_outputs(10108) <= a or b;
    layer0_outputs(10109) <= not b;
    layer0_outputs(10110) <= not a or b;
    layer0_outputs(10111) <= 1'b1;
    layer0_outputs(10112) <= not a;
    layer0_outputs(10113) <= a;
    layer0_outputs(10114) <= not (a and b);
    layer0_outputs(10115) <= a and b;
    layer0_outputs(10116) <= a xor b;
    layer0_outputs(10117) <= not (a and b);
    layer0_outputs(10118) <= not (a xor b);
    layer0_outputs(10119) <= 1'b1;
    layer0_outputs(10120) <= b;
    layer0_outputs(10121) <= not b;
    layer0_outputs(10122) <= not a or b;
    layer0_outputs(10123) <= not b;
    layer0_outputs(10124) <= not b;
    layer0_outputs(10125) <= a and not b;
    layer0_outputs(10126) <= a and not b;
    layer0_outputs(10127) <= 1'b1;
    layer0_outputs(10128) <= not b;
    layer0_outputs(10129) <= a and not b;
    layer0_outputs(10130) <= not b or a;
    layer0_outputs(10131) <= 1'b1;
    layer0_outputs(10132) <= b;
    layer0_outputs(10133) <= a or b;
    layer0_outputs(10134) <= a and not b;
    layer0_outputs(10135) <= 1'b1;
    layer0_outputs(10136) <= not a;
    layer0_outputs(10137) <= a or b;
    layer0_outputs(10138) <= a;
    layer0_outputs(10139) <= b and not a;
    layer0_outputs(10140) <= not (a xor b);
    layer0_outputs(10141) <= a or b;
    layer0_outputs(10142) <= not b;
    layer0_outputs(10143) <= a and not b;
    layer0_outputs(10144) <= not (a or b);
    layer0_outputs(10145) <= not a or b;
    layer0_outputs(10146) <= not (a xor b);
    layer0_outputs(10147) <= not (a and b);
    layer0_outputs(10148) <= a and b;
    layer0_outputs(10149) <= a;
    layer0_outputs(10150) <= a and b;
    layer0_outputs(10151) <= a or b;
    layer0_outputs(10152) <= a;
    layer0_outputs(10153) <= b and not a;
    layer0_outputs(10154) <= not (a and b);
    layer0_outputs(10155) <= not (a and b);
    layer0_outputs(10156) <= not b or a;
    layer0_outputs(10157) <= not b or a;
    layer0_outputs(10158) <= not b;
    layer0_outputs(10159) <= a or b;
    layer0_outputs(10160) <= b and not a;
    layer0_outputs(10161) <= not a;
    layer0_outputs(10162) <= 1'b0;
    layer0_outputs(10163) <= a;
    layer0_outputs(10164) <= b;
    layer0_outputs(10165) <= b;
    layer0_outputs(10166) <= a and not b;
    layer0_outputs(10167) <= not a or b;
    layer0_outputs(10168) <= not a or b;
    layer0_outputs(10169) <= not a;
    layer0_outputs(10170) <= 1'b1;
    layer0_outputs(10171) <= not (a and b);
    layer0_outputs(10172) <= not (a xor b);
    layer0_outputs(10173) <= not b or a;
    layer0_outputs(10174) <= not (a or b);
    layer0_outputs(10175) <= a;
    layer0_outputs(10176) <= not b;
    layer0_outputs(10177) <= not (a xor b);
    layer0_outputs(10178) <= not a;
    layer0_outputs(10179) <= a and not b;
    layer0_outputs(10180) <= a;
    layer0_outputs(10181) <= not a;
    layer0_outputs(10182) <= not (a xor b);
    layer0_outputs(10183) <= not a or b;
    layer0_outputs(10184) <= not a or b;
    layer0_outputs(10185) <= not a or b;
    layer0_outputs(10186) <= 1'b1;
    layer0_outputs(10187) <= not b;
    layer0_outputs(10188) <= a and not b;
    layer0_outputs(10189) <= not b;
    layer0_outputs(10190) <= not (a or b);
    layer0_outputs(10191) <= not (a or b);
    layer0_outputs(10192) <= not b;
    layer0_outputs(10193) <= not a or b;
    layer0_outputs(10194) <= not a;
    layer0_outputs(10195) <= a and b;
    layer0_outputs(10196) <= 1'b0;
    layer0_outputs(10197) <= a xor b;
    layer0_outputs(10198) <= not b or a;
    layer0_outputs(10199) <= not b;
    layer0_outputs(10200) <= not a;
    layer0_outputs(10201) <= not (a or b);
    layer0_outputs(10202) <= 1'b0;
    layer0_outputs(10203) <= 1'b1;
    layer0_outputs(10204) <= not (a and b);
    layer0_outputs(10205) <= a and b;
    layer0_outputs(10206) <= a xor b;
    layer0_outputs(10207) <= a;
    layer0_outputs(10208) <= b and not a;
    layer0_outputs(10209) <= not (a or b);
    layer0_outputs(10210) <= 1'b1;
    layer0_outputs(10211) <= not b;
    layer0_outputs(10212) <= 1'b0;
    layer0_outputs(10213) <= not (a or b);
    layer0_outputs(10214) <= not (a or b);
    layer0_outputs(10215) <= not b or a;
    layer0_outputs(10216) <= not b;
    layer0_outputs(10217) <= a and b;
    layer0_outputs(10218) <= 1'b0;
    layer0_outputs(10219) <= a;
    layer0_outputs(10220) <= a and not b;
    layer0_outputs(10221) <= a and b;
    layer0_outputs(10222) <= a and b;
    layer0_outputs(10223) <= not b;
    layer0_outputs(10224) <= not (a or b);
    layer0_outputs(10225) <= not (a or b);
    layer0_outputs(10226) <= a or b;
    layer0_outputs(10227) <= a xor b;
    layer0_outputs(10228) <= b;
    layer0_outputs(10229) <= not b or a;
    layer0_outputs(10230) <= b and not a;
    layer0_outputs(10231) <= 1'b1;
    layer0_outputs(10232) <= not a;
    layer0_outputs(10233) <= b;
    layer0_outputs(10234) <= not a;
    layer0_outputs(10235) <= a or b;
    layer0_outputs(10236) <= 1'b0;
    layer0_outputs(10237) <= b and not a;
    layer0_outputs(10238) <= 1'b1;
    layer0_outputs(10239) <= a and not b;
    layer1_outputs(0) <= not (a and b);
    layer1_outputs(1) <= a and not b;
    layer1_outputs(2) <= a;
    layer1_outputs(3) <= 1'b1;
    layer1_outputs(4) <= 1'b1;
    layer1_outputs(5) <= 1'b0;
    layer1_outputs(6) <= a xor b;
    layer1_outputs(7) <= not b;
    layer1_outputs(8) <= 1'b1;
    layer1_outputs(9) <= not (a xor b);
    layer1_outputs(10) <= not (a and b);
    layer1_outputs(11) <= not a;
    layer1_outputs(12) <= not b;
    layer1_outputs(13) <= a or b;
    layer1_outputs(14) <= a or b;
    layer1_outputs(15) <= b and not a;
    layer1_outputs(16) <= a or b;
    layer1_outputs(17) <= 1'b1;
    layer1_outputs(18) <= 1'b0;
    layer1_outputs(19) <= not b;
    layer1_outputs(20) <= a;
    layer1_outputs(21) <= a xor b;
    layer1_outputs(22) <= 1'b0;
    layer1_outputs(23) <= 1'b0;
    layer1_outputs(24) <= a or b;
    layer1_outputs(25) <= not (a and b);
    layer1_outputs(26) <= a or b;
    layer1_outputs(27) <= a xor b;
    layer1_outputs(28) <= b and not a;
    layer1_outputs(29) <= not a;
    layer1_outputs(30) <= a and not b;
    layer1_outputs(31) <= not b or a;
    layer1_outputs(32) <= not b;
    layer1_outputs(33) <= not (a or b);
    layer1_outputs(34) <= not b or a;
    layer1_outputs(35) <= not a or b;
    layer1_outputs(36) <= b;
    layer1_outputs(37) <= a and b;
    layer1_outputs(38) <= not (a or b);
    layer1_outputs(39) <= not (a or b);
    layer1_outputs(40) <= b;
    layer1_outputs(41) <= a and not b;
    layer1_outputs(42) <= a xor b;
    layer1_outputs(43) <= b;
    layer1_outputs(44) <= not (a and b);
    layer1_outputs(45) <= not (a or b);
    layer1_outputs(46) <= 1'b1;
    layer1_outputs(47) <= 1'b1;
    layer1_outputs(48) <= a or b;
    layer1_outputs(49) <= a;
    layer1_outputs(50) <= a xor b;
    layer1_outputs(51) <= a;
    layer1_outputs(52) <= a;
    layer1_outputs(53) <= not b or a;
    layer1_outputs(54) <= b and not a;
    layer1_outputs(55) <= not b;
    layer1_outputs(56) <= 1'b1;
    layer1_outputs(57) <= a and b;
    layer1_outputs(58) <= not (a xor b);
    layer1_outputs(59) <= not (a xor b);
    layer1_outputs(60) <= b and not a;
    layer1_outputs(61) <= b;
    layer1_outputs(62) <= not b;
    layer1_outputs(63) <= not b or a;
    layer1_outputs(64) <= not b or a;
    layer1_outputs(65) <= not b or a;
    layer1_outputs(66) <= b and not a;
    layer1_outputs(67) <= a or b;
    layer1_outputs(68) <= not a or b;
    layer1_outputs(69) <= not (a or b);
    layer1_outputs(70) <= b;
    layer1_outputs(71) <= not (a and b);
    layer1_outputs(72) <= a or b;
    layer1_outputs(73) <= not a or b;
    layer1_outputs(74) <= not a;
    layer1_outputs(75) <= not (a or b);
    layer1_outputs(76) <= a and b;
    layer1_outputs(77) <= a;
    layer1_outputs(78) <= not (a and b);
    layer1_outputs(79) <= a and not b;
    layer1_outputs(80) <= b and not a;
    layer1_outputs(81) <= 1'b0;
    layer1_outputs(82) <= not (a or b);
    layer1_outputs(83) <= not (a or b);
    layer1_outputs(84) <= not a;
    layer1_outputs(85) <= not (a and b);
    layer1_outputs(86) <= a and not b;
    layer1_outputs(87) <= a xor b;
    layer1_outputs(88) <= a and b;
    layer1_outputs(89) <= a xor b;
    layer1_outputs(90) <= a or b;
    layer1_outputs(91) <= not b;
    layer1_outputs(92) <= 1'b0;
    layer1_outputs(93) <= not a or b;
    layer1_outputs(94) <= b and not a;
    layer1_outputs(95) <= not b;
    layer1_outputs(96) <= not (a or b);
    layer1_outputs(97) <= b;
    layer1_outputs(98) <= not (a or b);
    layer1_outputs(99) <= a and not b;
    layer1_outputs(100) <= not a;
    layer1_outputs(101) <= 1'b0;
    layer1_outputs(102) <= not (a and b);
    layer1_outputs(103) <= a xor b;
    layer1_outputs(104) <= not b;
    layer1_outputs(105) <= a;
    layer1_outputs(106) <= not (a or b);
    layer1_outputs(107) <= not a or b;
    layer1_outputs(108) <= a or b;
    layer1_outputs(109) <= a and not b;
    layer1_outputs(110) <= b and not a;
    layer1_outputs(111) <= not b;
    layer1_outputs(112) <= not b;
    layer1_outputs(113) <= not a;
    layer1_outputs(114) <= not (a xor b);
    layer1_outputs(115) <= not b;
    layer1_outputs(116) <= not (a or b);
    layer1_outputs(117) <= a;
    layer1_outputs(118) <= not b or a;
    layer1_outputs(119) <= a and b;
    layer1_outputs(120) <= 1'b1;
    layer1_outputs(121) <= 1'b1;
    layer1_outputs(122) <= not (a or b);
    layer1_outputs(123) <= not (a or b);
    layer1_outputs(124) <= not b or a;
    layer1_outputs(125) <= a and not b;
    layer1_outputs(126) <= not b or a;
    layer1_outputs(127) <= a and b;
    layer1_outputs(128) <= b;
    layer1_outputs(129) <= 1'b1;
    layer1_outputs(130) <= a;
    layer1_outputs(131) <= b and not a;
    layer1_outputs(132) <= a or b;
    layer1_outputs(133) <= a and not b;
    layer1_outputs(134) <= not (a or b);
    layer1_outputs(135) <= 1'b1;
    layer1_outputs(136) <= a and b;
    layer1_outputs(137) <= not (a and b);
    layer1_outputs(138) <= a or b;
    layer1_outputs(139) <= not (a xor b);
    layer1_outputs(140) <= a and not b;
    layer1_outputs(141) <= not b or a;
    layer1_outputs(142) <= a;
    layer1_outputs(143) <= 1'b0;
    layer1_outputs(144) <= 1'b1;
    layer1_outputs(145) <= 1'b1;
    layer1_outputs(146) <= b;
    layer1_outputs(147) <= not (a or b);
    layer1_outputs(148) <= not a;
    layer1_outputs(149) <= a and b;
    layer1_outputs(150) <= a and b;
    layer1_outputs(151) <= a;
    layer1_outputs(152) <= 1'b0;
    layer1_outputs(153) <= not b or a;
    layer1_outputs(154) <= a or b;
    layer1_outputs(155) <= 1'b1;
    layer1_outputs(156) <= not (a xor b);
    layer1_outputs(157) <= not (a and b);
    layer1_outputs(158) <= a;
    layer1_outputs(159) <= a and not b;
    layer1_outputs(160) <= a and not b;
    layer1_outputs(161) <= 1'b0;
    layer1_outputs(162) <= not (a and b);
    layer1_outputs(163) <= not a or b;
    layer1_outputs(164) <= not a or b;
    layer1_outputs(165) <= not (a and b);
    layer1_outputs(166) <= 1'b1;
    layer1_outputs(167) <= not b;
    layer1_outputs(168) <= b and not a;
    layer1_outputs(169) <= not b;
    layer1_outputs(170) <= not b;
    layer1_outputs(171) <= a or b;
    layer1_outputs(172) <= a or b;
    layer1_outputs(173) <= 1'b1;
    layer1_outputs(174) <= not (a xor b);
    layer1_outputs(175) <= 1'b1;
    layer1_outputs(176) <= not a or b;
    layer1_outputs(177) <= not (a or b);
    layer1_outputs(178) <= b and not a;
    layer1_outputs(179) <= a and not b;
    layer1_outputs(180) <= a and b;
    layer1_outputs(181) <= a or b;
    layer1_outputs(182) <= not a;
    layer1_outputs(183) <= b and not a;
    layer1_outputs(184) <= b and not a;
    layer1_outputs(185) <= a;
    layer1_outputs(186) <= 1'b1;
    layer1_outputs(187) <= not (a and b);
    layer1_outputs(188) <= b;
    layer1_outputs(189) <= a;
    layer1_outputs(190) <= not b;
    layer1_outputs(191) <= not b or a;
    layer1_outputs(192) <= a;
    layer1_outputs(193) <= b and not a;
    layer1_outputs(194) <= a or b;
    layer1_outputs(195) <= a or b;
    layer1_outputs(196) <= b;
    layer1_outputs(197) <= a;
    layer1_outputs(198) <= not (a or b);
    layer1_outputs(199) <= not a or b;
    layer1_outputs(200) <= b and not a;
    layer1_outputs(201) <= 1'b1;
    layer1_outputs(202) <= 1'b0;
    layer1_outputs(203) <= a and b;
    layer1_outputs(204) <= not b or a;
    layer1_outputs(205) <= a;
    layer1_outputs(206) <= b;
    layer1_outputs(207) <= not a;
    layer1_outputs(208) <= a or b;
    layer1_outputs(209) <= not a or b;
    layer1_outputs(210) <= not (a or b);
    layer1_outputs(211) <= not b or a;
    layer1_outputs(212) <= not a or b;
    layer1_outputs(213) <= a and not b;
    layer1_outputs(214) <= a or b;
    layer1_outputs(215) <= a;
    layer1_outputs(216) <= 1'b0;
    layer1_outputs(217) <= b;
    layer1_outputs(218) <= not b;
    layer1_outputs(219) <= a and b;
    layer1_outputs(220) <= a or b;
    layer1_outputs(221) <= not b;
    layer1_outputs(222) <= a and not b;
    layer1_outputs(223) <= not (a and b);
    layer1_outputs(224) <= a and not b;
    layer1_outputs(225) <= 1'b0;
    layer1_outputs(226) <= b;
    layer1_outputs(227) <= a;
    layer1_outputs(228) <= 1'b1;
    layer1_outputs(229) <= a xor b;
    layer1_outputs(230) <= not (a xor b);
    layer1_outputs(231) <= b and not a;
    layer1_outputs(232) <= 1'b0;
    layer1_outputs(233) <= 1'b0;
    layer1_outputs(234) <= 1'b1;
    layer1_outputs(235) <= a and b;
    layer1_outputs(236) <= 1'b1;
    layer1_outputs(237) <= not (a xor b);
    layer1_outputs(238) <= a and b;
    layer1_outputs(239) <= not (a or b);
    layer1_outputs(240) <= a;
    layer1_outputs(241) <= not a;
    layer1_outputs(242) <= a;
    layer1_outputs(243) <= not b;
    layer1_outputs(244) <= a;
    layer1_outputs(245) <= not b or a;
    layer1_outputs(246) <= a and b;
    layer1_outputs(247) <= 1'b0;
    layer1_outputs(248) <= 1'b0;
    layer1_outputs(249) <= not a;
    layer1_outputs(250) <= not (a and b);
    layer1_outputs(251) <= not a;
    layer1_outputs(252) <= b;
    layer1_outputs(253) <= 1'b1;
    layer1_outputs(254) <= not (a or b);
    layer1_outputs(255) <= a;
    layer1_outputs(256) <= a or b;
    layer1_outputs(257) <= not b;
    layer1_outputs(258) <= b;
    layer1_outputs(259) <= not (a and b);
    layer1_outputs(260) <= not (a or b);
    layer1_outputs(261) <= 1'b1;
    layer1_outputs(262) <= not a;
    layer1_outputs(263) <= b and not a;
    layer1_outputs(264) <= not b or a;
    layer1_outputs(265) <= not a or b;
    layer1_outputs(266) <= a;
    layer1_outputs(267) <= a or b;
    layer1_outputs(268) <= 1'b1;
    layer1_outputs(269) <= not b;
    layer1_outputs(270) <= a and b;
    layer1_outputs(271) <= not a or b;
    layer1_outputs(272) <= 1'b1;
    layer1_outputs(273) <= a and not b;
    layer1_outputs(274) <= not a or b;
    layer1_outputs(275) <= not a or b;
    layer1_outputs(276) <= 1'b0;
    layer1_outputs(277) <= not a;
    layer1_outputs(278) <= not b;
    layer1_outputs(279) <= a or b;
    layer1_outputs(280) <= not b;
    layer1_outputs(281) <= not b or a;
    layer1_outputs(282) <= not b or a;
    layer1_outputs(283) <= a and not b;
    layer1_outputs(284) <= a;
    layer1_outputs(285) <= 1'b0;
    layer1_outputs(286) <= not a;
    layer1_outputs(287) <= not (a xor b);
    layer1_outputs(288) <= 1'b0;
    layer1_outputs(289) <= not b or a;
    layer1_outputs(290) <= 1'b0;
    layer1_outputs(291) <= 1'b0;
    layer1_outputs(292) <= 1'b1;
    layer1_outputs(293) <= a or b;
    layer1_outputs(294) <= not a;
    layer1_outputs(295) <= a;
    layer1_outputs(296) <= a and not b;
    layer1_outputs(297) <= b;
    layer1_outputs(298) <= a and not b;
    layer1_outputs(299) <= not a;
    layer1_outputs(300) <= 1'b1;
    layer1_outputs(301) <= b and not a;
    layer1_outputs(302) <= 1'b0;
    layer1_outputs(303) <= a and not b;
    layer1_outputs(304) <= not (a or b);
    layer1_outputs(305) <= 1'b0;
    layer1_outputs(306) <= a and b;
    layer1_outputs(307) <= not b or a;
    layer1_outputs(308) <= 1'b0;
    layer1_outputs(309) <= a;
    layer1_outputs(310) <= a and b;
    layer1_outputs(311) <= not a;
    layer1_outputs(312) <= a and not b;
    layer1_outputs(313) <= a xor b;
    layer1_outputs(314) <= not a or b;
    layer1_outputs(315) <= not (a or b);
    layer1_outputs(316) <= b;
    layer1_outputs(317) <= b and not a;
    layer1_outputs(318) <= not a or b;
    layer1_outputs(319) <= not a or b;
    layer1_outputs(320) <= not a;
    layer1_outputs(321) <= 1'b1;
    layer1_outputs(322) <= a or b;
    layer1_outputs(323) <= 1'b0;
    layer1_outputs(324) <= a xor b;
    layer1_outputs(325) <= not (a or b);
    layer1_outputs(326) <= b;
    layer1_outputs(327) <= not (a or b);
    layer1_outputs(328) <= b and not a;
    layer1_outputs(329) <= a and b;
    layer1_outputs(330) <= a and b;
    layer1_outputs(331) <= a and not b;
    layer1_outputs(332) <= a or b;
    layer1_outputs(333) <= not (a and b);
    layer1_outputs(334) <= a and b;
    layer1_outputs(335) <= a or b;
    layer1_outputs(336) <= a and b;
    layer1_outputs(337) <= not b or a;
    layer1_outputs(338) <= not a;
    layer1_outputs(339) <= b and not a;
    layer1_outputs(340) <= b;
    layer1_outputs(341) <= a or b;
    layer1_outputs(342) <= a and not b;
    layer1_outputs(343) <= b and not a;
    layer1_outputs(344) <= not a;
    layer1_outputs(345) <= b and not a;
    layer1_outputs(346) <= not b;
    layer1_outputs(347) <= 1'b1;
    layer1_outputs(348) <= 1'b0;
    layer1_outputs(349) <= a;
    layer1_outputs(350) <= not b or a;
    layer1_outputs(351) <= not a or b;
    layer1_outputs(352) <= not (a and b);
    layer1_outputs(353) <= 1'b0;
    layer1_outputs(354) <= not b or a;
    layer1_outputs(355) <= not b or a;
    layer1_outputs(356) <= not (a and b);
    layer1_outputs(357) <= 1'b1;
    layer1_outputs(358) <= not b or a;
    layer1_outputs(359) <= not b or a;
    layer1_outputs(360) <= a and not b;
    layer1_outputs(361) <= not (a and b);
    layer1_outputs(362) <= 1'b0;
    layer1_outputs(363) <= not b or a;
    layer1_outputs(364) <= not (a and b);
    layer1_outputs(365) <= b;
    layer1_outputs(366) <= 1'b0;
    layer1_outputs(367) <= not (a xor b);
    layer1_outputs(368) <= a xor b;
    layer1_outputs(369) <= not a;
    layer1_outputs(370) <= not (a or b);
    layer1_outputs(371) <= not a;
    layer1_outputs(372) <= 1'b0;
    layer1_outputs(373) <= not a or b;
    layer1_outputs(374) <= a and not b;
    layer1_outputs(375) <= not a or b;
    layer1_outputs(376) <= 1'b0;
    layer1_outputs(377) <= not (a and b);
    layer1_outputs(378) <= not b or a;
    layer1_outputs(379) <= a and b;
    layer1_outputs(380) <= not (a or b);
    layer1_outputs(381) <= not (a or b);
    layer1_outputs(382) <= a and not b;
    layer1_outputs(383) <= not (a and b);
    layer1_outputs(384) <= a or b;
    layer1_outputs(385) <= b;
    layer1_outputs(386) <= not a or b;
    layer1_outputs(387) <= not a;
    layer1_outputs(388) <= a or b;
    layer1_outputs(389) <= a or b;
    layer1_outputs(390) <= not b;
    layer1_outputs(391) <= a;
    layer1_outputs(392) <= not a;
    layer1_outputs(393) <= not (a or b);
    layer1_outputs(394) <= not a;
    layer1_outputs(395) <= b;
    layer1_outputs(396) <= not b;
    layer1_outputs(397) <= 1'b0;
    layer1_outputs(398) <= 1'b1;
    layer1_outputs(399) <= not a or b;
    layer1_outputs(400) <= 1'b0;
    layer1_outputs(401) <= not a or b;
    layer1_outputs(402) <= 1'b0;
    layer1_outputs(403) <= a;
    layer1_outputs(404) <= a and not b;
    layer1_outputs(405) <= 1'b0;
    layer1_outputs(406) <= 1'b0;
    layer1_outputs(407) <= not a;
    layer1_outputs(408) <= not (a and b);
    layer1_outputs(409) <= not (a or b);
    layer1_outputs(410) <= a or b;
    layer1_outputs(411) <= b;
    layer1_outputs(412) <= a or b;
    layer1_outputs(413) <= 1'b0;
    layer1_outputs(414) <= b and not a;
    layer1_outputs(415) <= 1'b1;
    layer1_outputs(416) <= 1'b1;
    layer1_outputs(417) <= not (a or b);
    layer1_outputs(418) <= a or b;
    layer1_outputs(419) <= not a or b;
    layer1_outputs(420) <= not (a and b);
    layer1_outputs(421) <= 1'b0;
    layer1_outputs(422) <= b;
    layer1_outputs(423) <= not (a or b);
    layer1_outputs(424) <= 1'b1;
    layer1_outputs(425) <= a;
    layer1_outputs(426) <= not (a or b);
    layer1_outputs(427) <= a xor b;
    layer1_outputs(428) <= 1'b0;
    layer1_outputs(429) <= a and b;
    layer1_outputs(430) <= not a;
    layer1_outputs(431) <= a and not b;
    layer1_outputs(432) <= a xor b;
    layer1_outputs(433) <= 1'b1;
    layer1_outputs(434) <= 1'b1;
    layer1_outputs(435) <= b and not a;
    layer1_outputs(436) <= not b or a;
    layer1_outputs(437) <= b and not a;
    layer1_outputs(438) <= not (a and b);
    layer1_outputs(439) <= a or b;
    layer1_outputs(440) <= b;
    layer1_outputs(441) <= not b;
    layer1_outputs(442) <= a and not b;
    layer1_outputs(443) <= a or b;
    layer1_outputs(444) <= not (a xor b);
    layer1_outputs(445) <= a;
    layer1_outputs(446) <= 1'b0;
    layer1_outputs(447) <= not a or b;
    layer1_outputs(448) <= not (a and b);
    layer1_outputs(449) <= not a or b;
    layer1_outputs(450) <= b and not a;
    layer1_outputs(451) <= a or b;
    layer1_outputs(452) <= a;
    layer1_outputs(453) <= not (a and b);
    layer1_outputs(454) <= 1'b1;
    layer1_outputs(455) <= a or b;
    layer1_outputs(456) <= b and not a;
    layer1_outputs(457) <= not b;
    layer1_outputs(458) <= 1'b0;
    layer1_outputs(459) <= not a or b;
    layer1_outputs(460) <= a or b;
    layer1_outputs(461) <= b and not a;
    layer1_outputs(462) <= not a or b;
    layer1_outputs(463) <= not (a and b);
    layer1_outputs(464) <= b and not a;
    layer1_outputs(465) <= a or b;
    layer1_outputs(466) <= 1'b1;
    layer1_outputs(467) <= 1'b1;
    layer1_outputs(468) <= b;
    layer1_outputs(469) <= a and not b;
    layer1_outputs(470) <= 1'b1;
    layer1_outputs(471) <= not b;
    layer1_outputs(472) <= a or b;
    layer1_outputs(473) <= a;
    layer1_outputs(474) <= a and b;
    layer1_outputs(475) <= not b or a;
    layer1_outputs(476) <= a or b;
    layer1_outputs(477) <= 1'b0;
    layer1_outputs(478) <= not a;
    layer1_outputs(479) <= 1'b1;
    layer1_outputs(480) <= b;
    layer1_outputs(481) <= not (a and b);
    layer1_outputs(482) <= not a;
    layer1_outputs(483) <= b;
    layer1_outputs(484) <= not (a or b);
    layer1_outputs(485) <= not (a and b);
    layer1_outputs(486) <= not (a or b);
    layer1_outputs(487) <= not (a and b);
    layer1_outputs(488) <= not a;
    layer1_outputs(489) <= 1'b0;
    layer1_outputs(490) <= 1'b1;
    layer1_outputs(491) <= a or b;
    layer1_outputs(492) <= b;
    layer1_outputs(493) <= 1'b0;
    layer1_outputs(494) <= not (a or b);
    layer1_outputs(495) <= 1'b1;
    layer1_outputs(496) <= a or b;
    layer1_outputs(497) <= a or b;
    layer1_outputs(498) <= 1'b0;
    layer1_outputs(499) <= b and not a;
    layer1_outputs(500) <= not (a and b);
    layer1_outputs(501) <= 1'b0;
    layer1_outputs(502) <= b and not a;
    layer1_outputs(503) <= a and b;
    layer1_outputs(504) <= not (a and b);
    layer1_outputs(505) <= 1'b1;
    layer1_outputs(506) <= not b or a;
    layer1_outputs(507) <= a and b;
    layer1_outputs(508) <= not (a and b);
    layer1_outputs(509) <= a;
    layer1_outputs(510) <= 1'b1;
    layer1_outputs(511) <= not b;
    layer1_outputs(512) <= b and not a;
    layer1_outputs(513) <= not (a or b);
    layer1_outputs(514) <= not b or a;
    layer1_outputs(515) <= not a or b;
    layer1_outputs(516) <= a;
    layer1_outputs(517) <= not a;
    layer1_outputs(518) <= a or b;
    layer1_outputs(519) <= not (a or b);
    layer1_outputs(520) <= a and not b;
    layer1_outputs(521) <= not (a or b);
    layer1_outputs(522) <= b and not a;
    layer1_outputs(523) <= not b or a;
    layer1_outputs(524) <= not a or b;
    layer1_outputs(525) <= 1'b0;
    layer1_outputs(526) <= not b or a;
    layer1_outputs(527) <= a or b;
    layer1_outputs(528) <= b;
    layer1_outputs(529) <= 1'b1;
    layer1_outputs(530) <= a or b;
    layer1_outputs(531) <= not b or a;
    layer1_outputs(532) <= 1'b1;
    layer1_outputs(533) <= b;
    layer1_outputs(534) <= b and not a;
    layer1_outputs(535) <= 1'b0;
    layer1_outputs(536) <= a;
    layer1_outputs(537) <= not a;
    layer1_outputs(538) <= b;
    layer1_outputs(539) <= b;
    layer1_outputs(540) <= not a or b;
    layer1_outputs(541) <= a and b;
    layer1_outputs(542) <= not a;
    layer1_outputs(543) <= not (a or b);
    layer1_outputs(544) <= not (a xor b);
    layer1_outputs(545) <= b;
    layer1_outputs(546) <= not a or b;
    layer1_outputs(547) <= a;
    layer1_outputs(548) <= not b or a;
    layer1_outputs(549) <= not (a and b);
    layer1_outputs(550) <= not (a or b);
    layer1_outputs(551) <= a and b;
    layer1_outputs(552) <= not (a and b);
    layer1_outputs(553) <= a and b;
    layer1_outputs(554) <= not (a or b);
    layer1_outputs(555) <= a or b;
    layer1_outputs(556) <= a;
    layer1_outputs(557) <= b;
    layer1_outputs(558) <= a and not b;
    layer1_outputs(559) <= 1'b1;
    layer1_outputs(560) <= a and b;
    layer1_outputs(561) <= not b;
    layer1_outputs(562) <= a and not b;
    layer1_outputs(563) <= b and not a;
    layer1_outputs(564) <= a xor b;
    layer1_outputs(565) <= not a or b;
    layer1_outputs(566) <= a and b;
    layer1_outputs(567) <= a and not b;
    layer1_outputs(568) <= a xor b;
    layer1_outputs(569) <= b and not a;
    layer1_outputs(570) <= not (a or b);
    layer1_outputs(571) <= not (a or b);
    layer1_outputs(572) <= a and b;
    layer1_outputs(573) <= a xor b;
    layer1_outputs(574) <= a or b;
    layer1_outputs(575) <= not b or a;
    layer1_outputs(576) <= not b;
    layer1_outputs(577) <= a;
    layer1_outputs(578) <= b;
    layer1_outputs(579) <= 1'b1;
    layer1_outputs(580) <= not (a and b);
    layer1_outputs(581) <= 1'b1;
    layer1_outputs(582) <= not (a or b);
    layer1_outputs(583) <= not a or b;
    layer1_outputs(584) <= not a;
    layer1_outputs(585) <= not b;
    layer1_outputs(586) <= 1'b1;
    layer1_outputs(587) <= a and not b;
    layer1_outputs(588) <= 1'b1;
    layer1_outputs(589) <= a and b;
    layer1_outputs(590) <= not a or b;
    layer1_outputs(591) <= a or b;
    layer1_outputs(592) <= a and not b;
    layer1_outputs(593) <= b;
    layer1_outputs(594) <= 1'b0;
    layer1_outputs(595) <= a and b;
    layer1_outputs(596) <= a and not b;
    layer1_outputs(597) <= 1'b0;
    layer1_outputs(598) <= not b or a;
    layer1_outputs(599) <= b;
    layer1_outputs(600) <= not (a and b);
    layer1_outputs(601) <= a xor b;
    layer1_outputs(602) <= b;
    layer1_outputs(603) <= a and b;
    layer1_outputs(604) <= a xor b;
    layer1_outputs(605) <= 1'b0;
    layer1_outputs(606) <= not b;
    layer1_outputs(607) <= 1'b0;
    layer1_outputs(608) <= b;
    layer1_outputs(609) <= a and not b;
    layer1_outputs(610) <= a or b;
    layer1_outputs(611) <= not b;
    layer1_outputs(612) <= 1'b1;
    layer1_outputs(613) <= not b;
    layer1_outputs(614) <= not b or a;
    layer1_outputs(615) <= b;
    layer1_outputs(616) <= a or b;
    layer1_outputs(617) <= 1'b0;
    layer1_outputs(618) <= a and b;
    layer1_outputs(619) <= a or b;
    layer1_outputs(620) <= b;
    layer1_outputs(621) <= not (a or b);
    layer1_outputs(622) <= a;
    layer1_outputs(623) <= not a;
    layer1_outputs(624) <= not (a and b);
    layer1_outputs(625) <= not (a and b);
    layer1_outputs(626) <= 1'b1;
    layer1_outputs(627) <= not b or a;
    layer1_outputs(628) <= not a;
    layer1_outputs(629) <= not b or a;
    layer1_outputs(630) <= not b;
    layer1_outputs(631) <= 1'b1;
    layer1_outputs(632) <= not b or a;
    layer1_outputs(633) <= b;
    layer1_outputs(634) <= a and b;
    layer1_outputs(635) <= 1'b0;
    layer1_outputs(636) <= a and not b;
    layer1_outputs(637) <= not b or a;
    layer1_outputs(638) <= 1'b1;
    layer1_outputs(639) <= not b;
    layer1_outputs(640) <= not a or b;
    layer1_outputs(641) <= not a;
    layer1_outputs(642) <= 1'b0;
    layer1_outputs(643) <= a and not b;
    layer1_outputs(644) <= not b or a;
    layer1_outputs(645) <= not a;
    layer1_outputs(646) <= not b or a;
    layer1_outputs(647) <= not (a and b);
    layer1_outputs(648) <= 1'b0;
    layer1_outputs(649) <= 1'b1;
    layer1_outputs(650) <= not (a and b);
    layer1_outputs(651) <= not b or a;
    layer1_outputs(652) <= a;
    layer1_outputs(653) <= not (a xor b);
    layer1_outputs(654) <= b;
    layer1_outputs(655) <= a or b;
    layer1_outputs(656) <= a;
    layer1_outputs(657) <= not (a or b);
    layer1_outputs(658) <= a;
    layer1_outputs(659) <= 1'b0;
    layer1_outputs(660) <= b and not a;
    layer1_outputs(661) <= 1'b1;
    layer1_outputs(662) <= not b;
    layer1_outputs(663) <= a or b;
    layer1_outputs(664) <= b and not a;
    layer1_outputs(665) <= a;
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= a or b;
    layer1_outputs(668) <= 1'b1;
    layer1_outputs(669) <= not a or b;
    layer1_outputs(670) <= not a;
    layer1_outputs(671) <= not a or b;
    layer1_outputs(672) <= a;
    layer1_outputs(673) <= not a or b;
    layer1_outputs(674) <= not b or a;
    layer1_outputs(675) <= not a;
    layer1_outputs(676) <= 1'b1;
    layer1_outputs(677) <= not b;
    layer1_outputs(678) <= b;
    layer1_outputs(679) <= not (a or b);
    layer1_outputs(680) <= not b or a;
    layer1_outputs(681) <= a;
    layer1_outputs(682) <= 1'b0;
    layer1_outputs(683) <= 1'b1;
    layer1_outputs(684) <= a xor b;
    layer1_outputs(685) <= 1'b1;
    layer1_outputs(686) <= a and not b;
    layer1_outputs(687) <= a or b;
    layer1_outputs(688) <= b;
    layer1_outputs(689) <= not a;
    layer1_outputs(690) <= 1'b0;
    layer1_outputs(691) <= 1'b1;
    layer1_outputs(692) <= a;
    layer1_outputs(693) <= not a;
    layer1_outputs(694) <= b;
    layer1_outputs(695) <= not (a or b);
    layer1_outputs(696) <= 1'b0;
    layer1_outputs(697) <= not a;
    layer1_outputs(698) <= 1'b1;
    layer1_outputs(699) <= not a;
    layer1_outputs(700) <= 1'b0;
    layer1_outputs(701) <= a;
    layer1_outputs(702) <= 1'b0;
    layer1_outputs(703) <= not a or b;
    layer1_outputs(704) <= 1'b0;
    layer1_outputs(705) <= a xor b;
    layer1_outputs(706) <= not b or a;
    layer1_outputs(707) <= a and not b;
    layer1_outputs(708) <= 1'b0;
    layer1_outputs(709) <= not a;
    layer1_outputs(710) <= a and not b;
    layer1_outputs(711) <= a or b;
    layer1_outputs(712) <= not (a or b);
    layer1_outputs(713) <= a xor b;
    layer1_outputs(714) <= 1'b1;
    layer1_outputs(715) <= b and not a;
    layer1_outputs(716) <= a or b;
    layer1_outputs(717) <= not b or a;
    layer1_outputs(718) <= not b or a;
    layer1_outputs(719) <= a and not b;
    layer1_outputs(720) <= a and not b;
    layer1_outputs(721) <= a;
    layer1_outputs(722) <= a and b;
    layer1_outputs(723) <= 1'b1;
    layer1_outputs(724) <= a and b;
    layer1_outputs(725) <= a xor b;
    layer1_outputs(726) <= not a or b;
    layer1_outputs(727) <= a;
    layer1_outputs(728) <= not a or b;
    layer1_outputs(729) <= a or b;
    layer1_outputs(730) <= a;
    layer1_outputs(731) <= a or b;
    layer1_outputs(732) <= not a or b;
    layer1_outputs(733) <= 1'b1;
    layer1_outputs(734) <= b;
    layer1_outputs(735) <= not b;
    layer1_outputs(736) <= a and not b;
    layer1_outputs(737) <= 1'b1;
    layer1_outputs(738) <= not a or b;
    layer1_outputs(739) <= a;
    layer1_outputs(740) <= 1'b0;
    layer1_outputs(741) <= a;
    layer1_outputs(742) <= b;
    layer1_outputs(743) <= not (a and b);
    layer1_outputs(744) <= 1'b0;
    layer1_outputs(745) <= not (a or b);
    layer1_outputs(746) <= b and not a;
    layer1_outputs(747) <= 1'b0;
    layer1_outputs(748) <= a;
    layer1_outputs(749) <= not b;
    layer1_outputs(750) <= 1'b1;
    layer1_outputs(751) <= 1'b0;
    layer1_outputs(752) <= not b or a;
    layer1_outputs(753) <= not (a or b);
    layer1_outputs(754) <= 1'b1;
    layer1_outputs(755) <= b;
    layer1_outputs(756) <= a and b;
    layer1_outputs(757) <= 1'b0;
    layer1_outputs(758) <= a;
    layer1_outputs(759) <= a and not b;
    layer1_outputs(760) <= a;
    layer1_outputs(761) <= not (a or b);
    layer1_outputs(762) <= not b or a;
    layer1_outputs(763) <= not b or a;
    layer1_outputs(764) <= not (a or b);
    layer1_outputs(765) <= a xor b;
    layer1_outputs(766) <= not (a xor b);
    layer1_outputs(767) <= not a or b;
    layer1_outputs(768) <= not (a and b);
    layer1_outputs(769) <= not (a and b);
    layer1_outputs(770) <= not a or b;
    layer1_outputs(771) <= a or b;
    layer1_outputs(772) <= not (a and b);
    layer1_outputs(773) <= not (a xor b);
    layer1_outputs(774) <= not a or b;
    layer1_outputs(775) <= not a;
    layer1_outputs(776) <= not b or a;
    layer1_outputs(777) <= a xor b;
    layer1_outputs(778) <= 1'b1;
    layer1_outputs(779) <= not (a and b);
    layer1_outputs(780) <= not b or a;
    layer1_outputs(781) <= a;
    layer1_outputs(782) <= b and not a;
    layer1_outputs(783) <= a and b;
    layer1_outputs(784) <= not b;
    layer1_outputs(785) <= not b or a;
    layer1_outputs(786) <= a;
    layer1_outputs(787) <= a;
    layer1_outputs(788) <= not a;
    layer1_outputs(789) <= a and not b;
    layer1_outputs(790) <= b and not a;
    layer1_outputs(791) <= b and not a;
    layer1_outputs(792) <= not a or b;
    layer1_outputs(793) <= a or b;
    layer1_outputs(794) <= not a or b;
    layer1_outputs(795) <= a;
    layer1_outputs(796) <= b;
    layer1_outputs(797) <= not (a and b);
    layer1_outputs(798) <= not a;
    layer1_outputs(799) <= 1'b0;
    layer1_outputs(800) <= not b;
    layer1_outputs(801) <= a or b;
    layer1_outputs(802) <= a;
    layer1_outputs(803) <= 1'b1;
    layer1_outputs(804) <= 1'b1;
    layer1_outputs(805) <= a;
    layer1_outputs(806) <= b;
    layer1_outputs(807) <= not a;
    layer1_outputs(808) <= b;
    layer1_outputs(809) <= a and b;
    layer1_outputs(810) <= 1'b0;
    layer1_outputs(811) <= not b or a;
    layer1_outputs(812) <= b and not a;
    layer1_outputs(813) <= not b;
    layer1_outputs(814) <= not (a xor b);
    layer1_outputs(815) <= a xor b;
    layer1_outputs(816) <= b and not a;
    layer1_outputs(817) <= a xor b;
    layer1_outputs(818) <= a and not b;
    layer1_outputs(819) <= not b or a;
    layer1_outputs(820) <= b;
    layer1_outputs(821) <= not a;
    layer1_outputs(822) <= a;
    layer1_outputs(823) <= not b;
    layer1_outputs(824) <= not b or a;
    layer1_outputs(825) <= not b;
    layer1_outputs(826) <= not a;
    layer1_outputs(827) <= not a or b;
    layer1_outputs(828) <= not (a or b);
    layer1_outputs(829) <= a and not b;
    layer1_outputs(830) <= a;
    layer1_outputs(831) <= 1'b0;
    layer1_outputs(832) <= b;
    layer1_outputs(833) <= not (a or b);
    layer1_outputs(834) <= a or b;
    layer1_outputs(835) <= not b;
    layer1_outputs(836) <= a;
    layer1_outputs(837) <= b and not a;
    layer1_outputs(838) <= not a or b;
    layer1_outputs(839) <= 1'b1;
    layer1_outputs(840) <= not b or a;
    layer1_outputs(841) <= b;
    layer1_outputs(842) <= not (a or b);
    layer1_outputs(843) <= not a or b;
    layer1_outputs(844) <= a and b;
    layer1_outputs(845) <= b;
    layer1_outputs(846) <= not a or b;
    layer1_outputs(847) <= 1'b1;
    layer1_outputs(848) <= 1'b1;
    layer1_outputs(849) <= not (a or b);
    layer1_outputs(850) <= b and not a;
    layer1_outputs(851) <= a and not b;
    layer1_outputs(852) <= not b;
    layer1_outputs(853) <= not (a or b);
    layer1_outputs(854) <= not a or b;
    layer1_outputs(855) <= 1'b0;
    layer1_outputs(856) <= b and not a;
    layer1_outputs(857) <= not (a and b);
    layer1_outputs(858) <= b and not a;
    layer1_outputs(859) <= 1'b1;
    layer1_outputs(860) <= not b or a;
    layer1_outputs(861) <= not (a or b);
    layer1_outputs(862) <= b;
    layer1_outputs(863) <= a and not b;
    layer1_outputs(864) <= a;
    layer1_outputs(865) <= not b or a;
    layer1_outputs(866) <= a and b;
    layer1_outputs(867) <= not (a or b);
    layer1_outputs(868) <= not a;
    layer1_outputs(869) <= a or b;
    layer1_outputs(870) <= 1'b1;
    layer1_outputs(871) <= not b or a;
    layer1_outputs(872) <= b and not a;
    layer1_outputs(873) <= a or b;
    layer1_outputs(874) <= not (a or b);
    layer1_outputs(875) <= 1'b1;
    layer1_outputs(876) <= a and not b;
    layer1_outputs(877) <= a xor b;
    layer1_outputs(878) <= not (a xor b);
    layer1_outputs(879) <= a and b;
    layer1_outputs(880) <= not b or a;
    layer1_outputs(881) <= 1'b0;
    layer1_outputs(882) <= not a;
    layer1_outputs(883) <= 1'b1;
    layer1_outputs(884) <= a or b;
    layer1_outputs(885) <= 1'b1;
    layer1_outputs(886) <= b and not a;
    layer1_outputs(887) <= 1'b0;
    layer1_outputs(888) <= not (a and b);
    layer1_outputs(889) <= a and b;
    layer1_outputs(890) <= a and b;
    layer1_outputs(891) <= not a or b;
    layer1_outputs(892) <= b;
    layer1_outputs(893) <= not (a xor b);
    layer1_outputs(894) <= 1'b1;
    layer1_outputs(895) <= b;
    layer1_outputs(896) <= not (a or b);
    layer1_outputs(897) <= not (a or b);
    layer1_outputs(898) <= b and not a;
    layer1_outputs(899) <= b;
    layer1_outputs(900) <= not a;
    layer1_outputs(901) <= not (a and b);
    layer1_outputs(902) <= a or b;
    layer1_outputs(903) <= b;
    layer1_outputs(904) <= 1'b1;
    layer1_outputs(905) <= not a;
    layer1_outputs(906) <= a and not b;
    layer1_outputs(907) <= not (a and b);
    layer1_outputs(908) <= a;
    layer1_outputs(909) <= not (a or b);
    layer1_outputs(910) <= 1'b1;
    layer1_outputs(911) <= 1'b1;
    layer1_outputs(912) <= not a;
    layer1_outputs(913) <= 1'b0;
    layer1_outputs(914) <= a or b;
    layer1_outputs(915) <= a;
    layer1_outputs(916) <= 1'b1;
    layer1_outputs(917) <= not (a and b);
    layer1_outputs(918) <= a and b;
    layer1_outputs(919) <= not (a or b);
    layer1_outputs(920) <= a;
    layer1_outputs(921) <= b and not a;
    layer1_outputs(922) <= a or b;
    layer1_outputs(923) <= a or b;
    layer1_outputs(924) <= not b;
    layer1_outputs(925) <= 1'b0;
    layer1_outputs(926) <= 1'b1;
    layer1_outputs(927) <= 1'b0;
    layer1_outputs(928) <= 1'b1;
    layer1_outputs(929) <= not b or a;
    layer1_outputs(930) <= a and not b;
    layer1_outputs(931) <= 1'b0;
    layer1_outputs(932) <= not (a and b);
    layer1_outputs(933) <= 1'b0;
    layer1_outputs(934) <= b;
    layer1_outputs(935) <= a;
    layer1_outputs(936) <= 1'b1;
    layer1_outputs(937) <= a and not b;
    layer1_outputs(938) <= 1'b0;
    layer1_outputs(939) <= not b;
    layer1_outputs(940) <= 1'b1;
    layer1_outputs(941) <= b;
    layer1_outputs(942) <= not b;
    layer1_outputs(943) <= not a;
    layer1_outputs(944) <= 1'b0;
    layer1_outputs(945) <= 1'b0;
    layer1_outputs(946) <= a or b;
    layer1_outputs(947) <= a or b;
    layer1_outputs(948) <= a;
    layer1_outputs(949) <= not (a and b);
    layer1_outputs(950) <= a and b;
    layer1_outputs(951) <= a;
    layer1_outputs(952) <= not a;
    layer1_outputs(953) <= not a;
    layer1_outputs(954) <= a and not b;
    layer1_outputs(955) <= a or b;
    layer1_outputs(956) <= not (a or b);
    layer1_outputs(957) <= 1'b1;
    layer1_outputs(958) <= 1'b1;
    layer1_outputs(959) <= a;
    layer1_outputs(960) <= a;
    layer1_outputs(961) <= not (a or b);
    layer1_outputs(962) <= b and not a;
    layer1_outputs(963) <= a xor b;
    layer1_outputs(964) <= not (a xor b);
    layer1_outputs(965) <= not (a or b);
    layer1_outputs(966) <= 1'b1;
    layer1_outputs(967) <= not (a and b);
    layer1_outputs(968) <= 1'b0;
    layer1_outputs(969) <= not b or a;
    layer1_outputs(970) <= b and not a;
    layer1_outputs(971) <= not (a or b);
    layer1_outputs(972) <= not (a or b);
    layer1_outputs(973) <= not (a and b);
    layer1_outputs(974) <= a and not b;
    layer1_outputs(975) <= 1'b0;
    layer1_outputs(976) <= a xor b;
    layer1_outputs(977) <= a and b;
    layer1_outputs(978) <= b;
    layer1_outputs(979) <= not b or a;
    layer1_outputs(980) <= 1'b1;
    layer1_outputs(981) <= a and b;
    layer1_outputs(982) <= not a;
    layer1_outputs(983) <= not a or b;
    layer1_outputs(984) <= a and not b;
    layer1_outputs(985) <= b and not a;
    layer1_outputs(986) <= not (a and b);
    layer1_outputs(987) <= a and not b;
    layer1_outputs(988) <= 1'b0;
    layer1_outputs(989) <= b;
    layer1_outputs(990) <= not (a and b);
    layer1_outputs(991) <= b and not a;
    layer1_outputs(992) <= not a or b;
    layer1_outputs(993) <= a and not b;
    layer1_outputs(994) <= b;
    layer1_outputs(995) <= b;
    layer1_outputs(996) <= a or b;
    layer1_outputs(997) <= 1'b0;
    layer1_outputs(998) <= a;
    layer1_outputs(999) <= not a or b;
    layer1_outputs(1000) <= not (a xor b);
    layer1_outputs(1001) <= a;
    layer1_outputs(1002) <= b and not a;
    layer1_outputs(1003) <= 1'b1;
    layer1_outputs(1004) <= not b;
    layer1_outputs(1005) <= a;
    layer1_outputs(1006) <= a or b;
    layer1_outputs(1007) <= a and b;
    layer1_outputs(1008) <= not (a xor b);
    layer1_outputs(1009) <= 1'b1;
    layer1_outputs(1010) <= not b;
    layer1_outputs(1011) <= not b;
    layer1_outputs(1012) <= not a;
    layer1_outputs(1013) <= not a or b;
    layer1_outputs(1014) <= not b or a;
    layer1_outputs(1015) <= b and not a;
    layer1_outputs(1016) <= not a or b;
    layer1_outputs(1017) <= b;
    layer1_outputs(1018) <= a and b;
    layer1_outputs(1019) <= a and not b;
    layer1_outputs(1020) <= a or b;
    layer1_outputs(1021) <= not b or a;
    layer1_outputs(1022) <= not (a and b);
    layer1_outputs(1023) <= not b;
    layer1_outputs(1024) <= not a;
    layer1_outputs(1025) <= not (a xor b);
    layer1_outputs(1026) <= not a or b;
    layer1_outputs(1027) <= not b;
    layer1_outputs(1028) <= not a;
    layer1_outputs(1029) <= 1'b0;
    layer1_outputs(1030) <= 1'b1;
    layer1_outputs(1031) <= not b or a;
    layer1_outputs(1032) <= 1'b0;
    layer1_outputs(1033) <= not (a and b);
    layer1_outputs(1034) <= not b;
    layer1_outputs(1035) <= 1'b0;
    layer1_outputs(1036) <= not (a or b);
    layer1_outputs(1037) <= not (a and b);
    layer1_outputs(1038) <= not (a or b);
    layer1_outputs(1039) <= not (a and b);
    layer1_outputs(1040) <= b;
    layer1_outputs(1041) <= a and not b;
    layer1_outputs(1042) <= 1'b0;
    layer1_outputs(1043) <= a xor b;
    layer1_outputs(1044) <= not a;
    layer1_outputs(1045) <= a and b;
    layer1_outputs(1046) <= not a;
    layer1_outputs(1047) <= not a or b;
    layer1_outputs(1048) <= a and b;
    layer1_outputs(1049) <= not a;
    layer1_outputs(1050) <= b;
    layer1_outputs(1051) <= a and b;
    layer1_outputs(1052) <= not a;
    layer1_outputs(1053) <= not (a or b);
    layer1_outputs(1054) <= not b or a;
    layer1_outputs(1055) <= 1'b1;
    layer1_outputs(1056) <= a;
    layer1_outputs(1057) <= not (a or b);
    layer1_outputs(1058) <= not (a and b);
    layer1_outputs(1059) <= not (a and b);
    layer1_outputs(1060) <= 1'b0;
    layer1_outputs(1061) <= not (a or b);
    layer1_outputs(1062) <= a and b;
    layer1_outputs(1063) <= 1'b1;
    layer1_outputs(1064) <= not b;
    layer1_outputs(1065) <= a;
    layer1_outputs(1066) <= a and not b;
    layer1_outputs(1067) <= not a;
    layer1_outputs(1068) <= not (a and b);
    layer1_outputs(1069) <= 1'b1;
    layer1_outputs(1070) <= a and not b;
    layer1_outputs(1071) <= a or b;
    layer1_outputs(1072) <= not (a and b);
    layer1_outputs(1073) <= b;
    layer1_outputs(1074) <= 1'b1;
    layer1_outputs(1075) <= not a;
    layer1_outputs(1076) <= 1'b1;
    layer1_outputs(1077) <= not (a and b);
    layer1_outputs(1078) <= b and not a;
    layer1_outputs(1079) <= not (a or b);
    layer1_outputs(1080) <= not (a or b);
    layer1_outputs(1081) <= not b or a;
    layer1_outputs(1082) <= b;
    layer1_outputs(1083) <= a or b;
    layer1_outputs(1084) <= 1'b0;
    layer1_outputs(1085) <= not b;
    layer1_outputs(1086) <= a;
    layer1_outputs(1087) <= b and not a;
    layer1_outputs(1088) <= a and b;
    layer1_outputs(1089) <= 1'b0;
    layer1_outputs(1090) <= not (a or b);
    layer1_outputs(1091) <= not a or b;
    layer1_outputs(1092) <= not b or a;
    layer1_outputs(1093) <= 1'b1;
    layer1_outputs(1094) <= not (a or b);
    layer1_outputs(1095) <= 1'b0;
    layer1_outputs(1096) <= a or b;
    layer1_outputs(1097) <= 1'b0;
    layer1_outputs(1098) <= 1'b0;
    layer1_outputs(1099) <= not (a xor b);
    layer1_outputs(1100) <= 1'b1;
    layer1_outputs(1101) <= a or b;
    layer1_outputs(1102) <= b and not a;
    layer1_outputs(1103) <= not (a or b);
    layer1_outputs(1104) <= a xor b;
    layer1_outputs(1105) <= 1'b0;
    layer1_outputs(1106) <= a and not b;
    layer1_outputs(1107) <= not b;
    layer1_outputs(1108) <= not (a or b);
    layer1_outputs(1109) <= 1'b0;
    layer1_outputs(1110) <= a and b;
    layer1_outputs(1111) <= 1'b0;
    layer1_outputs(1112) <= not a or b;
    layer1_outputs(1113) <= 1'b0;
    layer1_outputs(1114) <= not (a or b);
    layer1_outputs(1115) <= a or b;
    layer1_outputs(1116) <= not a or b;
    layer1_outputs(1117) <= not (a and b);
    layer1_outputs(1118) <= a xor b;
    layer1_outputs(1119) <= b;
    layer1_outputs(1120) <= a and b;
    layer1_outputs(1121) <= not (a or b);
    layer1_outputs(1122) <= 1'b1;
    layer1_outputs(1123) <= not a or b;
    layer1_outputs(1124) <= a xor b;
    layer1_outputs(1125) <= not a or b;
    layer1_outputs(1126) <= a;
    layer1_outputs(1127) <= b and not a;
    layer1_outputs(1128) <= not b or a;
    layer1_outputs(1129) <= not (a and b);
    layer1_outputs(1130) <= a;
    layer1_outputs(1131) <= not (a or b);
    layer1_outputs(1132) <= a and b;
    layer1_outputs(1133) <= a and not b;
    layer1_outputs(1134) <= not (a and b);
    layer1_outputs(1135) <= b and not a;
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= not a;
    layer1_outputs(1138) <= 1'b0;
    layer1_outputs(1139) <= b;
    layer1_outputs(1140) <= b and not a;
    layer1_outputs(1141) <= not (a and b);
    layer1_outputs(1142) <= not b;
    layer1_outputs(1143) <= a and not b;
    layer1_outputs(1144) <= a and b;
    layer1_outputs(1145) <= 1'b1;
    layer1_outputs(1146) <= a and b;
    layer1_outputs(1147) <= not (a and b);
    layer1_outputs(1148) <= not (a and b);
    layer1_outputs(1149) <= not (a or b);
    layer1_outputs(1150) <= b;
    layer1_outputs(1151) <= a and not b;
    layer1_outputs(1152) <= 1'b1;
    layer1_outputs(1153) <= not b;
    layer1_outputs(1154) <= a and not b;
    layer1_outputs(1155) <= 1'b1;
    layer1_outputs(1156) <= not b or a;
    layer1_outputs(1157) <= not (a xor b);
    layer1_outputs(1158) <= a and not b;
    layer1_outputs(1159) <= a or b;
    layer1_outputs(1160) <= a;
    layer1_outputs(1161) <= 1'b1;
    layer1_outputs(1162) <= 1'b1;
    layer1_outputs(1163) <= not (a or b);
    layer1_outputs(1164) <= 1'b1;
    layer1_outputs(1165) <= 1'b0;
    layer1_outputs(1166) <= a;
    layer1_outputs(1167) <= a;
    layer1_outputs(1168) <= a;
    layer1_outputs(1169) <= a and not b;
    layer1_outputs(1170) <= not a or b;
    layer1_outputs(1171) <= not (a xor b);
    layer1_outputs(1172) <= not a or b;
    layer1_outputs(1173) <= not a;
    layer1_outputs(1174) <= b;
    layer1_outputs(1175) <= a xor b;
    layer1_outputs(1176) <= not (a or b);
    layer1_outputs(1177) <= not (a and b);
    layer1_outputs(1178) <= not a;
    layer1_outputs(1179) <= a and b;
    layer1_outputs(1180) <= not (a and b);
    layer1_outputs(1181) <= a;
    layer1_outputs(1182) <= a xor b;
    layer1_outputs(1183) <= a or b;
    layer1_outputs(1184) <= 1'b1;
    layer1_outputs(1185) <= not b;
    layer1_outputs(1186) <= 1'b1;
    layer1_outputs(1187) <= not (a xor b);
    layer1_outputs(1188) <= a;
    layer1_outputs(1189) <= not b or a;
    layer1_outputs(1190) <= 1'b1;
    layer1_outputs(1191) <= b;
    layer1_outputs(1192) <= b;
    layer1_outputs(1193) <= 1'b0;
    layer1_outputs(1194) <= a;
    layer1_outputs(1195) <= not (a or b);
    layer1_outputs(1196) <= not b;
    layer1_outputs(1197) <= 1'b1;
    layer1_outputs(1198) <= b;
    layer1_outputs(1199) <= b and not a;
    layer1_outputs(1200) <= a;
    layer1_outputs(1201) <= not b or a;
    layer1_outputs(1202) <= a;
    layer1_outputs(1203) <= a and not b;
    layer1_outputs(1204) <= a and b;
    layer1_outputs(1205) <= 1'b0;
    layer1_outputs(1206) <= b;
    layer1_outputs(1207) <= not a;
    layer1_outputs(1208) <= not (a and b);
    layer1_outputs(1209) <= a xor b;
    layer1_outputs(1210) <= not a;
    layer1_outputs(1211) <= not a or b;
    layer1_outputs(1212) <= a and b;
    layer1_outputs(1213) <= 1'b0;
    layer1_outputs(1214) <= b and not a;
    layer1_outputs(1215) <= a;
    layer1_outputs(1216) <= not (a or b);
    layer1_outputs(1217) <= not (a xor b);
    layer1_outputs(1218) <= not b or a;
    layer1_outputs(1219) <= 1'b0;
    layer1_outputs(1220) <= a;
    layer1_outputs(1221) <= b;
    layer1_outputs(1222) <= a and not b;
    layer1_outputs(1223) <= 1'b1;
    layer1_outputs(1224) <= 1'b1;
    layer1_outputs(1225) <= not a;
    layer1_outputs(1226) <= not a;
    layer1_outputs(1227) <= not (a and b);
    layer1_outputs(1228) <= a;
    layer1_outputs(1229) <= 1'b1;
    layer1_outputs(1230) <= not b;
    layer1_outputs(1231) <= a or b;
    layer1_outputs(1232) <= not b or a;
    layer1_outputs(1233) <= 1'b0;
    layer1_outputs(1234) <= not b;
    layer1_outputs(1235) <= a and not b;
    layer1_outputs(1236) <= a and not b;
    layer1_outputs(1237) <= a xor b;
    layer1_outputs(1238) <= a;
    layer1_outputs(1239) <= a and b;
    layer1_outputs(1240) <= not a or b;
    layer1_outputs(1241) <= not a or b;
    layer1_outputs(1242) <= not (a or b);
    layer1_outputs(1243) <= not (a or b);
    layer1_outputs(1244) <= not b or a;
    layer1_outputs(1245) <= a and b;
    layer1_outputs(1246) <= not (a xor b);
    layer1_outputs(1247) <= a and not b;
    layer1_outputs(1248) <= not (a or b);
    layer1_outputs(1249) <= not a;
    layer1_outputs(1250) <= not b;
    layer1_outputs(1251) <= a;
    layer1_outputs(1252) <= not b;
    layer1_outputs(1253) <= b and not a;
    layer1_outputs(1254) <= b and not a;
    layer1_outputs(1255) <= b and not a;
    layer1_outputs(1256) <= a and b;
    layer1_outputs(1257) <= not a or b;
    layer1_outputs(1258) <= not (a xor b);
    layer1_outputs(1259) <= 1'b0;
    layer1_outputs(1260) <= not (a xor b);
    layer1_outputs(1261) <= a and b;
    layer1_outputs(1262) <= not (a and b);
    layer1_outputs(1263) <= not (a or b);
    layer1_outputs(1264) <= 1'b0;
    layer1_outputs(1265) <= a and b;
    layer1_outputs(1266) <= not a or b;
    layer1_outputs(1267) <= a and not b;
    layer1_outputs(1268) <= 1'b0;
    layer1_outputs(1269) <= a and b;
    layer1_outputs(1270) <= not a;
    layer1_outputs(1271) <= not a;
    layer1_outputs(1272) <= not (a and b);
    layer1_outputs(1273) <= 1'b0;
    layer1_outputs(1274) <= a;
    layer1_outputs(1275) <= not (a or b);
    layer1_outputs(1276) <= a;
    layer1_outputs(1277) <= not a or b;
    layer1_outputs(1278) <= not (a xor b);
    layer1_outputs(1279) <= not b or a;
    layer1_outputs(1280) <= b;
    layer1_outputs(1281) <= 1'b0;
    layer1_outputs(1282) <= not a or b;
    layer1_outputs(1283) <= not (a or b);
    layer1_outputs(1284) <= a;
    layer1_outputs(1285) <= a or b;
    layer1_outputs(1286) <= a and not b;
    layer1_outputs(1287) <= not (a xor b);
    layer1_outputs(1288) <= not (a or b);
    layer1_outputs(1289) <= a;
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= not b or a;
    layer1_outputs(1292) <= a and not b;
    layer1_outputs(1293) <= b;
    layer1_outputs(1294) <= 1'b1;
    layer1_outputs(1295) <= not (a or b);
    layer1_outputs(1296) <= a and not b;
    layer1_outputs(1297) <= not b;
    layer1_outputs(1298) <= not a;
    layer1_outputs(1299) <= a;
    layer1_outputs(1300) <= 1'b0;
    layer1_outputs(1301) <= not b;
    layer1_outputs(1302) <= a and b;
    layer1_outputs(1303) <= not b;
    layer1_outputs(1304) <= b and not a;
    layer1_outputs(1305) <= 1'b0;
    layer1_outputs(1306) <= not a or b;
    layer1_outputs(1307) <= not (a xor b);
    layer1_outputs(1308) <= not a or b;
    layer1_outputs(1309) <= not b;
    layer1_outputs(1310) <= 1'b0;
    layer1_outputs(1311) <= a or b;
    layer1_outputs(1312) <= not (a or b);
    layer1_outputs(1313) <= 1'b0;
    layer1_outputs(1314) <= not (a and b);
    layer1_outputs(1315) <= b;
    layer1_outputs(1316) <= a or b;
    layer1_outputs(1317) <= not (a or b);
    layer1_outputs(1318) <= a and not b;
    layer1_outputs(1319) <= b and not a;
    layer1_outputs(1320) <= 1'b1;
    layer1_outputs(1321) <= b and not a;
    layer1_outputs(1322) <= not (a and b);
    layer1_outputs(1323) <= 1'b0;
    layer1_outputs(1324) <= 1'b1;
    layer1_outputs(1325) <= not b;
    layer1_outputs(1326) <= not (a or b);
    layer1_outputs(1327) <= 1'b1;
    layer1_outputs(1328) <= b and not a;
    layer1_outputs(1329) <= 1'b1;
    layer1_outputs(1330) <= not (a xor b);
    layer1_outputs(1331) <= not a;
    layer1_outputs(1332) <= a xor b;
    layer1_outputs(1333) <= a;
    layer1_outputs(1334) <= b;
    layer1_outputs(1335) <= a or b;
    layer1_outputs(1336) <= not (a or b);
    layer1_outputs(1337) <= a or b;
    layer1_outputs(1338) <= 1'b1;
    layer1_outputs(1339) <= b;
    layer1_outputs(1340) <= not b;
    layer1_outputs(1341) <= not (a xor b);
    layer1_outputs(1342) <= a and not b;
    layer1_outputs(1343) <= not (a or b);
    layer1_outputs(1344) <= not (a or b);
    layer1_outputs(1345) <= b;
    layer1_outputs(1346) <= not b;
    layer1_outputs(1347) <= a or b;
    layer1_outputs(1348) <= not a;
    layer1_outputs(1349) <= a or b;
    layer1_outputs(1350) <= b and not a;
    layer1_outputs(1351) <= not (a and b);
    layer1_outputs(1352) <= not (a or b);
    layer1_outputs(1353) <= not a or b;
    layer1_outputs(1354) <= not b;
    layer1_outputs(1355) <= not a or b;
    layer1_outputs(1356) <= 1'b0;
    layer1_outputs(1357) <= b and not a;
    layer1_outputs(1358) <= 1'b0;
    layer1_outputs(1359) <= a xor b;
    layer1_outputs(1360) <= not (a and b);
    layer1_outputs(1361) <= a and not b;
    layer1_outputs(1362) <= 1'b0;
    layer1_outputs(1363) <= a or b;
    layer1_outputs(1364) <= not (a or b);
    layer1_outputs(1365) <= not (a xor b);
    layer1_outputs(1366) <= a and b;
    layer1_outputs(1367) <= not a or b;
    layer1_outputs(1368) <= 1'b1;
    layer1_outputs(1369) <= 1'b0;
    layer1_outputs(1370) <= a or b;
    layer1_outputs(1371) <= not (a xor b);
    layer1_outputs(1372) <= b and not a;
    layer1_outputs(1373) <= b and not a;
    layer1_outputs(1374) <= not b;
    layer1_outputs(1375) <= a or b;
    layer1_outputs(1376) <= 1'b1;
    layer1_outputs(1377) <= not b or a;
    layer1_outputs(1378) <= a and b;
    layer1_outputs(1379) <= not (a and b);
    layer1_outputs(1380) <= b and not a;
    layer1_outputs(1381) <= 1'b0;
    layer1_outputs(1382) <= not (a and b);
    layer1_outputs(1383) <= not a or b;
    layer1_outputs(1384) <= not b or a;
    layer1_outputs(1385) <= a;
    layer1_outputs(1386) <= not a or b;
    layer1_outputs(1387) <= 1'b1;
    layer1_outputs(1388) <= a and not b;
    layer1_outputs(1389) <= a and b;
    layer1_outputs(1390) <= not (a and b);
    layer1_outputs(1391) <= not (a and b);
    layer1_outputs(1392) <= a or b;
    layer1_outputs(1393) <= a xor b;
    layer1_outputs(1394) <= 1'b0;
    layer1_outputs(1395) <= 1'b0;
    layer1_outputs(1396) <= not (a or b);
    layer1_outputs(1397) <= 1'b0;
    layer1_outputs(1398) <= 1'b1;
    layer1_outputs(1399) <= a and b;
    layer1_outputs(1400) <= not (a or b);
    layer1_outputs(1401) <= 1'b0;
    layer1_outputs(1402) <= not a or b;
    layer1_outputs(1403) <= 1'b0;
    layer1_outputs(1404) <= not (a xor b);
    layer1_outputs(1405) <= a and not b;
    layer1_outputs(1406) <= 1'b0;
    layer1_outputs(1407) <= a and b;
    layer1_outputs(1408) <= not a or b;
    layer1_outputs(1409) <= a and not b;
    layer1_outputs(1410) <= b and not a;
    layer1_outputs(1411) <= a and not b;
    layer1_outputs(1412) <= not a;
    layer1_outputs(1413) <= not a;
    layer1_outputs(1414) <= 1'b1;
    layer1_outputs(1415) <= 1'b1;
    layer1_outputs(1416) <= not a or b;
    layer1_outputs(1417) <= 1'b0;
    layer1_outputs(1418) <= not a;
    layer1_outputs(1419) <= b;
    layer1_outputs(1420) <= not b or a;
    layer1_outputs(1421) <= 1'b0;
    layer1_outputs(1422) <= b;
    layer1_outputs(1423) <= a and b;
    layer1_outputs(1424) <= a and not b;
    layer1_outputs(1425) <= not (a and b);
    layer1_outputs(1426) <= not (a or b);
    layer1_outputs(1427) <= 1'b1;
    layer1_outputs(1428) <= not a or b;
    layer1_outputs(1429) <= not a;
    layer1_outputs(1430) <= not b or a;
    layer1_outputs(1431) <= a;
    layer1_outputs(1432) <= not (a or b);
    layer1_outputs(1433) <= not b;
    layer1_outputs(1434) <= a and b;
    layer1_outputs(1435) <= b;
    layer1_outputs(1436) <= not (a xor b);
    layer1_outputs(1437) <= not b;
    layer1_outputs(1438) <= not (a and b);
    layer1_outputs(1439) <= b;
    layer1_outputs(1440) <= not (a xor b);
    layer1_outputs(1441) <= a and b;
    layer1_outputs(1442) <= not (a and b);
    layer1_outputs(1443) <= a xor b;
    layer1_outputs(1444) <= a or b;
    layer1_outputs(1445) <= a;
    layer1_outputs(1446) <= not a;
    layer1_outputs(1447) <= 1'b0;
    layer1_outputs(1448) <= a or b;
    layer1_outputs(1449) <= a;
    layer1_outputs(1450) <= not a or b;
    layer1_outputs(1451) <= a and not b;
    layer1_outputs(1452) <= b;
    layer1_outputs(1453) <= 1'b0;
    layer1_outputs(1454) <= a and b;
    layer1_outputs(1455) <= not (a or b);
    layer1_outputs(1456) <= b;
    layer1_outputs(1457) <= a xor b;
    layer1_outputs(1458) <= 1'b1;
    layer1_outputs(1459) <= a or b;
    layer1_outputs(1460) <= 1'b1;
    layer1_outputs(1461) <= not (a or b);
    layer1_outputs(1462) <= b;
    layer1_outputs(1463) <= not (a and b);
    layer1_outputs(1464) <= b and not a;
    layer1_outputs(1465) <= not (a or b);
    layer1_outputs(1466) <= not b;
    layer1_outputs(1467) <= not b or a;
    layer1_outputs(1468) <= 1'b1;
    layer1_outputs(1469) <= not b or a;
    layer1_outputs(1470) <= a or b;
    layer1_outputs(1471) <= b and not a;
    layer1_outputs(1472) <= b and not a;
    layer1_outputs(1473) <= a;
    layer1_outputs(1474) <= a and not b;
    layer1_outputs(1475) <= not b or a;
    layer1_outputs(1476) <= a and not b;
    layer1_outputs(1477) <= not (a or b);
    layer1_outputs(1478) <= 1'b1;
    layer1_outputs(1479) <= b;
    layer1_outputs(1480) <= a and b;
    layer1_outputs(1481) <= b and not a;
    layer1_outputs(1482) <= a or b;
    layer1_outputs(1483) <= a and b;
    layer1_outputs(1484) <= a or b;
    layer1_outputs(1485) <= a;
    layer1_outputs(1486) <= not (a and b);
    layer1_outputs(1487) <= not (a or b);
    layer1_outputs(1488) <= not a or b;
    layer1_outputs(1489) <= not (a or b);
    layer1_outputs(1490) <= a and not b;
    layer1_outputs(1491) <= 1'b0;
    layer1_outputs(1492) <= not a;
    layer1_outputs(1493) <= b;
    layer1_outputs(1494) <= a and not b;
    layer1_outputs(1495) <= not a or b;
    layer1_outputs(1496) <= not (a or b);
    layer1_outputs(1497) <= b and not a;
    layer1_outputs(1498) <= not (a or b);
    layer1_outputs(1499) <= not (a xor b);
    layer1_outputs(1500) <= a and b;
    layer1_outputs(1501) <= 1'b0;
    layer1_outputs(1502) <= 1'b1;
    layer1_outputs(1503) <= a and not b;
    layer1_outputs(1504) <= not a;
    layer1_outputs(1505) <= b;
    layer1_outputs(1506) <= a and b;
    layer1_outputs(1507) <= not (a and b);
    layer1_outputs(1508) <= not b or a;
    layer1_outputs(1509) <= b;
    layer1_outputs(1510) <= 1'b0;
    layer1_outputs(1511) <= 1'b1;
    layer1_outputs(1512) <= a xor b;
    layer1_outputs(1513) <= b;
    layer1_outputs(1514) <= a xor b;
    layer1_outputs(1515) <= a and b;
    layer1_outputs(1516) <= not b;
    layer1_outputs(1517) <= 1'b1;
    layer1_outputs(1518) <= not b or a;
    layer1_outputs(1519) <= 1'b1;
    layer1_outputs(1520) <= 1'b0;
    layer1_outputs(1521) <= a and not b;
    layer1_outputs(1522) <= a and b;
    layer1_outputs(1523) <= not (a and b);
    layer1_outputs(1524) <= b and not a;
    layer1_outputs(1525) <= 1'b0;
    layer1_outputs(1526) <= 1'b0;
    layer1_outputs(1527) <= a or b;
    layer1_outputs(1528) <= not (a or b);
    layer1_outputs(1529) <= a xor b;
    layer1_outputs(1530) <= not (a and b);
    layer1_outputs(1531) <= not (a or b);
    layer1_outputs(1532) <= not a;
    layer1_outputs(1533) <= 1'b1;
    layer1_outputs(1534) <= a and not b;
    layer1_outputs(1535) <= a;
    layer1_outputs(1536) <= not a or b;
    layer1_outputs(1537) <= not b or a;
    layer1_outputs(1538) <= a and b;
    layer1_outputs(1539) <= a and not b;
    layer1_outputs(1540) <= 1'b0;
    layer1_outputs(1541) <= not (a and b);
    layer1_outputs(1542) <= a or b;
    layer1_outputs(1543) <= not a;
    layer1_outputs(1544) <= 1'b1;
    layer1_outputs(1545) <= a and not b;
    layer1_outputs(1546) <= 1'b0;
    layer1_outputs(1547) <= 1'b0;
    layer1_outputs(1548) <= not (a and b);
    layer1_outputs(1549) <= 1'b1;
    layer1_outputs(1550) <= b;
    layer1_outputs(1551) <= a and b;
    layer1_outputs(1552) <= b;
    layer1_outputs(1553) <= 1'b1;
    layer1_outputs(1554) <= 1'b0;
    layer1_outputs(1555) <= a and b;
    layer1_outputs(1556) <= a or b;
    layer1_outputs(1557) <= a and not b;
    layer1_outputs(1558) <= a and not b;
    layer1_outputs(1559) <= not (a or b);
    layer1_outputs(1560) <= not b;
    layer1_outputs(1561) <= not b;
    layer1_outputs(1562) <= 1'b1;
    layer1_outputs(1563) <= not (a xor b);
    layer1_outputs(1564) <= a and not b;
    layer1_outputs(1565) <= not b or a;
    layer1_outputs(1566) <= not (a or b);
    layer1_outputs(1567) <= 1'b0;
    layer1_outputs(1568) <= a or b;
    layer1_outputs(1569) <= not b or a;
    layer1_outputs(1570) <= 1'b0;
    layer1_outputs(1571) <= a or b;
    layer1_outputs(1572) <= a or b;
    layer1_outputs(1573) <= a and not b;
    layer1_outputs(1574) <= not b;
    layer1_outputs(1575) <= not (a xor b);
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= 1'b0;
    layer1_outputs(1578) <= b;
    layer1_outputs(1579) <= b and not a;
    layer1_outputs(1580) <= not b;
    layer1_outputs(1581) <= 1'b1;
    layer1_outputs(1582) <= 1'b0;
    layer1_outputs(1583) <= not a or b;
    layer1_outputs(1584) <= not b;
    layer1_outputs(1585) <= not b;
    layer1_outputs(1586) <= a and b;
    layer1_outputs(1587) <= a and not b;
    layer1_outputs(1588) <= not (a and b);
    layer1_outputs(1589) <= not a;
    layer1_outputs(1590) <= not b;
    layer1_outputs(1591) <= a;
    layer1_outputs(1592) <= a xor b;
    layer1_outputs(1593) <= a and not b;
    layer1_outputs(1594) <= b;
    layer1_outputs(1595) <= b;
    layer1_outputs(1596) <= a and not b;
    layer1_outputs(1597) <= a and not b;
    layer1_outputs(1598) <= not (a and b);
    layer1_outputs(1599) <= a and not b;
    layer1_outputs(1600) <= not (a and b);
    layer1_outputs(1601) <= not b or a;
    layer1_outputs(1602) <= b and not a;
    layer1_outputs(1603) <= not b or a;
    layer1_outputs(1604) <= 1'b0;
    layer1_outputs(1605) <= 1'b1;
    layer1_outputs(1606) <= a;
    layer1_outputs(1607) <= not b or a;
    layer1_outputs(1608) <= not (a or b);
    layer1_outputs(1609) <= b and not a;
    layer1_outputs(1610) <= not b or a;
    layer1_outputs(1611) <= 1'b1;
    layer1_outputs(1612) <= not b;
    layer1_outputs(1613) <= not b;
    layer1_outputs(1614) <= not (a and b);
    layer1_outputs(1615) <= not (a and b);
    layer1_outputs(1616) <= not a;
    layer1_outputs(1617) <= a or b;
    layer1_outputs(1618) <= 1'b0;
    layer1_outputs(1619) <= not (a or b);
    layer1_outputs(1620) <= 1'b0;
    layer1_outputs(1621) <= b and not a;
    layer1_outputs(1622) <= a and b;
    layer1_outputs(1623) <= a and b;
    layer1_outputs(1624) <= not a;
    layer1_outputs(1625) <= 1'b0;
    layer1_outputs(1626) <= a xor b;
    layer1_outputs(1627) <= not a or b;
    layer1_outputs(1628) <= not b;
    layer1_outputs(1629) <= not b or a;
    layer1_outputs(1630) <= a and not b;
    layer1_outputs(1631) <= a and not b;
    layer1_outputs(1632) <= 1'b1;
    layer1_outputs(1633) <= a or b;
    layer1_outputs(1634) <= a;
    layer1_outputs(1635) <= a or b;
    layer1_outputs(1636) <= not (a or b);
    layer1_outputs(1637) <= a and b;
    layer1_outputs(1638) <= not a or b;
    layer1_outputs(1639) <= not b;
    layer1_outputs(1640) <= b;
    layer1_outputs(1641) <= a or b;
    layer1_outputs(1642) <= a and not b;
    layer1_outputs(1643) <= a;
    layer1_outputs(1644) <= a and b;
    layer1_outputs(1645) <= 1'b0;
    layer1_outputs(1646) <= not (a or b);
    layer1_outputs(1647) <= a and not b;
    layer1_outputs(1648) <= 1'b1;
    layer1_outputs(1649) <= a;
    layer1_outputs(1650) <= not (a or b);
    layer1_outputs(1651) <= a;
    layer1_outputs(1652) <= 1'b1;
    layer1_outputs(1653) <= a xor b;
    layer1_outputs(1654) <= not a;
    layer1_outputs(1655) <= not (a and b);
    layer1_outputs(1656) <= b and not a;
    layer1_outputs(1657) <= a and not b;
    layer1_outputs(1658) <= 1'b1;
    layer1_outputs(1659) <= not a or b;
    layer1_outputs(1660) <= a;
    layer1_outputs(1661) <= not (a and b);
    layer1_outputs(1662) <= a;
    layer1_outputs(1663) <= not b;
    layer1_outputs(1664) <= a xor b;
    layer1_outputs(1665) <= not (a or b);
    layer1_outputs(1666) <= 1'b0;
    layer1_outputs(1667) <= a and not b;
    layer1_outputs(1668) <= b and not a;
    layer1_outputs(1669) <= not (a and b);
    layer1_outputs(1670) <= not b;
    layer1_outputs(1671) <= not b or a;
    layer1_outputs(1672) <= b;
    layer1_outputs(1673) <= not b;
    layer1_outputs(1674) <= not b;
    layer1_outputs(1675) <= b;
    layer1_outputs(1676) <= 1'b1;
    layer1_outputs(1677) <= a and b;
    layer1_outputs(1678) <= 1'b0;
    layer1_outputs(1679) <= b and not a;
    layer1_outputs(1680) <= a;
    layer1_outputs(1681) <= a and b;
    layer1_outputs(1682) <= a or b;
    layer1_outputs(1683) <= b and not a;
    layer1_outputs(1684) <= 1'b0;
    layer1_outputs(1685) <= not b;
    layer1_outputs(1686) <= 1'b1;
    layer1_outputs(1687) <= a or b;
    layer1_outputs(1688) <= not (a or b);
    layer1_outputs(1689) <= not a;
    layer1_outputs(1690) <= not (a or b);
    layer1_outputs(1691) <= not b;
    layer1_outputs(1692) <= not a;
    layer1_outputs(1693) <= b;
    layer1_outputs(1694) <= a and b;
    layer1_outputs(1695) <= a;
    layer1_outputs(1696) <= a or b;
    layer1_outputs(1697) <= b;
    layer1_outputs(1698) <= a or b;
    layer1_outputs(1699) <= not b;
    layer1_outputs(1700) <= not b or a;
    layer1_outputs(1701) <= a or b;
    layer1_outputs(1702) <= b and not a;
    layer1_outputs(1703) <= b;
    layer1_outputs(1704) <= not (a and b);
    layer1_outputs(1705) <= not a or b;
    layer1_outputs(1706) <= not (a and b);
    layer1_outputs(1707) <= not a or b;
    layer1_outputs(1708) <= not b or a;
    layer1_outputs(1709) <= a or b;
    layer1_outputs(1710) <= a and not b;
    layer1_outputs(1711) <= 1'b0;
    layer1_outputs(1712) <= a;
    layer1_outputs(1713) <= not b;
    layer1_outputs(1714) <= a and not b;
    layer1_outputs(1715) <= a and b;
    layer1_outputs(1716) <= 1'b1;
    layer1_outputs(1717) <= b;
    layer1_outputs(1718) <= not a;
    layer1_outputs(1719) <= not (a xor b);
    layer1_outputs(1720) <= not b;
    layer1_outputs(1721) <= a and not b;
    layer1_outputs(1722) <= a;
    layer1_outputs(1723) <= a and not b;
    layer1_outputs(1724) <= not a;
    layer1_outputs(1725) <= 1'b0;
    layer1_outputs(1726) <= 1'b1;
    layer1_outputs(1727) <= not b;
    layer1_outputs(1728) <= b and not a;
    layer1_outputs(1729) <= a or b;
    layer1_outputs(1730) <= 1'b0;
    layer1_outputs(1731) <= 1'b0;
    layer1_outputs(1732) <= not b;
    layer1_outputs(1733) <= a xor b;
    layer1_outputs(1734) <= not a;
    layer1_outputs(1735) <= not (a xor b);
    layer1_outputs(1736) <= not b or a;
    layer1_outputs(1737) <= a and not b;
    layer1_outputs(1738) <= not (a or b);
    layer1_outputs(1739) <= not b or a;
    layer1_outputs(1740) <= b;
    layer1_outputs(1741) <= b;
    layer1_outputs(1742) <= 1'b1;
    layer1_outputs(1743) <= a or b;
    layer1_outputs(1744) <= not b;
    layer1_outputs(1745) <= a and b;
    layer1_outputs(1746) <= 1'b1;
    layer1_outputs(1747) <= not b;
    layer1_outputs(1748) <= a;
    layer1_outputs(1749) <= 1'b1;
    layer1_outputs(1750) <= 1'b1;
    layer1_outputs(1751) <= not b or a;
    layer1_outputs(1752) <= not a;
    layer1_outputs(1753) <= not a or b;
    layer1_outputs(1754) <= not (a and b);
    layer1_outputs(1755) <= b and not a;
    layer1_outputs(1756) <= a xor b;
    layer1_outputs(1757) <= a or b;
    layer1_outputs(1758) <= 1'b0;
    layer1_outputs(1759) <= b and not a;
    layer1_outputs(1760) <= b and not a;
    layer1_outputs(1761) <= a and b;
    layer1_outputs(1762) <= a and b;
    layer1_outputs(1763) <= a and b;
    layer1_outputs(1764) <= not (a and b);
    layer1_outputs(1765) <= not (a and b);
    layer1_outputs(1766) <= a or b;
    layer1_outputs(1767) <= not b or a;
    layer1_outputs(1768) <= a xor b;
    layer1_outputs(1769) <= a and b;
    layer1_outputs(1770) <= not b or a;
    layer1_outputs(1771) <= not (a xor b);
    layer1_outputs(1772) <= not (a and b);
    layer1_outputs(1773) <= not (a or b);
    layer1_outputs(1774) <= b and not a;
    layer1_outputs(1775) <= a or b;
    layer1_outputs(1776) <= not (a or b);
    layer1_outputs(1777) <= not (a or b);
    layer1_outputs(1778) <= not a;
    layer1_outputs(1779) <= 1'b1;
    layer1_outputs(1780) <= b;
    layer1_outputs(1781) <= not (a and b);
    layer1_outputs(1782) <= b and not a;
    layer1_outputs(1783) <= b;
    layer1_outputs(1784) <= not b or a;
    layer1_outputs(1785) <= 1'b0;
    layer1_outputs(1786) <= not (a xor b);
    layer1_outputs(1787) <= not b or a;
    layer1_outputs(1788) <= b and not a;
    layer1_outputs(1789) <= 1'b1;
    layer1_outputs(1790) <= a and not b;
    layer1_outputs(1791) <= 1'b1;
    layer1_outputs(1792) <= not a or b;
    layer1_outputs(1793) <= not a;
    layer1_outputs(1794) <= not b;
    layer1_outputs(1795) <= not (a and b);
    layer1_outputs(1796) <= a and not b;
    layer1_outputs(1797) <= a;
    layer1_outputs(1798) <= b and not a;
    layer1_outputs(1799) <= 1'b0;
    layer1_outputs(1800) <= b and not a;
    layer1_outputs(1801) <= not (a and b);
    layer1_outputs(1802) <= b and not a;
    layer1_outputs(1803) <= a and not b;
    layer1_outputs(1804) <= not (a or b);
    layer1_outputs(1805) <= a xor b;
    layer1_outputs(1806) <= not b;
    layer1_outputs(1807) <= not (a and b);
    layer1_outputs(1808) <= a or b;
    layer1_outputs(1809) <= not a or b;
    layer1_outputs(1810) <= 1'b0;
    layer1_outputs(1811) <= 1'b0;
    layer1_outputs(1812) <= a or b;
    layer1_outputs(1813) <= not (a and b);
    layer1_outputs(1814) <= b;
    layer1_outputs(1815) <= 1'b1;
    layer1_outputs(1816) <= b;
    layer1_outputs(1817) <= not (a and b);
    layer1_outputs(1818) <= b;
    layer1_outputs(1819) <= not (a and b);
    layer1_outputs(1820) <= a or b;
    layer1_outputs(1821) <= not (a or b);
    layer1_outputs(1822) <= not (a or b);
    layer1_outputs(1823) <= 1'b1;
    layer1_outputs(1824) <= a;
    layer1_outputs(1825) <= b;
    layer1_outputs(1826) <= a and not b;
    layer1_outputs(1827) <= not (a or b);
    layer1_outputs(1828) <= not b;
    layer1_outputs(1829) <= not a or b;
    layer1_outputs(1830) <= not (a and b);
    layer1_outputs(1831) <= a;
    layer1_outputs(1832) <= 1'b0;
    layer1_outputs(1833) <= a or b;
    layer1_outputs(1834) <= not (a or b);
    layer1_outputs(1835) <= a and not b;
    layer1_outputs(1836) <= a and not b;
    layer1_outputs(1837) <= 1'b1;
    layer1_outputs(1838) <= a;
    layer1_outputs(1839) <= b and not a;
    layer1_outputs(1840) <= a and b;
    layer1_outputs(1841) <= not b or a;
    layer1_outputs(1842) <= a;
    layer1_outputs(1843) <= not (a or b);
    layer1_outputs(1844) <= a and not b;
    layer1_outputs(1845) <= b;
    layer1_outputs(1846) <= a;
    layer1_outputs(1847) <= not (a or b);
    layer1_outputs(1848) <= 1'b0;
    layer1_outputs(1849) <= 1'b1;
    layer1_outputs(1850) <= a;
    layer1_outputs(1851) <= a and b;
    layer1_outputs(1852) <= not b or a;
    layer1_outputs(1853) <= a;
    layer1_outputs(1854) <= b;
    layer1_outputs(1855) <= a xor b;
    layer1_outputs(1856) <= not (a or b);
    layer1_outputs(1857) <= a;
    layer1_outputs(1858) <= b;
    layer1_outputs(1859) <= b and not a;
    layer1_outputs(1860) <= a and not b;
    layer1_outputs(1861) <= b;
    layer1_outputs(1862) <= not a;
    layer1_outputs(1863) <= b;
    layer1_outputs(1864) <= b and not a;
    layer1_outputs(1865) <= a and b;
    layer1_outputs(1866) <= b;
    layer1_outputs(1867) <= 1'b1;
    layer1_outputs(1868) <= not a or b;
    layer1_outputs(1869) <= not (a and b);
    layer1_outputs(1870) <= 1'b1;
    layer1_outputs(1871) <= not a;
    layer1_outputs(1872) <= a;
    layer1_outputs(1873) <= 1'b0;
    layer1_outputs(1874) <= a or b;
    layer1_outputs(1875) <= not (a xor b);
    layer1_outputs(1876) <= 1'b1;
    layer1_outputs(1877) <= not a;
    layer1_outputs(1878) <= a and not b;
    layer1_outputs(1879) <= not (a or b);
    layer1_outputs(1880) <= b and not a;
    layer1_outputs(1881) <= not b;
    layer1_outputs(1882) <= a and b;
    layer1_outputs(1883) <= a and not b;
    layer1_outputs(1884) <= not (a or b);
    layer1_outputs(1885) <= a xor b;
    layer1_outputs(1886) <= not a;
    layer1_outputs(1887) <= not b;
    layer1_outputs(1888) <= not b;
    layer1_outputs(1889) <= b and not a;
    layer1_outputs(1890) <= a or b;
    layer1_outputs(1891) <= not a or b;
    layer1_outputs(1892) <= 1'b0;
    layer1_outputs(1893) <= not b or a;
    layer1_outputs(1894) <= not (a and b);
    layer1_outputs(1895) <= 1'b0;
    layer1_outputs(1896) <= a;
    layer1_outputs(1897) <= a and b;
    layer1_outputs(1898) <= not b or a;
    layer1_outputs(1899) <= a and not b;
    layer1_outputs(1900) <= a and b;
    layer1_outputs(1901) <= b and not a;
    layer1_outputs(1902) <= not (a xor b);
    layer1_outputs(1903) <= a xor b;
    layer1_outputs(1904) <= b;
    layer1_outputs(1905) <= 1'b0;
    layer1_outputs(1906) <= 1'b0;
    layer1_outputs(1907) <= a or b;
    layer1_outputs(1908) <= not a or b;
    layer1_outputs(1909) <= 1'b0;
    layer1_outputs(1910) <= 1'b0;
    layer1_outputs(1911) <= 1'b0;
    layer1_outputs(1912) <= not b or a;
    layer1_outputs(1913) <= not a or b;
    layer1_outputs(1914) <= a;
    layer1_outputs(1915) <= a and not b;
    layer1_outputs(1916) <= not (a or b);
    layer1_outputs(1917) <= a;
    layer1_outputs(1918) <= 1'b0;
    layer1_outputs(1919) <= 1'b0;
    layer1_outputs(1920) <= not a;
    layer1_outputs(1921) <= not b or a;
    layer1_outputs(1922) <= 1'b0;
    layer1_outputs(1923) <= not b;
    layer1_outputs(1924) <= b;
    layer1_outputs(1925) <= b;
    layer1_outputs(1926) <= b and not a;
    layer1_outputs(1927) <= a or b;
    layer1_outputs(1928) <= a and not b;
    layer1_outputs(1929) <= not a or b;
    layer1_outputs(1930) <= a and not b;
    layer1_outputs(1931) <= a and not b;
    layer1_outputs(1932) <= a xor b;
    layer1_outputs(1933) <= a or b;
    layer1_outputs(1934) <= a;
    layer1_outputs(1935) <= not (a or b);
    layer1_outputs(1936) <= not (a or b);
    layer1_outputs(1937) <= not a;
    layer1_outputs(1938) <= not (a or b);
    layer1_outputs(1939) <= 1'b1;
    layer1_outputs(1940) <= not b or a;
    layer1_outputs(1941) <= not b;
    layer1_outputs(1942) <= 1'b1;
    layer1_outputs(1943) <= b;
    layer1_outputs(1944) <= a and not b;
    layer1_outputs(1945) <= a;
    layer1_outputs(1946) <= not (a or b);
    layer1_outputs(1947) <= b;
    layer1_outputs(1948) <= a and not b;
    layer1_outputs(1949) <= not a or b;
    layer1_outputs(1950) <= a or b;
    layer1_outputs(1951) <= not a or b;
    layer1_outputs(1952) <= b and not a;
    layer1_outputs(1953) <= not (a or b);
    layer1_outputs(1954) <= 1'b0;
    layer1_outputs(1955) <= b and not a;
    layer1_outputs(1956) <= not b;
    layer1_outputs(1957) <= not (a or b);
    layer1_outputs(1958) <= not a;
    layer1_outputs(1959) <= 1'b0;
    layer1_outputs(1960) <= b;
    layer1_outputs(1961) <= not b;
    layer1_outputs(1962) <= not b or a;
    layer1_outputs(1963) <= a or b;
    layer1_outputs(1964) <= 1'b1;
    layer1_outputs(1965) <= not b;
    layer1_outputs(1966) <= a xor b;
    layer1_outputs(1967) <= 1'b1;
    layer1_outputs(1968) <= b;
    layer1_outputs(1969) <= b;
    layer1_outputs(1970) <= a and not b;
    layer1_outputs(1971) <= a or b;
    layer1_outputs(1972) <= not (a or b);
    layer1_outputs(1973) <= not (a xor b);
    layer1_outputs(1974) <= not a or b;
    layer1_outputs(1975) <= a xor b;
    layer1_outputs(1976) <= 1'b0;
    layer1_outputs(1977) <= not (a or b);
    layer1_outputs(1978) <= 1'b0;
    layer1_outputs(1979) <= a or b;
    layer1_outputs(1980) <= b;
    layer1_outputs(1981) <= a;
    layer1_outputs(1982) <= 1'b1;
    layer1_outputs(1983) <= b;
    layer1_outputs(1984) <= 1'b0;
    layer1_outputs(1985) <= not (a and b);
    layer1_outputs(1986) <= a or b;
    layer1_outputs(1987) <= not b;
    layer1_outputs(1988) <= not b or a;
    layer1_outputs(1989) <= not (a and b);
    layer1_outputs(1990) <= b and not a;
    layer1_outputs(1991) <= 1'b1;
    layer1_outputs(1992) <= not b or a;
    layer1_outputs(1993) <= not (a and b);
    layer1_outputs(1994) <= not a or b;
    layer1_outputs(1995) <= a and not b;
    layer1_outputs(1996) <= 1'b1;
    layer1_outputs(1997) <= a and b;
    layer1_outputs(1998) <= not b;
    layer1_outputs(1999) <= 1'b1;
    layer1_outputs(2000) <= 1'b1;
    layer1_outputs(2001) <= b and not a;
    layer1_outputs(2002) <= not (a xor b);
    layer1_outputs(2003) <= not (a or b);
    layer1_outputs(2004) <= 1'b0;
    layer1_outputs(2005) <= not b;
    layer1_outputs(2006) <= not a or b;
    layer1_outputs(2007) <= not a;
    layer1_outputs(2008) <= not b or a;
    layer1_outputs(2009) <= a and b;
    layer1_outputs(2010) <= b;
    layer1_outputs(2011) <= a and b;
    layer1_outputs(2012) <= 1'b0;
    layer1_outputs(2013) <= not a;
    layer1_outputs(2014) <= not (a xor b);
    layer1_outputs(2015) <= 1'b1;
    layer1_outputs(2016) <= b;
    layer1_outputs(2017) <= not (a xor b);
    layer1_outputs(2018) <= not a;
    layer1_outputs(2019) <= 1'b0;
    layer1_outputs(2020) <= not b;
    layer1_outputs(2021) <= not a;
    layer1_outputs(2022) <= not b;
    layer1_outputs(2023) <= not a or b;
    layer1_outputs(2024) <= a and b;
    layer1_outputs(2025) <= not a or b;
    layer1_outputs(2026) <= b and not a;
    layer1_outputs(2027) <= not (a or b);
    layer1_outputs(2028) <= 1'b1;
    layer1_outputs(2029) <= not a;
    layer1_outputs(2030) <= a and not b;
    layer1_outputs(2031) <= not b;
    layer1_outputs(2032) <= 1'b0;
    layer1_outputs(2033) <= a and b;
    layer1_outputs(2034) <= 1'b1;
    layer1_outputs(2035) <= a and not b;
    layer1_outputs(2036) <= not b or a;
    layer1_outputs(2037) <= a;
    layer1_outputs(2038) <= 1'b0;
    layer1_outputs(2039) <= not b or a;
    layer1_outputs(2040) <= a;
    layer1_outputs(2041) <= not b or a;
    layer1_outputs(2042) <= a or b;
    layer1_outputs(2043) <= 1'b1;
    layer1_outputs(2044) <= a and not b;
    layer1_outputs(2045) <= 1'b0;
    layer1_outputs(2046) <= 1'b0;
    layer1_outputs(2047) <= not a;
    layer1_outputs(2048) <= b;
    layer1_outputs(2049) <= not a;
    layer1_outputs(2050) <= b;
    layer1_outputs(2051) <= not (a and b);
    layer1_outputs(2052) <= a and b;
    layer1_outputs(2053) <= 1'b0;
    layer1_outputs(2054) <= a and not b;
    layer1_outputs(2055) <= b;
    layer1_outputs(2056) <= a or b;
    layer1_outputs(2057) <= not b;
    layer1_outputs(2058) <= 1'b1;
    layer1_outputs(2059) <= not b;
    layer1_outputs(2060) <= not a or b;
    layer1_outputs(2061) <= a;
    layer1_outputs(2062) <= b;
    layer1_outputs(2063) <= a;
    layer1_outputs(2064) <= 1'b1;
    layer1_outputs(2065) <= not a or b;
    layer1_outputs(2066) <= not b;
    layer1_outputs(2067) <= a;
    layer1_outputs(2068) <= b;
    layer1_outputs(2069) <= a and b;
    layer1_outputs(2070) <= a or b;
    layer1_outputs(2071) <= not (a or b);
    layer1_outputs(2072) <= 1'b1;
    layer1_outputs(2073) <= not (a or b);
    layer1_outputs(2074) <= a and b;
    layer1_outputs(2075) <= not b or a;
    layer1_outputs(2076) <= not a;
    layer1_outputs(2077) <= 1'b1;
    layer1_outputs(2078) <= a xor b;
    layer1_outputs(2079) <= a and not b;
    layer1_outputs(2080) <= not (a and b);
    layer1_outputs(2081) <= 1'b0;
    layer1_outputs(2082) <= not (a or b);
    layer1_outputs(2083) <= a and not b;
    layer1_outputs(2084) <= not a;
    layer1_outputs(2085) <= b;
    layer1_outputs(2086) <= not b or a;
    layer1_outputs(2087) <= not a;
    layer1_outputs(2088) <= not a;
    layer1_outputs(2089) <= 1'b1;
    layer1_outputs(2090) <= b and not a;
    layer1_outputs(2091) <= a;
    layer1_outputs(2092) <= not (a and b);
    layer1_outputs(2093) <= a;
    layer1_outputs(2094) <= not (a and b);
    layer1_outputs(2095) <= not (a or b);
    layer1_outputs(2096) <= 1'b0;
    layer1_outputs(2097) <= 1'b0;
    layer1_outputs(2098) <= not b or a;
    layer1_outputs(2099) <= not (a or b);
    layer1_outputs(2100) <= b;
    layer1_outputs(2101) <= not a;
    layer1_outputs(2102) <= a xor b;
    layer1_outputs(2103) <= not a or b;
    layer1_outputs(2104) <= 1'b0;
    layer1_outputs(2105) <= 1'b1;
    layer1_outputs(2106) <= not b;
    layer1_outputs(2107) <= a or b;
    layer1_outputs(2108) <= b;
    layer1_outputs(2109) <= not a;
    layer1_outputs(2110) <= not a or b;
    layer1_outputs(2111) <= 1'b1;
    layer1_outputs(2112) <= not b;
    layer1_outputs(2113) <= b and not a;
    layer1_outputs(2114) <= a or b;
    layer1_outputs(2115) <= a;
    layer1_outputs(2116) <= not a or b;
    layer1_outputs(2117) <= 1'b1;
    layer1_outputs(2118) <= not a;
    layer1_outputs(2119) <= a or b;
    layer1_outputs(2120) <= not a;
    layer1_outputs(2121) <= not b;
    layer1_outputs(2122) <= b and not a;
    layer1_outputs(2123) <= not a;
    layer1_outputs(2124) <= not (a and b);
    layer1_outputs(2125) <= not (a and b);
    layer1_outputs(2126) <= not a;
    layer1_outputs(2127) <= not b or a;
    layer1_outputs(2128) <= 1'b1;
    layer1_outputs(2129) <= b and not a;
    layer1_outputs(2130) <= a and not b;
    layer1_outputs(2131) <= not a or b;
    layer1_outputs(2132) <= not b or a;
    layer1_outputs(2133) <= b;
    layer1_outputs(2134) <= a or b;
    layer1_outputs(2135) <= not (a and b);
    layer1_outputs(2136) <= not (a or b);
    layer1_outputs(2137) <= not (a xor b);
    layer1_outputs(2138) <= not (a or b);
    layer1_outputs(2139) <= a;
    layer1_outputs(2140) <= a;
    layer1_outputs(2141) <= not (a and b);
    layer1_outputs(2142) <= b;
    layer1_outputs(2143) <= 1'b1;
    layer1_outputs(2144) <= a and b;
    layer1_outputs(2145) <= not a;
    layer1_outputs(2146) <= a and not b;
    layer1_outputs(2147) <= a or b;
    layer1_outputs(2148) <= a and not b;
    layer1_outputs(2149) <= not (a or b);
    layer1_outputs(2150) <= a and b;
    layer1_outputs(2151) <= a or b;
    layer1_outputs(2152) <= not b or a;
    layer1_outputs(2153) <= not (a xor b);
    layer1_outputs(2154) <= not (a and b);
    layer1_outputs(2155) <= not (a and b);
    layer1_outputs(2156) <= 1'b1;
    layer1_outputs(2157) <= a;
    layer1_outputs(2158) <= a xor b;
    layer1_outputs(2159) <= 1'b0;
    layer1_outputs(2160) <= not b;
    layer1_outputs(2161) <= not b;
    layer1_outputs(2162) <= a and not b;
    layer1_outputs(2163) <= 1'b1;
    layer1_outputs(2164) <= not a or b;
    layer1_outputs(2165) <= a xor b;
    layer1_outputs(2166) <= a and not b;
    layer1_outputs(2167) <= 1'b1;
    layer1_outputs(2168) <= b and not a;
    layer1_outputs(2169) <= a;
    layer1_outputs(2170) <= not b;
    layer1_outputs(2171) <= not (a xor b);
    layer1_outputs(2172) <= not a;
    layer1_outputs(2173) <= not b;
    layer1_outputs(2174) <= b;
    layer1_outputs(2175) <= a;
    layer1_outputs(2176) <= not (a and b);
    layer1_outputs(2177) <= a or b;
    layer1_outputs(2178) <= a xor b;
    layer1_outputs(2179) <= not (a or b);
    layer1_outputs(2180) <= a and not b;
    layer1_outputs(2181) <= a;
    layer1_outputs(2182) <= not a;
    layer1_outputs(2183) <= a and not b;
    layer1_outputs(2184) <= a or b;
    layer1_outputs(2185) <= 1'b0;
    layer1_outputs(2186) <= not (a or b);
    layer1_outputs(2187) <= a and not b;
    layer1_outputs(2188) <= not (a and b);
    layer1_outputs(2189) <= not b or a;
    layer1_outputs(2190) <= 1'b0;
    layer1_outputs(2191) <= not b or a;
    layer1_outputs(2192) <= 1'b0;
    layer1_outputs(2193) <= 1'b0;
    layer1_outputs(2194) <= a and not b;
    layer1_outputs(2195) <= not (a or b);
    layer1_outputs(2196) <= 1'b0;
    layer1_outputs(2197) <= b and not a;
    layer1_outputs(2198) <= b and not a;
    layer1_outputs(2199) <= a;
    layer1_outputs(2200) <= b;
    layer1_outputs(2201) <= b;
    layer1_outputs(2202) <= a;
    layer1_outputs(2203) <= a and not b;
    layer1_outputs(2204) <= not b or a;
    layer1_outputs(2205) <= a and b;
    layer1_outputs(2206) <= not (a and b);
    layer1_outputs(2207) <= not b;
    layer1_outputs(2208) <= b and not a;
    layer1_outputs(2209) <= not a;
    layer1_outputs(2210) <= b;
    layer1_outputs(2211) <= not a;
    layer1_outputs(2212) <= a and not b;
    layer1_outputs(2213) <= not (a and b);
    layer1_outputs(2214) <= not a or b;
    layer1_outputs(2215) <= 1'b1;
    layer1_outputs(2216) <= b;
    layer1_outputs(2217) <= not b;
    layer1_outputs(2218) <= not (a or b);
    layer1_outputs(2219) <= b;
    layer1_outputs(2220) <= 1'b1;
    layer1_outputs(2221) <= not b;
    layer1_outputs(2222) <= a or b;
    layer1_outputs(2223) <= 1'b1;
    layer1_outputs(2224) <= a xor b;
    layer1_outputs(2225) <= 1'b0;
    layer1_outputs(2226) <= a;
    layer1_outputs(2227) <= not a or b;
    layer1_outputs(2228) <= not (a xor b);
    layer1_outputs(2229) <= a;
    layer1_outputs(2230) <= b and not a;
    layer1_outputs(2231) <= not b;
    layer1_outputs(2232) <= a xor b;
    layer1_outputs(2233) <= 1'b0;
    layer1_outputs(2234) <= 1'b1;
    layer1_outputs(2235) <= not (a and b);
    layer1_outputs(2236) <= b;
    layer1_outputs(2237) <= not a or b;
    layer1_outputs(2238) <= 1'b1;
    layer1_outputs(2239) <= not a;
    layer1_outputs(2240) <= not b or a;
    layer1_outputs(2241) <= 1'b1;
    layer1_outputs(2242) <= 1'b0;
    layer1_outputs(2243) <= 1'b1;
    layer1_outputs(2244) <= 1'b1;
    layer1_outputs(2245) <= a or b;
    layer1_outputs(2246) <= a and not b;
    layer1_outputs(2247) <= a and b;
    layer1_outputs(2248) <= not (a and b);
    layer1_outputs(2249) <= not (a and b);
    layer1_outputs(2250) <= 1'b0;
    layer1_outputs(2251) <= not a or b;
    layer1_outputs(2252) <= 1'b1;
    layer1_outputs(2253) <= not (a or b);
    layer1_outputs(2254) <= a and not b;
    layer1_outputs(2255) <= not (a or b);
    layer1_outputs(2256) <= not b or a;
    layer1_outputs(2257) <= not b or a;
    layer1_outputs(2258) <= b;
    layer1_outputs(2259) <= a;
    layer1_outputs(2260) <= not a or b;
    layer1_outputs(2261) <= a and b;
    layer1_outputs(2262) <= 1'b1;
    layer1_outputs(2263) <= a and not b;
    layer1_outputs(2264) <= not b or a;
    layer1_outputs(2265) <= 1'b0;
    layer1_outputs(2266) <= a or b;
    layer1_outputs(2267) <= a and not b;
    layer1_outputs(2268) <= 1'b1;
    layer1_outputs(2269) <= a and not b;
    layer1_outputs(2270) <= a and b;
    layer1_outputs(2271) <= not (a and b);
    layer1_outputs(2272) <= a;
    layer1_outputs(2273) <= 1'b0;
    layer1_outputs(2274) <= not (a xor b);
    layer1_outputs(2275) <= not b;
    layer1_outputs(2276) <= 1'b1;
    layer1_outputs(2277) <= b and not a;
    layer1_outputs(2278) <= a and not b;
    layer1_outputs(2279) <= b and not a;
    layer1_outputs(2280) <= not a or b;
    layer1_outputs(2281) <= a and b;
    layer1_outputs(2282) <= not a or b;
    layer1_outputs(2283) <= not (a and b);
    layer1_outputs(2284) <= not a or b;
    layer1_outputs(2285) <= b;
    layer1_outputs(2286) <= a and b;
    layer1_outputs(2287) <= not (a or b);
    layer1_outputs(2288) <= b and not a;
    layer1_outputs(2289) <= 1'b1;
    layer1_outputs(2290) <= not b;
    layer1_outputs(2291) <= not b or a;
    layer1_outputs(2292) <= 1'b1;
    layer1_outputs(2293) <= b and not a;
    layer1_outputs(2294) <= not a;
    layer1_outputs(2295) <= not b;
    layer1_outputs(2296) <= not (a or b);
    layer1_outputs(2297) <= 1'b1;
    layer1_outputs(2298) <= b;
    layer1_outputs(2299) <= a;
    layer1_outputs(2300) <= a and b;
    layer1_outputs(2301) <= a and not b;
    layer1_outputs(2302) <= not b or a;
    layer1_outputs(2303) <= a and not b;
    layer1_outputs(2304) <= not (a or b);
    layer1_outputs(2305) <= not b or a;
    layer1_outputs(2306) <= a and not b;
    layer1_outputs(2307) <= not (a and b);
    layer1_outputs(2308) <= 1'b1;
    layer1_outputs(2309) <= a xor b;
    layer1_outputs(2310) <= 1'b0;
    layer1_outputs(2311) <= not a or b;
    layer1_outputs(2312) <= not b;
    layer1_outputs(2313) <= not (a and b);
    layer1_outputs(2314) <= not b;
    layer1_outputs(2315) <= not a;
    layer1_outputs(2316) <= not a or b;
    layer1_outputs(2317) <= a and b;
    layer1_outputs(2318) <= b;
    layer1_outputs(2319) <= 1'b0;
    layer1_outputs(2320) <= a and b;
    layer1_outputs(2321) <= 1'b0;
    layer1_outputs(2322) <= a and not b;
    layer1_outputs(2323) <= not b;
    layer1_outputs(2324) <= a and not b;
    layer1_outputs(2325) <= b and not a;
    layer1_outputs(2326) <= a xor b;
    layer1_outputs(2327) <= b;
    layer1_outputs(2328) <= b;
    layer1_outputs(2329) <= not (a and b);
    layer1_outputs(2330) <= not (a and b);
    layer1_outputs(2331) <= not b or a;
    layer1_outputs(2332) <= b and not a;
    layer1_outputs(2333) <= not a;
    layer1_outputs(2334) <= b;
    layer1_outputs(2335) <= a and not b;
    layer1_outputs(2336) <= 1'b1;
    layer1_outputs(2337) <= a and not b;
    layer1_outputs(2338) <= 1'b0;
    layer1_outputs(2339) <= not a;
    layer1_outputs(2340) <= 1'b0;
    layer1_outputs(2341) <= not b;
    layer1_outputs(2342) <= 1'b0;
    layer1_outputs(2343) <= 1'b1;
    layer1_outputs(2344) <= a or b;
    layer1_outputs(2345) <= b and not a;
    layer1_outputs(2346) <= not a;
    layer1_outputs(2347) <= 1'b1;
    layer1_outputs(2348) <= 1'b0;
    layer1_outputs(2349) <= a and b;
    layer1_outputs(2350) <= a xor b;
    layer1_outputs(2351) <= 1'b0;
    layer1_outputs(2352) <= not b;
    layer1_outputs(2353) <= not (a xor b);
    layer1_outputs(2354) <= not b or a;
    layer1_outputs(2355) <= not a;
    layer1_outputs(2356) <= 1'b0;
    layer1_outputs(2357) <= 1'b1;
    layer1_outputs(2358) <= a or b;
    layer1_outputs(2359) <= not b or a;
    layer1_outputs(2360) <= not b;
    layer1_outputs(2361) <= a;
    layer1_outputs(2362) <= b and not a;
    layer1_outputs(2363) <= 1'b0;
    layer1_outputs(2364) <= a and not b;
    layer1_outputs(2365) <= 1'b1;
    layer1_outputs(2366) <= not b;
    layer1_outputs(2367) <= not b or a;
    layer1_outputs(2368) <= a or b;
    layer1_outputs(2369) <= a and not b;
    layer1_outputs(2370) <= not b;
    layer1_outputs(2371) <= a xor b;
    layer1_outputs(2372) <= not b or a;
    layer1_outputs(2373) <= 1'b0;
    layer1_outputs(2374) <= a and not b;
    layer1_outputs(2375) <= b;
    layer1_outputs(2376) <= a;
    layer1_outputs(2377) <= 1'b1;
    layer1_outputs(2378) <= a and not b;
    layer1_outputs(2379) <= a or b;
    layer1_outputs(2380) <= a or b;
    layer1_outputs(2381) <= a and not b;
    layer1_outputs(2382) <= a or b;
    layer1_outputs(2383) <= a and b;
    layer1_outputs(2384) <= not (a and b);
    layer1_outputs(2385) <= a or b;
    layer1_outputs(2386) <= not a;
    layer1_outputs(2387) <= a and b;
    layer1_outputs(2388) <= not a or b;
    layer1_outputs(2389) <= not b;
    layer1_outputs(2390) <= not (a or b);
    layer1_outputs(2391) <= 1'b1;
    layer1_outputs(2392) <= not (a and b);
    layer1_outputs(2393) <= 1'b1;
    layer1_outputs(2394) <= a and not b;
    layer1_outputs(2395) <= b;
    layer1_outputs(2396) <= b;
    layer1_outputs(2397) <= 1'b0;
    layer1_outputs(2398) <= not (a and b);
    layer1_outputs(2399) <= not (a and b);
    layer1_outputs(2400) <= a or b;
    layer1_outputs(2401) <= a or b;
    layer1_outputs(2402) <= a;
    layer1_outputs(2403) <= b and not a;
    layer1_outputs(2404) <= a and not b;
    layer1_outputs(2405) <= a and b;
    layer1_outputs(2406) <= not b or a;
    layer1_outputs(2407) <= not b;
    layer1_outputs(2408) <= not b or a;
    layer1_outputs(2409) <= a and b;
    layer1_outputs(2410) <= b;
    layer1_outputs(2411) <= a or b;
    layer1_outputs(2412) <= not a or b;
    layer1_outputs(2413) <= a xor b;
    layer1_outputs(2414) <= not a or b;
    layer1_outputs(2415) <= 1'b0;
    layer1_outputs(2416) <= b and not a;
    layer1_outputs(2417) <= a xor b;
    layer1_outputs(2418) <= not (a and b);
    layer1_outputs(2419) <= a and b;
    layer1_outputs(2420) <= b;
    layer1_outputs(2421) <= b;
    layer1_outputs(2422) <= a or b;
    layer1_outputs(2423) <= a and not b;
    layer1_outputs(2424) <= not b or a;
    layer1_outputs(2425) <= not b;
    layer1_outputs(2426) <= 1'b1;
    layer1_outputs(2427) <= b and not a;
    layer1_outputs(2428) <= not b or a;
    layer1_outputs(2429) <= 1'b0;
    layer1_outputs(2430) <= not (a and b);
    layer1_outputs(2431) <= a xor b;
    layer1_outputs(2432) <= b and not a;
    layer1_outputs(2433) <= a;
    layer1_outputs(2434) <= not a or b;
    layer1_outputs(2435) <= 1'b0;
    layer1_outputs(2436) <= b;
    layer1_outputs(2437) <= not (a or b);
    layer1_outputs(2438) <= b and not a;
    layer1_outputs(2439) <= a and b;
    layer1_outputs(2440) <= b;
    layer1_outputs(2441) <= 1'b1;
    layer1_outputs(2442) <= b and not a;
    layer1_outputs(2443) <= not (a and b);
    layer1_outputs(2444) <= a and b;
    layer1_outputs(2445) <= not a;
    layer1_outputs(2446) <= 1'b1;
    layer1_outputs(2447) <= not b or a;
    layer1_outputs(2448) <= a or b;
    layer1_outputs(2449) <= not a or b;
    layer1_outputs(2450) <= 1'b1;
    layer1_outputs(2451) <= b;
    layer1_outputs(2452) <= 1'b0;
    layer1_outputs(2453) <= b and not a;
    layer1_outputs(2454) <= a and not b;
    layer1_outputs(2455) <= a and b;
    layer1_outputs(2456) <= 1'b0;
    layer1_outputs(2457) <= a;
    layer1_outputs(2458) <= 1'b0;
    layer1_outputs(2459) <= a and b;
    layer1_outputs(2460) <= not (a or b);
    layer1_outputs(2461) <= a xor b;
    layer1_outputs(2462) <= 1'b0;
    layer1_outputs(2463) <= not (a or b);
    layer1_outputs(2464) <= 1'b0;
    layer1_outputs(2465) <= 1'b1;
    layer1_outputs(2466) <= 1'b0;
    layer1_outputs(2467) <= 1'b1;
    layer1_outputs(2468) <= not (a xor b);
    layer1_outputs(2469) <= not (a xor b);
    layer1_outputs(2470) <= 1'b1;
    layer1_outputs(2471) <= not (a or b);
    layer1_outputs(2472) <= not (a and b);
    layer1_outputs(2473) <= not (a and b);
    layer1_outputs(2474) <= a;
    layer1_outputs(2475) <= 1'b0;
    layer1_outputs(2476) <= 1'b1;
    layer1_outputs(2477) <= b;
    layer1_outputs(2478) <= 1'b0;
    layer1_outputs(2479) <= not (a xor b);
    layer1_outputs(2480) <= not a;
    layer1_outputs(2481) <= not b;
    layer1_outputs(2482) <= a xor b;
    layer1_outputs(2483) <= not a or b;
    layer1_outputs(2484) <= b;
    layer1_outputs(2485) <= 1'b0;
    layer1_outputs(2486) <= not b;
    layer1_outputs(2487) <= 1'b0;
    layer1_outputs(2488) <= not b or a;
    layer1_outputs(2489) <= not (a and b);
    layer1_outputs(2490) <= 1'b1;
    layer1_outputs(2491) <= 1'b1;
    layer1_outputs(2492) <= a and b;
    layer1_outputs(2493) <= 1'b0;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= not b;
    layer1_outputs(2496) <= not b;
    layer1_outputs(2497) <= b;
    layer1_outputs(2498) <= b;
    layer1_outputs(2499) <= not (a and b);
    layer1_outputs(2500) <= not b;
    layer1_outputs(2501) <= 1'b1;
    layer1_outputs(2502) <= a;
    layer1_outputs(2503) <= 1'b0;
    layer1_outputs(2504) <= not (a or b);
    layer1_outputs(2505) <= not (a and b);
    layer1_outputs(2506) <= not a or b;
    layer1_outputs(2507) <= a and not b;
    layer1_outputs(2508) <= not b;
    layer1_outputs(2509) <= not (a or b);
    layer1_outputs(2510) <= not b or a;
    layer1_outputs(2511) <= not b;
    layer1_outputs(2512) <= 1'b1;
    layer1_outputs(2513) <= not a or b;
    layer1_outputs(2514) <= a;
    layer1_outputs(2515) <= not (a xor b);
    layer1_outputs(2516) <= b;
    layer1_outputs(2517) <= not a;
    layer1_outputs(2518) <= not (a and b);
    layer1_outputs(2519) <= not (a and b);
    layer1_outputs(2520) <= a xor b;
    layer1_outputs(2521) <= a or b;
    layer1_outputs(2522) <= not b or a;
    layer1_outputs(2523) <= a;
    layer1_outputs(2524) <= a and b;
    layer1_outputs(2525) <= 1'b0;
    layer1_outputs(2526) <= not b;
    layer1_outputs(2527) <= 1'b1;
    layer1_outputs(2528) <= not a or b;
    layer1_outputs(2529) <= not (a or b);
    layer1_outputs(2530) <= not b or a;
    layer1_outputs(2531) <= a and b;
    layer1_outputs(2532) <= not (a or b);
    layer1_outputs(2533) <= b;
    layer1_outputs(2534) <= not (a and b);
    layer1_outputs(2535) <= b and not a;
    layer1_outputs(2536) <= not (a and b);
    layer1_outputs(2537) <= not a;
    layer1_outputs(2538) <= 1'b0;
    layer1_outputs(2539) <= not b or a;
    layer1_outputs(2540) <= 1'b0;
    layer1_outputs(2541) <= not b or a;
    layer1_outputs(2542) <= not a;
    layer1_outputs(2543) <= b and not a;
    layer1_outputs(2544) <= b;
    layer1_outputs(2545) <= not b;
    layer1_outputs(2546) <= 1'b1;
    layer1_outputs(2547) <= 1'b1;
    layer1_outputs(2548) <= 1'b0;
    layer1_outputs(2549) <= not b or a;
    layer1_outputs(2550) <= not b or a;
    layer1_outputs(2551) <= not (a or b);
    layer1_outputs(2552) <= a and not b;
    layer1_outputs(2553) <= not (a xor b);
    layer1_outputs(2554) <= not a;
    layer1_outputs(2555) <= a and not b;
    layer1_outputs(2556) <= a and not b;
    layer1_outputs(2557) <= b;
    layer1_outputs(2558) <= not b;
    layer1_outputs(2559) <= 1'b1;
    layer1_outputs(2560) <= 1'b0;
    layer1_outputs(2561) <= a or b;
    layer1_outputs(2562) <= a or b;
    layer1_outputs(2563) <= b;
    layer1_outputs(2564) <= not (a and b);
    layer1_outputs(2565) <= not (a and b);
    layer1_outputs(2566) <= not b;
    layer1_outputs(2567) <= 1'b0;
    layer1_outputs(2568) <= 1'b1;
    layer1_outputs(2569) <= not b or a;
    layer1_outputs(2570) <= a;
    layer1_outputs(2571) <= a;
    layer1_outputs(2572) <= not b;
    layer1_outputs(2573) <= 1'b0;
    layer1_outputs(2574) <= not b;
    layer1_outputs(2575) <= not (a and b);
    layer1_outputs(2576) <= not a or b;
    layer1_outputs(2577) <= not a;
    layer1_outputs(2578) <= not b or a;
    layer1_outputs(2579) <= not a;
    layer1_outputs(2580) <= 1'b0;
    layer1_outputs(2581) <= b and not a;
    layer1_outputs(2582) <= not (a xor b);
    layer1_outputs(2583) <= b;
    layer1_outputs(2584) <= not b;
    layer1_outputs(2585) <= 1'b1;
    layer1_outputs(2586) <= a and b;
    layer1_outputs(2587) <= b and not a;
    layer1_outputs(2588) <= a or b;
    layer1_outputs(2589) <= a and b;
    layer1_outputs(2590) <= a and not b;
    layer1_outputs(2591) <= not a or b;
    layer1_outputs(2592) <= 1'b1;
    layer1_outputs(2593) <= not b or a;
    layer1_outputs(2594) <= 1'b0;
    layer1_outputs(2595) <= not a or b;
    layer1_outputs(2596) <= not a;
    layer1_outputs(2597) <= 1'b0;
    layer1_outputs(2598) <= b and not a;
    layer1_outputs(2599) <= 1'b1;
    layer1_outputs(2600) <= not (a and b);
    layer1_outputs(2601) <= a or b;
    layer1_outputs(2602) <= a and not b;
    layer1_outputs(2603) <= not (a or b);
    layer1_outputs(2604) <= a and b;
    layer1_outputs(2605) <= not a;
    layer1_outputs(2606) <= not (a xor b);
    layer1_outputs(2607) <= a or b;
    layer1_outputs(2608) <= not (a and b);
    layer1_outputs(2609) <= not a or b;
    layer1_outputs(2610) <= 1'b1;
    layer1_outputs(2611) <= a or b;
    layer1_outputs(2612) <= 1'b0;
    layer1_outputs(2613) <= a and b;
    layer1_outputs(2614) <= b;
    layer1_outputs(2615) <= b;
    layer1_outputs(2616) <= not a;
    layer1_outputs(2617) <= 1'b0;
    layer1_outputs(2618) <= a;
    layer1_outputs(2619) <= not b;
    layer1_outputs(2620) <= a xor b;
    layer1_outputs(2621) <= not b or a;
    layer1_outputs(2622) <= a and not b;
    layer1_outputs(2623) <= not (a or b);
    layer1_outputs(2624) <= b;
    layer1_outputs(2625) <= not a or b;
    layer1_outputs(2626) <= a or b;
    layer1_outputs(2627) <= 1'b0;
    layer1_outputs(2628) <= a and b;
    layer1_outputs(2629) <= 1'b1;
    layer1_outputs(2630) <= not (a or b);
    layer1_outputs(2631) <= a or b;
    layer1_outputs(2632) <= not (a or b);
    layer1_outputs(2633) <= a and not b;
    layer1_outputs(2634) <= not a or b;
    layer1_outputs(2635) <= not (a xor b);
    layer1_outputs(2636) <= not b or a;
    layer1_outputs(2637) <= 1'b0;
    layer1_outputs(2638) <= not b or a;
    layer1_outputs(2639) <= a and not b;
    layer1_outputs(2640) <= 1'b0;
    layer1_outputs(2641) <= not (a and b);
    layer1_outputs(2642) <= b;
    layer1_outputs(2643) <= not b;
    layer1_outputs(2644) <= not (a and b);
    layer1_outputs(2645) <= not b;
    layer1_outputs(2646) <= a;
    layer1_outputs(2647) <= 1'b0;
    layer1_outputs(2648) <= a;
    layer1_outputs(2649) <= b and not a;
    layer1_outputs(2650) <= not b;
    layer1_outputs(2651) <= a;
    layer1_outputs(2652) <= b and not a;
    layer1_outputs(2653) <= not b;
    layer1_outputs(2654) <= not (a and b);
    layer1_outputs(2655) <= b and not a;
    layer1_outputs(2656) <= not (a and b);
    layer1_outputs(2657) <= b;
    layer1_outputs(2658) <= a and not b;
    layer1_outputs(2659) <= not a or b;
    layer1_outputs(2660) <= a;
    layer1_outputs(2661) <= not b or a;
    layer1_outputs(2662) <= a and b;
    layer1_outputs(2663) <= not (a xor b);
    layer1_outputs(2664) <= b;
    layer1_outputs(2665) <= not a;
    layer1_outputs(2666) <= not a;
    layer1_outputs(2667) <= not a or b;
    layer1_outputs(2668) <= not a or b;
    layer1_outputs(2669) <= 1'b1;
    layer1_outputs(2670) <= not (a and b);
    layer1_outputs(2671) <= not a;
    layer1_outputs(2672) <= b and not a;
    layer1_outputs(2673) <= not (a and b);
    layer1_outputs(2674) <= not b or a;
    layer1_outputs(2675) <= not b;
    layer1_outputs(2676) <= not a or b;
    layer1_outputs(2677) <= not b or a;
    layer1_outputs(2678) <= not (a and b);
    layer1_outputs(2679) <= not a or b;
    layer1_outputs(2680) <= 1'b0;
    layer1_outputs(2681) <= 1'b1;
    layer1_outputs(2682) <= not b or a;
    layer1_outputs(2683) <= not a;
    layer1_outputs(2684) <= a;
    layer1_outputs(2685) <= 1'b0;
    layer1_outputs(2686) <= a and b;
    layer1_outputs(2687) <= not (a or b);
    layer1_outputs(2688) <= a and not b;
    layer1_outputs(2689) <= a;
    layer1_outputs(2690) <= not b or a;
    layer1_outputs(2691) <= not b;
    layer1_outputs(2692) <= not (a and b);
    layer1_outputs(2693) <= a;
    layer1_outputs(2694) <= 1'b0;
    layer1_outputs(2695) <= not a or b;
    layer1_outputs(2696) <= 1'b1;
    layer1_outputs(2697) <= a and not b;
    layer1_outputs(2698) <= not (a and b);
    layer1_outputs(2699) <= not a or b;
    layer1_outputs(2700) <= a or b;
    layer1_outputs(2701) <= 1'b0;
    layer1_outputs(2702) <= not (a or b);
    layer1_outputs(2703) <= not a or b;
    layer1_outputs(2704) <= b and not a;
    layer1_outputs(2705) <= 1'b0;
    layer1_outputs(2706) <= 1'b0;
    layer1_outputs(2707) <= 1'b0;
    layer1_outputs(2708) <= not b or a;
    layer1_outputs(2709) <= b;
    layer1_outputs(2710) <= 1'b0;
    layer1_outputs(2711) <= not a;
    layer1_outputs(2712) <= a or b;
    layer1_outputs(2713) <= 1'b0;
    layer1_outputs(2714) <= not a or b;
    layer1_outputs(2715) <= b and not a;
    layer1_outputs(2716) <= not (a xor b);
    layer1_outputs(2717) <= not b or a;
    layer1_outputs(2718) <= a and not b;
    layer1_outputs(2719) <= b and not a;
    layer1_outputs(2720) <= not a or b;
    layer1_outputs(2721) <= a and b;
    layer1_outputs(2722) <= a and not b;
    layer1_outputs(2723) <= a;
    layer1_outputs(2724) <= not b;
    layer1_outputs(2725) <= a;
    layer1_outputs(2726) <= not a;
    layer1_outputs(2727) <= not b;
    layer1_outputs(2728) <= not (a and b);
    layer1_outputs(2729) <= b and not a;
    layer1_outputs(2730) <= not a;
    layer1_outputs(2731) <= not b or a;
    layer1_outputs(2732) <= not b;
    layer1_outputs(2733) <= not (a or b);
    layer1_outputs(2734) <= 1'b0;
    layer1_outputs(2735) <= not a or b;
    layer1_outputs(2736) <= 1'b1;
    layer1_outputs(2737) <= not (a and b);
    layer1_outputs(2738) <= not a or b;
    layer1_outputs(2739) <= not a;
    layer1_outputs(2740) <= a;
    layer1_outputs(2741) <= a and not b;
    layer1_outputs(2742) <= not (a or b);
    layer1_outputs(2743) <= 1'b1;
    layer1_outputs(2744) <= not b;
    layer1_outputs(2745) <= not a;
    layer1_outputs(2746) <= not a or b;
    layer1_outputs(2747) <= 1'b1;
    layer1_outputs(2748) <= not (a or b);
    layer1_outputs(2749) <= a;
    layer1_outputs(2750) <= b and not a;
    layer1_outputs(2751) <= 1'b1;
    layer1_outputs(2752) <= not b or a;
    layer1_outputs(2753) <= not a;
    layer1_outputs(2754) <= not a;
    layer1_outputs(2755) <= not a or b;
    layer1_outputs(2756) <= a or b;
    layer1_outputs(2757) <= not (a and b);
    layer1_outputs(2758) <= a;
    layer1_outputs(2759) <= a and not b;
    layer1_outputs(2760) <= 1'b0;
    layer1_outputs(2761) <= b and not a;
    layer1_outputs(2762) <= b;
    layer1_outputs(2763) <= a and b;
    layer1_outputs(2764) <= b and not a;
    layer1_outputs(2765) <= not a or b;
    layer1_outputs(2766) <= not a;
    layer1_outputs(2767) <= b;
    layer1_outputs(2768) <= 1'b1;
    layer1_outputs(2769) <= not b;
    layer1_outputs(2770) <= b;
    layer1_outputs(2771) <= not b;
    layer1_outputs(2772) <= a xor b;
    layer1_outputs(2773) <= not b or a;
    layer1_outputs(2774) <= not a;
    layer1_outputs(2775) <= a or b;
    layer1_outputs(2776) <= a;
    layer1_outputs(2777) <= a;
    layer1_outputs(2778) <= a and b;
    layer1_outputs(2779) <= a or b;
    layer1_outputs(2780) <= a or b;
    layer1_outputs(2781) <= not b;
    layer1_outputs(2782) <= not (a and b);
    layer1_outputs(2783) <= 1'b0;
    layer1_outputs(2784) <= not (a and b);
    layer1_outputs(2785) <= not (a and b);
    layer1_outputs(2786) <= a or b;
    layer1_outputs(2787) <= not a or b;
    layer1_outputs(2788) <= b and not a;
    layer1_outputs(2789) <= not b;
    layer1_outputs(2790) <= not a;
    layer1_outputs(2791) <= not (a xor b);
    layer1_outputs(2792) <= not (a or b);
    layer1_outputs(2793) <= 1'b0;
    layer1_outputs(2794) <= a and not b;
    layer1_outputs(2795) <= a and not b;
    layer1_outputs(2796) <= b and not a;
    layer1_outputs(2797) <= a or b;
    layer1_outputs(2798) <= not b or a;
    layer1_outputs(2799) <= not (a or b);
    layer1_outputs(2800) <= a;
    layer1_outputs(2801) <= not b;
    layer1_outputs(2802) <= a and not b;
    layer1_outputs(2803) <= not b;
    layer1_outputs(2804) <= a and not b;
    layer1_outputs(2805) <= a and b;
    layer1_outputs(2806) <= 1'b1;
    layer1_outputs(2807) <= b and not a;
    layer1_outputs(2808) <= a and b;
    layer1_outputs(2809) <= 1'b0;
    layer1_outputs(2810) <= 1'b0;
    layer1_outputs(2811) <= a xor b;
    layer1_outputs(2812) <= b and not a;
    layer1_outputs(2813) <= 1'b1;
    layer1_outputs(2814) <= a;
    layer1_outputs(2815) <= a;
    layer1_outputs(2816) <= not b or a;
    layer1_outputs(2817) <= not a;
    layer1_outputs(2818) <= not (a and b);
    layer1_outputs(2819) <= b and not a;
    layer1_outputs(2820) <= not b or a;
    layer1_outputs(2821) <= not (a or b);
    layer1_outputs(2822) <= not a or b;
    layer1_outputs(2823) <= not (a and b);
    layer1_outputs(2824) <= a or b;
    layer1_outputs(2825) <= not b;
    layer1_outputs(2826) <= b;
    layer1_outputs(2827) <= a or b;
    layer1_outputs(2828) <= not (a xor b);
    layer1_outputs(2829) <= a;
    layer1_outputs(2830) <= a;
    layer1_outputs(2831) <= not (a or b);
    layer1_outputs(2832) <= b;
    layer1_outputs(2833) <= 1'b0;
    layer1_outputs(2834) <= a and not b;
    layer1_outputs(2835) <= a or b;
    layer1_outputs(2836) <= b and not a;
    layer1_outputs(2837) <= 1'b1;
    layer1_outputs(2838) <= not b;
    layer1_outputs(2839) <= not a;
    layer1_outputs(2840) <= b and not a;
    layer1_outputs(2841) <= 1'b1;
    layer1_outputs(2842) <= a and not b;
    layer1_outputs(2843) <= b and not a;
    layer1_outputs(2844) <= not (a or b);
    layer1_outputs(2845) <= 1'b1;
    layer1_outputs(2846) <= a or b;
    layer1_outputs(2847) <= a or b;
    layer1_outputs(2848) <= 1'b0;
    layer1_outputs(2849) <= not a;
    layer1_outputs(2850) <= b;
    layer1_outputs(2851) <= 1'b0;
    layer1_outputs(2852) <= not (a and b);
    layer1_outputs(2853) <= not (a or b);
    layer1_outputs(2854) <= b;
    layer1_outputs(2855) <= not (a or b);
    layer1_outputs(2856) <= 1'b1;
    layer1_outputs(2857) <= not b;
    layer1_outputs(2858) <= not (a or b);
    layer1_outputs(2859) <= not b or a;
    layer1_outputs(2860) <= not (a xor b);
    layer1_outputs(2861) <= not a or b;
    layer1_outputs(2862) <= not b;
    layer1_outputs(2863) <= a or b;
    layer1_outputs(2864) <= 1'b0;
    layer1_outputs(2865) <= not a or b;
    layer1_outputs(2866) <= b and not a;
    layer1_outputs(2867) <= b;
    layer1_outputs(2868) <= b;
    layer1_outputs(2869) <= not b;
    layer1_outputs(2870) <= a;
    layer1_outputs(2871) <= a and not b;
    layer1_outputs(2872) <= a and b;
    layer1_outputs(2873) <= not a or b;
    layer1_outputs(2874) <= not (a or b);
    layer1_outputs(2875) <= a and b;
    layer1_outputs(2876) <= not a;
    layer1_outputs(2877) <= not (a and b);
    layer1_outputs(2878) <= 1'b0;
    layer1_outputs(2879) <= a and b;
    layer1_outputs(2880) <= not (a or b);
    layer1_outputs(2881) <= not b;
    layer1_outputs(2882) <= a and not b;
    layer1_outputs(2883) <= not (a and b);
    layer1_outputs(2884) <= b;
    layer1_outputs(2885) <= not (a or b);
    layer1_outputs(2886) <= a and not b;
    layer1_outputs(2887) <= a and not b;
    layer1_outputs(2888) <= a and not b;
    layer1_outputs(2889) <= not a or b;
    layer1_outputs(2890) <= 1'b1;
    layer1_outputs(2891) <= not (a xor b);
    layer1_outputs(2892) <= not (a or b);
    layer1_outputs(2893) <= a and not b;
    layer1_outputs(2894) <= a and b;
    layer1_outputs(2895) <= a or b;
    layer1_outputs(2896) <= 1'b0;
    layer1_outputs(2897) <= a;
    layer1_outputs(2898) <= not a;
    layer1_outputs(2899) <= b and not a;
    layer1_outputs(2900) <= not a;
    layer1_outputs(2901) <= b;
    layer1_outputs(2902) <= a and b;
    layer1_outputs(2903) <= b and not a;
    layer1_outputs(2904) <= not (a or b);
    layer1_outputs(2905) <= a and b;
    layer1_outputs(2906) <= a or b;
    layer1_outputs(2907) <= not a;
    layer1_outputs(2908) <= a or b;
    layer1_outputs(2909) <= 1'b1;
    layer1_outputs(2910) <= not a or b;
    layer1_outputs(2911) <= not b;
    layer1_outputs(2912) <= a and b;
    layer1_outputs(2913) <= 1'b0;
    layer1_outputs(2914) <= a and b;
    layer1_outputs(2915) <= a or b;
    layer1_outputs(2916) <= not b;
    layer1_outputs(2917) <= 1'b0;
    layer1_outputs(2918) <= not a or b;
    layer1_outputs(2919) <= not (a or b);
    layer1_outputs(2920) <= not (a xor b);
    layer1_outputs(2921) <= not a;
    layer1_outputs(2922) <= not (a and b);
    layer1_outputs(2923) <= 1'b1;
    layer1_outputs(2924) <= not (a and b);
    layer1_outputs(2925) <= not a;
    layer1_outputs(2926) <= b;
    layer1_outputs(2927) <= a and not b;
    layer1_outputs(2928) <= not (a and b);
    layer1_outputs(2929) <= a;
    layer1_outputs(2930) <= b and not a;
    layer1_outputs(2931) <= a and not b;
    layer1_outputs(2932) <= b;
    layer1_outputs(2933) <= a and b;
    layer1_outputs(2934) <= a;
    layer1_outputs(2935) <= 1'b1;
    layer1_outputs(2936) <= a and not b;
    layer1_outputs(2937) <= 1'b0;
    layer1_outputs(2938) <= a or b;
    layer1_outputs(2939) <= not (a and b);
    layer1_outputs(2940) <= not a;
    layer1_outputs(2941) <= not b or a;
    layer1_outputs(2942) <= b and not a;
    layer1_outputs(2943) <= not (a xor b);
    layer1_outputs(2944) <= not (a or b);
    layer1_outputs(2945) <= 1'b1;
    layer1_outputs(2946) <= not (a and b);
    layer1_outputs(2947) <= b;
    layer1_outputs(2948) <= b;
    layer1_outputs(2949) <= a and not b;
    layer1_outputs(2950) <= not b;
    layer1_outputs(2951) <= a or b;
    layer1_outputs(2952) <= not a;
    layer1_outputs(2953) <= not (a and b);
    layer1_outputs(2954) <= a or b;
    layer1_outputs(2955) <= a and not b;
    layer1_outputs(2956) <= not b;
    layer1_outputs(2957) <= a or b;
    layer1_outputs(2958) <= b;
    layer1_outputs(2959) <= not b or a;
    layer1_outputs(2960) <= not (a or b);
    layer1_outputs(2961) <= not a or b;
    layer1_outputs(2962) <= a;
    layer1_outputs(2963) <= b and not a;
    layer1_outputs(2964) <= not (a and b);
    layer1_outputs(2965) <= not b or a;
    layer1_outputs(2966) <= b;
    layer1_outputs(2967) <= a and b;
    layer1_outputs(2968) <= not a or b;
    layer1_outputs(2969) <= a or b;
    layer1_outputs(2970) <= b and not a;
    layer1_outputs(2971) <= not a;
    layer1_outputs(2972) <= not (a or b);
    layer1_outputs(2973) <= not a;
    layer1_outputs(2974) <= 1'b1;
    layer1_outputs(2975) <= not (a xor b);
    layer1_outputs(2976) <= not b;
    layer1_outputs(2977) <= b;
    layer1_outputs(2978) <= not (a xor b);
    layer1_outputs(2979) <= not b;
    layer1_outputs(2980) <= a or b;
    layer1_outputs(2981) <= b and not a;
    layer1_outputs(2982) <= a and b;
    layer1_outputs(2983) <= not b or a;
    layer1_outputs(2984) <= b and not a;
    layer1_outputs(2985) <= a and not b;
    layer1_outputs(2986) <= b;
    layer1_outputs(2987) <= 1'b1;
    layer1_outputs(2988) <= a and b;
    layer1_outputs(2989) <= not (a or b);
    layer1_outputs(2990) <= not b or a;
    layer1_outputs(2991) <= a;
    layer1_outputs(2992) <= not (a and b);
    layer1_outputs(2993) <= not (a and b);
    layer1_outputs(2994) <= not (a xor b);
    layer1_outputs(2995) <= 1'b1;
    layer1_outputs(2996) <= not (a or b);
    layer1_outputs(2997) <= a and not b;
    layer1_outputs(2998) <= not (a or b);
    layer1_outputs(2999) <= not (a xor b);
    layer1_outputs(3000) <= not b or a;
    layer1_outputs(3001) <= a and not b;
    layer1_outputs(3002) <= a;
    layer1_outputs(3003) <= a and not b;
    layer1_outputs(3004) <= a;
    layer1_outputs(3005) <= a and b;
    layer1_outputs(3006) <= not b;
    layer1_outputs(3007) <= 1'b1;
    layer1_outputs(3008) <= a or b;
    layer1_outputs(3009) <= a xor b;
    layer1_outputs(3010) <= 1'b0;
    layer1_outputs(3011) <= not b or a;
    layer1_outputs(3012) <= not (a and b);
    layer1_outputs(3013) <= b;
    layer1_outputs(3014) <= a;
    layer1_outputs(3015) <= not a or b;
    layer1_outputs(3016) <= not (a and b);
    layer1_outputs(3017) <= 1'b1;
    layer1_outputs(3018) <= b and not a;
    layer1_outputs(3019) <= 1'b1;
    layer1_outputs(3020) <= not (a and b);
    layer1_outputs(3021) <= not b;
    layer1_outputs(3022) <= not (a or b);
    layer1_outputs(3023) <= 1'b0;
    layer1_outputs(3024) <= a or b;
    layer1_outputs(3025) <= not (a and b);
    layer1_outputs(3026) <= 1'b1;
    layer1_outputs(3027) <= 1'b1;
    layer1_outputs(3028) <= 1'b0;
    layer1_outputs(3029) <= not b;
    layer1_outputs(3030) <= 1'b1;
    layer1_outputs(3031) <= not b;
    layer1_outputs(3032) <= 1'b1;
    layer1_outputs(3033) <= not b;
    layer1_outputs(3034) <= a;
    layer1_outputs(3035) <= 1'b1;
    layer1_outputs(3036) <= a and b;
    layer1_outputs(3037) <= 1'b0;
    layer1_outputs(3038) <= a or b;
    layer1_outputs(3039) <= not (a and b);
    layer1_outputs(3040) <= 1'b0;
    layer1_outputs(3041) <= 1'b0;
    layer1_outputs(3042) <= 1'b1;
    layer1_outputs(3043) <= a or b;
    layer1_outputs(3044) <= 1'b1;
    layer1_outputs(3045) <= a;
    layer1_outputs(3046) <= a or b;
    layer1_outputs(3047) <= a xor b;
    layer1_outputs(3048) <= a and not b;
    layer1_outputs(3049) <= a and b;
    layer1_outputs(3050) <= not (a and b);
    layer1_outputs(3051) <= not (a and b);
    layer1_outputs(3052) <= a and b;
    layer1_outputs(3053) <= not b or a;
    layer1_outputs(3054) <= not (a or b);
    layer1_outputs(3055) <= not (a or b);
    layer1_outputs(3056) <= not b;
    layer1_outputs(3057) <= not a or b;
    layer1_outputs(3058) <= 1'b0;
    layer1_outputs(3059) <= b and not a;
    layer1_outputs(3060) <= a and b;
    layer1_outputs(3061) <= 1'b0;
    layer1_outputs(3062) <= not (a and b);
    layer1_outputs(3063) <= not a;
    layer1_outputs(3064) <= b;
    layer1_outputs(3065) <= a or b;
    layer1_outputs(3066) <= 1'b1;
    layer1_outputs(3067) <= 1'b1;
    layer1_outputs(3068) <= not (a and b);
    layer1_outputs(3069) <= a or b;
    layer1_outputs(3070) <= a or b;
    layer1_outputs(3071) <= b and not a;
    layer1_outputs(3072) <= a and b;
    layer1_outputs(3073) <= a;
    layer1_outputs(3074) <= not (a or b);
    layer1_outputs(3075) <= not a;
    layer1_outputs(3076) <= a and not b;
    layer1_outputs(3077) <= not b or a;
    layer1_outputs(3078) <= a or b;
    layer1_outputs(3079) <= 1'b1;
    layer1_outputs(3080) <= b and not a;
    layer1_outputs(3081) <= not b;
    layer1_outputs(3082) <= 1'b0;
    layer1_outputs(3083) <= not a;
    layer1_outputs(3084) <= a;
    layer1_outputs(3085) <= a and b;
    layer1_outputs(3086) <= b;
    layer1_outputs(3087) <= not b;
    layer1_outputs(3088) <= not a;
    layer1_outputs(3089) <= not b;
    layer1_outputs(3090) <= b and not a;
    layer1_outputs(3091) <= 1'b0;
    layer1_outputs(3092) <= a;
    layer1_outputs(3093) <= a xor b;
    layer1_outputs(3094) <= 1'b1;
    layer1_outputs(3095) <= a;
    layer1_outputs(3096) <= not b;
    layer1_outputs(3097) <= a xor b;
    layer1_outputs(3098) <= not a;
    layer1_outputs(3099) <= not a;
    layer1_outputs(3100) <= b and not a;
    layer1_outputs(3101) <= not a;
    layer1_outputs(3102) <= b;
    layer1_outputs(3103) <= a and not b;
    layer1_outputs(3104) <= a and b;
    layer1_outputs(3105) <= b and not a;
    layer1_outputs(3106) <= not b or a;
    layer1_outputs(3107) <= not (a or b);
    layer1_outputs(3108) <= not (a or b);
    layer1_outputs(3109) <= 1'b0;
    layer1_outputs(3110) <= not (a and b);
    layer1_outputs(3111) <= 1'b1;
    layer1_outputs(3112) <= b;
    layer1_outputs(3113) <= b and not a;
    layer1_outputs(3114) <= not b or a;
    layer1_outputs(3115) <= a xor b;
    layer1_outputs(3116) <= not b;
    layer1_outputs(3117) <= 1'b0;
    layer1_outputs(3118) <= not a or b;
    layer1_outputs(3119) <= a and b;
    layer1_outputs(3120) <= b;
    layer1_outputs(3121) <= b;
    layer1_outputs(3122) <= a and not b;
    layer1_outputs(3123) <= not (a and b);
    layer1_outputs(3124) <= not (a and b);
    layer1_outputs(3125) <= b and not a;
    layer1_outputs(3126) <= 1'b1;
    layer1_outputs(3127) <= not b or a;
    layer1_outputs(3128) <= 1'b1;
    layer1_outputs(3129) <= a and not b;
    layer1_outputs(3130) <= not a;
    layer1_outputs(3131) <= 1'b1;
    layer1_outputs(3132) <= not b or a;
    layer1_outputs(3133) <= not a or b;
    layer1_outputs(3134) <= not (a and b);
    layer1_outputs(3135) <= a;
    layer1_outputs(3136) <= 1'b0;
    layer1_outputs(3137) <= not (a and b);
    layer1_outputs(3138) <= b;
    layer1_outputs(3139) <= b;
    layer1_outputs(3140) <= not a or b;
    layer1_outputs(3141) <= not a;
    layer1_outputs(3142) <= 1'b0;
    layer1_outputs(3143) <= 1'b1;
    layer1_outputs(3144) <= not a or b;
    layer1_outputs(3145) <= a and not b;
    layer1_outputs(3146) <= a;
    layer1_outputs(3147) <= a xor b;
    layer1_outputs(3148) <= not b;
    layer1_outputs(3149) <= a and b;
    layer1_outputs(3150) <= a and b;
    layer1_outputs(3151) <= not a;
    layer1_outputs(3152) <= b;
    layer1_outputs(3153) <= 1'b1;
    layer1_outputs(3154) <= b and not a;
    layer1_outputs(3155) <= b;
    layer1_outputs(3156) <= a or b;
    layer1_outputs(3157) <= not (a and b);
    layer1_outputs(3158) <= not (a xor b);
    layer1_outputs(3159) <= b;
    layer1_outputs(3160) <= a or b;
    layer1_outputs(3161) <= 1'b0;
    layer1_outputs(3162) <= a or b;
    layer1_outputs(3163) <= not b or a;
    layer1_outputs(3164) <= b;
    layer1_outputs(3165) <= 1'b1;
    layer1_outputs(3166) <= not b or a;
    layer1_outputs(3167) <= not (a or b);
    layer1_outputs(3168) <= a or b;
    layer1_outputs(3169) <= a xor b;
    layer1_outputs(3170) <= a and b;
    layer1_outputs(3171) <= not (a and b);
    layer1_outputs(3172) <= 1'b0;
    layer1_outputs(3173) <= a and b;
    layer1_outputs(3174) <= a and not b;
    layer1_outputs(3175) <= a or b;
    layer1_outputs(3176) <= not b or a;
    layer1_outputs(3177) <= a and not b;
    layer1_outputs(3178) <= a xor b;
    layer1_outputs(3179) <= not b or a;
    layer1_outputs(3180) <= not a or b;
    layer1_outputs(3181) <= b and not a;
    layer1_outputs(3182) <= not a or b;
    layer1_outputs(3183) <= not (a and b);
    layer1_outputs(3184) <= a and b;
    layer1_outputs(3185) <= b;
    layer1_outputs(3186) <= a;
    layer1_outputs(3187) <= not (a or b);
    layer1_outputs(3188) <= b;
    layer1_outputs(3189) <= a or b;
    layer1_outputs(3190) <= a;
    layer1_outputs(3191) <= a;
    layer1_outputs(3192) <= not (a and b);
    layer1_outputs(3193) <= not (a or b);
    layer1_outputs(3194) <= not b or a;
    layer1_outputs(3195) <= a;
    layer1_outputs(3196) <= a xor b;
    layer1_outputs(3197) <= not a;
    layer1_outputs(3198) <= 1'b0;
    layer1_outputs(3199) <= a or b;
    layer1_outputs(3200) <= a or b;
    layer1_outputs(3201) <= not b;
    layer1_outputs(3202) <= 1'b0;
    layer1_outputs(3203) <= a;
    layer1_outputs(3204) <= 1'b1;
    layer1_outputs(3205) <= not b;
    layer1_outputs(3206) <= not (a or b);
    layer1_outputs(3207) <= b and not a;
    layer1_outputs(3208) <= a or b;
    layer1_outputs(3209) <= 1'b0;
    layer1_outputs(3210) <= b and not a;
    layer1_outputs(3211) <= 1'b1;
    layer1_outputs(3212) <= 1'b1;
    layer1_outputs(3213) <= not (a and b);
    layer1_outputs(3214) <= a or b;
    layer1_outputs(3215) <= a xor b;
    layer1_outputs(3216) <= a and b;
    layer1_outputs(3217) <= not b;
    layer1_outputs(3218) <= 1'b0;
    layer1_outputs(3219) <= 1'b1;
    layer1_outputs(3220) <= not a;
    layer1_outputs(3221) <= b and not a;
    layer1_outputs(3222) <= a;
    layer1_outputs(3223) <= a;
    layer1_outputs(3224) <= b;
    layer1_outputs(3225) <= 1'b0;
    layer1_outputs(3226) <= a or b;
    layer1_outputs(3227) <= a or b;
    layer1_outputs(3228) <= not (a or b);
    layer1_outputs(3229) <= not (a or b);
    layer1_outputs(3230) <= not a or b;
    layer1_outputs(3231) <= a or b;
    layer1_outputs(3232) <= not b;
    layer1_outputs(3233) <= 1'b1;
    layer1_outputs(3234) <= not (a or b);
    layer1_outputs(3235) <= not b or a;
    layer1_outputs(3236) <= 1'b1;
    layer1_outputs(3237) <= not b or a;
    layer1_outputs(3238) <= not (a or b);
    layer1_outputs(3239) <= not (a and b);
    layer1_outputs(3240) <= b;
    layer1_outputs(3241) <= not a;
    layer1_outputs(3242) <= a;
    layer1_outputs(3243) <= b;
    layer1_outputs(3244) <= not b or a;
    layer1_outputs(3245) <= not a or b;
    layer1_outputs(3246) <= not b;
    layer1_outputs(3247) <= not a or b;
    layer1_outputs(3248) <= a and not b;
    layer1_outputs(3249) <= 1'b1;
    layer1_outputs(3250) <= a or b;
    layer1_outputs(3251) <= 1'b0;
    layer1_outputs(3252) <= not b;
    layer1_outputs(3253) <= not (a or b);
    layer1_outputs(3254) <= 1'b1;
    layer1_outputs(3255) <= a xor b;
    layer1_outputs(3256) <= a;
    layer1_outputs(3257) <= not (a and b);
    layer1_outputs(3258) <= not (a and b);
    layer1_outputs(3259) <= b;
    layer1_outputs(3260) <= 1'b0;
    layer1_outputs(3261) <= not (a xor b);
    layer1_outputs(3262) <= not (a or b);
    layer1_outputs(3263) <= b;
    layer1_outputs(3264) <= a and not b;
    layer1_outputs(3265) <= b and not a;
    layer1_outputs(3266) <= not (a or b);
    layer1_outputs(3267) <= not (a and b);
    layer1_outputs(3268) <= b and not a;
    layer1_outputs(3269) <= 1'b0;
    layer1_outputs(3270) <= a and not b;
    layer1_outputs(3271) <= b and not a;
    layer1_outputs(3272) <= b;
    layer1_outputs(3273) <= 1'b0;
    layer1_outputs(3274) <= b;
    layer1_outputs(3275) <= 1'b1;
    layer1_outputs(3276) <= b and not a;
    layer1_outputs(3277) <= a or b;
    layer1_outputs(3278) <= not b or a;
    layer1_outputs(3279) <= b;
    layer1_outputs(3280) <= a or b;
    layer1_outputs(3281) <= not (a xor b);
    layer1_outputs(3282) <= not (a xor b);
    layer1_outputs(3283) <= b;
    layer1_outputs(3284) <= a or b;
    layer1_outputs(3285) <= a or b;
    layer1_outputs(3286) <= a;
    layer1_outputs(3287) <= a and not b;
    layer1_outputs(3288) <= a and not b;
    layer1_outputs(3289) <= not (a and b);
    layer1_outputs(3290) <= b and not a;
    layer1_outputs(3291) <= not b or a;
    layer1_outputs(3292) <= a and not b;
    layer1_outputs(3293) <= a and not b;
    layer1_outputs(3294) <= a and not b;
    layer1_outputs(3295) <= 1'b1;
    layer1_outputs(3296) <= not (a and b);
    layer1_outputs(3297) <= not (a xor b);
    layer1_outputs(3298) <= not a;
    layer1_outputs(3299) <= not a or b;
    layer1_outputs(3300) <= b and not a;
    layer1_outputs(3301) <= not (a or b);
    layer1_outputs(3302) <= not a or b;
    layer1_outputs(3303) <= 1'b0;
    layer1_outputs(3304) <= not b or a;
    layer1_outputs(3305) <= not (a xor b);
    layer1_outputs(3306) <= a and b;
    layer1_outputs(3307) <= b;
    layer1_outputs(3308) <= not (a and b);
    layer1_outputs(3309) <= not (a or b);
    layer1_outputs(3310) <= a and not b;
    layer1_outputs(3311) <= not a;
    layer1_outputs(3312) <= not b;
    layer1_outputs(3313) <= not a;
    layer1_outputs(3314) <= b and not a;
    layer1_outputs(3315) <= not (a xor b);
    layer1_outputs(3316) <= b and not a;
    layer1_outputs(3317) <= not a or b;
    layer1_outputs(3318) <= not (a or b);
    layer1_outputs(3319) <= not b or a;
    layer1_outputs(3320) <= not (a or b);
    layer1_outputs(3321) <= b and not a;
    layer1_outputs(3322) <= a;
    layer1_outputs(3323) <= not b or a;
    layer1_outputs(3324) <= a and not b;
    layer1_outputs(3325) <= a or b;
    layer1_outputs(3326) <= b;
    layer1_outputs(3327) <= not (a or b);
    layer1_outputs(3328) <= b and not a;
    layer1_outputs(3329) <= a and not b;
    layer1_outputs(3330) <= a;
    layer1_outputs(3331) <= not a;
    layer1_outputs(3332) <= not (a and b);
    layer1_outputs(3333) <= a or b;
    layer1_outputs(3334) <= a and not b;
    layer1_outputs(3335) <= not (a xor b);
    layer1_outputs(3336) <= not (a xor b);
    layer1_outputs(3337) <= 1'b1;
    layer1_outputs(3338) <= not b;
    layer1_outputs(3339) <= not (a or b);
    layer1_outputs(3340) <= not b;
    layer1_outputs(3341) <= not b;
    layer1_outputs(3342) <= 1'b0;
    layer1_outputs(3343) <= a and not b;
    layer1_outputs(3344) <= not (a xor b);
    layer1_outputs(3345) <= a or b;
    layer1_outputs(3346) <= not (a and b);
    layer1_outputs(3347) <= 1'b0;
    layer1_outputs(3348) <= a and not b;
    layer1_outputs(3349) <= not b or a;
    layer1_outputs(3350) <= not a or b;
    layer1_outputs(3351) <= b and not a;
    layer1_outputs(3352) <= not (a or b);
    layer1_outputs(3353) <= not (a and b);
    layer1_outputs(3354) <= not b or a;
    layer1_outputs(3355) <= not a or b;
    layer1_outputs(3356) <= not (a and b);
    layer1_outputs(3357) <= a;
    layer1_outputs(3358) <= not b or a;
    layer1_outputs(3359) <= a;
    layer1_outputs(3360) <= a and b;
    layer1_outputs(3361) <= not a or b;
    layer1_outputs(3362) <= a;
    layer1_outputs(3363) <= b;
    layer1_outputs(3364) <= not (a xor b);
    layer1_outputs(3365) <= a;
    layer1_outputs(3366) <= 1'b0;
    layer1_outputs(3367) <= a and b;
    layer1_outputs(3368) <= b;
    layer1_outputs(3369) <= a or b;
    layer1_outputs(3370) <= a or b;
    layer1_outputs(3371) <= a or b;
    layer1_outputs(3372) <= not b;
    layer1_outputs(3373) <= 1'b1;
    layer1_outputs(3374) <= not b or a;
    layer1_outputs(3375) <= 1'b0;
    layer1_outputs(3376) <= not b or a;
    layer1_outputs(3377) <= a and b;
    layer1_outputs(3378) <= 1'b0;
    layer1_outputs(3379) <= a xor b;
    layer1_outputs(3380) <= a;
    layer1_outputs(3381) <= not b or a;
    layer1_outputs(3382) <= a;
    layer1_outputs(3383) <= not a;
    layer1_outputs(3384) <= not (a or b);
    layer1_outputs(3385) <= b and not a;
    layer1_outputs(3386) <= not (a or b);
    layer1_outputs(3387) <= not b or a;
    layer1_outputs(3388) <= not b;
    layer1_outputs(3389) <= a and b;
    layer1_outputs(3390) <= 1'b0;
    layer1_outputs(3391) <= not b or a;
    layer1_outputs(3392) <= a or b;
    layer1_outputs(3393) <= not b;
    layer1_outputs(3394) <= a;
    layer1_outputs(3395) <= 1'b0;
    layer1_outputs(3396) <= not a;
    layer1_outputs(3397) <= not a or b;
    layer1_outputs(3398) <= 1'b1;
    layer1_outputs(3399) <= not b or a;
    layer1_outputs(3400) <= a or b;
    layer1_outputs(3401) <= not a;
    layer1_outputs(3402) <= 1'b0;
    layer1_outputs(3403) <= not b or a;
    layer1_outputs(3404) <= b and not a;
    layer1_outputs(3405) <= a and not b;
    layer1_outputs(3406) <= b;
    layer1_outputs(3407) <= b;
    layer1_outputs(3408) <= not a or b;
    layer1_outputs(3409) <= not b or a;
    layer1_outputs(3410) <= a or b;
    layer1_outputs(3411) <= a or b;
    layer1_outputs(3412) <= not (a xor b);
    layer1_outputs(3413) <= 1'b1;
    layer1_outputs(3414) <= b and not a;
    layer1_outputs(3415) <= not b or a;
    layer1_outputs(3416) <= not a;
    layer1_outputs(3417) <= 1'b0;
    layer1_outputs(3418) <= b;
    layer1_outputs(3419) <= 1'b1;
    layer1_outputs(3420) <= not (a and b);
    layer1_outputs(3421) <= not b or a;
    layer1_outputs(3422) <= not (a xor b);
    layer1_outputs(3423) <= b and not a;
    layer1_outputs(3424) <= not (a or b);
    layer1_outputs(3425) <= a and b;
    layer1_outputs(3426) <= not a or b;
    layer1_outputs(3427) <= 1'b1;
    layer1_outputs(3428) <= not a or b;
    layer1_outputs(3429) <= not a;
    layer1_outputs(3430) <= a and not b;
    layer1_outputs(3431) <= not a or b;
    layer1_outputs(3432) <= a and b;
    layer1_outputs(3433) <= a or b;
    layer1_outputs(3434) <= not b or a;
    layer1_outputs(3435) <= not (a xor b);
    layer1_outputs(3436) <= b and not a;
    layer1_outputs(3437) <= a and not b;
    layer1_outputs(3438) <= b and not a;
    layer1_outputs(3439) <= a and not b;
    layer1_outputs(3440) <= 1'b1;
    layer1_outputs(3441) <= 1'b0;
    layer1_outputs(3442) <= b;
    layer1_outputs(3443) <= not b or a;
    layer1_outputs(3444) <= a or b;
    layer1_outputs(3445) <= 1'b0;
    layer1_outputs(3446) <= not (a or b);
    layer1_outputs(3447) <= not a;
    layer1_outputs(3448) <= a or b;
    layer1_outputs(3449) <= 1'b0;
    layer1_outputs(3450) <= a xor b;
    layer1_outputs(3451) <= a and not b;
    layer1_outputs(3452) <= not b or a;
    layer1_outputs(3453) <= not (a and b);
    layer1_outputs(3454) <= b;
    layer1_outputs(3455) <= a and not b;
    layer1_outputs(3456) <= not b or a;
    layer1_outputs(3457) <= not (a and b);
    layer1_outputs(3458) <= not b or a;
    layer1_outputs(3459) <= not a or b;
    layer1_outputs(3460) <= a and b;
    layer1_outputs(3461) <= not (a or b);
    layer1_outputs(3462) <= a;
    layer1_outputs(3463) <= not (a xor b);
    layer1_outputs(3464) <= not b;
    layer1_outputs(3465) <= not b;
    layer1_outputs(3466) <= not b;
    layer1_outputs(3467) <= b;
    layer1_outputs(3468) <= not b or a;
    layer1_outputs(3469) <= a and b;
    layer1_outputs(3470) <= not b or a;
    layer1_outputs(3471) <= a and b;
    layer1_outputs(3472) <= a and not b;
    layer1_outputs(3473) <= a or b;
    layer1_outputs(3474) <= 1'b1;
    layer1_outputs(3475) <= a and not b;
    layer1_outputs(3476) <= a and b;
    layer1_outputs(3477) <= a and not b;
    layer1_outputs(3478) <= not b or a;
    layer1_outputs(3479) <= 1'b0;
    layer1_outputs(3480) <= a and not b;
    layer1_outputs(3481) <= b;
    layer1_outputs(3482) <= not (a or b);
    layer1_outputs(3483) <= b;
    layer1_outputs(3484) <= not b;
    layer1_outputs(3485) <= a and not b;
    layer1_outputs(3486) <= b and not a;
    layer1_outputs(3487) <= not a or b;
    layer1_outputs(3488) <= a or b;
    layer1_outputs(3489) <= b;
    layer1_outputs(3490) <= not a;
    layer1_outputs(3491) <= 1'b0;
    layer1_outputs(3492) <= b and not a;
    layer1_outputs(3493) <= not (a or b);
    layer1_outputs(3494) <= not (a or b);
    layer1_outputs(3495) <= a;
    layer1_outputs(3496) <= not a;
    layer1_outputs(3497) <= a and not b;
    layer1_outputs(3498) <= b;
    layer1_outputs(3499) <= not (a or b);
    layer1_outputs(3500) <= a xor b;
    layer1_outputs(3501) <= not (a xor b);
    layer1_outputs(3502) <= a and b;
    layer1_outputs(3503) <= b and not a;
    layer1_outputs(3504) <= not (a and b);
    layer1_outputs(3505) <= not b;
    layer1_outputs(3506) <= b;
    layer1_outputs(3507) <= not a or b;
    layer1_outputs(3508) <= a xor b;
    layer1_outputs(3509) <= a and b;
    layer1_outputs(3510) <= a or b;
    layer1_outputs(3511) <= not (a and b);
    layer1_outputs(3512) <= not (a and b);
    layer1_outputs(3513) <= not a;
    layer1_outputs(3514) <= a and not b;
    layer1_outputs(3515) <= b and not a;
    layer1_outputs(3516) <= not (a or b);
    layer1_outputs(3517) <= 1'b1;
    layer1_outputs(3518) <= not (a and b);
    layer1_outputs(3519) <= 1'b1;
    layer1_outputs(3520) <= a;
    layer1_outputs(3521) <= not (a and b);
    layer1_outputs(3522) <= not (a or b);
    layer1_outputs(3523) <= not (a or b);
    layer1_outputs(3524) <= not b or a;
    layer1_outputs(3525) <= not a or b;
    layer1_outputs(3526) <= a;
    layer1_outputs(3527) <= not (a and b);
    layer1_outputs(3528) <= b and not a;
    layer1_outputs(3529) <= a and b;
    layer1_outputs(3530) <= 1'b0;
    layer1_outputs(3531) <= 1'b0;
    layer1_outputs(3532) <= b;
    layer1_outputs(3533) <= not b;
    layer1_outputs(3534) <= b;
    layer1_outputs(3535) <= not b;
    layer1_outputs(3536) <= a and b;
    layer1_outputs(3537) <= b and not a;
    layer1_outputs(3538) <= a and not b;
    layer1_outputs(3539) <= not (a or b);
    layer1_outputs(3540) <= 1'b0;
    layer1_outputs(3541) <= b;
    layer1_outputs(3542) <= not b;
    layer1_outputs(3543) <= b and not a;
    layer1_outputs(3544) <= 1'b0;
    layer1_outputs(3545) <= not b or a;
    layer1_outputs(3546) <= not (a and b);
    layer1_outputs(3547) <= not (a and b);
    layer1_outputs(3548) <= not b or a;
    layer1_outputs(3549) <= not (a and b);
    layer1_outputs(3550) <= not a;
    layer1_outputs(3551) <= not b;
    layer1_outputs(3552) <= a and not b;
    layer1_outputs(3553) <= not b;
    layer1_outputs(3554) <= not (a and b);
    layer1_outputs(3555) <= b and not a;
    layer1_outputs(3556) <= not b or a;
    layer1_outputs(3557) <= not a or b;
    layer1_outputs(3558) <= b;
    layer1_outputs(3559) <= b and not a;
    layer1_outputs(3560) <= 1'b1;
    layer1_outputs(3561) <= a and not b;
    layer1_outputs(3562) <= not (a and b);
    layer1_outputs(3563) <= not b;
    layer1_outputs(3564) <= b and not a;
    layer1_outputs(3565) <= not (a xor b);
    layer1_outputs(3566) <= not a;
    layer1_outputs(3567) <= 1'b0;
    layer1_outputs(3568) <= not (a and b);
    layer1_outputs(3569) <= a xor b;
    layer1_outputs(3570) <= not (a xor b);
    layer1_outputs(3571) <= a;
    layer1_outputs(3572) <= not (a or b);
    layer1_outputs(3573) <= not (a or b);
    layer1_outputs(3574) <= not (a and b);
    layer1_outputs(3575) <= a and b;
    layer1_outputs(3576) <= a and b;
    layer1_outputs(3577) <= a or b;
    layer1_outputs(3578) <= 1'b1;
    layer1_outputs(3579) <= not a or b;
    layer1_outputs(3580) <= b and not a;
    layer1_outputs(3581) <= not b or a;
    layer1_outputs(3582) <= a;
    layer1_outputs(3583) <= a and b;
    layer1_outputs(3584) <= 1'b0;
    layer1_outputs(3585) <= not a or b;
    layer1_outputs(3586) <= a and not b;
    layer1_outputs(3587) <= a;
    layer1_outputs(3588) <= b and not a;
    layer1_outputs(3589) <= b and not a;
    layer1_outputs(3590) <= not (a and b);
    layer1_outputs(3591) <= a and b;
    layer1_outputs(3592) <= a and b;
    layer1_outputs(3593) <= a and b;
    layer1_outputs(3594) <= not (a or b);
    layer1_outputs(3595) <= a or b;
    layer1_outputs(3596) <= a or b;
    layer1_outputs(3597) <= not a or b;
    layer1_outputs(3598) <= b;
    layer1_outputs(3599) <= b and not a;
    layer1_outputs(3600) <= b;
    layer1_outputs(3601) <= not (a and b);
    layer1_outputs(3602) <= a and b;
    layer1_outputs(3603) <= not a or b;
    layer1_outputs(3604) <= not b;
    layer1_outputs(3605) <= not a or b;
    layer1_outputs(3606) <= 1'b1;
    layer1_outputs(3607) <= b and not a;
    layer1_outputs(3608) <= not (a and b);
    layer1_outputs(3609) <= not (a or b);
    layer1_outputs(3610) <= 1'b1;
    layer1_outputs(3611) <= 1'b0;
    layer1_outputs(3612) <= not (a or b);
    layer1_outputs(3613) <= 1'b0;
    layer1_outputs(3614) <= not a;
    layer1_outputs(3615) <= b;
    layer1_outputs(3616) <= b and not a;
    layer1_outputs(3617) <= not b;
    layer1_outputs(3618) <= 1'b1;
    layer1_outputs(3619) <= not b or a;
    layer1_outputs(3620) <= a or b;
    layer1_outputs(3621) <= not a or b;
    layer1_outputs(3622) <= 1'b0;
    layer1_outputs(3623) <= b;
    layer1_outputs(3624) <= not (a or b);
    layer1_outputs(3625) <= not a;
    layer1_outputs(3626) <= a and b;
    layer1_outputs(3627) <= not (a and b);
    layer1_outputs(3628) <= not a or b;
    layer1_outputs(3629) <= 1'b1;
    layer1_outputs(3630) <= not (a xor b);
    layer1_outputs(3631) <= not (a or b);
    layer1_outputs(3632) <= not a;
    layer1_outputs(3633) <= 1'b0;
    layer1_outputs(3634) <= not (a or b);
    layer1_outputs(3635) <= a xor b;
    layer1_outputs(3636) <= 1'b1;
    layer1_outputs(3637) <= 1'b0;
    layer1_outputs(3638) <= a or b;
    layer1_outputs(3639) <= not b;
    layer1_outputs(3640) <= not (a and b);
    layer1_outputs(3641) <= not (a xor b);
    layer1_outputs(3642) <= not (a or b);
    layer1_outputs(3643) <= a and not b;
    layer1_outputs(3644) <= b;
    layer1_outputs(3645) <= not a;
    layer1_outputs(3646) <= not a or b;
    layer1_outputs(3647) <= b;
    layer1_outputs(3648) <= a and not b;
    layer1_outputs(3649) <= not b;
    layer1_outputs(3650) <= a and b;
    layer1_outputs(3651) <= a and b;
    layer1_outputs(3652) <= not b;
    layer1_outputs(3653) <= 1'b1;
    layer1_outputs(3654) <= 1'b1;
    layer1_outputs(3655) <= a and b;
    layer1_outputs(3656) <= not b or a;
    layer1_outputs(3657) <= b;
    layer1_outputs(3658) <= not a;
    layer1_outputs(3659) <= not a;
    layer1_outputs(3660) <= b;
    layer1_outputs(3661) <= not (a or b);
    layer1_outputs(3662) <= not b or a;
    layer1_outputs(3663) <= not (a or b);
    layer1_outputs(3664) <= not b;
    layer1_outputs(3665) <= a;
    layer1_outputs(3666) <= not a;
    layer1_outputs(3667) <= 1'b1;
    layer1_outputs(3668) <= 1'b1;
    layer1_outputs(3669) <= 1'b0;
    layer1_outputs(3670) <= a and b;
    layer1_outputs(3671) <= not (a or b);
    layer1_outputs(3672) <= 1'b1;
    layer1_outputs(3673) <= a and not b;
    layer1_outputs(3674) <= a or b;
    layer1_outputs(3675) <= not a;
    layer1_outputs(3676) <= not b or a;
    layer1_outputs(3677) <= a or b;
    layer1_outputs(3678) <= not (a and b);
    layer1_outputs(3679) <= a;
    layer1_outputs(3680) <= a or b;
    layer1_outputs(3681) <= not (a and b);
    layer1_outputs(3682) <= a and not b;
    layer1_outputs(3683) <= not (a and b);
    layer1_outputs(3684) <= a and not b;
    layer1_outputs(3685) <= 1'b1;
    layer1_outputs(3686) <= a;
    layer1_outputs(3687) <= not (a or b);
    layer1_outputs(3688) <= b and not a;
    layer1_outputs(3689) <= 1'b1;
    layer1_outputs(3690) <= not b;
    layer1_outputs(3691) <= a xor b;
    layer1_outputs(3692) <= b;
    layer1_outputs(3693) <= not b or a;
    layer1_outputs(3694) <= not b or a;
    layer1_outputs(3695) <= not (a or b);
    layer1_outputs(3696) <= 1'b0;
    layer1_outputs(3697) <= not a or b;
    layer1_outputs(3698) <= not (a xor b);
    layer1_outputs(3699) <= a and b;
    layer1_outputs(3700) <= 1'b0;
    layer1_outputs(3701) <= not (a and b);
    layer1_outputs(3702) <= not a;
    layer1_outputs(3703) <= not (a or b);
    layer1_outputs(3704) <= a xor b;
    layer1_outputs(3705) <= not (a or b);
    layer1_outputs(3706) <= a and b;
    layer1_outputs(3707) <= 1'b1;
    layer1_outputs(3708) <= a;
    layer1_outputs(3709) <= 1'b0;
    layer1_outputs(3710) <= not b;
    layer1_outputs(3711) <= not (a xor b);
    layer1_outputs(3712) <= a and b;
    layer1_outputs(3713) <= a and not b;
    layer1_outputs(3714) <= 1'b1;
    layer1_outputs(3715) <= not b;
    layer1_outputs(3716) <= not a;
    layer1_outputs(3717) <= not (a or b);
    layer1_outputs(3718) <= a and not b;
    layer1_outputs(3719) <= not b;
    layer1_outputs(3720) <= 1'b0;
    layer1_outputs(3721) <= 1'b0;
    layer1_outputs(3722) <= not (a and b);
    layer1_outputs(3723) <= not b or a;
    layer1_outputs(3724) <= not (a or b);
    layer1_outputs(3725) <= not b or a;
    layer1_outputs(3726) <= a;
    layer1_outputs(3727) <= not a;
    layer1_outputs(3728) <= a and b;
    layer1_outputs(3729) <= a and not b;
    layer1_outputs(3730) <= a or b;
    layer1_outputs(3731) <= not a;
    layer1_outputs(3732) <= not (a and b);
    layer1_outputs(3733) <= not (a xor b);
    layer1_outputs(3734) <= b;
    layer1_outputs(3735) <= not b;
    layer1_outputs(3736) <= a xor b;
    layer1_outputs(3737) <= a or b;
    layer1_outputs(3738) <= b;
    layer1_outputs(3739) <= b;
    layer1_outputs(3740) <= a and b;
    layer1_outputs(3741) <= a and b;
    layer1_outputs(3742) <= not (a or b);
    layer1_outputs(3743) <= not b;
    layer1_outputs(3744) <= 1'b1;
    layer1_outputs(3745) <= b;
    layer1_outputs(3746) <= b and not a;
    layer1_outputs(3747) <= b;
    layer1_outputs(3748) <= not (a or b);
    layer1_outputs(3749) <= not a;
    layer1_outputs(3750) <= 1'b1;
    layer1_outputs(3751) <= 1'b0;
    layer1_outputs(3752) <= b and not a;
    layer1_outputs(3753) <= a and not b;
    layer1_outputs(3754) <= not (a or b);
    layer1_outputs(3755) <= a xor b;
    layer1_outputs(3756) <= not (a xor b);
    layer1_outputs(3757) <= not b;
    layer1_outputs(3758) <= not b or a;
    layer1_outputs(3759) <= a;
    layer1_outputs(3760) <= not a or b;
    layer1_outputs(3761) <= a;
    layer1_outputs(3762) <= not a or b;
    layer1_outputs(3763) <= not b;
    layer1_outputs(3764) <= not a;
    layer1_outputs(3765) <= 1'b1;
    layer1_outputs(3766) <= a;
    layer1_outputs(3767) <= a and not b;
    layer1_outputs(3768) <= 1'b0;
    layer1_outputs(3769) <= 1'b0;
    layer1_outputs(3770) <= a;
    layer1_outputs(3771) <= not (a or b);
    layer1_outputs(3772) <= not (a or b);
    layer1_outputs(3773) <= not a;
    layer1_outputs(3774) <= not a;
    layer1_outputs(3775) <= not a;
    layer1_outputs(3776) <= b and not a;
    layer1_outputs(3777) <= not b;
    layer1_outputs(3778) <= not (a and b);
    layer1_outputs(3779) <= a;
    layer1_outputs(3780) <= b;
    layer1_outputs(3781) <= not a;
    layer1_outputs(3782) <= a and b;
    layer1_outputs(3783) <= 1'b0;
    layer1_outputs(3784) <= 1'b0;
    layer1_outputs(3785) <= a and not b;
    layer1_outputs(3786) <= 1'b1;
    layer1_outputs(3787) <= 1'b1;
    layer1_outputs(3788) <= a or b;
    layer1_outputs(3789) <= not (a xor b);
    layer1_outputs(3790) <= a and not b;
    layer1_outputs(3791) <= not (a or b);
    layer1_outputs(3792) <= a and b;
    layer1_outputs(3793) <= b;
    layer1_outputs(3794) <= not b;
    layer1_outputs(3795) <= a or b;
    layer1_outputs(3796) <= a;
    layer1_outputs(3797) <= a xor b;
    layer1_outputs(3798) <= a or b;
    layer1_outputs(3799) <= 1'b0;
    layer1_outputs(3800) <= not (a or b);
    layer1_outputs(3801) <= a and b;
    layer1_outputs(3802) <= not a;
    layer1_outputs(3803) <= 1'b1;
    layer1_outputs(3804) <= b;
    layer1_outputs(3805) <= 1'b0;
    layer1_outputs(3806) <= b and not a;
    layer1_outputs(3807) <= not (a xor b);
    layer1_outputs(3808) <= 1'b0;
    layer1_outputs(3809) <= 1'b0;
    layer1_outputs(3810) <= 1'b0;
    layer1_outputs(3811) <= 1'b1;
    layer1_outputs(3812) <= not a;
    layer1_outputs(3813) <= not (a or b);
    layer1_outputs(3814) <= 1'b1;
    layer1_outputs(3815) <= not a or b;
    layer1_outputs(3816) <= b;
    layer1_outputs(3817) <= not (a and b);
    layer1_outputs(3818) <= a;
    layer1_outputs(3819) <= not b;
    layer1_outputs(3820) <= a and b;
    layer1_outputs(3821) <= not (a or b);
    layer1_outputs(3822) <= b and not a;
    layer1_outputs(3823) <= 1'b1;
    layer1_outputs(3824) <= a and not b;
    layer1_outputs(3825) <= a and not b;
    layer1_outputs(3826) <= not b or a;
    layer1_outputs(3827) <= a and b;
    layer1_outputs(3828) <= a and b;
    layer1_outputs(3829) <= 1'b1;
    layer1_outputs(3830) <= a;
    layer1_outputs(3831) <= 1'b0;
    layer1_outputs(3832) <= not b;
    layer1_outputs(3833) <= a;
    layer1_outputs(3834) <= a and b;
    layer1_outputs(3835) <= a xor b;
    layer1_outputs(3836) <= a and b;
    layer1_outputs(3837) <= not (a or b);
    layer1_outputs(3838) <= not (a or b);
    layer1_outputs(3839) <= a and not b;
    layer1_outputs(3840) <= b;
    layer1_outputs(3841) <= not b;
    layer1_outputs(3842) <= not (a and b);
    layer1_outputs(3843) <= a and not b;
    layer1_outputs(3844) <= 1'b0;
    layer1_outputs(3845) <= not b;
    layer1_outputs(3846) <= not b;
    layer1_outputs(3847) <= b;
    layer1_outputs(3848) <= a and b;
    layer1_outputs(3849) <= not b or a;
    layer1_outputs(3850) <= a;
    layer1_outputs(3851) <= a and b;
    layer1_outputs(3852) <= not a;
    layer1_outputs(3853) <= not (a and b);
    layer1_outputs(3854) <= a and not b;
    layer1_outputs(3855) <= not (a or b);
    layer1_outputs(3856) <= b;
    layer1_outputs(3857) <= not b or a;
    layer1_outputs(3858) <= not b or a;
    layer1_outputs(3859) <= a or b;
    layer1_outputs(3860) <= b and not a;
    layer1_outputs(3861) <= not b;
    layer1_outputs(3862) <= not a or b;
    layer1_outputs(3863) <= 1'b0;
    layer1_outputs(3864) <= not a or b;
    layer1_outputs(3865) <= not b;
    layer1_outputs(3866) <= 1'b0;
    layer1_outputs(3867) <= not (a xor b);
    layer1_outputs(3868) <= a or b;
    layer1_outputs(3869) <= 1'b0;
    layer1_outputs(3870) <= 1'b0;
    layer1_outputs(3871) <= not b or a;
    layer1_outputs(3872) <= a;
    layer1_outputs(3873) <= b;
    layer1_outputs(3874) <= a;
    layer1_outputs(3875) <= a or b;
    layer1_outputs(3876) <= 1'b1;
    layer1_outputs(3877) <= b and not a;
    layer1_outputs(3878) <= 1'b0;
    layer1_outputs(3879) <= b;
    layer1_outputs(3880) <= 1'b0;
    layer1_outputs(3881) <= a or b;
    layer1_outputs(3882) <= a or b;
    layer1_outputs(3883) <= 1'b0;
    layer1_outputs(3884) <= a and not b;
    layer1_outputs(3885) <= not (a or b);
    layer1_outputs(3886) <= not (a or b);
    layer1_outputs(3887) <= a or b;
    layer1_outputs(3888) <= a;
    layer1_outputs(3889) <= b and not a;
    layer1_outputs(3890) <= not a or b;
    layer1_outputs(3891) <= a or b;
    layer1_outputs(3892) <= a;
    layer1_outputs(3893) <= not (a and b);
    layer1_outputs(3894) <= 1'b0;
    layer1_outputs(3895) <= 1'b0;
    layer1_outputs(3896) <= b and not a;
    layer1_outputs(3897) <= a;
    layer1_outputs(3898) <= not b;
    layer1_outputs(3899) <= b and not a;
    layer1_outputs(3900) <= not (a and b);
    layer1_outputs(3901) <= not b;
    layer1_outputs(3902) <= not b;
    layer1_outputs(3903) <= 1'b0;
    layer1_outputs(3904) <= 1'b1;
    layer1_outputs(3905) <= not a or b;
    layer1_outputs(3906) <= not a or b;
    layer1_outputs(3907) <= not (a or b);
    layer1_outputs(3908) <= 1'b1;
    layer1_outputs(3909) <= not b;
    layer1_outputs(3910) <= not a;
    layer1_outputs(3911) <= not a;
    layer1_outputs(3912) <= not (a xor b);
    layer1_outputs(3913) <= not (a or b);
    layer1_outputs(3914) <= a and not b;
    layer1_outputs(3915) <= a and b;
    layer1_outputs(3916) <= a;
    layer1_outputs(3917) <= a;
    layer1_outputs(3918) <= not a or b;
    layer1_outputs(3919) <= a and b;
    layer1_outputs(3920) <= b;
    layer1_outputs(3921) <= not a or b;
    layer1_outputs(3922) <= b;
    layer1_outputs(3923) <= not b or a;
    layer1_outputs(3924) <= b and not a;
    layer1_outputs(3925) <= not (a or b);
    layer1_outputs(3926) <= not b;
    layer1_outputs(3927) <= 1'b1;
    layer1_outputs(3928) <= b and not a;
    layer1_outputs(3929) <= b and not a;
    layer1_outputs(3930) <= not b;
    layer1_outputs(3931) <= not b;
    layer1_outputs(3932) <= 1'b0;
    layer1_outputs(3933) <= not (a xor b);
    layer1_outputs(3934) <= a xor b;
    layer1_outputs(3935) <= not b;
    layer1_outputs(3936) <= not b;
    layer1_outputs(3937) <= not (a or b);
    layer1_outputs(3938) <= a or b;
    layer1_outputs(3939) <= a and b;
    layer1_outputs(3940) <= 1'b0;
    layer1_outputs(3941) <= a or b;
    layer1_outputs(3942) <= b;
    layer1_outputs(3943) <= a xor b;
    layer1_outputs(3944) <= not (a and b);
    layer1_outputs(3945) <= a and not b;
    layer1_outputs(3946) <= 1'b0;
    layer1_outputs(3947) <= 1'b1;
    layer1_outputs(3948) <= a and not b;
    layer1_outputs(3949) <= not b or a;
    layer1_outputs(3950) <= not (a or b);
    layer1_outputs(3951) <= a xor b;
    layer1_outputs(3952) <= a and not b;
    layer1_outputs(3953) <= not a;
    layer1_outputs(3954) <= a;
    layer1_outputs(3955) <= b and not a;
    layer1_outputs(3956) <= b and not a;
    layer1_outputs(3957) <= 1'b1;
    layer1_outputs(3958) <= not (a xor b);
    layer1_outputs(3959) <= a and b;
    layer1_outputs(3960) <= a;
    layer1_outputs(3961) <= not a;
    layer1_outputs(3962) <= a and b;
    layer1_outputs(3963) <= a and b;
    layer1_outputs(3964) <= not a;
    layer1_outputs(3965) <= a and not b;
    layer1_outputs(3966) <= b;
    layer1_outputs(3967) <= not a;
    layer1_outputs(3968) <= a and not b;
    layer1_outputs(3969) <= 1'b0;
    layer1_outputs(3970) <= 1'b0;
    layer1_outputs(3971) <= not a;
    layer1_outputs(3972) <= a and b;
    layer1_outputs(3973) <= not (a and b);
    layer1_outputs(3974) <= b;
    layer1_outputs(3975) <= not (a or b);
    layer1_outputs(3976) <= not a;
    layer1_outputs(3977) <= b and not a;
    layer1_outputs(3978) <= not (a or b);
    layer1_outputs(3979) <= b;
    layer1_outputs(3980) <= a xor b;
    layer1_outputs(3981) <= a and not b;
    layer1_outputs(3982) <= a;
    layer1_outputs(3983) <= a and not b;
    layer1_outputs(3984) <= not (a or b);
    layer1_outputs(3985) <= not (a xor b);
    layer1_outputs(3986) <= not b;
    layer1_outputs(3987) <= a and not b;
    layer1_outputs(3988) <= a xor b;
    layer1_outputs(3989) <= not a;
    layer1_outputs(3990) <= a or b;
    layer1_outputs(3991) <= not (a or b);
    layer1_outputs(3992) <= not a;
    layer1_outputs(3993) <= not a;
    layer1_outputs(3994) <= b;
    layer1_outputs(3995) <= not b or a;
    layer1_outputs(3996) <= not b;
    layer1_outputs(3997) <= not a or b;
    layer1_outputs(3998) <= not b;
    layer1_outputs(3999) <= not (a or b);
    layer1_outputs(4000) <= a and b;
    layer1_outputs(4001) <= not (a and b);
    layer1_outputs(4002) <= a and not b;
    layer1_outputs(4003) <= a or b;
    layer1_outputs(4004) <= not a or b;
    layer1_outputs(4005) <= not a;
    layer1_outputs(4006) <= a or b;
    layer1_outputs(4007) <= not a or b;
    layer1_outputs(4008) <= b;
    layer1_outputs(4009) <= 1'b0;
    layer1_outputs(4010) <= 1'b1;
    layer1_outputs(4011) <= not a;
    layer1_outputs(4012) <= b and not a;
    layer1_outputs(4013) <= not (a or b);
    layer1_outputs(4014) <= not a or b;
    layer1_outputs(4015) <= not a;
    layer1_outputs(4016) <= a and not b;
    layer1_outputs(4017) <= a and b;
    layer1_outputs(4018) <= b;
    layer1_outputs(4019) <= a;
    layer1_outputs(4020) <= not (a or b);
    layer1_outputs(4021) <= not a;
    layer1_outputs(4022) <= not b or a;
    layer1_outputs(4023) <= not a or b;
    layer1_outputs(4024) <= a and not b;
    layer1_outputs(4025) <= not (a and b);
    layer1_outputs(4026) <= a xor b;
    layer1_outputs(4027) <= 1'b1;
    layer1_outputs(4028) <= a or b;
    layer1_outputs(4029) <= b;
    layer1_outputs(4030) <= not b or a;
    layer1_outputs(4031) <= a and b;
    layer1_outputs(4032) <= a;
    layer1_outputs(4033) <= not a;
    layer1_outputs(4034) <= a xor b;
    layer1_outputs(4035) <= a and b;
    layer1_outputs(4036) <= not b or a;
    layer1_outputs(4037) <= not b;
    layer1_outputs(4038) <= not b;
    layer1_outputs(4039) <= not (a or b);
    layer1_outputs(4040) <= not (a or b);
    layer1_outputs(4041) <= a and b;
    layer1_outputs(4042) <= b and not a;
    layer1_outputs(4043) <= 1'b1;
    layer1_outputs(4044) <= b;
    layer1_outputs(4045) <= b;
    layer1_outputs(4046) <= a and b;
    layer1_outputs(4047) <= 1'b1;
    layer1_outputs(4048) <= not (a and b);
    layer1_outputs(4049) <= a;
    layer1_outputs(4050) <= 1'b1;
    layer1_outputs(4051) <= a and b;
    layer1_outputs(4052) <= not a;
    layer1_outputs(4053) <= 1'b1;
    layer1_outputs(4054) <= a;
    layer1_outputs(4055) <= 1'b1;
    layer1_outputs(4056) <= not (a or b);
    layer1_outputs(4057) <= b;
    layer1_outputs(4058) <= not a or b;
    layer1_outputs(4059) <= 1'b0;
    layer1_outputs(4060) <= b and not a;
    layer1_outputs(4061) <= a;
    layer1_outputs(4062) <= not a or b;
    layer1_outputs(4063) <= a or b;
    layer1_outputs(4064) <= 1'b1;
    layer1_outputs(4065) <= 1'b1;
    layer1_outputs(4066) <= a;
    layer1_outputs(4067) <= not (a or b);
    layer1_outputs(4068) <= not (a or b);
    layer1_outputs(4069) <= not b or a;
    layer1_outputs(4070) <= a xor b;
    layer1_outputs(4071) <= 1'b1;
    layer1_outputs(4072) <= a and b;
    layer1_outputs(4073) <= not (a or b);
    layer1_outputs(4074) <= not (a or b);
    layer1_outputs(4075) <= a or b;
    layer1_outputs(4076) <= a and not b;
    layer1_outputs(4077) <= a and b;
    layer1_outputs(4078) <= not a;
    layer1_outputs(4079) <= not (a xor b);
    layer1_outputs(4080) <= not a;
    layer1_outputs(4081) <= a or b;
    layer1_outputs(4082) <= not (a and b);
    layer1_outputs(4083) <= 1'b1;
    layer1_outputs(4084) <= a;
    layer1_outputs(4085) <= a or b;
    layer1_outputs(4086) <= a;
    layer1_outputs(4087) <= b and not a;
    layer1_outputs(4088) <= not b or a;
    layer1_outputs(4089) <= not a;
    layer1_outputs(4090) <= not b;
    layer1_outputs(4091) <= not a;
    layer1_outputs(4092) <= not b or a;
    layer1_outputs(4093) <= b;
    layer1_outputs(4094) <= a xor b;
    layer1_outputs(4095) <= b;
    layer1_outputs(4096) <= not a or b;
    layer1_outputs(4097) <= 1'b0;
    layer1_outputs(4098) <= b;
    layer1_outputs(4099) <= not b or a;
    layer1_outputs(4100) <= not b or a;
    layer1_outputs(4101) <= 1'b0;
    layer1_outputs(4102) <= a or b;
    layer1_outputs(4103) <= 1'b0;
    layer1_outputs(4104) <= not (a or b);
    layer1_outputs(4105) <= not a;
    layer1_outputs(4106) <= a;
    layer1_outputs(4107) <= 1'b1;
    layer1_outputs(4108) <= 1'b1;
    layer1_outputs(4109) <= not (a and b);
    layer1_outputs(4110) <= 1'b1;
    layer1_outputs(4111) <= 1'b0;
    layer1_outputs(4112) <= a;
    layer1_outputs(4113) <= 1'b1;
    layer1_outputs(4114) <= not a or b;
    layer1_outputs(4115) <= a or b;
    layer1_outputs(4116) <= not b;
    layer1_outputs(4117) <= not a or b;
    layer1_outputs(4118) <= b;
    layer1_outputs(4119) <= not a or b;
    layer1_outputs(4120) <= b and not a;
    layer1_outputs(4121) <= not a or b;
    layer1_outputs(4122) <= not (a or b);
    layer1_outputs(4123) <= 1'b0;
    layer1_outputs(4124) <= not a;
    layer1_outputs(4125) <= not b or a;
    layer1_outputs(4126) <= 1'b1;
    layer1_outputs(4127) <= not a;
    layer1_outputs(4128) <= not (a and b);
    layer1_outputs(4129) <= a and not b;
    layer1_outputs(4130) <= not b or a;
    layer1_outputs(4131) <= a or b;
    layer1_outputs(4132) <= a;
    layer1_outputs(4133) <= a and b;
    layer1_outputs(4134) <= b and not a;
    layer1_outputs(4135) <= not (a xor b);
    layer1_outputs(4136) <= not (a or b);
    layer1_outputs(4137) <= a xor b;
    layer1_outputs(4138) <= 1'b1;
    layer1_outputs(4139) <= not a;
    layer1_outputs(4140) <= not a;
    layer1_outputs(4141) <= b and not a;
    layer1_outputs(4142) <= a and not b;
    layer1_outputs(4143) <= 1'b0;
    layer1_outputs(4144) <= a or b;
    layer1_outputs(4145) <= a or b;
    layer1_outputs(4146) <= 1'b0;
    layer1_outputs(4147) <= not b or a;
    layer1_outputs(4148) <= not (a and b);
    layer1_outputs(4149) <= a and not b;
    layer1_outputs(4150) <= not a;
    layer1_outputs(4151) <= a xor b;
    layer1_outputs(4152) <= a;
    layer1_outputs(4153) <= not b;
    layer1_outputs(4154) <= not b or a;
    layer1_outputs(4155) <= a;
    layer1_outputs(4156) <= b and not a;
    layer1_outputs(4157) <= 1'b0;
    layer1_outputs(4158) <= a;
    layer1_outputs(4159) <= a;
    layer1_outputs(4160) <= not (a or b);
    layer1_outputs(4161) <= not (a xor b);
    layer1_outputs(4162) <= a and b;
    layer1_outputs(4163) <= not b or a;
    layer1_outputs(4164) <= not a;
    layer1_outputs(4165) <= not b or a;
    layer1_outputs(4166) <= a;
    layer1_outputs(4167) <= not b;
    layer1_outputs(4168) <= 1'b0;
    layer1_outputs(4169) <= a xor b;
    layer1_outputs(4170) <= 1'b1;
    layer1_outputs(4171) <= a and not b;
    layer1_outputs(4172) <= not a or b;
    layer1_outputs(4173) <= a and b;
    layer1_outputs(4174) <= b and not a;
    layer1_outputs(4175) <= not b;
    layer1_outputs(4176) <= b and not a;
    layer1_outputs(4177) <= b and not a;
    layer1_outputs(4178) <= 1'b1;
    layer1_outputs(4179) <= not a or b;
    layer1_outputs(4180) <= 1'b0;
    layer1_outputs(4181) <= not b;
    layer1_outputs(4182) <= a and not b;
    layer1_outputs(4183) <= a and b;
    layer1_outputs(4184) <= b and not a;
    layer1_outputs(4185) <= not (a or b);
    layer1_outputs(4186) <= b and not a;
    layer1_outputs(4187) <= b;
    layer1_outputs(4188) <= b;
    layer1_outputs(4189) <= not a or b;
    layer1_outputs(4190) <= b and not a;
    layer1_outputs(4191) <= b and not a;
    layer1_outputs(4192) <= not a;
    layer1_outputs(4193) <= not b or a;
    layer1_outputs(4194) <= a or b;
    layer1_outputs(4195) <= not (a xor b);
    layer1_outputs(4196) <= b;
    layer1_outputs(4197) <= a;
    layer1_outputs(4198) <= not (a or b);
    layer1_outputs(4199) <= b;
    layer1_outputs(4200) <= not a or b;
    layer1_outputs(4201) <= a;
    layer1_outputs(4202) <= not b;
    layer1_outputs(4203) <= not a;
    layer1_outputs(4204) <= not (a or b);
    layer1_outputs(4205) <= a;
    layer1_outputs(4206) <= not a or b;
    layer1_outputs(4207) <= 1'b0;
    layer1_outputs(4208) <= not b;
    layer1_outputs(4209) <= b and not a;
    layer1_outputs(4210) <= 1'b1;
    layer1_outputs(4211) <= 1'b0;
    layer1_outputs(4212) <= 1'b1;
    layer1_outputs(4213) <= not b;
    layer1_outputs(4214) <= a and not b;
    layer1_outputs(4215) <= b and not a;
    layer1_outputs(4216) <= not b or a;
    layer1_outputs(4217) <= not (a or b);
    layer1_outputs(4218) <= not a;
    layer1_outputs(4219) <= b;
    layer1_outputs(4220) <= b and not a;
    layer1_outputs(4221) <= 1'b1;
    layer1_outputs(4222) <= 1'b0;
    layer1_outputs(4223) <= a and b;
    layer1_outputs(4224) <= 1'b0;
    layer1_outputs(4225) <= not (a or b);
    layer1_outputs(4226) <= a or b;
    layer1_outputs(4227) <= 1'b0;
    layer1_outputs(4228) <= a or b;
    layer1_outputs(4229) <= a or b;
    layer1_outputs(4230) <= b and not a;
    layer1_outputs(4231) <= b;
    layer1_outputs(4232) <= a;
    layer1_outputs(4233) <= not (a or b);
    layer1_outputs(4234) <= not a or b;
    layer1_outputs(4235) <= not a;
    layer1_outputs(4236) <= b and not a;
    layer1_outputs(4237) <= not a or b;
    layer1_outputs(4238) <= not b;
    layer1_outputs(4239) <= not a or b;
    layer1_outputs(4240) <= a and b;
    layer1_outputs(4241) <= b and not a;
    layer1_outputs(4242) <= not b;
    layer1_outputs(4243) <= b;
    layer1_outputs(4244) <= not (a and b);
    layer1_outputs(4245) <= not a or b;
    layer1_outputs(4246) <= not (a xor b);
    layer1_outputs(4247) <= 1'b0;
    layer1_outputs(4248) <= not a or b;
    layer1_outputs(4249) <= a and not b;
    layer1_outputs(4250) <= a and not b;
    layer1_outputs(4251) <= 1'b1;
    layer1_outputs(4252) <= not b or a;
    layer1_outputs(4253) <= b and not a;
    layer1_outputs(4254) <= not a;
    layer1_outputs(4255) <= not (a xor b);
    layer1_outputs(4256) <= 1'b0;
    layer1_outputs(4257) <= not (a or b);
    layer1_outputs(4258) <= a;
    layer1_outputs(4259) <= a and b;
    layer1_outputs(4260) <= 1'b1;
    layer1_outputs(4261) <= b and not a;
    layer1_outputs(4262) <= 1'b0;
    layer1_outputs(4263) <= 1'b1;
    layer1_outputs(4264) <= a and not b;
    layer1_outputs(4265) <= not (a and b);
    layer1_outputs(4266) <= 1'b0;
    layer1_outputs(4267) <= not b;
    layer1_outputs(4268) <= a or b;
    layer1_outputs(4269) <= 1'b0;
    layer1_outputs(4270) <= b and not a;
    layer1_outputs(4271) <= a and not b;
    layer1_outputs(4272) <= 1'b1;
    layer1_outputs(4273) <= a;
    layer1_outputs(4274) <= not b or a;
    layer1_outputs(4275) <= not (a and b);
    layer1_outputs(4276) <= a;
    layer1_outputs(4277) <= 1'b0;
    layer1_outputs(4278) <= not b or a;
    layer1_outputs(4279) <= not (a and b);
    layer1_outputs(4280) <= a or b;
    layer1_outputs(4281) <= not (a or b);
    layer1_outputs(4282) <= a and not b;
    layer1_outputs(4283) <= a;
    layer1_outputs(4284) <= not b or a;
    layer1_outputs(4285) <= a and not b;
    layer1_outputs(4286) <= a or b;
    layer1_outputs(4287) <= a;
    layer1_outputs(4288) <= not (a and b);
    layer1_outputs(4289) <= not (a xor b);
    layer1_outputs(4290) <= a and b;
    layer1_outputs(4291) <= a and not b;
    layer1_outputs(4292) <= a xor b;
    layer1_outputs(4293) <= 1'b1;
    layer1_outputs(4294) <= 1'b0;
    layer1_outputs(4295) <= not (a and b);
    layer1_outputs(4296) <= 1'b1;
    layer1_outputs(4297) <= b and not a;
    layer1_outputs(4298) <= a and not b;
    layer1_outputs(4299) <= 1'b0;
    layer1_outputs(4300) <= a and b;
    layer1_outputs(4301) <= not a;
    layer1_outputs(4302) <= not a;
    layer1_outputs(4303) <= not b or a;
    layer1_outputs(4304) <= not b or a;
    layer1_outputs(4305) <= not (a or b);
    layer1_outputs(4306) <= a or b;
    layer1_outputs(4307) <= 1'b1;
    layer1_outputs(4308) <= not b;
    layer1_outputs(4309) <= b and not a;
    layer1_outputs(4310) <= a and not b;
    layer1_outputs(4311) <= not a;
    layer1_outputs(4312) <= b and not a;
    layer1_outputs(4313) <= a;
    layer1_outputs(4314) <= not b or a;
    layer1_outputs(4315) <= a or b;
    layer1_outputs(4316) <= a and not b;
    layer1_outputs(4317) <= not (a and b);
    layer1_outputs(4318) <= not (a or b);
    layer1_outputs(4319) <= 1'b1;
    layer1_outputs(4320) <= not a;
    layer1_outputs(4321) <= a and b;
    layer1_outputs(4322) <= not b;
    layer1_outputs(4323) <= a and b;
    layer1_outputs(4324) <= b;
    layer1_outputs(4325) <= 1'b0;
    layer1_outputs(4326) <= a;
    layer1_outputs(4327) <= not a;
    layer1_outputs(4328) <= not b or a;
    layer1_outputs(4329) <= not a;
    layer1_outputs(4330) <= not (a and b);
    layer1_outputs(4331) <= a;
    layer1_outputs(4332) <= 1'b1;
    layer1_outputs(4333) <= not b or a;
    layer1_outputs(4334) <= a and b;
    layer1_outputs(4335) <= not a;
    layer1_outputs(4336) <= not (a xor b);
    layer1_outputs(4337) <= not b or a;
    layer1_outputs(4338) <= 1'b0;
    layer1_outputs(4339) <= 1'b1;
    layer1_outputs(4340) <= 1'b0;
    layer1_outputs(4341) <= a and b;
    layer1_outputs(4342) <= 1'b1;
    layer1_outputs(4343) <= a and not b;
    layer1_outputs(4344) <= 1'b1;
    layer1_outputs(4345) <= not b;
    layer1_outputs(4346) <= not a;
    layer1_outputs(4347) <= a and b;
    layer1_outputs(4348) <= b and not a;
    layer1_outputs(4349) <= not a;
    layer1_outputs(4350) <= not (a and b);
    layer1_outputs(4351) <= 1'b1;
    layer1_outputs(4352) <= a and b;
    layer1_outputs(4353) <= not b or a;
    layer1_outputs(4354) <= 1'b0;
    layer1_outputs(4355) <= 1'b0;
    layer1_outputs(4356) <= not a or b;
    layer1_outputs(4357) <= b and not a;
    layer1_outputs(4358) <= a or b;
    layer1_outputs(4359) <= b;
    layer1_outputs(4360) <= b and not a;
    layer1_outputs(4361) <= b;
    layer1_outputs(4362) <= not (a xor b);
    layer1_outputs(4363) <= not a or b;
    layer1_outputs(4364) <= b;
    layer1_outputs(4365) <= a;
    layer1_outputs(4366) <= 1'b0;
    layer1_outputs(4367) <= not (a or b);
    layer1_outputs(4368) <= a and not b;
    layer1_outputs(4369) <= not a;
    layer1_outputs(4370) <= 1'b1;
    layer1_outputs(4371) <= b and not a;
    layer1_outputs(4372) <= b;
    layer1_outputs(4373) <= not (a and b);
    layer1_outputs(4374) <= a and b;
    layer1_outputs(4375) <= 1'b1;
    layer1_outputs(4376) <= not a or b;
    layer1_outputs(4377) <= not (a and b);
    layer1_outputs(4378) <= b and not a;
    layer1_outputs(4379) <= not b;
    layer1_outputs(4380) <= a;
    layer1_outputs(4381) <= a and b;
    layer1_outputs(4382) <= b and not a;
    layer1_outputs(4383) <= not a or b;
    layer1_outputs(4384) <= not b or a;
    layer1_outputs(4385) <= not (a or b);
    layer1_outputs(4386) <= a and b;
    layer1_outputs(4387) <= 1'b0;
    layer1_outputs(4388) <= a;
    layer1_outputs(4389) <= 1'b0;
    layer1_outputs(4390) <= a and not b;
    layer1_outputs(4391) <= a and not b;
    layer1_outputs(4392) <= b and not a;
    layer1_outputs(4393) <= not b or a;
    layer1_outputs(4394) <= a;
    layer1_outputs(4395) <= a;
    layer1_outputs(4396) <= b;
    layer1_outputs(4397) <= a;
    layer1_outputs(4398) <= 1'b0;
    layer1_outputs(4399) <= 1'b1;
    layer1_outputs(4400) <= not b or a;
    layer1_outputs(4401) <= 1'b1;
    layer1_outputs(4402) <= not a;
    layer1_outputs(4403) <= not a or b;
    layer1_outputs(4404) <= not (a or b);
    layer1_outputs(4405) <= a;
    layer1_outputs(4406) <= b and not a;
    layer1_outputs(4407) <= b;
    layer1_outputs(4408) <= 1'b0;
    layer1_outputs(4409) <= a and not b;
    layer1_outputs(4410) <= not a;
    layer1_outputs(4411) <= not a;
    layer1_outputs(4412) <= a;
    layer1_outputs(4413) <= not (a or b);
    layer1_outputs(4414) <= not (a or b);
    layer1_outputs(4415) <= not (a xor b);
    layer1_outputs(4416) <= a;
    layer1_outputs(4417) <= not a;
    layer1_outputs(4418) <= not b or a;
    layer1_outputs(4419) <= not a;
    layer1_outputs(4420) <= not (a or b);
    layer1_outputs(4421) <= not a or b;
    layer1_outputs(4422) <= not (a and b);
    layer1_outputs(4423) <= not b;
    layer1_outputs(4424) <= b and not a;
    layer1_outputs(4425) <= a xor b;
    layer1_outputs(4426) <= 1'b0;
    layer1_outputs(4427) <= 1'b1;
    layer1_outputs(4428) <= not b;
    layer1_outputs(4429) <= 1'b0;
    layer1_outputs(4430) <= b;
    layer1_outputs(4431) <= a;
    layer1_outputs(4432) <= not a or b;
    layer1_outputs(4433) <= a and not b;
    layer1_outputs(4434) <= b and not a;
    layer1_outputs(4435) <= a xor b;
    layer1_outputs(4436) <= not b or a;
    layer1_outputs(4437) <= 1'b1;
    layer1_outputs(4438) <= 1'b0;
    layer1_outputs(4439) <= not (a and b);
    layer1_outputs(4440) <= not b;
    layer1_outputs(4441) <= not b;
    layer1_outputs(4442) <= a and b;
    layer1_outputs(4443) <= b and not a;
    layer1_outputs(4444) <= not a;
    layer1_outputs(4445) <= a;
    layer1_outputs(4446) <= b and not a;
    layer1_outputs(4447) <= a;
    layer1_outputs(4448) <= not (a or b);
    layer1_outputs(4449) <= a and not b;
    layer1_outputs(4450) <= a and b;
    layer1_outputs(4451) <= not b or a;
    layer1_outputs(4452) <= not (a and b);
    layer1_outputs(4453) <= b and not a;
    layer1_outputs(4454) <= b;
    layer1_outputs(4455) <= a and not b;
    layer1_outputs(4456) <= a and not b;
    layer1_outputs(4457) <= not (a and b);
    layer1_outputs(4458) <= not (a and b);
    layer1_outputs(4459) <= a and not b;
    layer1_outputs(4460) <= b;
    layer1_outputs(4461) <= not (a or b);
    layer1_outputs(4462) <= b;
    layer1_outputs(4463) <= 1'b0;
    layer1_outputs(4464) <= a and not b;
    layer1_outputs(4465) <= not a or b;
    layer1_outputs(4466) <= not (a or b);
    layer1_outputs(4467) <= a or b;
    layer1_outputs(4468) <= a and not b;
    layer1_outputs(4469) <= 1'b0;
    layer1_outputs(4470) <= a;
    layer1_outputs(4471) <= not (a or b);
    layer1_outputs(4472) <= not (a or b);
    layer1_outputs(4473) <= a and b;
    layer1_outputs(4474) <= 1'b0;
    layer1_outputs(4475) <= not a or b;
    layer1_outputs(4476) <= 1'b1;
    layer1_outputs(4477) <= a or b;
    layer1_outputs(4478) <= a and not b;
    layer1_outputs(4479) <= not (a and b);
    layer1_outputs(4480) <= a xor b;
    layer1_outputs(4481) <= not a;
    layer1_outputs(4482) <= a and not b;
    layer1_outputs(4483) <= a and b;
    layer1_outputs(4484) <= a;
    layer1_outputs(4485) <= a or b;
    layer1_outputs(4486) <= b;
    layer1_outputs(4487) <= not a;
    layer1_outputs(4488) <= not a;
    layer1_outputs(4489) <= not a or b;
    layer1_outputs(4490) <= not a;
    layer1_outputs(4491) <= a and b;
    layer1_outputs(4492) <= a;
    layer1_outputs(4493) <= a and not b;
    layer1_outputs(4494) <= a or b;
    layer1_outputs(4495) <= not (a or b);
    layer1_outputs(4496) <= a and b;
    layer1_outputs(4497) <= a or b;
    layer1_outputs(4498) <= not b or a;
    layer1_outputs(4499) <= not b or a;
    layer1_outputs(4500) <= not b;
    layer1_outputs(4501) <= a and b;
    layer1_outputs(4502) <= 1'b0;
    layer1_outputs(4503) <= not (a or b);
    layer1_outputs(4504) <= b and not a;
    layer1_outputs(4505) <= b and not a;
    layer1_outputs(4506) <= not b or a;
    layer1_outputs(4507) <= 1'b0;
    layer1_outputs(4508) <= not b;
    layer1_outputs(4509) <= not a or b;
    layer1_outputs(4510) <= a;
    layer1_outputs(4511) <= not (a xor b);
    layer1_outputs(4512) <= not (a and b);
    layer1_outputs(4513) <= not b;
    layer1_outputs(4514) <= not (a and b);
    layer1_outputs(4515) <= not a or b;
    layer1_outputs(4516) <= b and not a;
    layer1_outputs(4517) <= 1'b0;
    layer1_outputs(4518) <= b and not a;
    layer1_outputs(4519) <= not (a xor b);
    layer1_outputs(4520) <= not a;
    layer1_outputs(4521) <= not (a and b);
    layer1_outputs(4522) <= b and not a;
    layer1_outputs(4523) <= 1'b0;
    layer1_outputs(4524) <= not b;
    layer1_outputs(4525) <= a;
    layer1_outputs(4526) <= b;
    layer1_outputs(4527) <= a or b;
    layer1_outputs(4528) <= a and not b;
    layer1_outputs(4529) <= not a;
    layer1_outputs(4530) <= not (a or b);
    layer1_outputs(4531) <= 1'b1;
    layer1_outputs(4532) <= not b;
    layer1_outputs(4533) <= 1'b0;
    layer1_outputs(4534) <= not a or b;
    layer1_outputs(4535) <= a xor b;
    layer1_outputs(4536) <= b and not a;
    layer1_outputs(4537) <= a or b;
    layer1_outputs(4538) <= b;
    layer1_outputs(4539) <= a;
    layer1_outputs(4540) <= a and b;
    layer1_outputs(4541) <= not a;
    layer1_outputs(4542) <= 1'b1;
    layer1_outputs(4543) <= not (a and b);
    layer1_outputs(4544) <= 1'b1;
    layer1_outputs(4545) <= b;
    layer1_outputs(4546) <= 1'b1;
    layer1_outputs(4547) <= not b;
    layer1_outputs(4548) <= not a or b;
    layer1_outputs(4549) <= b;
    layer1_outputs(4550) <= a and b;
    layer1_outputs(4551) <= a;
    layer1_outputs(4552) <= not a or b;
    layer1_outputs(4553) <= not a or b;
    layer1_outputs(4554) <= 1'b0;
    layer1_outputs(4555) <= a and not b;
    layer1_outputs(4556) <= a or b;
    layer1_outputs(4557) <= a and b;
    layer1_outputs(4558) <= a and not b;
    layer1_outputs(4559) <= not (a xor b);
    layer1_outputs(4560) <= b;
    layer1_outputs(4561) <= not b;
    layer1_outputs(4562) <= a;
    layer1_outputs(4563) <= not b;
    layer1_outputs(4564) <= a and not b;
    layer1_outputs(4565) <= not a;
    layer1_outputs(4566) <= not (a or b);
    layer1_outputs(4567) <= 1'b1;
    layer1_outputs(4568) <= not b;
    layer1_outputs(4569) <= not a or b;
    layer1_outputs(4570) <= b and not a;
    layer1_outputs(4571) <= 1'b0;
    layer1_outputs(4572) <= not (a or b);
    layer1_outputs(4573) <= b and not a;
    layer1_outputs(4574) <= not a or b;
    layer1_outputs(4575) <= a and b;
    layer1_outputs(4576) <= not b or a;
    layer1_outputs(4577) <= not b or a;
    layer1_outputs(4578) <= not b;
    layer1_outputs(4579) <= a;
    layer1_outputs(4580) <= not a;
    layer1_outputs(4581) <= a and b;
    layer1_outputs(4582) <= not (a xor b);
    layer1_outputs(4583) <= not (a xor b);
    layer1_outputs(4584) <= a and b;
    layer1_outputs(4585) <= not b or a;
    layer1_outputs(4586) <= 1'b0;
    layer1_outputs(4587) <= a or b;
    layer1_outputs(4588) <= a and not b;
    layer1_outputs(4589) <= 1'b1;
    layer1_outputs(4590) <= a or b;
    layer1_outputs(4591) <= a or b;
    layer1_outputs(4592) <= a;
    layer1_outputs(4593) <= not (a or b);
    layer1_outputs(4594) <= 1'b1;
    layer1_outputs(4595) <= not a;
    layer1_outputs(4596) <= not (a xor b);
    layer1_outputs(4597) <= a xor b;
    layer1_outputs(4598) <= a and not b;
    layer1_outputs(4599) <= a;
    layer1_outputs(4600) <= not b or a;
    layer1_outputs(4601) <= a;
    layer1_outputs(4602) <= not a;
    layer1_outputs(4603) <= not (a or b);
    layer1_outputs(4604) <= b;
    layer1_outputs(4605) <= a or b;
    layer1_outputs(4606) <= not b;
    layer1_outputs(4607) <= a or b;
    layer1_outputs(4608) <= b;
    layer1_outputs(4609) <= a;
    layer1_outputs(4610) <= a and b;
    layer1_outputs(4611) <= 1'b0;
    layer1_outputs(4612) <= a and b;
    layer1_outputs(4613) <= 1'b0;
    layer1_outputs(4614) <= not b or a;
    layer1_outputs(4615) <= 1'b1;
    layer1_outputs(4616) <= not a;
    layer1_outputs(4617) <= not b or a;
    layer1_outputs(4618) <= 1'b1;
    layer1_outputs(4619) <= not (a or b);
    layer1_outputs(4620) <= not b or a;
    layer1_outputs(4621) <= not a;
    layer1_outputs(4622) <= not (a or b);
    layer1_outputs(4623) <= not b or a;
    layer1_outputs(4624) <= not a;
    layer1_outputs(4625) <= not (a or b);
    layer1_outputs(4626) <= 1'b1;
    layer1_outputs(4627) <= not (a or b);
    layer1_outputs(4628) <= not b;
    layer1_outputs(4629) <= b;
    layer1_outputs(4630) <= a or b;
    layer1_outputs(4631) <= not a or b;
    layer1_outputs(4632) <= 1'b0;
    layer1_outputs(4633) <= 1'b1;
    layer1_outputs(4634) <= b;
    layer1_outputs(4635) <= not a or b;
    layer1_outputs(4636) <= not a;
    layer1_outputs(4637) <= b and not a;
    layer1_outputs(4638) <= not a or b;
    layer1_outputs(4639) <= not (a or b);
    layer1_outputs(4640) <= not a or b;
    layer1_outputs(4641) <= b and not a;
    layer1_outputs(4642) <= 1'b0;
    layer1_outputs(4643) <= not (a or b);
    layer1_outputs(4644) <= a;
    layer1_outputs(4645) <= not a;
    layer1_outputs(4646) <= not b;
    layer1_outputs(4647) <= not b;
    layer1_outputs(4648) <= a;
    layer1_outputs(4649) <= a and not b;
    layer1_outputs(4650) <= not (a or b);
    layer1_outputs(4651) <= not b or a;
    layer1_outputs(4652) <= not b;
    layer1_outputs(4653) <= not (a and b);
    layer1_outputs(4654) <= a xor b;
    layer1_outputs(4655) <= not (a or b);
    layer1_outputs(4656) <= not a;
    layer1_outputs(4657) <= not b;
    layer1_outputs(4658) <= not (a and b);
    layer1_outputs(4659) <= a xor b;
    layer1_outputs(4660) <= a and not b;
    layer1_outputs(4661) <= b;
    layer1_outputs(4662) <= a xor b;
    layer1_outputs(4663) <= a;
    layer1_outputs(4664) <= not (a and b);
    layer1_outputs(4665) <= b and not a;
    layer1_outputs(4666) <= a and b;
    layer1_outputs(4667) <= a and not b;
    layer1_outputs(4668) <= b and not a;
    layer1_outputs(4669) <= not (a or b);
    layer1_outputs(4670) <= not a;
    layer1_outputs(4671) <= not (a and b);
    layer1_outputs(4672) <= a and not b;
    layer1_outputs(4673) <= not (a or b);
    layer1_outputs(4674) <= a;
    layer1_outputs(4675) <= 1'b0;
    layer1_outputs(4676) <= 1'b1;
    layer1_outputs(4677) <= not a;
    layer1_outputs(4678) <= a or b;
    layer1_outputs(4679) <= a and b;
    layer1_outputs(4680) <= not a;
    layer1_outputs(4681) <= 1'b0;
    layer1_outputs(4682) <= not a or b;
    layer1_outputs(4683) <= 1'b1;
    layer1_outputs(4684) <= not a or b;
    layer1_outputs(4685) <= not (a or b);
    layer1_outputs(4686) <= a or b;
    layer1_outputs(4687) <= not a or b;
    layer1_outputs(4688) <= not a or b;
    layer1_outputs(4689) <= a or b;
    layer1_outputs(4690) <= 1'b0;
    layer1_outputs(4691) <= 1'b0;
    layer1_outputs(4692) <= a or b;
    layer1_outputs(4693) <= not (a and b);
    layer1_outputs(4694) <= not a or b;
    layer1_outputs(4695) <= a;
    layer1_outputs(4696) <= a;
    layer1_outputs(4697) <= a or b;
    layer1_outputs(4698) <= 1'b0;
    layer1_outputs(4699) <= b and not a;
    layer1_outputs(4700) <= a and not b;
    layer1_outputs(4701) <= not (a and b);
    layer1_outputs(4702) <= not a or b;
    layer1_outputs(4703) <= not (a xor b);
    layer1_outputs(4704) <= not a;
    layer1_outputs(4705) <= not a or b;
    layer1_outputs(4706) <= b and not a;
    layer1_outputs(4707) <= not a or b;
    layer1_outputs(4708) <= 1'b1;
    layer1_outputs(4709) <= not b;
    layer1_outputs(4710) <= b and not a;
    layer1_outputs(4711) <= 1'b1;
    layer1_outputs(4712) <= 1'b0;
    layer1_outputs(4713) <= not (a or b);
    layer1_outputs(4714) <= 1'b0;
    layer1_outputs(4715) <= b and not a;
    layer1_outputs(4716) <= not a or b;
    layer1_outputs(4717) <= b;
    layer1_outputs(4718) <= not (a and b);
    layer1_outputs(4719) <= 1'b0;
    layer1_outputs(4720) <= 1'b1;
    layer1_outputs(4721) <= a and not b;
    layer1_outputs(4722) <= a and b;
    layer1_outputs(4723) <= not b or a;
    layer1_outputs(4724) <= b and not a;
    layer1_outputs(4725) <= not a;
    layer1_outputs(4726) <= not a or b;
    layer1_outputs(4727) <= a and not b;
    layer1_outputs(4728) <= 1'b1;
    layer1_outputs(4729) <= b;
    layer1_outputs(4730) <= not a;
    layer1_outputs(4731) <= not b;
    layer1_outputs(4732) <= 1'b0;
    layer1_outputs(4733) <= a and b;
    layer1_outputs(4734) <= a and not b;
    layer1_outputs(4735) <= 1'b1;
    layer1_outputs(4736) <= b;
    layer1_outputs(4737) <= not b or a;
    layer1_outputs(4738) <= 1'b1;
    layer1_outputs(4739) <= b and not a;
    layer1_outputs(4740) <= a;
    layer1_outputs(4741) <= a xor b;
    layer1_outputs(4742) <= b;
    layer1_outputs(4743) <= a or b;
    layer1_outputs(4744) <= not b;
    layer1_outputs(4745) <= b;
    layer1_outputs(4746) <= 1'b1;
    layer1_outputs(4747) <= a and not b;
    layer1_outputs(4748) <= a and b;
    layer1_outputs(4749) <= not a or b;
    layer1_outputs(4750) <= 1'b1;
    layer1_outputs(4751) <= a;
    layer1_outputs(4752) <= a or b;
    layer1_outputs(4753) <= 1'b0;
    layer1_outputs(4754) <= not a or b;
    layer1_outputs(4755) <= not a;
    layer1_outputs(4756) <= b;
    layer1_outputs(4757) <= 1'b0;
    layer1_outputs(4758) <= 1'b0;
    layer1_outputs(4759) <= not b or a;
    layer1_outputs(4760) <= b and not a;
    layer1_outputs(4761) <= not (a or b);
    layer1_outputs(4762) <= b;
    layer1_outputs(4763) <= not a or b;
    layer1_outputs(4764) <= a or b;
    layer1_outputs(4765) <= not (a and b);
    layer1_outputs(4766) <= not b;
    layer1_outputs(4767) <= 1'b0;
    layer1_outputs(4768) <= a or b;
    layer1_outputs(4769) <= a;
    layer1_outputs(4770) <= 1'b0;
    layer1_outputs(4771) <= not a or b;
    layer1_outputs(4772) <= not b;
    layer1_outputs(4773) <= not (a xor b);
    layer1_outputs(4774) <= not a or b;
    layer1_outputs(4775) <= a and b;
    layer1_outputs(4776) <= a and b;
    layer1_outputs(4777) <= 1'b0;
    layer1_outputs(4778) <= 1'b1;
    layer1_outputs(4779) <= 1'b0;
    layer1_outputs(4780) <= not a;
    layer1_outputs(4781) <= not a or b;
    layer1_outputs(4782) <= 1'b1;
    layer1_outputs(4783) <= b;
    layer1_outputs(4784) <= a xor b;
    layer1_outputs(4785) <= not b or a;
    layer1_outputs(4786) <= 1'b0;
    layer1_outputs(4787) <= a and not b;
    layer1_outputs(4788) <= a and not b;
    layer1_outputs(4789) <= a and b;
    layer1_outputs(4790) <= 1'b0;
    layer1_outputs(4791) <= a or b;
    layer1_outputs(4792) <= 1'b0;
    layer1_outputs(4793) <= not (a and b);
    layer1_outputs(4794) <= not a;
    layer1_outputs(4795) <= not a;
    layer1_outputs(4796) <= a and b;
    layer1_outputs(4797) <= not b;
    layer1_outputs(4798) <= not (a xor b);
    layer1_outputs(4799) <= not (a xor b);
    layer1_outputs(4800) <= a and not b;
    layer1_outputs(4801) <= a and not b;
    layer1_outputs(4802) <= a or b;
    layer1_outputs(4803) <= not a;
    layer1_outputs(4804) <= not (a and b);
    layer1_outputs(4805) <= 1'b0;
    layer1_outputs(4806) <= not (a or b);
    layer1_outputs(4807) <= not a or b;
    layer1_outputs(4808) <= not b;
    layer1_outputs(4809) <= a or b;
    layer1_outputs(4810) <= not (a and b);
    layer1_outputs(4811) <= not (a or b);
    layer1_outputs(4812) <= 1'b0;
    layer1_outputs(4813) <= not (a and b);
    layer1_outputs(4814) <= not a;
    layer1_outputs(4815) <= a and b;
    layer1_outputs(4816) <= not a;
    layer1_outputs(4817) <= not (a or b);
    layer1_outputs(4818) <= not b;
    layer1_outputs(4819) <= b;
    layer1_outputs(4820) <= not b or a;
    layer1_outputs(4821) <= b;
    layer1_outputs(4822) <= a xor b;
    layer1_outputs(4823) <= b and not a;
    layer1_outputs(4824) <= a and not b;
    layer1_outputs(4825) <= b;
    layer1_outputs(4826) <= not b;
    layer1_outputs(4827) <= a and not b;
    layer1_outputs(4828) <= not a or b;
    layer1_outputs(4829) <= a;
    layer1_outputs(4830) <= not b;
    layer1_outputs(4831) <= not a;
    layer1_outputs(4832) <= 1'b1;
    layer1_outputs(4833) <= 1'b0;
    layer1_outputs(4834) <= 1'b0;
    layer1_outputs(4835) <= not (a or b);
    layer1_outputs(4836) <= not a or b;
    layer1_outputs(4837) <= a and not b;
    layer1_outputs(4838) <= 1'b0;
    layer1_outputs(4839) <= a xor b;
    layer1_outputs(4840) <= 1'b0;
    layer1_outputs(4841) <= a and b;
    layer1_outputs(4842) <= a and b;
    layer1_outputs(4843) <= not a;
    layer1_outputs(4844) <= 1'b0;
    layer1_outputs(4845) <= 1'b1;
    layer1_outputs(4846) <= b and not a;
    layer1_outputs(4847) <= b and not a;
    layer1_outputs(4848) <= not (a or b);
    layer1_outputs(4849) <= a;
    layer1_outputs(4850) <= not (a or b);
    layer1_outputs(4851) <= b and not a;
    layer1_outputs(4852) <= not (a and b);
    layer1_outputs(4853) <= 1'b0;
    layer1_outputs(4854) <= 1'b1;
    layer1_outputs(4855) <= a;
    layer1_outputs(4856) <= 1'b0;
    layer1_outputs(4857) <= not b or a;
    layer1_outputs(4858) <= a xor b;
    layer1_outputs(4859) <= not b or a;
    layer1_outputs(4860) <= not a;
    layer1_outputs(4861) <= not b or a;
    layer1_outputs(4862) <= 1'b0;
    layer1_outputs(4863) <= 1'b1;
    layer1_outputs(4864) <= b and not a;
    layer1_outputs(4865) <= a and b;
    layer1_outputs(4866) <= a and b;
    layer1_outputs(4867) <= 1'b1;
    layer1_outputs(4868) <= a;
    layer1_outputs(4869) <= not (a xor b);
    layer1_outputs(4870) <= a xor b;
    layer1_outputs(4871) <= not b;
    layer1_outputs(4872) <= not (a xor b);
    layer1_outputs(4873) <= b and not a;
    layer1_outputs(4874) <= not (a and b);
    layer1_outputs(4875) <= not a or b;
    layer1_outputs(4876) <= a;
    layer1_outputs(4877) <= not (a or b);
    layer1_outputs(4878) <= 1'b0;
    layer1_outputs(4879) <= not (a and b);
    layer1_outputs(4880) <= a;
    layer1_outputs(4881) <= not b or a;
    layer1_outputs(4882) <= b;
    layer1_outputs(4883) <= not a or b;
    layer1_outputs(4884) <= b and not a;
    layer1_outputs(4885) <= 1'b0;
    layer1_outputs(4886) <= b and not a;
    layer1_outputs(4887) <= not (a and b);
    layer1_outputs(4888) <= a or b;
    layer1_outputs(4889) <= b;
    layer1_outputs(4890) <= b and not a;
    layer1_outputs(4891) <= a xor b;
    layer1_outputs(4892) <= 1'b0;
    layer1_outputs(4893) <= 1'b0;
    layer1_outputs(4894) <= b and not a;
    layer1_outputs(4895) <= 1'b1;
    layer1_outputs(4896) <= 1'b0;
    layer1_outputs(4897) <= b;
    layer1_outputs(4898) <= not (a and b);
    layer1_outputs(4899) <= b;
    layer1_outputs(4900) <= not (a or b);
    layer1_outputs(4901) <= b;
    layer1_outputs(4902) <= a;
    layer1_outputs(4903) <= 1'b0;
    layer1_outputs(4904) <= a or b;
    layer1_outputs(4905) <= a;
    layer1_outputs(4906) <= 1'b0;
    layer1_outputs(4907) <= a or b;
    layer1_outputs(4908) <= not (a and b);
    layer1_outputs(4909) <= not b;
    layer1_outputs(4910) <= 1'b0;
    layer1_outputs(4911) <= b and not a;
    layer1_outputs(4912) <= a or b;
    layer1_outputs(4913) <= a xor b;
    layer1_outputs(4914) <= not b or a;
    layer1_outputs(4915) <= b;
    layer1_outputs(4916) <= a and b;
    layer1_outputs(4917) <= not (a and b);
    layer1_outputs(4918) <= not (a and b);
    layer1_outputs(4919) <= b;
    layer1_outputs(4920) <= not a;
    layer1_outputs(4921) <= 1'b1;
    layer1_outputs(4922) <= not a;
    layer1_outputs(4923) <= not b;
    layer1_outputs(4924) <= not a or b;
    layer1_outputs(4925) <= not b;
    layer1_outputs(4926) <= a and not b;
    layer1_outputs(4927) <= a and not b;
    layer1_outputs(4928) <= a;
    layer1_outputs(4929) <= a or b;
    layer1_outputs(4930) <= not (a or b);
    layer1_outputs(4931) <= not (a xor b);
    layer1_outputs(4932) <= 1'b1;
    layer1_outputs(4933) <= 1'b0;
    layer1_outputs(4934) <= not a;
    layer1_outputs(4935) <= a or b;
    layer1_outputs(4936) <= 1'b0;
    layer1_outputs(4937) <= a;
    layer1_outputs(4938) <= a and not b;
    layer1_outputs(4939) <= a and b;
    layer1_outputs(4940) <= not (a and b);
    layer1_outputs(4941) <= not b;
    layer1_outputs(4942) <= 1'b1;
    layer1_outputs(4943) <= 1'b0;
    layer1_outputs(4944) <= a and not b;
    layer1_outputs(4945) <= not a or b;
    layer1_outputs(4946) <= a and b;
    layer1_outputs(4947) <= a;
    layer1_outputs(4948) <= a and b;
    layer1_outputs(4949) <= not a or b;
    layer1_outputs(4950) <= 1'b1;
    layer1_outputs(4951) <= a or b;
    layer1_outputs(4952) <= a and b;
    layer1_outputs(4953) <= a or b;
    layer1_outputs(4954) <= b;
    layer1_outputs(4955) <= a and not b;
    layer1_outputs(4956) <= 1'b0;
    layer1_outputs(4957) <= not a;
    layer1_outputs(4958) <= a and not b;
    layer1_outputs(4959) <= a or b;
    layer1_outputs(4960) <= not (a or b);
    layer1_outputs(4961) <= not b;
    layer1_outputs(4962) <= not a or b;
    layer1_outputs(4963) <= a xor b;
    layer1_outputs(4964) <= a;
    layer1_outputs(4965) <= a xor b;
    layer1_outputs(4966) <= a or b;
    layer1_outputs(4967) <= a and b;
    layer1_outputs(4968) <= 1'b1;
    layer1_outputs(4969) <= a and b;
    layer1_outputs(4970) <= not b or a;
    layer1_outputs(4971) <= 1'b1;
    layer1_outputs(4972) <= not a;
    layer1_outputs(4973) <= 1'b0;
    layer1_outputs(4974) <= 1'b0;
    layer1_outputs(4975) <= 1'b1;
    layer1_outputs(4976) <= not b or a;
    layer1_outputs(4977) <= not (a and b);
    layer1_outputs(4978) <= b;
    layer1_outputs(4979) <= b and not a;
    layer1_outputs(4980) <= 1'b1;
    layer1_outputs(4981) <= b and not a;
    layer1_outputs(4982) <= a or b;
    layer1_outputs(4983) <= b;
    layer1_outputs(4984) <= a and not b;
    layer1_outputs(4985) <= not b;
    layer1_outputs(4986) <= not b or a;
    layer1_outputs(4987) <= a xor b;
    layer1_outputs(4988) <= b and not a;
    layer1_outputs(4989) <= not b or a;
    layer1_outputs(4990) <= not a or b;
    layer1_outputs(4991) <= not b or a;
    layer1_outputs(4992) <= 1'b1;
    layer1_outputs(4993) <= a and not b;
    layer1_outputs(4994) <= b and not a;
    layer1_outputs(4995) <= a or b;
    layer1_outputs(4996) <= a and not b;
    layer1_outputs(4997) <= not a;
    layer1_outputs(4998) <= not b;
    layer1_outputs(4999) <= not a;
    layer1_outputs(5000) <= 1'b1;
    layer1_outputs(5001) <= 1'b1;
    layer1_outputs(5002) <= not a or b;
    layer1_outputs(5003) <= 1'b1;
    layer1_outputs(5004) <= a or b;
    layer1_outputs(5005) <= a and not b;
    layer1_outputs(5006) <= 1'b1;
    layer1_outputs(5007) <= a and not b;
    layer1_outputs(5008) <= b;
    layer1_outputs(5009) <= not (a or b);
    layer1_outputs(5010) <= a;
    layer1_outputs(5011) <= not b or a;
    layer1_outputs(5012) <= a xor b;
    layer1_outputs(5013) <= 1'b1;
    layer1_outputs(5014) <= not b;
    layer1_outputs(5015) <= a;
    layer1_outputs(5016) <= not (a and b);
    layer1_outputs(5017) <= b;
    layer1_outputs(5018) <= a or b;
    layer1_outputs(5019) <= a and b;
    layer1_outputs(5020) <= not (a or b);
    layer1_outputs(5021) <= not b;
    layer1_outputs(5022) <= 1'b0;
    layer1_outputs(5023) <= 1'b1;
    layer1_outputs(5024) <= b and not a;
    layer1_outputs(5025) <= not a;
    layer1_outputs(5026) <= 1'b0;
    layer1_outputs(5027) <= a;
    layer1_outputs(5028) <= 1'b1;
    layer1_outputs(5029) <= 1'b0;
    layer1_outputs(5030) <= not b;
    layer1_outputs(5031) <= 1'b1;
    layer1_outputs(5032) <= a or b;
    layer1_outputs(5033) <= a and b;
    layer1_outputs(5034) <= not a;
    layer1_outputs(5035) <= not (a and b);
    layer1_outputs(5036) <= 1'b0;
    layer1_outputs(5037) <= 1'b1;
    layer1_outputs(5038) <= not b;
    layer1_outputs(5039) <= 1'b0;
    layer1_outputs(5040) <= b and not a;
    layer1_outputs(5041) <= a;
    layer1_outputs(5042) <= b and not a;
    layer1_outputs(5043) <= a;
    layer1_outputs(5044) <= b;
    layer1_outputs(5045) <= a;
    layer1_outputs(5046) <= a or b;
    layer1_outputs(5047) <= not b;
    layer1_outputs(5048) <= a and not b;
    layer1_outputs(5049) <= not b;
    layer1_outputs(5050) <= b and not a;
    layer1_outputs(5051) <= not a or b;
    layer1_outputs(5052) <= b;
    layer1_outputs(5053) <= not (a or b);
    layer1_outputs(5054) <= not b;
    layer1_outputs(5055) <= b and not a;
    layer1_outputs(5056) <= 1'b1;
    layer1_outputs(5057) <= not b or a;
    layer1_outputs(5058) <= not a;
    layer1_outputs(5059) <= a and b;
    layer1_outputs(5060) <= a or b;
    layer1_outputs(5061) <= not (a and b);
    layer1_outputs(5062) <= not b;
    layer1_outputs(5063) <= 1'b1;
    layer1_outputs(5064) <= not b or a;
    layer1_outputs(5065) <= b and not a;
    layer1_outputs(5066) <= not b or a;
    layer1_outputs(5067) <= 1'b0;
    layer1_outputs(5068) <= not b;
    layer1_outputs(5069) <= b;
    layer1_outputs(5070) <= not (a or b);
    layer1_outputs(5071) <= a and b;
    layer1_outputs(5072) <= not a;
    layer1_outputs(5073) <= a and not b;
    layer1_outputs(5074) <= not a or b;
    layer1_outputs(5075) <= not a;
    layer1_outputs(5076) <= b and not a;
    layer1_outputs(5077) <= not b;
    layer1_outputs(5078) <= 1'b0;
    layer1_outputs(5079) <= not a;
    layer1_outputs(5080) <= a xor b;
    layer1_outputs(5081) <= not a;
    layer1_outputs(5082) <= not (a or b);
    layer1_outputs(5083) <= not (a or b);
    layer1_outputs(5084) <= not b or a;
    layer1_outputs(5085) <= a and b;
    layer1_outputs(5086) <= b;
    layer1_outputs(5087) <= a;
    layer1_outputs(5088) <= a or b;
    layer1_outputs(5089) <= a or b;
    layer1_outputs(5090) <= not a;
    layer1_outputs(5091) <= b;
    layer1_outputs(5092) <= not (a xor b);
    layer1_outputs(5093) <= a or b;
    layer1_outputs(5094) <= not a;
    layer1_outputs(5095) <= b;
    layer1_outputs(5096) <= 1'b1;
    layer1_outputs(5097) <= not a or b;
    layer1_outputs(5098) <= a and b;
    layer1_outputs(5099) <= b;
    layer1_outputs(5100) <= not a or b;
    layer1_outputs(5101) <= b;
    layer1_outputs(5102) <= not (a or b);
    layer1_outputs(5103) <= not a or b;
    layer1_outputs(5104) <= not (a and b);
    layer1_outputs(5105) <= a and b;
    layer1_outputs(5106) <= not a;
    layer1_outputs(5107) <= not (a xor b);
    layer1_outputs(5108) <= 1'b0;
    layer1_outputs(5109) <= a or b;
    layer1_outputs(5110) <= a or b;
    layer1_outputs(5111) <= not (a and b);
    layer1_outputs(5112) <= a and b;
    layer1_outputs(5113) <= not (a xor b);
    layer1_outputs(5114) <= a and not b;
    layer1_outputs(5115) <= not b;
    layer1_outputs(5116) <= a and b;
    layer1_outputs(5117) <= 1'b0;
    layer1_outputs(5118) <= 1'b0;
    layer1_outputs(5119) <= a and b;
    layer1_outputs(5120) <= 1'b0;
    layer1_outputs(5121) <= b and not a;
    layer1_outputs(5122) <= not a or b;
    layer1_outputs(5123) <= not b or a;
    layer1_outputs(5124) <= not b or a;
    layer1_outputs(5125) <= not a;
    layer1_outputs(5126) <= a xor b;
    layer1_outputs(5127) <= 1'b1;
    layer1_outputs(5128) <= b and not a;
    layer1_outputs(5129) <= not (a or b);
    layer1_outputs(5130) <= 1'b0;
    layer1_outputs(5131) <= not (a and b);
    layer1_outputs(5132) <= not (a and b);
    layer1_outputs(5133) <= 1'b1;
    layer1_outputs(5134) <= not a;
    layer1_outputs(5135) <= 1'b1;
    layer1_outputs(5136) <= 1'b1;
    layer1_outputs(5137) <= a and b;
    layer1_outputs(5138) <= not b or a;
    layer1_outputs(5139) <= not a or b;
    layer1_outputs(5140) <= not a or b;
    layer1_outputs(5141) <= b and not a;
    layer1_outputs(5142) <= not a;
    layer1_outputs(5143) <= a and not b;
    layer1_outputs(5144) <= a and b;
    layer1_outputs(5145) <= not b;
    layer1_outputs(5146) <= not a or b;
    layer1_outputs(5147) <= 1'b0;
    layer1_outputs(5148) <= not (a xor b);
    layer1_outputs(5149) <= a and not b;
    layer1_outputs(5150) <= 1'b1;
    layer1_outputs(5151) <= a and b;
    layer1_outputs(5152) <= not (a and b);
    layer1_outputs(5153) <= not a or b;
    layer1_outputs(5154) <= 1'b0;
    layer1_outputs(5155) <= not (a and b);
    layer1_outputs(5156) <= a or b;
    layer1_outputs(5157) <= not b or a;
    layer1_outputs(5158) <= not b;
    layer1_outputs(5159) <= a and b;
    layer1_outputs(5160) <= b and not a;
    layer1_outputs(5161) <= 1'b0;
    layer1_outputs(5162) <= 1'b0;
    layer1_outputs(5163) <= b and not a;
    layer1_outputs(5164) <= 1'b1;
    layer1_outputs(5165) <= 1'b0;
    layer1_outputs(5166) <= a;
    layer1_outputs(5167) <= not (a or b);
    layer1_outputs(5168) <= not a or b;
    layer1_outputs(5169) <= not (a or b);
    layer1_outputs(5170) <= 1'b1;
    layer1_outputs(5171) <= a;
    layer1_outputs(5172) <= 1'b0;
    layer1_outputs(5173) <= not a or b;
    layer1_outputs(5174) <= not a;
    layer1_outputs(5175) <= a and b;
    layer1_outputs(5176) <= 1'b0;
    layer1_outputs(5177) <= not b or a;
    layer1_outputs(5178) <= 1'b1;
    layer1_outputs(5179) <= not (a xor b);
    layer1_outputs(5180) <= not b;
    layer1_outputs(5181) <= not (a or b);
    layer1_outputs(5182) <= a or b;
    layer1_outputs(5183) <= 1'b0;
    layer1_outputs(5184) <= a xor b;
    layer1_outputs(5185) <= 1'b1;
    layer1_outputs(5186) <= not (a xor b);
    layer1_outputs(5187) <= not (a and b);
    layer1_outputs(5188) <= a;
    layer1_outputs(5189) <= b and not a;
    layer1_outputs(5190) <= not (a or b);
    layer1_outputs(5191) <= a or b;
    layer1_outputs(5192) <= a;
    layer1_outputs(5193) <= not (a and b);
    layer1_outputs(5194) <= not (a and b);
    layer1_outputs(5195) <= a xor b;
    layer1_outputs(5196) <= not (a and b);
    layer1_outputs(5197) <= not a or b;
    layer1_outputs(5198) <= not (a and b);
    layer1_outputs(5199) <= a xor b;
    layer1_outputs(5200) <= a;
    layer1_outputs(5201) <= not (a or b);
    layer1_outputs(5202) <= not (a xor b);
    layer1_outputs(5203) <= not (a xor b);
    layer1_outputs(5204) <= a or b;
    layer1_outputs(5205) <= not b;
    layer1_outputs(5206) <= not (a and b);
    layer1_outputs(5207) <= a;
    layer1_outputs(5208) <= not b;
    layer1_outputs(5209) <= not b or a;
    layer1_outputs(5210) <= a and b;
    layer1_outputs(5211) <= not a;
    layer1_outputs(5212) <= 1'b0;
    layer1_outputs(5213) <= not (a and b);
    layer1_outputs(5214) <= not (a and b);
    layer1_outputs(5215) <= not b or a;
    layer1_outputs(5216) <= 1'b0;
    layer1_outputs(5217) <= 1'b1;
    layer1_outputs(5218) <= 1'b1;
    layer1_outputs(5219) <= 1'b1;
    layer1_outputs(5220) <= not (a and b);
    layer1_outputs(5221) <= 1'b0;
    layer1_outputs(5222) <= not (a and b);
    layer1_outputs(5223) <= not b;
    layer1_outputs(5224) <= not (a xor b);
    layer1_outputs(5225) <= not (a xor b);
    layer1_outputs(5226) <= a and not b;
    layer1_outputs(5227) <= a and b;
    layer1_outputs(5228) <= a and not b;
    layer1_outputs(5229) <= 1'b1;
    layer1_outputs(5230) <= not (a and b);
    layer1_outputs(5231) <= a and b;
    layer1_outputs(5232) <= not a;
    layer1_outputs(5233) <= 1'b0;
    layer1_outputs(5234) <= a xor b;
    layer1_outputs(5235) <= a;
    layer1_outputs(5236) <= not a;
    layer1_outputs(5237) <= b and not a;
    layer1_outputs(5238) <= b;
    layer1_outputs(5239) <= b;
    layer1_outputs(5240) <= 1'b0;
    layer1_outputs(5241) <= b;
    layer1_outputs(5242) <= 1'b0;
    layer1_outputs(5243) <= not b;
    layer1_outputs(5244) <= a and not b;
    layer1_outputs(5245) <= b;
    layer1_outputs(5246) <= b;
    layer1_outputs(5247) <= a;
    layer1_outputs(5248) <= a;
    layer1_outputs(5249) <= not a or b;
    layer1_outputs(5250) <= a and not b;
    layer1_outputs(5251) <= not (a or b);
    layer1_outputs(5252) <= a;
    layer1_outputs(5253) <= not b;
    layer1_outputs(5254) <= 1'b0;
    layer1_outputs(5255) <= not b or a;
    layer1_outputs(5256) <= not a or b;
    layer1_outputs(5257) <= a and b;
    layer1_outputs(5258) <= a and b;
    layer1_outputs(5259) <= not (a or b);
    layer1_outputs(5260) <= 1'b0;
    layer1_outputs(5261) <= b and not a;
    layer1_outputs(5262) <= a or b;
    layer1_outputs(5263) <= a or b;
    layer1_outputs(5264) <= a and b;
    layer1_outputs(5265) <= b;
    layer1_outputs(5266) <= not a or b;
    layer1_outputs(5267) <= 1'b1;
    layer1_outputs(5268) <= a and not b;
    layer1_outputs(5269) <= a and b;
    layer1_outputs(5270) <= 1'b0;
    layer1_outputs(5271) <= a xor b;
    layer1_outputs(5272) <= a;
    layer1_outputs(5273) <= b;
    layer1_outputs(5274) <= 1'b1;
    layer1_outputs(5275) <= 1'b0;
    layer1_outputs(5276) <= a and not b;
    layer1_outputs(5277) <= not (a or b);
    layer1_outputs(5278) <= 1'b0;
    layer1_outputs(5279) <= a and b;
    layer1_outputs(5280) <= a xor b;
    layer1_outputs(5281) <= a;
    layer1_outputs(5282) <= b;
    layer1_outputs(5283) <= not a or b;
    layer1_outputs(5284) <= 1'b0;
    layer1_outputs(5285) <= not (a and b);
    layer1_outputs(5286) <= not b or a;
    layer1_outputs(5287) <= not (a and b);
    layer1_outputs(5288) <= a or b;
    layer1_outputs(5289) <= b;
    layer1_outputs(5290) <= not (a and b);
    layer1_outputs(5291) <= not b or a;
    layer1_outputs(5292) <= not b;
    layer1_outputs(5293) <= a;
    layer1_outputs(5294) <= not a or b;
    layer1_outputs(5295) <= 1'b0;
    layer1_outputs(5296) <= a and b;
    layer1_outputs(5297) <= not b or a;
    layer1_outputs(5298) <= not a;
    layer1_outputs(5299) <= not (a or b);
    layer1_outputs(5300) <= not (a or b);
    layer1_outputs(5301) <= a xor b;
    layer1_outputs(5302) <= a and b;
    layer1_outputs(5303) <= not b or a;
    layer1_outputs(5304) <= not b or a;
    layer1_outputs(5305) <= a or b;
    layer1_outputs(5306) <= b;
    layer1_outputs(5307) <= not a;
    layer1_outputs(5308) <= not a;
    layer1_outputs(5309) <= not (a and b);
    layer1_outputs(5310) <= not b or a;
    layer1_outputs(5311) <= not b or a;
    layer1_outputs(5312) <= not b;
    layer1_outputs(5313) <= not a;
    layer1_outputs(5314) <= a xor b;
    layer1_outputs(5315) <= 1'b1;
    layer1_outputs(5316) <= a and b;
    layer1_outputs(5317) <= 1'b0;
    layer1_outputs(5318) <= not b or a;
    layer1_outputs(5319) <= a or b;
    layer1_outputs(5320) <= 1'b1;
    layer1_outputs(5321) <= a or b;
    layer1_outputs(5322) <= not a or b;
    layer1_outputs(5323) <= not (a and b);
    layer1_outputs(5324) <= not b or a;
    layer1_outputs(5325) <= a or b;
    layer1_outputs(5326) <= a xor b;
    layer1_outputs(5327) <= b;
    layer1_outputs(5328) <= a xor b;
    layer1_outputs(5329) <= 1'b1;
    layer1_outputs(5330) <= a or b;
    layer1_outputs(5331) <= a and b;
    layer1_outputs(5332) <= not b;
    layer1_outputs(5333) <= not (a or b);
    layer1_outputs(5334) <= 1'b1;
    layer1_outputs(5335) <= b;
    layer1_outputs(5336) <= not b or a;
    layer1_outputs(5337) <= 1'b1;
    layer1_outputs(5338) <= not a or b;
    layer1_outputs(5339) <= 1'b0;
    layer1_outputs(5340) <= not (a and b);
    layer1_outputs(5341) <= not (a or b);
    layer1_outputs(5342) <= 1'b0;
    layer1_outputs(5343) <= a and not b;
    layer1_outputs(5344) <= not (a xor b);
    layer1_outputs(5345) <= a or b;
    layer1_outputs(5346) <= not b;
    layer1_outputs(5347) <= 1'b0;
    layer1_outputs(5348) <= not a or b;
    layer1_outputs(5349) <= a;
    layer1_outputs(5350) <= b;
    layer1_outputs(5351) <= a and not b;
    layer1_outputs(5352) <= 1'b0;
    layer1_outputs(5353) <= 1'b0;
    layer1_outputs(5354) <= not (a and b);
    layer1_outputs(5355) <= not a;
    layer1_outputs(5356) <= a;
    layer1_outputs(5357) <= b and not a;
    layer1_outputs(5358) <= not (a or b);
    layer1_outputs(5359) <= 1'b0;
    layer1_outputs(5360) <= b and not a;
    layer1_outputs(5361) <= 1'b1;
    layer1_outputs(5362) <= not (a and b);
    layer1_outputs(5363) <= not (a or b);
    layer1_outputs(5364) <= not (a and b);
    layer1_outputs(5365) <= not a or b;
    layer1_outputs(5366) <= b and not a;
    layer1_outputs(5367) <= not (a and b);
    layer1_outputs(5368) <= a and b;
    layer1_outputs(5369) <= a and b;
    layer1_outputs(5370) <= 1'b0;
    layer1_outputs(5371) <= not (a and b);
    layer1_outputs(5372) <= 1'b0;
    layer1_outputs(5373) <= not a;
    layer1_outputs(5374) <= a and not b;
    layer1_outputs(5375) <= a;
    layer1_outputs(5376) <= a or b;
    layer1_outputs(5377) <= a xor b;
    layer1_outputs(5378) <= not a;
    layer1_outputs(5379) <= 1'b0;
    layer1_outputs(5380) <= not (a or b);
    layer1_outputs(5381) <= 1'b0;
    layer1_outputs(5382) <= 1'b0;
    layer1_outputs(5383) <= not (a xor b);
    layer1_outputs(5384) <= b and not a;
    layer1_outputs(5385) <= 1'b0;
    layer1_outputs(5386) <= not a or b;
    layer1_outputs(5387) <= a;
    layer1_outputs(5388) <= not a;
    layer1_outputs(5389) <= not (a or b);
    layer1_outputs(5390) <= not b or a;
    layer1_outputs(5391) <= not b;
    layer1_outputs(5392) <= 1'b0;
    layer1_outputs(5393) <= b and not a;
    layer1_outputs(5394) <= 1'b1;
    layer1_outputs(5395) <= not (a or b);
    layer1_outputs(5396) <= 1'b1;
    layer1_outputs(5397) <= not (a or b);
    layer1_outputs(5398) <= a and not b;
    layer1_outputs(5399) <= b and not a;
    layer1_outputs(5400) <= 1'b1;
    layer1_outputs(5401) <= not (a or b);
    layer1_outputs(5402) <= 1'b1;
    layer1_outputs(5403) <= 1'b1;
    layer1_outputs(5404) <= not a or b;
    layer1_outputs(5405) <= b;
    layer1_outputs(5406) <= a and not b;
    layer1_outputs(5407) <= not a;
    layer1_outputs(5408) <= b and not a;
    layer1_outputs(5409) <= a and not b;
    layer1_outputs(5410) <= not a or b;
    layer1_outputs(5411) <= b and not a;
    layer1_outputs(5412) <= a xor b;
    layer1_outputs(5413) <= not (a and b);
    layer1_outputs(5414) <= not a or b;
    layer1_outputs(5415) <= not a;
    layer1_outputs(5416) <= not b;
    layer1_outputs(5417) <= b;
    layer1_outputs(5418) <= not b or a;
    layer1_outputs(5419) <= a;
    layer1_outputs(5420) <= not (a and b);
    layer1_outputs(5421) <= not a;
    layer1_outputs(5422) <= a and b;
    layer1_outputs(5423) <= a;
    layer1_outputs(5424) <= not (a xor b);
    layer1_outputs(5425) <= b;
    layer1_outputs(5426) <= not a;
    layer1_outputs(5427) <= not (a or b);
    layer1_outputs(5428) <= not a or b;
    layer1_outputs(5429) <= b and not a;
    layer1_outputs(5430) <= not (a or b);
    layer1_outputs(5431) <= b and not a;
    layer1_outputs(5432) <= a and not b;
    layer1_outputs(5433) <= b and not a;
    layer1_outputs(5434) <= not (a or b);
    layer1_outputs(5435) <= 1'b0;
    layer1_outputs(5436) <= a and b;
    layer1_outputs(5437) <= 1'b0;
    layer1_outputs(5438) <= 1'b0;
    layer1_outputs(5439) <= 1'b0;
    layer1_outputs(5440) <= 1'b0;
    layer1_outputs(5441) <= not b;
    layer1_outputs(5442) <= not (a or b);
    layer1_outputs(5443) <= not (a and b);
    layer1_outputs(5444) <= not a;
    layer1_outputs(5445) <= a;
    layer1_outputs(5446) <= b and not a;
    layer1_outputs(5447) <= not b or a;
    layer1_outputs(5448) <= not a;
    layer1_outputs(5449) <= a xor b;
    layer1_outputs(5450) <= 1'b1;
    layer1_outputs(5451) <= b;
    layer1_outputs(5452) <= 1'b1;
    layer1_outputs(5453) <= not (a and b);
    layer1_outputs(5454) <= a or b;
    layer1_outputs(5455) <= a;
    layer1_outputs(5456) <= not a;
    layer1_outputs(5457) <= 1'b0;
    layer1_outputs(5458) <= not (a xor b);
    layer1_outputs(5459) <= a or b;
    layer1_outputs(5460) <= not b;
    layer1_outputs(5461) <= not (a or b);
    layer1_outputs(5462) <= not (a and b);
    layer1_outputs(5463) <= not a;
    layer1_outputs(5464) <= not a or b;
    layer1_outputs(5465) <= a xor b;
    layer1_outputs(5466) <= not a;
    layer1_outputs(5467) <= not a or b;
    layer1_outputs(5468) <= not b;
    layer1_outputs(5469) <= not b;
    layer1_outputs(5470) <= not (a and b);
    layer1_outputs(5471) <= not a or b;
    layer1_outputs(5472) <= a or b;
    layer1_outputs(5473) <= not b or a;
    layer1_outputs(5474) <= not (a and b);
    layer1_outputs(5475) <= not (a and b);
    layer1_outputs(5476) <= not a;
    layer1_outputs(5477) <= a and b;
    layer1_outputs(5478) <= not (a or b);
    layer1_outputs(5479) <= 1'b1;
    layer1_outputs(5480) <= 1'b1;
    layer1_outputs(5481) <= a or b;
    layer1_outputs(5482) <= a xor b;
    layer1_outputs(5483) <= a;
    layer1_outputs(5484) <= 1'b1;
    layer1_outputs(5485) <= not b;
    layer1_outputs(5486) <= b;
    layer1_outputs(5487) <= a;
    layer1_outputs(5488) <= not (a or b);
    layer1_outputs(5489) <= 1'b1;
    layer1_outputs(5490) <= not a;
    layer1_outputs(5491) <= a;
    layer1_outputs(5492) <= 1'b0;
    layer1_outputs(5493) <= a and b;
    layer1_outputs(5494) <= b and not a;
    layer1_outputs(5495) <= 1'b0;
    layer1_outputs(5496) <= not (a and b);
    layer1_outputs(5497) <= 1'b0;
    layer1_outputs(5498) <= 1'b0;
    layer1_outputs(5499) <= 1'b0;
    layer1_outputs(5500) <= not a;
    layer1_outputs(5501) <= b and not a;
    layer1_outputs(5502) <= not a or b;
    layer1_outputs(5503) <= not (a or b);
    layer1_outputs(5504) <= not b or a;
    layer1_outputs(5505) <= a and not b;
    layer1_outputs(5506) <= 1'b0;
    layer1_outputs(5507) <= 1'b0;
    layer1_outputs(5508) <= a or b;
    layer1_outputs(5509) <= not a or b;
    layer1_outputs(5510) <= 1'b0;
    layer1_outputs(5511) <= not b or a;
    layer1_outputs(5512) <= not (a and b);
    layer1_outputs(5513) <= not (a or b);
    layer1_outputs(5514) <= not a;
    layer1_outputs(5515) <= a;
    layer1_outputs(5516) <= not (a and b);
    layer1_outputs(5517) <= not a or b;
    layer1_outputs(5518) <= a;
    layer1_outputs(5519) <= a;
    layer1_outputs(5520) <= a and not b;
    layer1_outputs(5521) <= not b or a;
    layer1_outputs(5522) <= 1'b1;
    layer1_outputs(5523) <= a;
    layer1_outputs(5524) <= a and b;
    layer1_outputs(5525) <= 1'b1;
    layer1_outputs(5526) <= 1'b1;
    layer1_outputs(5527) <= 1'b0;
    layer1_outputs(5528) <= a or b;
    layer1_outputs(5529) <= a and not b;
    layer1_outputs(5530) <= a or b;
    layer1_outputs(5531) <= 1'b1;
    layer1_outputs(5532) <= not a or b;
    layer1_outputs(5533) <= not b;
    layer1_outputs(5534) <= a and b;
    layer1_outputs(5535) <= a or b;
    layer1_outputs(5536) <= a;
    layer1_outputs(5537) <= a or b;
    layer1_outputs(5538) <= not (a or b);
    layer1_outputs(5539) <= not (a or b);
    layer1_outputs(5540) <= not a or b;
    layer1_outputs(5541) <= 1'b0;
    layer1_outputs(5542) <= 1'b0;
    layer1_outputs(5543) <= not b;
    layer1_outputs(5544) <= not b or a;
    layer1_outputs(5545) <= not a or b;
    layer1_outputs(5546) <= 1'b0;
    layer1_outputs(5547) <= a;
    layer1_outputs(5548) <= 1'b0;
    layer1_outputs(5549) <= not b or a;
    layer1_outputs(5550) <= a or b;
    layer1_outputs(5551) <= 1'b1;
    layer1_outputs(5552) <= a and b;
    layer1_outputs(5553) <= not a;
    layer1_outputs(5554) <= not (a or b);
    layer1_outputs(5555) <= not (a or b);
    layer1_outputs(5556) <= b and not a;
    layer1_outputs(5557) <= b;
    layer1_outputs(5558) <= a and b;
    layer1_outputs(5559) <= not b or a;
    layer1_outputs(5560) <= not b;
    layer1_outputs(5561) <= not a or b;
    layer1_outputs(5562) <= 1'b0;
    layer1_outputs(5563) <= not (a and b);
    layer1_outputs(5564) <= a and b;
    layer1_outputs(5565) <= b and not a;
    layer1_outputs(5566) <= a xor b;
    layer1_outputs(5567) <= a or b;
    layer1_outputs(5568) <= not b or a;
    layer1_outputs(5569) <= 1'b0;
    layer1_outputs(5570) <= not (a and b);
    layer1_outputs(5571) <= not a;
    layer1_outputs(5572) <= 1'b1;
    layer1_outputs(5573) <= not b;
    layer1_outputs(5574) <= not (a or b);
    layer1_outputs(5575) <= a or b;
    layer1_outputs(5576) <= a;
    layer1_outputs(5577) <= not a or b;
    layer1_outputs(5578) <= not (a and b);
    layer1_outputs(5579) <= a and not b;
    layer1_outputs(5580) <= not (a or b);
    layer1_outputs(5581) <= a or b;
    layer1_outputs(5582) <= a and b;
    layer1_outputs(5583) <= not (a and b);
    layer1_outputs(5584) <= not b;
    layer1_outputs(5585) <= not (a or b);
    layer1_outputs(5586) <= a xor b;
    layer1_outputs(5587) <= b;
    layer1_outputs(5588) <= 1'b0;
    layer1_outputs(5589) <= not b;
    layer1_outputs(5590) <= 1'b0;
    layer1_outputs(5591) <= 1'b0;
    layer1_outputs(5592) <= not a or b;
    layer1_outputs(5593) <= not a;
    layer1_outputs(5594) <= a or b;
    layer1_outputs(5595) <= 1'b1;
    layer1_outputs(5596) <= 1'b1;
    layer1_outputs(5597) <= not a or b;
    layer1_outputs(5598) <= a and b;
    layer1_outputs(5599) <= a and not b;
    layer1_outputs(5600) <= not b or a;
    layer1_outputs(5601) <= a and b;
    layer1_outputs(5602) <= 1'b0;
    layer1_outputs(5603) <= a xor b;
    layer1_outputs(5604) <= not (a and b);
    layer1_outputs(5605) <= not a or b;
    layer1_outputs(5606) <= a and b;
    layer1_outputs(5607) <= 1'b0;
    layer1_outputs(5608) <= a or b;
    layer1_outputs(5609) <= not b;
    layer1_outputs(5610) <= 1'b1;
    layer1_outputs(5611) <= 1'b0;
    layer1_outputs(5612) <= not (a and b);
    layer1_outputs(5613) <= a and b;
    layer1_outputs(5614) <= not (a or b);
    layer1_outputs(5615) <= b;
    layer1_outputs(5616) <= b and not a;
    layer1_outputs(5617) <= 1'b0;
    layer1_outputs(5618) <= 1'b0;
    layer1_outputs(5619) <= a and b;
    layer1_outputs(5620) <= not b;
    layer1_outputs(5621) <= a xor b;
    layer1_outputs(5622) <= not b or a;
    layer1_outputs(5623) <= a;
    layer1_outputs(5624) <= a or b;
    layer1_outputs(5625) <= a xor b;
    layer1_outputs(5626) <= b;
    layer1_outputs(5627) <= 1'b1;
    layer1_outputs(5628) <= not (a and b);
    layer1_outputs(5629) <= not (a and b);
    layer1_outputs(5630) <= not (a and b);
    layer1_outputs(5631) <= not b or a;
    layer1_outputs(5632) <= not (a and b);
    layer1_outputs(5633) <= a xor b;
    layer1_outputs(5634) <= a or b;
    layer1_outputs(5635) <= not a or b;
    layer1_outputs(5636) <= a and not b;
    layer1_outputs(5637) <= not (a and b);
    layer1_outputs(5638) <= 1'b1;
    layer1_outputs(5639) <= a and not b;
    layer1_outputs(5640) <= 1'b0;
    layer1_outputs(5641) <= a or b;
    layer1_outputs(5642) <= not (a or b);
    layer1_outputs(5643) <= a or b;
    layer1_outputs(5644) <= not (a xor b);
    layer1_outputs(5645) <= b and not a;
    layer1_outputs(5646) <= not a;
    layer1_outputs(5647) <= 1'b1;
    layer1_outputs(5648) <= 1'b1;
    layer1_outputs(5649) <= not (a xor b);
    layer1_outputs(5650) <= b and not a;
    layer1_outputs(5651) <= a and b;
    layer1_outputs(5652) <= a or b;
    layer1_outputs(5653) <= a and not b;
    layer1_outputs(5654) <= 1'b0;
    layer1_outputs(5655) <= b;
    layer1_outputs(5656) <= a and b;
    layer1_outputs(5657) <= b;
    layer1_outputs(5658) <= 1'b1;
    layer1_outputs(5659) <= not b;
    layer1_outputs(5660) <= not a;
    layer1_outputs(5661) <= not a or b;
    layer1_outputs(5662) <= not b;
    layer1_outputs(5663) <= not a or b;
    layer1_outputs(5664) <= not b or a;
    layer1_outputs(5665) <= a;
    layer1_outputs(5666) <= not a or b;
    layer1_outputs(5667) <= not a;
    layer1_outputs(5668) <= b;
    layer1_outputs(5669) <= a and b;
    layer1_outputs(5670) <= a or b;
    layer1_outputs(5671) <= 1'b1;
    layer1_outputs(5672) <= b;
    layer1_outputs(5673) <= 1'b0;
    layer1_outputs(5674) <= a;
    layer1_outputs(5675) <= a and b;
    layer1_outputs(5676) <= a and b;
    layer1_outputs(5677) <= not a;
    layer1_outputs(5678) <= a xor b;
    layer1_outputs(5679) <= not a;
    layer1_outputs(5680) <= a;
    layer1_outputs(5681) <= 1'b0;
    layer1_outputs(5682) <= b and not a;
    layer1_outputs(5683) <= 1'b1;
    layer1_outputs(5684) <= not b;
    layer1_outputs(5685) <= not b or a;
    layer1_outputs(5686) <= not a or b;
    layer1_outputs(5687) <= not a or b;
    layer1_outputs(5688) <= b and not a;
    layer1_outputs(5689) <= a and not b;
    layer1_outputs(5690) <= 1'b1;
    layer1_outputs(5691) <= not a or b;
    layer1_outputs(5692) <= not (a or b);
    layer1_outputs(5693) <= not b;
    layer1_outputs(5694) <= not (a or b);
    layer1_outputs(5695) <= b;
    layer1_outputs(5696) <= not a or b;
    layer1_outputs(5697) <= a and b;
    layer1_outputs(5698) <= a or b;
    layer1_outputs(5699) <= 1'b0;
    layer1_outputs(5700) <= 1'b1;
    layer1_outputs(5701) <= 1'b0;
    layer1_outputs(5702) <= not b or a;
    layer1_outputs(5703) <= b;
    layer1_outputs(5704) <= a and b;
    layer1_outputs(5705) <= not a or b;
    layer1_outputs(5706) <= b and not a;
    layer1_outputs(5707) <= not b or a;
    layer1_outputs(5708) <= not (a and b);
    layer1_outputs(5709) <= not b;
    layer1_outputs(5710) <= a and not b;
    layer1_outputs(5711) <= a and b;
    layer1_outputs(5712) <= a;
    layer1_outputs(5713) <= a or b;
    layer1_outputs(5714) <= b;
    layer1_outputs(5715) <= not b;
    layer1_outputs(5716) <= not (a or b);
    layer1_outputs(5717) <= 1'b0;
    layer1_outputs(5718) <= a and not b;
    layer1_outputs(5719) <= not a;
    layer1_outputs(5720) <= a and not b;
    layer1_outputs(5721) <= 1'b0;
    layer1_outputs(5722) <= a and not b;
    layer1_outputs(5723) <= not (a or b);
    layer1_outputs(5724) <= a and not b;
    layer1_outputs(5725) <= not a;
    layer1_outputs(5726) <= a;
    layer1_outputs(5727) <= 1'b0;
    layer1_outputs(5728) <= not b;
    layer1_outputs(5729) <= not b;
    layer1_outputs(5730) <= not (a xor b);
    layer1_outputs(5731) <= not (a or b);
    layer1_outputs(5732) <= a and not b;
    layer1_outputs(5733) <= b;
    layer1_outputs(5734) <= b;
    layer1_outputs(5735) <= not a or b;
    layer1_outputs(5736) <= 1'b1;
    layer1_outputs(5737) <= a;
    layer1_outputs(5738) <= a and not b;
    layer1_outputs(5739) <= a and b;
    layer1_outputs(5740) <= not (a and b);
    layer1_outputs(5741) <= 1'b1;
    layer1_outputs(5742) <= a and not b;
    layer1_outputs(5743) <= a or b;
    layer1_outputs(5744) <= not b;
    layer1_outputs(5745) <= not (a and b);
    layer1_outputs(5746) <= a;
    layer1_outputs(5747) <= b;
    layer1_outputs(5748) <= not (a or b);
    layer1_outputs(5749) <= not (a or b);
    layer1_outputs(5750) <= 1'b1;
    layer1_outputs(5751) <= b and not a;
    layer1_outputs(5752) <= a xor b;
    layer1_outputs(5753) <= a or b;
    layer1_outputs(5754) <= a and not b;
    layer1_outputs(5755) <= 1'b1;
    layer1_outputs(5756) <= not (a and b);
    layer1_outputs(5757) <= not a;
    layer1_outputs(5758) <= not a;
    layer1_outputs(5759) <= a;
    layer1_outputs(5760) <= not a;
    layer1_outputs(5761) <= not (a or b);
    layer1_outputs(5762) <= a;
    layer1_outputs(5763) <= not b or a;
    layer1_outputs(5764) <= a and b;
    layer1_outputs(5765) <= a;
    layer1_outputs(5766) <= a;
    layer1_outputs(5767) <= not (a or b);
    layer1_outputs(5768) <= 1'b0;
    layer1_outputs(5769) <= 1'b0;
    layer1_outputs(5770) <= not (a or b);
    layer1_outputs(5771) <= 1'b1;
    layer1_outputs(5772) <= a or b;
    layer1_outputs(5773) <= not (a or b);
    layer1_outputs(5774) <= b;
    layer1_outputs(5775) <= not a or b;
    layer1_outputs(5776) <= not (a or b);
    layer1_outputs(5777) <= b and not a;
    layer1_outputs(5778) <= a and not b;
    layer1_outputs(5779) <= a and b;
    layer1_outputs(5780) <= a and b;
    layer1_outputs(5781) <= a;
    layer1_outputs(5782) <= not (a or b);
    layer1_outputs(5783) <= b and not a;
    layer1_outputs(5784) <= not (a and b);
    layer1_outputs(5785) <= a;
    layer1_outputs(5786) <= 1'b1;
    layer1_outputs(5787) <= 1'b1;
    layer1_outputs(5788) <= 1'b0;
    layer1_outputs(5789) <= not a;
    layer1_outputs(5790) <= not a or b;
    layer1_outputs(5791) <= b;
    layer1_outputs(5792) <= not b or a;
    layer1_outputs(5793) <= not (a and b);
    layer1_outputs(5794) <= a or b;
    layer1_outputs(5795) <= 1'b1;
    layer1_outputs(5796) <= not b;
    layer1_outputs(5797) <= a;
    layer1_outputs(5798) <= not (a and b);
    layer1_outputs(5799) <= a and b;
    layer1_outputs(5800) <= a or b;
    layer1_outputs(5801) <= 1'b0;
    layer1_outputs(5802) <= a and not b;
    layer1_outputs(5803) <= b and not a;
    layer1_outputs(5804) <= b;
    layer1_outputs(5805) <= b and not a;
    layer1_outputs(5806) <= 1'b0;
    layer1_outputs(5807) <= not (a or b);
    layer1_outputs(5808) <= a or b;
    layer1_outputs(5809) <= not b;
    layer1_outputs(5810) <= 1'b1;
    layer1_outputs(5811) <= not b or a;
    layer1_outputs(5812) <= not a;
    layer1_outputs(5813) <= b and not a;
    layer1_outputs(5814) <= not (a or b);
    layer1_outputs(5815) <= 1'b0;
    layer1_outputs(5816) <= not b or a;
    layer1_outputs(5817) <= not (a and b);
    layer1_outputs(5818) <= a;
    layer1_outputs(5819) <= not b or a;
    layer1_outputs(5820) <= a or b;
    layer1_outputs(5821) <= not a or b;
    layer1_outputs(5822) <= a and b;
    layer1_outputs(5823) <= not a;
    layer1_outputs(5824) <= 1'b0;
    layer1_outputs(5825) <= not a;
    layer1_outputs(5826) <= b;
    layer1_outputs(5827) <= not a or b;
    layer1_outputs(5828) <= not b or a;
    layer1_outputs(5829) <= b;
    layer1_outputs(5830) <= not b or a;
    layer1_outputs(5831) <= not b or a;
    layer1_outputs(5832) <= a or b;
    layer1_outputs(5833) <= b;
    layer1_outputs(5834) <= b and not a;
    layer1_outputs(5835) <= not (a and b);
    layer1_outputs(5836) <= a;
    layer1_outputs(5837) <= a and not b;
    layer1_outputs(5838) <= a;
    layer1_outputs(5839) <= 1'b0;
    layer1_outputs(5840) <= 1'b1;
    layer1_outputs(5841) <= not a;
    layer1_outputs(5842) <= a;
    layer1_outputs(5843) <= 1'b1;
    layer1_outputs(5844) <= 1'b0;
    layer1_outputs(5845) <= 1'b1;
    layer1_outputs(5846) <= a xor b;
    layer1_outputs(5847) <= a or b;
    layer1_outputs(5848) <= b and not a;
    layer1_outputs(5849) <= 1'b1;
    layer1_outputs(5850) <= a xor b;
    layer1_outputs(5851) <= a or b;
    layer1_outputs(5852) <= 1'b0;
    layer1_outputs(5853) <= not a;
    layer1_outputs(5854) <= 1'b0;
    layer1_outputs(5855) <= 1'b1;
    layer1_outputs(5856) <= not a or b;
    layer1_outputs(5857) <= 1'b1;
    layer1_outputs(5858) <= a and b;
    layer1_outputs(5859) <= b and not a;
    layer1_outputs(5860) <= not a;
    layer1_outputs(5861) <= not a;
    layer1_outputs(5862) <= a and not b;
    layer1_outputs(5863) <= a and not b;
    layer1_outputs(5864) <= a or b;
    layer1_outputs(5865) <= b and not a;
    layer1_outputs(5866) <= a or b;
    layer1_outputs(5867) <= a or b;
    layer1_outputs(5868) <= not a;
    layer1_outputs(5869) <= 1'b1;
    layer1_outputs(5870) <= b and not a;
    layer1_outputs(5871) <= b and not a;
    layer1_outputs(5872) <= not (a or b);
    layer1_outputs(5873) <= 1'b0;
    layer1_outputs(5874) <= b;
    layer1_outputs(5875) <= not (a and b);
    layer1_outputs(5876) <= a or b;
    layer1_outputs(5877) <= a;
    layer1_outputs(5878) <= not a;
    layer1_outputs(5879) <= 1'b0;
    layer1_outputs(5880) <= not a;
    layer1_outputs(5881) <= a or b;
    layer1_outputs(5882) <= 1'b0;
    layer1_outputs(5883) <= not (a or b);
    layer1_outputs(5884) <= not (a and b);
    layer1_outputs(5885) <= not b;
    layer1_outputs(5886) <= 1'b1;
    layer1_outputs(5887) <= a or b;
    layer1_outputs(5888) <= a and not b;
    layer1_outputs(5889) <= a xor b;
    layer1_outputs(5890) <= not a or b;
    layer1_outputs(5891) <= not (a and b);
    layer1_outputs(5892) <= 1'b1;
    layer1_outputs(5893) <= not (a or b);
    layer1_outputs(5894) <= not (a or b);
    layer1_outputs(5895) <= b and not a;
    layer1_outputs(5896) <= not a;
    layer1_outputs(5897) <= not (a or b);
    layer1_outputs(5898) <= a;
    layer1_outputs(5899) <= not b;
    layer1_outputs(5900) <= a or b;
    layer1_outputs(5901) <= not b;
    layer1_outputs(5902) <= not a;
    layer1_outputs(5903) <= b;
    layer1_outputs(5904) <= a;
    layer1_outputs(5905) <= not b or a;
    layer1_outputs(5906) <= a and b;
    layer1_outputs(5907) <= not (a or b);
    layer1_outputs(5908) <= a and not b;
    layer1_outputs(5909) <= a and b;
    layer1_outputs(5910) <= not (a or b);
    layer1_outputs(5911) <= 1'b1;
    layer1_outputs(5912) <= b;
    layer1_outputs(5913) <= not (a or b);
    layer1_outputs(5914) <= a and b;
    layer1_outputs(5915) <= 1'b0;
    layer1_outputs(5916) <= not (a xor b);
    layer1_outputs(5917) <= a and b;
    layer1_outputs(5918) <= a or b;
    layer1_outputs(5919) <= not (a and b);
    layer1_outputs(5920) <= a or b;
    layer1_outputs(5921) <= a and not b;
    layer1_outputs(5922) <= not b;
    layer1_outputs(5923) <= not (a or b);
    layer1_outputs(5924) <= not (a and b);
    layer1_outputs(5925) <= not b or a;
    layer1_outputs(5926) <= b;
    layer1_outputs(5927) <= a and not b;
    layer1_outputs(5928) <= not (a or b);
    layer1_outputs(5929) <= not (a and b);
    layer1_outputs(5930) <= a and b;
    layer1_outputs(5931) <= not b;
    layer1_outputs(5932) <= a;
    layer1_outputs(5933) <= not (a or b);
    layer1_outputs(5934) <= a and b;
    layer1_outputs(5935) <= 1'b1;
    layer1_outputs(5936) <= a and b;
    layer1_outputs(5937) <= 1'b1;
    layer1_outputs(5938) <= a or b;
    layer1_outputs(5939) <= not b;
    layer1_outputs(5940) <= not (a or b);
    layer1_outputs(5941) <= 1'b0;
    layer1_outputs(5942) <= not b;
    layer1_outputs(5943) <= not a or b;
    layer1_outputs(5944) <= not b;
    layer1_outputs(5945) <= 1'b1;
    layer1_outputs(5946) <= a or b;
    layer1_outputs(5947) <= not (a or b);
    layer1_outputs(5948) <= a or b;
    layer1_outputs(5949) <= b and not a;
    layer1_outputs(5950) <= 1'b1;
    layer1_outputs(5951) <= not a or b;
    layer1_outputs(5952) <= a;
    layer1_outputs(5953) <= 1'b0;
    layer1_outputs(5954) <= 1'b0;
    layer1_outputs(5955) <= not (a or b);
    layer1_outputs(5956) <= b and not a;
    layer1_outputs(5957) <= 1'b1;
    layer1_outputs(5958) <= a and not b;
    layer1_outputs(5959) <= not a;
    layer1_outputs(5960) <= a or b;
    layer1_outputs(5961) <= a and not b;
    layer1_outputs(5962) <= not (a or b);
    layer1_outputs(5963) <= not b;
    layer1_outputs(5964) <= a;
    layer1_outputs(5965) <= a and b;
    layer1_outputs(5966) <= not (a or b);
    layer1_outputs(5967) <= 1'b0;
    layer1_outputs(5968) <= not (a or b);
    layer1_outputs(5969) <= a and b;
    layer1_outputs(5970) <= 1'b1;
    layer1_outputs(5971) <= not a or b;
    layer1_outputs(5972) <= not (a and b);
    layer1_outputs(5973) <= not (a or b);
    layer1_outputs(5974) <= not a;
    layer1_outputs(5975) <= not b;
    layer1_outputs(5976) <= not (a xor b);
    layer1_outputs(5977) <= not a or b;
    layer1_outputs(5978) <= not (a and b);
    layer1_outputs(5979) <= b;
    layer1_outputs(5980) <= a xor b;
    layer1_outputs(5981) <= not (a xor b);
    layer1_outputs(5982) <= not a or b;
    layer1_outputs(5983) <= not b or a;
    layer1_outputs(5984) <= a xor b;
    layer1_outputs(5985) <= not a or b;
    layer1_outputs(5986) <= a and b;
    layer1_outputs(5987) <= not (a xor b);
    layer1_outputs(5988) <= a xor b;
    layer1_outputs(5989) <= a and not b;
    layer1_outputs(5990) <= a and not b;
    layer1_outputs(5991) <= a and not b;
    layer1_outputs(5992) <= not (a or b);
    layer1_outputs(5993) <= a xor b;
    layer1_outputs(5994) <= a and b;
    layer1_outputs(5995) <= b and not a;
    layer1_outputs(5996) <= b and not a;
    layer1_outputs(5997) <= not (a and b);
    layer1_outputs(5998) <= 1'b0;
    layer1_outputs(5999) <= a or b;
    layer1_outputs(6000) <= not b or a;
    layer1_outputs(6001) <= not (a or b);
    layer1_outputs(6002) <= not (a and b);
    layer1_outputs(6003) <= 1'b0;
    layer1_outputs(6004) <= b;
    layer1_outputs(6005) <= not b or a;
    layer1_outputs(6006) <= not b or a;
    layer1_outputs(6007) <= a and not b;
    layer1_outputs(6008) <= 1'b1;
    layer1_outputs(6009) <= a or b;
    layer1_outputs(6010) <= not b;
    layer1_outputs(6011) <= a and not b;
    layer1_outputs(6012) <= not (a and b);
    layer1_outputs(6013) <= not a or b;
    layer1_outputs(6014) <= a and b;
    layer1_outputs(6015) <= a and b;
    layer1_outputs(6016) <= a and b;
    layer1_outputs(6017) <= not b;
    layer1_outputs(6018) <= not (a or b);
    layer1_outputs(6019) <= a or b;
    layer1_outputs(6020) <= a and not b;
    layer1_outputs(6021) <= b and not a;
    layer1_outputs(6022) <= a and not b;
    layer1_outputs(6023) <= 1'b0;
    layer1_outputs(6024) <= 1'b0;
    layer1_outputs(6025) <= not a;
    layer1_outputs(6026) <= 1'b1;
    layer1_outputs(6027) <= not (a or b);
    layer1_outputs(6028) <= 1'b1;
    layer1_outputs(6029) <= 1'b0;
    layer1_outputs(6030) <= a or b;
    layer1_outputs(6031) <= a;
    layer1_outputs(6032) <= a;
    layer1_outputs(6033) <= b and not a;
    layer1_outputs(6034) <= b;
    layer1_outputs(6035) <= a;
    layer1_outputs(6036) <= b;
    layer1_outputs(6037) <= not a;
    layer1_outputs(6038) <= not b;
    layer1_outputs(6039) <= 1'b0;
    layer1_outputs(6040) <= a;
    layer1_outputs(6041) <= not (a and b);
    layer1_outputs(6042) <= a and b;
    layer1_outputs(6043) <= not (a and b);
    layer1_outputs(6044) <= a and not b;
    layer1_outputs(6045) <= not (a and b);
    layer1_outputs(6046) <= a;
    layer1_outputs(6047) <= a;
    layer1_outputs(6048) <= not (a and b);
    layer1_outputs(6049) <= a xor b;
    layer1_outputs(6050) <= not b or a;
    layer1_outputs(6051) <= not b;
    layer1_outputs(6052) <= a and b;
    layer1_outputs(6053) <= 1'b0;
    layer1_outputs(6054) <= a and not b;
    layer1_outputs(6055) <= not b or a;
    layer1_outputs(6056) <= not (a and b);
    layer1_outputs(6057) <= a and b;
    layer1_outputs(6058) <= a and b;
    layer1_outputs(6059) <= 1'b1;
    layer1_outputs(6060) <= not b;
    layer1_outputs(6061) <= a and not b;
    layer1_outputs(6062) <= not a or b;
    layer1_outputs(6063) <= not b or a;
    layer1_outputs(6064) <= not a;
    layer1_outputs(6065) <= not a or b;
    layer1_outputs(6066) <= not a;
    layer1_outputs(6067) <= not (a and b);
    layer1_outputs(6068) <= a or b;
    layer1_outputs(6069) <= b;
    layer1_outputs(6070) <= not a or b;
    layer1_outputs(6071) <= 1'b0;
    layer1_outputs(6072) <= not (a and b);
    layer1_outputs(6073) <= b and not a;
    layer1_outputs(6074) <= not (a or b);
    layer1_outputs(6075) <= not (a xor b);
    layer1_outputs(6076) <= b;
    layer1_outputs(6077) <= not a;
    layer1_outputs(6078) <= 1'b1;
    layer1_outputs(6079) <= b and not a;
    layer1_outputs(6080) <= a and b;
    layer1_outputs(6081) <= b;
    layer1_outputs(6082) <= b and not a;
    layer1_outputs(6083) <= b and not a;
    layer1_outputs(6084) <= not b or a;
    layer1_outputs(6085) <= a or b;
    layer1_outputs(6086) <= b and not a;
    layer1_outputs(6087) <= not a or b;
    layer1_outputs(6088) <= 1'b1;
    layer1_outputs(6089) <= 1'b1;
    layer1_outputs(6090) <= not a;
    layer1_outputs(6091) <= not (a or b);
    layer1_outputs(6092) <= b and not a;
    layer1_outputs(6093) <= a and b;
    layer1_outputs(6094) <= 1'b0;
    layer1_outputs(6095) <= not b;
    layer1_outputs(6096) <= not a;
    layer1_outputs(6097) <= a and not b;
    layer1_outputs(6098) <= b;
    layer1_outputs(6099) <= b;
    layer1_outputs(6100) <= not a;
    layer1_outputs(6101) <= not a;
    layer1_outputs(6102) <= 1'b0;
    layer1_outputs(6103) <= a or b;
    layer1_outputs(6104) <= not a or b;
    layer1_outputs(6105) <= 1'b0;
    layer1_outputs(6106) <= 1'b0;
    layer1_outputs(6107) <= not b;
    layer1_outputs(6108) <= not a or b;
    layer1_outputs(6109) <= b and not a;
    layer1_outputs(6110) <= not a;
    layer1_outputs(6111) <= b;
    layer1_outputs(6112) <= not b or a;
    layer1_outputs(6113) <= b;
    layer1_outputs(6114) <= not a or b;
    layer1_outputs(6115) <= b and not a;
    layer1_outputs(6116) <= a and not b;
    layer1_outputs(6117) <= not a or b;
    layer1_outputs(6118) <= a and not b;
    layer1_outputs(6119) <= not (a or b);
    layer1_outputs(6120) <= not b or a;
    layer1_outputs(6121) <= b;
    layer1_outputs(6122) <= a or b;
    layer1_outputs(6123) <= a xor b;
    layer1_outputs(6124) <= 1'b0;
    layer1_outputs(6125) <= not b;
    layer1_outputs(6126) <= not (a xor b);
    layer1_outputs(6127) <= 1'b0;
    layer1_outputs(6128) <= not (a and b);
    layer1_outputs(6129) <= not (a or b);
    layer1_outputs(6130) <= a;
    layer1_outputs(6131) <= not a or b;
    layer1_outputs(6132) <= not (a or b);
    layer1_outputs(6133) <= a and b;
    layer1_outputs(6134) <= 1'b1;
    layer1_outputs(6135) <= b and not a;
    layer1_outputs(6136) <= a and not b;
    layer1_outputs(6137) <= a or b;
    layer1_outputs(6138) <= not a or b;
    layer1_outputs(6139) <= not (a and b);
    layer1_outputs(6140) <= a xor b;
    layer1_outputs(6141) <= 1'b1;
    layer1_outputs(6142) <= a or b;
    layer1_outputs(6143) <= not b or a;
    layer1_outputs(6144) <= 1'b1;
    layer1_outputs(6145) <= not a;
    layer1_outputs(6146) <= a xor b;
    layer1_outputs(6147) <= a or b;
    layer1_outputs(6148) <= b;
    layer1_outputs(6149) <= not a;
    layer1_outputs(6150) <= not (a and b);
    layer1_outputs(6151) <= b and not a;
    layer1_outputs(6152) <= not (a and b);
    layer1_outputs(6153) <= not a or b;
    layer1_outputs(6154) <= not b;
    layer1_outputs(6155) <= a and b;
    layer1_outputs(6156) <= b and not a;
    layer1_outputs(6157) <= a or b;
    layer1_outputs(6158) <= b and not a;
    layer1_outputs(6159) <= not b or a;
    layer1_outputs(6160) <= b and not a;
    layer1_outputs(6161) <= 1'b1;
    layer1_outputs(6162) <= not (a and b);
    layer1_outputs(6163) <= not (a and b);
    layer1_outputs(6164) <= a;
    layer1_outputs(6165) <= a or b;
    layer1_outputs(6166) <= not (a xor b);
    layer1_outputs(6167) <= not b or a;
    layer1_outputs(6168) <= b;
    layer1_outputs(6169) <= 1'b1;
    layer1_outputs(6170) <= not b;
    layer1_outputs(6171) <= 1'b1;
    layer1_outputs(6172) <= a;
    layer1_outputs(6173) <= not (a and b);
    layer1_outputs(6174) <= 1'b1;
    layer1_outputs(6175) <= b;
    layer1_outputs(6176) <= 1'b1;
    layer1_outputs(6177) <= 1'b0;
    layer1_outputs(6178) <= not a or b;
    layer1_outputs(6179) <= a;
    layer1_outputs(6180) <= a and not b;
    layer1_outputs(6181) <= 1'b0;
    layer1_outputs(6182) <= not (a xor b);
    layer1_outputs(6183) <= a xor b;
    layer1_outputs(6184) <= a xor b;
    layer1_outputs(6185) <= a xor b;
    layer1_outputs(6186) <= a and b;
    layer1_outputs(6187) <= not b;
    layer1_outputs(6188) <= a and not b;
    layer1_outputs(6189) <= a or b;
    layer1_outputs(6190) <= a or b;
    layer1_outputs(6191) <= a;
    layer1_outputs(6192) <= a and b;
    layer1_outputs(6193) <= 1'b1;
    layer1_outputs(6194) <= a and not b;
    layer1_outputs(6195) <= 1'b1;
    layer1_outputs(6196) <= 1'b1;
    layer1_outputs(6197) <= a and not b;
    layer1_outputs(6198) <= not (a or b);
    layer1_outputs(6199) <= not b;
    layer1_outputs(6200) <= b;
    layer1_outputs(6201) <= not (a xor b);
    layer1_outputs(6202) <= not (a and b);
    layer1_outputs(6203) <= not b;
    layer1_outputs(6204) <= a or b;
    layer1_outputs(6205) <= b and not a;
    layer1_outputs(6206) <= not (a and b);
    layer1_outputs(6207) <= b and not a;
    layer1_outputs(6208) <= not a;
    layer1_outputs(6209) <= 1'b1;
    layer1_outputs(6210) <= not a or b;
    layer1_outputs(6211) <= b;
    layer1_outputs(6212) <= a and b;
    layer1_outputs(6213) <= not a;
    layer1_outputs(6214) <= not (a and b);
    layer1_outputs(6215) <= a xor b;
    layer1_outputs(6216) <= a;
    layer1_outputs(6217) <= not b or a;
    layer1_outputs(6218) <= b and not a;
    layer1_outputs(6219) <= not a or b;
    layer1_outputs(6220) <= a;
    layer1_outputs(6221) <= a;
    layer1_outputs(6222) <= not (a or b);
    layer1_outputs(6223) <= b and not a;
    layer1_outputs(6224) <= a xor b;
    layer1_outputs(6225) <= not b or a;
    layer1_outputs(6226) <= 1'b0;
    layer1_outputs(6227) <= 1'b0;
    layer1_outputs(6228) <= not (a or b);
    layer1_outputs(6229) <= not a or b;
    layer1_outputs(6230) <= 1'b1;
    layer1_outputs(6231) <= 1'b0;
    layer1_outputs(6232) <= not a;
    layer1_outputs(6233) <= a or b;
    layer1_outputs(6234) <= not a or b;
    layer1_outputs(6235) <= not a or b;
    layer1_outputs(6236) <= not (a and b);
    layer1_outputs(6237) <= not a;
    layer1_outputs(6238) <= not (a and b);
    layer1_outputs(6239) <= not (a and b);
    layer1_outputs(6240) <= a or b;
    layer1_outputs(6241) <= not (a and b);
    layer1_outputs(6242) <= b and not a;
    layer1_outputs(6243) <= not a;
    layer1_outputs(6244) <= a and not b;
    layer1_outputs(6245) <= b;
    layer1_outputs(6246) <= b;
    layer1_outputs(6247) <= 1'b1;
    layer1_outputs(6248) <= not (a and b);
    layer1_outputs(6249) <= b;
    layer1_outputs(6250) <= not (a and b);
    layer1_outputs(6251) <= b;
    layer1_outputs(6252) <= not (a or b);
    layer1_outputs(6253) <= a;
    layer1_outputs(6254) <= not (a and b);
    layer1_outputs(6255) <= a and b;
    layer1_outputs(6256) <= 1'b1;
    layer1_outputs(6257) <= a and not b;
    layer1_outputs(6258) <= a and b;
    layer1_outputs(6259) <= a and not b;
    layer1_outputs(6260) <= a xor b;
    layer1_outputs(6261) <= a and not b;
    layer1_outputs(6262) <= b;
    layer1_outputs(6263) <= a and not b;
    layer1_outputs(6264) <= 1'b1;
    layer1_outputs(6265) <= a;
    layer1_outputs(6266) <= a;
    layer1_outputs(6267) <= b and not a;
    layer1_outputs(6268) <= b;
    layer1_outputs(6269) <= not (a xor b);
    layer1_outputs(6270) <= not (a xor b);
    layer1_outputs(6271) <= b and not a;
    layer1_outputs(6272) <= not (a or b);
    layer1_outputs(6273) <= not (a or b);
    layer1_outputs(6274) <= a and not b;
    layer1_outputs(6275) <= b and not a;
    layer1_outputs(6276) <= 1'b0;
    layer1_outputs(6277) <= a;
    layer1_outputs(6278) <= a or b;
    layer1_outputs(6279) <= a;
    layer1_outputs(6280) <= a and b;
    layer1_outputs(6281) <= not b or a;
    layer1_outputs(6282) <= a or b;
    layer1_outputs(6283) <= not b or a;
    layer1_outputs(6284) <= 1'b1;
    layer1_outputs(6285) <= 1'b0;
    layer1_outputs(6286) <= 1'b1;
    layer1_outputs(6287) <= 1'b0;
    layer1_outputs(6288) <= 1'b0;
    layer1_outputs(6289) <= 1'b1;
    layer1_outputs(6290) <= 1'b1;
    layer1_outputs(6291) <= a and not b;
    layer1_outputs(6292) <= a and b;
    layer1_outputs(6293) <= b and not a;
    layer1_outputs(6294) <= not a or b;
    layer1_outputs(6295) <= not b or a;
    layer1_outputs(6296) <= 1'b1;
    layer1_outputs(6297) <= not b;
    layer1_outputs(6298) <= a and b;
    layer1_outputs(6299) <= not a;
    layer1_outputs(6300) <= a;
    layer1_outputs(6301) <= a xor b;
    layer1_outputs(6302) <= not (a and b);
    layer1_outputs(6303) <= a and not b;
    layer1_outputs(6304) <= b and not a;
    layer1_outputs(6305) <= 1'b0;
    layer1_outputs(6306) <= not a;
    layer1_outputs(6307) <= a and not b;
    layer1_outputs(6308) <= a xor b;
    layer1_outputs(6309) <= a;
    layer1_outputs(6310) <= 1'b0;
    layer1_outputs(6311) <= not b;
    layer1_outputs(6312) <= 1'b0;
    layer1_outputs(6313) <= a and not b;
    layer1_outputs(6314) <= not a or b;
    layer1_outputs(6315) <= not a or b;
    layer1_outputs(6316) <= not a;
    layer1_outputs(6317) <= a and not b;
    layer1_outputs(6318) <= not (a xor b);
    layer1_outputs(6319) <= a;
    layer1_outputs(6320) <= 1'b0;
    layer1_outputs(6321) <= not b or a;
    layer1_outputs(6322) <= not b;
    layer1_outputs(6323) <= 1'b1;
    layer1_outputs(6324) <= a and b;
    layer1_outputs(6325) <= not b;
    layer1_outputs(6326) <= a and b;
    layer1_outputs(6327) <= not b or a;
    layer1_outputs(6328) <= not (a xor b);
    layer1_outputs(6329) <= not (a and b);
    layer1_outputs(6330) <= not a or b;
    layer1_outputs(6331) <= not (a xor b);
    layer1_outputs(6332) <= a and b;
    layer1_outputs(6333) <= not b or a;
    layer1_outputs(6334) <= not b or a;
    layer1_outputs(6335) <= not b or a;
    layer1_outputs(6336) <= not a or b;
    layer1_outputs(6337) <= 1'b1;
    layer1_outputs(6338) <= a and not b;
    layer1_outputs(6339) <= b and not a;
    layer1_outputs(6340) <= not b or a;
    layer1_outputs(6341) <= a and not b;
    layer1_outputs(6342) <= b;
    layer1_outputs(6343) <= 1'b0;
    layer1_outputs(6344) <= b and not a;
    layer1_outputs(6345) <= a or b;
    layer1_outputs(6346) <= a and b;
    layer1_outputs(6347) <= not b;
    layer1_outputs(6348) <= not (a and b);
    layer1_outputs(6349) <= not a;
    layer1_outputs(6350) <= not a;
    layer1_outputs(6351) <= not (a or b);
    layer1_outputs(6352) <= a and b;
    layer1_outputs(6353) <= not (a and b);
    layer1_outputs(6354) <= not b or a;
    layer1_outputs(6355) <= a and not b;
    layer1_outputs(6356) <= 1'b1;
    layer1_outputs(6357) <= b and not a;
    layer1_outputs(6358) <= a and not b;
    layer1_outputs(6359) <= not (a and b);
    layer1_outputs(6360) <= not (a xor b);
    layer1_outputs(6361) <= 1'b0;
    layer1_outputs(6362) <= 1'b1;
    layer1_outputs(6363) <= a and not b;
    layer1_outputs(6364) <= not (a or b);
    layer1_outputs(6365) <= 1'b1;
    layer1_outputs(6366) <= 1'b0;
    layer1_outputs(6367) <= a and b;
    layer1_outputs(6368) <= a and b;
    layer1_outputs(6369) <= not b or a;
    layer1_outputs(6370) <= b;
    layer1_outputs(6371) <= b;
    layer1_outputs(6372) <= 1'b1;
    layer1_outputs(6373) <= a and b;
    layer1_outputs(6374) <= not (a xor b);
    layer1_outputs(6375) <= a xor b;
    layer1_outputs(6376) <= b and not a;
    layer1_outputs(6377) <= a or b;
    layer1_outputs(6378) <= b;
    layer1_outputs(6379) <= b and not a;
    layer1_outputs(6380) <= a;
    layer1_outputs(6381) <= 1'b0;
    layer1_outputs(6382) <= not (a xor b);
    layer1_outputs(6383) <= not a or b;
    layer1_outputs(6384) <= a;
    layer1_outputs(6385) <= b;
    layer1_outputs(6386) <= a;
    layer1_outputs(6387) <= 1'b1;
    layer1_outputs(6388) <= b and not a;
    layer1_outputs(6389) <= a and not b;
    layer1_outputs(6390) <= not a or b;
    layer1_outputs(6391) <= not b;
    layer1_outputs(6392) <= not (a and b);
    layer1_outputs(6393) <= 1'b1;
    layer1_outputs(6394) <= a xor b;
    layer1_outputs(6395) <= a;
    layer1_outputs(6396) <= a;
    layer1_outputs(6397) <= a and not b;
    layer1_outputs(6398) <= 1'b1;
    layer1_outputs(6399) <= not (a or b);
    layer1_outputs(6400) <= 1'b1;
    layer1_outputs(6401) <= not b;
    layer1_outputs(6402) <= b and not a;
    layer1_outputs(6403) <= not b;
    layer1_outputs(6404) <= not b or a;
    layer1_outputs(6405) <= not b or a;
    layer1_outputs(6406) <= a xor b;
    layer1_outputs(6407) <= a and not b;
    layer1_outputs(6408) <= a and b;
    layer1_outputs(6409) <= a xor b;
    layer1_outputs(6410) <= not b;
    layer1_outputs(6411) <= 1'b0;
    layer1_outputs(6412) <= 1'b0;
    layer1_outputs(6413) <= a;
    layer1_outputs(6414) <= not b or a;
    layer1_outputs(6415) <= b and not a;
    layer1_outputs(6416) <= a and not b;
    layer1_outputs(6417) <= 1'b1;
    layer1_outputs(6418) <= not a;
    layer1_outputs(6419) <= not (a or b);
    layer1_outputs(6420) <= a and b;
    layer1_outputs(6421) <= b and not a;
    layer1_outputs(6422) <= b;
    layer1_outputs(6423) <= not a or b;
    layer1_outputs(6424) <= 1'b0;
    layer1_outputs(6425) <= a and not b;
    layer1_outputs(6426) <= not (a or b);
    layer1_outputs(6427) <= a and b;
    layer1_outputs(6428) <= not (a and b);
    layer1_outputs(6429) <= b;
    layer1_outputs(6430) <= not a;
    layer1_outputs(6431) <= b;
    layer1_outputs(6432) <= b and not a;
    layer1_outputs(6433) <= 1'b1;
    layer1_outputs(6434) <= 1'b1;
    layer1_outputs(6435) <= not a;
    layer1_outputs(6436) <= a or b;
    layer1_outputs(6437) <= b and not a;
    layer1_outputs(6438) <= 1'b1;
    layer1_outputs(6439) <= 1'b1;
    layer1_outputs(6440) <= 1'b0;
    layer1_outputs(6441) <= b;
    layer1_outputs(6442) <= a and not b;
    layer1_outputs(6443) <= a and b;
    layer1_outputs(6444) <= not (a or b);
    layer1_outputs(6445) <= not a;
    layer1_outputs(6446) <= b and not a;
    layer1_outputs(6447) <= b;
    layer1_outputs(6448) <= 1'b0;
    layer1_outputs(6449) <= not a;
    layer1_outputs(6450) <= a and b;
    layer1_outputs(6451) <= a;
    layer1_outputs(6452) <= b and not a;
    layer1_outputs(6453) <= not a or b;
    layer1_outputs(6454) <= b and not a;
    layer1_outputs(6455) <= a and not b;
    layer1_outputs(6456) <= a and not b;
    layer1_outputs(6457) <= not (a xor b);
    layer1_outputs(6458) <= a xor b;
    layer1_outputs(6459) <= 1'b1;
    layer1_outputs(6460) <= a or b;
    layer1_outputs(6461) <= not b;
    layer1_outputs(6462) <= 1'b0;
    layer1_outputs(6463) <= not b;
    layer1_outputs(6464) <= a or b;
    layer1_outputs(6465) <= not (a and b);
    layer1_outputs(6466) <= b;
    layer1_outputs(6467) <= not (a or b);
    layer1_outputs(6468) <= not a;
    layer1_outputs(6469) <= a xor b;
    layer1_outputs(6470) <= not b or a;
    layer1_outputs(6471) <= a or b;
    layer1_outputs(6472) <= 1'b0;
    layer1_outputs(6473) <= a or b;
    layer1_outputs(6474) <= not (a and b);
    layer1_outputs(6475) <= a and not b;
    layer1_outputs(6476) <= b and not a;
    layer1_outputs(6477) <= 1'b0;
    layer1_outputs(6478) <= not (a or b);
    layer1_outputs(6479) <= a;
    layer1_outputs(6480) <= 1'b1;
    layer1_outputs(6481) <= b;
    layer1_outputs(6482) <= not a or b;
    layer1_outputs(6483) <= 1'b0;
    layer1_outputs(6484) <= not b;
    layer1_outputs(6485) <= not (a or b);
    layer1_outputs(6486) <= a;
    layer1_outputs(6487) <= b and not a;
    layer1_outputs(6488) <= 1'b0;
    layer1_outputs(6489) <= b and not a;
    layer1_outputs(6490) <= a and not b;
    layer1_outputs(6491) <= not b;
    layer1_outputs(6492) <= a and not b;
    layer1_outputs(6493) <= b and not a;
    layer1_outputs(6494) <= 1'b1;
    layer1_outputs(6495) <= not a;
    layer1_outputs(6496) <= not b or a;
    layer1_outputs(6497) <= b and not a;
    layer1_outputs(6498) <= b and not a;
    layer1_outputs(6499) <= b;
    layer1_outputs(6500) <= not a;
    layer1_outputs(6501) <= not a or b;
    layer1_outputs(6502) <= 1'b0;
    layer1_outputs(6503) <= not (a and b);
    layer1_outputs(6504) <= 1'b1;
    layer1_outputs(6505) <= a;
    layer1_outputs(6506) <= not a or b;
    layer1_outputs(6507) <= a and not b;
    layer1_outputs(6508) <= a;
    layer1_outputs(6509) <= 1'b0;
    layer1_outputs(6510) <= 1'b0;
    layer1_outputs(6511) <= 1'b0;
    layer1_outputs(6512) <= not a or b;
    layer1_outputs(6513) <= b and not a;
    layer1_outputs(6514) <= a xor b;
    layer1_outputs(6515) <= not a;
    layer1_outputs(6516) <= 1'b1;
    layer1_outputs(6517) <= a;
    layer1_outputs(6518) <= a and not b;
    layer1_outputs(6519) <= a and b;
    layer1_outputs(6520) <= not b or a;
    layer1_outputs(6521) <= 1'b1;
    layer1_outputs(6522) <= a;
    layer1_outputs(6523) <= a xor b;
    layer1_outputs(6524) <= b and not a;
    layer1_outputs(6525) <= a;
    layer1_outputs(6526) <= not a;
    layer1_outputs(6527) <= not a or b;
    layer1_outputs(6528) <= 1'b0;
    layer1_outputs(6529) <= not a or b;
    layer1_outputs(6530) <= a or b;
    layer1_outputs(6531) <= not b or a;
    layer1_outputs(6532) <= a and b;
    layer1_outputs(6533) <= a and not b;
    layer1_outputs(6534) <= a and not b;
    layer1_outputs(6535) <= b and not a;
    layer1_outputs(6536) <= not a;
    layer1_outputs(6537) <= b;
    layer1_outputs(6538) <= 1'b0;
    layer1_outputs(6539) <= b and not a;
    layer1_outputs(6540) <= b and not a;
    layer1_outputs(6541) <= not b or a;
    layer1_outputs(6542) <= not (a or b);
    layer1_outputs(6543) <= b;
    layer1_outputs(6544) <= 1'b1;
    layer1_outputs(6545) <= a and not b;
    layer1_outputs(6546) <= a and b;
    layer1_outputs(6547) <= not (a and b);
    layer1_outputs(6548) <= b;
    layer1_outputs(6549) <= not (a xor b);
    layer1_outputs(6550) <= a;
    layer1_outputs(6551) <= a;
    layer1_outputs(6552) <= not (a and b);
    layer1_outputs(6553) <= not (a or b);
    layer1_outputs(6554) <= not (a and b);
    layer1_outputs(6555) <= a;
    layer1_outputs(6556) <= not (a xor b);
    layer1_outputs(6557) <= a and not b;
    layer1_outputs(6558) <= a;
    layer1_outputs(6559) <= 1'b1;
    layer1_outputs(6560) <= a;
    layer1_outputs(6561) <= 1'b1;
    layer1_outputs(6562) <= a and not b;
    layer1_outputs(6563) <= 1'b0;
    layer1_outputs(6564) <= a and b;
    layer1_outputs(6565) <= not (a and b);
    layer1_outputs(6566) <= not (a or b);
    layer1_outputs(6567) <= not a or b;
    layer1_outputs(6568) <= b and not a;
    layer1_outputs(6569) <= 1'b0;
    layer1_outputs(6570) <= not b;
    layer1_outputs(6571) <= a xor b;
    layer1_outputs(6572) <= 1'b1;
    layer1_outputs(6573) <= not (a or b);
    layer1_outputs(6574) <= not a;
    layer1_outputs(6575) <= a or b;
    layer1_outputs(6576) <= a and not b;
    layer1_outputs(6577) <= not b or a;
    layer1_outputs(6578) <= a;
    layer1_outputs(6579) <= not b or a;
    layer1_outputs(6580) <= a and b;
    layer1_outputs(6581) <= not (a or b);
    layer1_outputs(6582) <= 1'b1;
    layer1_outputs(6583) <= 1'b1;
    layer1_outputs(6584) <= a;
    layer1_outputs(6585) <= b;
    layer1_outputs(6586) <= 1'b1;
    layer1_outputs(6587) <= a xor b;
    layer1_outputs(6588) <= not a;
    layer1_outputs(6589) <= not a;
    layer1_outputs(6590) <= not (a and b);
    layer1_outputs(6591) <= not (a and b);
    layer1_outputs(6592) <= 1'b0;
    layer1_outputs(6593) <= a and not b;
    layer1_outputs(6594) <= a and not b;
    layer1_outputs(6595) <= not a;
    layer1_outputs(6596) <= not a;
    layer1_outputs(6597) <= not b or a;
    layer1_outputs(6598) <= a or b;
    layer1_outputs(6599) <= a and b;
    layer1_outputs(6600) <= 1'b1;
    layer1_outputs(6601) <= b and not a;
    layer1_outputs(6602) <= a and b;
    layer1_outputs(6603) <= not a or b;
    layer1_outputs(6604) <= b;
    layer1_outputs(6605) <= 1'b0;
    layer1_outputs(6606) <= a or b;
    layer1_outputs(6607) <= 1'b1;
    layer1_outputs(6608) <= not b or a;
    layer1_outputs(6609) <= not (a or b);
    layer1_outputs(6610) <= a and b;
    layer1_outputs(6611) <= not (a and b);
    layer1_outputs(6612) <= a xor b;
    layer1_outputs(6613) <= not a;
    layer1_outputs(6614) <= not a or b;
    layer1_outputs(6615) <= a xor b;
    layer1_outputs(6616) <= 1'b0;
    layer1_outputs(6617) <= a;
    layer1_outputs(6618) <= a and not b;
    layer1_outputs(6619) <= a and not b;
    layer1_outputs(6620) <= not (a or b);
    layer1_outputs(6621) <= a;
    layer1_outputs(6622) <= 1'b0;
    layer1_outputs(6623) <= 1'b0;
    layer1_outputs(6624) <= not (a or b);
    layer1_outputs(6625) <= 1'b0;
    layer1_outputs(6626) <= a xor b;
    layer1_outputs(6627) <= not a;
    layer1_outputs(6628) <= not a;
    layer1_outputs(6629) <= not (a or b);
    layer1_outputs(6630) <= not a or b;
    layer1_outputs(6631) <= b and not a;
    layer1_outputs(6632) <= not a;
    layer1_outputs(6633) <= a xor b;
    layer1_outputs(6634) <= 1'b0;
    layer1_outputs(6635) <= not (a xor b);
    layer1_outputs(6636) <= not a;
    layer1_outputs(6637) <= not (a or b);
    layer1_outputs(6638) <= not a;
    layer1_outputs(6639) <= not a or b;
    layer1_outputs(6640) <= a;
    layer1_outputs(6641) <= 1'b1;
    layer1_outputs(6642) <= a and b;
    layer1_outputs(6643) <= a or b;
    layer1_outputs(6644) <= not (a or b);
    layer1_outputs(6645) <= 1'b1;
    layer1_outputs(6646) <= a and not b;
    layer1_outputs(6647) <= b;
    layer1_outputs(6648) <= not a;
    layer1_outputs(6649) <= not b;
    layer1_outputs(6650) <= 1'b1;
    layer1_outputs(6651) <= a and b;
    layer1_outputs(6652) <= a and b;
    layer1_outputs(6653) <= 1'b0;
    layer1_outputs(6654) <= not a or b;
    layer1_outputs(6655) <= a and b;
    layer1_outputs(6656) <= not (a or b);
    layer1_outputs(6657) <= not a or b;
    layer1_outputs(6658) <= 1'b0;
    layer1_outputs(6659) <= not a;
    layer1_outputs(6660) <= not (a or b);
    layer1_outputs(6661) <= not (a or b);
    layer1_outputs(6662) <= b;
    layer1_outputs(6663) <= a and b;
    layer1_outputs(6664) <= a;
    layer1_outputs(6665) <= not (a or b);
    layer1_outputs(6666) <= a and b;
    layer1_outputs(6667) <= not b;
    layer1_outputs(6668) <= a or b;
    layer1_outputs(6669) <= a and not b;
    layer1_outputs(6670) <= 1'b0;
    layer1_outputs(6671) <= b;
    layer1_outputs(6672) <= 1'b0;
    layer1_outputs(6673) <= not a or b;
    layer1_outputs(6674) <= a;
    layer1_outputs(6675) <= b and not a;
    layer1_outputs(6676) <= a or b;
    layer1_outputs(6677) <= not b or a;
    layer1_outputs(6678) <= a and not b;
    layer1_outputs(6679) <= not (a or b);
    layer1_outputs(6680) <= not b or a;
    layer1_outputs(6681) <= not b;
    layer1_outputs(6682) <= not b or a;
    layer1_outputs(6683) <= not b or a;
    layer1_outputs(6684) <= b;
    layer1_outputs(6685) <= not a or b;
    layer1_outputs(6686) <= a and not b;
    layer1_outputs(6687) <= a and b;
    layer1_outputs(6688) <= not (a xor b);
    layer1_outputs(6689) <= b and not a;
    layer1_outputs(6690) <= 1'b0;
    layer1_outputs(6691) <= not a or b;
    layer1_outputs(6692) <= not a or b;
    layer1_outputs(6693) <= not b;
    layer1_outputs(6694) <= a xor b;
    layer1_outputs(6695) <= a or b;
    layer1_outputs(6696) <= a and not b;
    layer1_outputs(6697) <= a and b;
    layer1_outputs(6698) <= a or b;
    layer1_outputs(6699) <= b;
    layer1_outputs(6700) <= a or b;
    layer1_outputs(6701) <= not (a and b);
    layer1_outputs(6702) <= not b or a;
    layer1_outputs(6703) <= a and b;
    layer1_outputs(6704) <= not b;
    layer1_outputs(6705) <= a or b;
    layer1_outputs(6706) <= b;
    layer1_outputs(6707) <= a or b;
    layer1_outputs(6708) <= a and b;
    layer1_outputs(6709) <= a and b;
    layer1_outputs(6710) <= a;
    layer1_outputs(6711) <= not b;
    layer1_outputs(6712) <= not a or b;
    layer1_outputs(6713) <= not a or b;
    layer1_outputs(6714) <= not a or b;
    layer1_outputs(6715) <= b and not a;
    layer1_outputs(6716) <= 1'b0;
    layer1_outputs(6717) <= not (a or b);
    layer1_outputs(6718) <= not (a xor b);
    layer1_outputs(6719) <= a xor b;
    layer1_outputs(6720) <= not (a or b);
    layer1_outputs(6721) <= b and not a;
    layer1_outputs(6722) <= b;
    layer1_outputs(6723) <= b;
    layer1_outputs(6724) <= a xor b;
    layer1_outputs(6725) <= a or b;
    layer1_outputs(6726) <= not (a or b);
    layer1_outputs(6727) <= b and not a;
    layer1_outputs(6728) <= a and not b;
    layer1_outputs(6729) <= b and not a;
    layer1_outputs(6730) <= a and not b;
    layer1_outputs(6731) <= a and not b;
    layer1_outputs(6732) <= not b;
    layer1_outputs(6733) <= not a;
    layer1_outputs(6734) <= b and not a;
    layer1_outputs(6735) <= a and b;
    layer1_outputs(6736) <= not (a and b);
    layer1_outputs(6737) <= not b or a;
    layer1_outputs(6738) <= 1'b0;
    layer1_outputs(6739) <= not a or b;
    layer1_outputs(6740) <= a xor b;
    layer1_outputs(6741) <= not a or b;
    layer1_outputs(6742) <= not (a and b);
    layer1_outputs(6743) <= not (a and b);
    layer1_outputs(6744) <= not a or b;
    layer1_outputs(6745) <= a and not b;
    layer1_outputs(6746) <= a and not b;
    layer1_outputs(6747) <= not b;
    layer1_outputs(6748) <= a xor b;
    layer1_outputs(6749) <= not a or b;
    layer1_outputs(6750) <= not a;
    layer1_outputs(6751) <= a and not b;
    layer1_outputs(6752) <= a;
    layer1_outputs(6753) <= not (a xor b);
    layer1_outputs(6754) <= not b or a;
    layer1_outputs(6755) <= not (a or b);
    layer1_outputs(6756) <= b and not a;
    layer1_outputs(6757) <= a and not b;
    layer1_outputs(6758) <= not (a and b);
    layer1_outputs(6759) <= not b;
    layer1_outputs(6760) <= 1'b1;
    layer1_outputs(6761) <= not a;
    layer1_outputs(6762) <= not b;
    layer1_outputs(6763) <= not a or b;
    layer1_outputs(6764) <= not (a and b);
    layer1_outputs(6765) <= a or b;
    layer1_outputs(6766) <= 1'b0;
    layer1_outputs(6767) <= not b;
    layer1_outputs(6768) <= not (a or b);
    layer1_outputs(6769) <= not (a and b);
    layer1_outputs(6770) <= a and b;
    layer1_outputs(6771) <= a and b;
    layer1_outputs(6772) <= 1'b0;
    layer1_outputs(6773) <= b and not a;
    layer1_outputs(6774) <= not (a and b);
    layer1_outputs(6775) <= not (a xor b);
    layer1_outputs(6776) <= not b or a;
    layer1_outputs(6777) <= a and b;
    layer1_outputs(6778) <= a;
    layer1_outputs(6779) <= 1'b1;
    layer1_outputs(6780) <= not (a or b);
    layer1_outputs(6781) <= not (a or b);
    layer1_outputs(6782) <= a xor b;
    layer1_outputs(6783) <= b and not a;
    layer1_outputs(6784) <= not a;
    layer1_outputs(6785) <= b and not a;
    layer1_outputs(6786) <= not a or b;
    layer1_outputs(6787) <= b and not a;
    layer1_outputs(6788) <= a and b;
    layer1_outputs(6789) <= not b;
    layer1_outputs(6790) <= a and not b;
    layer1_outputs(6791) <= a or b;
    layer1_outputs(6792) <= not b;
    layer1_outputs(6793) <= 1'b0;
    layer1_outputs(6794) <= 1'b1;
    layer1_outputs(6795) <= a or b;
    layer1_outputs(6796) <= not a;
    layer1_outputs(6797) <= b and not a;
    layer1_outputs(6798) <= a or b;
    layer1_outputs(6799) <= not b;
    layer1_outputs(6800) <= not b;
    layer1_outputs(6801) <= b and not a;
    layer1_outputs(6802) <= 1'b0;
    layer1_outputs(6803) <= not b or a;
    layer1_outputs(6804) <= a or b;
    layer1_outputs(6805) <= not (a or b);
    layer1_outputs(6806) <= not a;
    layer1_outputs(6807) <= not b or a;
    layer1_outputs(6808) <= not (a and b);
    layer1_outputs(6809) <= not b or a;
    layer1_outputs(6810) <= not a or b;
    layer1_outputs(6811) <= not b;
    layer1_outputs(6812) <= 1'b1;
    layer1_outputs(6813) <= a or b;
    layer1_outputs(6814) <= not (a and b);
    layer1_outputs(6815) <= not b or a;
    layer1_outputs(6816) <= not b or a;
    layer1_outputs(6817) <= a and not b;
    layer1_outputs(6818) <= not (a or b);
    layer1_outputs(6819) <= b;
    layer1_outputs(6820) <= not a or b;
    layer1_outputs(6821) <= not (a and b);
    layer1_outputs(6822) <= not (a xor b);
    layer1_outputs(6823) <= a or b;
    layer1_outputs(6824) <= b;
    layer1_outputs(6825) <= 1'b1;
    layer1_outputs(6826) <= a xor b;
    layer1_outputs(6827) <= 1'b1;
    layer1_outputs(6828) <= not (a or b);
    layer1_outputs(6829) <= not b or a;
    layer1_outputs(6830) <= b and not a;
    layer1_outputs(6831) <= a and not b;
    layer1_outputs(6832) <= 1'b0;
    layer1_outputs(6833) <= 1'b1;
    layer1_outputs(6834) <= a and not b;
    layer1_outputs(6835) <= b and not a;
    layer1_outputs(6836) <= not b;
    layer1_outputs(6837) <= not (a xor b);
    layer1_outputs(6838) <= not a;
    layer1_outputs(6839) <= a and not b;
    layer1_outputs(6840) <= not a;
    layer1_outputs(6841) <= 1'b0;
    layer1_outputs(6842) <= b;
    layer1_outputs(6843) <= not b;
    layer1_outputs(6844) <= not b;
    layer1_outputs(6845) <= a or b;
    layer1_outputs(6846) <= 1'b1;
    layer1_outputs(6847) <= not (a and b);
    layer1_outputs(6848) <= not a or b;
    layer1_outputs(6849) <= not b;
    layer1_outputs(6850) <= 1'b1;
    layer1_outputs(6851) <= a and not b;
    layer1_outputs(6852) <= a xor b;
    layer1_outputs(6853) <= not (a xor b);
    layer1_outputs(6854) <= not a or b;
    layer1_outputs(6855) <= not (a or b);
    layer1_outputs(6856) <= a or b;
    layer1_outputs(6857) <= not b;
    layer1_outputs(6858) <= not (a and b);
    layer1_outputs(6859) <= a and b;
    layer1_outputs(6860) <= not (a or b);
    layer1_outputs(6861) <= a xor b;
    layer1_outputs(6862) <= not (a and b);
    layer1_outputs(6863) <= not b or a;
    layer1_outputs(6864) <= not a or b;
    layer1_outputs(6865) <= not a;
    layer1_outputs(6866) <= a and not b;
    layer1_outputs(6867) <= not a;
    layer1_outputs(6868) <= 1'b1;
    layer1_outputs(6869) <= b;
    layer1_outputs(6870) <= a;
    layer1_outputs(6871) <= not (a or b);
    layer1_outputs(6872) <= a and b;
    layer1_outputs(6873) <= not b or a;
    layer1_outputs(6874) <= not (a and b);
    layer1_outputs(6875) <= 1'b1;
    layer1_outputs(6876) <= not a or b;
    layer1_outputs(6877) <= a and not b;
    layer1_outputs(6878) <= a and b;
    layer1_outputs(6879) <= not (a or b);
    layer1_outputs(6880) <= not a;
    layer1_outputs(6881) <= a and b;
    layer1_outputs(6882) <= not a;
    layer1_outputs(6883) <= not b or a;
    layer1_outputs(6884) <= a or b;
    layer1_outputs(6885) <= a and not b;
    layer1_outputs(6886) <= b and not a;
    layer1_outputs(6887) <= not a or b;
    layer1_outputs(6888) <= a and not b;
    layer1_outputs(6889) <= 1'b1;
    layer1_outputs(6890) <= 1'b0;
    layer1_outputs(6891) <= b and not a;
    layer1_outputs(6892) <= not (a or b);
    layer1_outputs(6893) <= 1'b1;
    layer1_outputs(6894) <= a;
    layer1_outputs(6895) <= 1'b1;
    layer1_outputs(6896) <= not (a and b);
    layer1_outputs(6897) <= b and not a;
    layer1_outputs(6898) <= not (a and b);
    layer1_outputs(6899) <= not b;
    layer1_outputs(6900) <= 1'b1;
    layer1_outputs(6901) <= a and not b;
    layer1_outputs(6902) <= not b;
    layer1_outputs(6903) <= 1'b0;
    layer1_outputs(6904) <= not a;
    layer1_outputs(6905) <= not b or a;
    layer1_outputs(6906) <= not (a xor b);
    layer1_outputs(6907) <= not b;
    layer1_outputs(6908) <= a and not b;
    layer1_outputs(6909) <= not a or b;
    layer1_outputs(6910) <= not (a or b);
    layer1_outputs(6911) <= not b;
    layer1_outputs(6912) <= 1'b0;
    layer1_outputs(6913) <= not b;
    layer1_outputs(6914) <= not (a or b);
    layer1_outputs(6915) <= a and not b;
    layer1_outputs(6916) <= a and b;
    layer1_outputs(6917) <= 1'b0;
    layer1_outputs(6918) <= 1'b1;
    layer1_outputs(6919) <= b and not a;
    layer1_outputs(6920) <= 1'b1;
    layer1_outputs(6921) <= 1'b1;
    layer1_outputs(6922) <= a and b;
    layer1_outputs(6923) <= a;
    layer1_outputs(6924) <= a and not b;
    layer1_outputs(6925) <= a and b;
    layer1_outputs(6926) <= not a or b;
    layer1_outputs(6927) <= 1'b0;
    layer1_outputs(6928) <= not b;
    layer1_outputs(6929) <= not a;
    layer1_outputs(6930) <= b;
    layer1_outputs(6931) <= a xor b;
    layer1_outputs(6932) <= a xor b;
    layer1_outputs(6933) <= not (a and b);
    layer1_outputs(6934) <= not a or b;
    layer1_outputs(6935) <= not b or a;
    layer1_outputs(6936) <= a;
    layer1_outputs(6937) <= 1'b1;
    layer1_outputs(6938) <= 1'b0;
    layer1_outputs(6939) <= a;
    layer1_outputs(6940) <= not (a and b);
    layer1_outputs(6941) <= not a;
    layer1_outputs(6942) <= not b;
    layer1_outputs(6943) <= not a or b;
    layer1_outputs(6944) <= a and not b;
    layer1_outputs(6945) <= not a or b;
    layer1_outputs(6946) <= a and b;
    layer1_outputs(6947) <= not a;
    layer1_outputs(6948) <= not b;
    layer1_outputs(6949) <= a and not b;
    layer1_outputs(6950) <= not b or a;
    layer1_outputs(6951) <= not b or a;
    layer1_outputs(6952) <= a and b;
    layer1_outputs(6953) <= b and not a;
    layer1_outputs(6954) <= not (a or b);
    layer1_outputs(6955) <= a;
    layer1_outputs(6956) <= not (a and b);
    layer1_outputs(6957) <= a and not b;
    layer1_outputs(6958) <= b;
    layer1_outputs(6959) <= not a;
    layer1_outputs(6960) <= not b;
    layer1_outputs(6961) <= not b or a;
    layer1_outputs(6962) <= not (a or b);
    layer1_outputs(6963) <= not b or a;
    layer1_outputs(6964) <= 1'b1;
    layer1_outputs(6965) <= not a or b;
    layer1_outputs(6966) <= b and not a;
    layer1_outputs(6967) <= 1'b0;
    layer1_outputs(6968) <= not (a or b);
    layer1_outputs(6969) <= not b or a;
    layer1_outputs(6970) <= 1'b1;
    layer1_outputs(6971) <= not a;
    layer1_outputs(6972) <= b and not a;
    layer1_outputs(6973) <= 1'b1;
    layer1_outputs(6974) <= b;
    layer1_outputs(6975) <= a or b;
    layer1_outputs(6976) <= b and not a;
    layer1_outputs(6977) <= not a or b;
    layer1_outputs(6978) <= not a or b;
    layer1_outputs(6979) <= not (a or b);
    layer1_outputs(6980) <= 1'b0;
    layer1_outputs(6981) <= 1'b1;
    layer1_outputs(6982) <= not (a and b);
    layer1_outputs(6983) <= 1'b1;
    layer1_outputs(6984) <= not (a and b);
    layer1_outputs(6985) <= b;
    layer1_outputs(6986) <= not (a xor b);
    layer1_outputs(6987) <= a and b;
    layer1_outputs(6988) <= a and not b;
    layer1_outputs(6989) <= 1'b0;
    layer1_outputs(6990) <= a;
    layer1_outputs(6991) <= 1'b1;
    layer1_outputs(6992) <= a or b;
    layer1_outputs(6993) <= a xor b;
    layer1_outputs(6994) <= 1'b1;
    layer1_outputs(6995) <= 1'b0;
    layer1_outputs(6996) <= 1'b0;
    layer1_outputs(6997) <= 1'b0;
    layer1_outputs(6998) <= not (a or b);
    layer1_outputs(6999) <= not b;
    layer1_outputs(7000) <= a and not b;
    layer1_outputs(7001) <= a and not b;
    layer1_outputs(7002) <= not b or a;
    layer1_outputs(7003) <= 1'b1;
    layer1_outputs(7004) <= a xor b;
    layer1_outputs(7005) <= b;
    layer1_outputs(7006) <= b and not a;
    layer1_outputs(7007) <= a and not b;
    layer1_outputs(7008) <= not a or b;
    layer1_outputs(7009) <= b;
    layer1_outputs(7010) <= 1'b0;
    layer1_outputs(7011) <= b;
    layer1_outputs(7012) <= 1'b1;
    layer1_outputs(7013) <= a and b;
    layer1_outputs(7014) <= a and b;
    layer1_outputs(7015) <= 1'b1;
    layer1_outputs(7016) <= not (a or b);
    layer1_outputs(7017) <= not (a or b);
    layer1_outputs(7018) <= not a;
    layer1_outputs(7019) <= not (a and b);
    layer1_outputs(7020) <= b and not a;
    layer1_outputs(7021) <= a or b;
    layer1_outputs(7022) <= not (a and b);
    layer1_outputs(7023) <= b;
    layer1_outputs(7024) <= b and not a;
    layer1_outputs(7025) <= b and not a;
    layer1_outputs(7026) <= a and b;
    layer1_outputs(7027) <= 1'b1;
    layer1_outputs(7028) <= a and b;
    layer1_outputs(7029) <= a or b;
    layer1_outputs(7030) <= not (a or b);
    layer1_outputs(7031) <= a or b;
    layer1_outputs(7032) <= 1'b0;
    layer1_outputs(7033) <= a xor b;
    layer1_outputs(7034) <= 1'b0;
    layer1_outputs(7035) <= not a;
    layer1_outputs(7036) <= not (a xor b);
    layer1_outputs(7037) <= 1'b0;
    layer1_outputs(7038) <= a;
    layer1_outputs(7039) <= 1'b0;
    layer1_outputs(7040) <= not (a and b);
    layer1_outputs(7041) <= 1'b1;
    layer1_outputs(7042) <= not (a or b);
    layer1_outputs(7043) <= b;
    layer1_outputs(7044) <= a and b;
    layer1_outputs(7045) <= not b or a;
    layer1_outputs(7046) <= 1'b0;
    layer1_outputs(7047) <= a or b;
    layer1_outputs(7048) <= not (a and b);
    layer1_outputs(7049) <= not (a and b);
    layer1_outputs(7050) <= b and not a;
    layer1_outputs(7051) <= a;
    layer1_outputs(7052) <= a xor b;
    layer1_outputs(7053) <= not a;
    layer1_outputs(7054) <= not (a or b);
    layer1_outputs(7055) <= not b;
    layer1_outputs(7056) <= a and b;
    layer1_outputs(7057) <= b;
    layer1_outputs(7058) <= a and b;
    layer1_outputs(7059) <= not b or a;
    layer1_outputs(7060) <= not (a xor b);
    layer1_outputs(7061) <= 1'b1;
    layer1_outputs(7062) <= not (a and b);
    layer1_outputs(7063) <= not b or a;
    layer1_outputs(7064) <= not a;
    layer1_outputs(7065) <= not b or a;
    layer1_outputs(7066) <= not a;
    layer1_outputs(7067) <= 1'b1;
    layer1_outputs(7068) <= not (a and b);
    layer1_outputs(7069) <= not (a or b);
    layer1_outputs(7070) <= b;
    layer1_outputs(7071) <= a and not b;
    layer1_outputs(7072) <= b;
    layer1_outputs(7073) <= b;
    layer1_outputs(7074) <= not b or a;
    layer1_outputs(7075) <= not (a and b);
    layer1_outputs(7076) <= not a or b;
    layer1_outputs(7077) <= 1'b0;
    layer1_outputs(7078) <= not a;
    layer1_outputs(7079) <= not b;
    layer1_outputs(7080) <= a and b;
    layer1_outputs(7081) <= not (a or b);
    layer1_outputs(7082) <= 1'b1;
    layer1_outputs(7083) <= b;
    layer1_outputs(7084) <= a or b;
    layer1_outputs(7085) <= not b;
    layer1_outputs(7086) <= b;
    layer1_outputs(7087) <= a or b;
    layer1_outputs(7088) <= not (a xor b);
    layer1_outputs(7089) <= a and not b;
    layer1_outputs(7090) <= b and not a;
    layer1_outputs(7091) <= not (a or b);
    layer1_outputs(7092) <= not a;
    layer1_outputs(7093) <= 1'b1;
    layer1_outputs(7094) <= not (a xor b);
    layer1_outputs(7095) <= not b;
    layer1_outputs(7096) <= not (a xor b);
    layer1_outputs(7097) <= b;
    layer1_outputs(7098) <= not a;
    layer1_outputs(7099) <= not a or b;
    layer1_outputs(7100) <= a and b;
    layer1_outputs(7101) <= a and not b;
    layer1_outputs(7102) <= a or b;
    layer1_outputs(7103) <= a;
    layer1_outputs(7104) <= a and not b;
    layer1_outputs(7105) <= not (a or b);
    layer1_outputs(7106) <= a or b;
    layer1_outputs(7107) <= b and not a;
    layer1_outputs(7108) <= b;
    layer1_outputs(7109) <= not a;
    layer1_outputs(7110) <= a xor b;
    layer1_outputs(7111) <= not b;
    layer1_outputs(7112) <= not (a or b);
    layer1_outputs(7113) <= 1'b1;
    layer1_outputs(7114) <= b and not a;
    layer1_outputs(7115) <= a or b;
    layer1_outputs(7116) <= not b or a;
    layer1_outputs(7117) <= not b or a;
    layer1_outputs(7118) <= not a or b;
    layer1_outputs(7119) <= not (a xor b);
    layer1_outputs(7120) <= a and not b;
    layer1_outputs(7121) <= b;
    layer1_outputs(7122) <= not (a or b);
    layer1_outputs(7123) <= not b;
    layer1_outputs(7124) <= a xor b;
    layer1_outputs(7125) <= 1'b1;
    layer1_outputs(7126) <= not a or b;
    layer1_outputs(7127) <= b and not a;
    layer1_outputs(7128) <= not b or a;
    layer1_outputs(7129) <= b;
    layer1_outputs(7130) <= a or b;
    layer1_outputs(7131) <= not b or a;
    layer1_outputs(7132) <= not b;
    layer1_outputs(7133) <= 1'b1;
    layer1_outputs(7134) <= b and not a;
    layer1_outputs(7135) <= 1'b1;
    layer1_outputs(7136) <= a or b;
    layer1_outputs(7137) <= not a;
    layer1_outputs(7138) <= not b or a;
    layer1_outputs(7139) <= b and not a;
    layer1_outputs(7140) <= b and not a;
    layer1_outputs(7141) <= not (a and b);
    layer1_outputs(7142) <= a or b;
    layer1_outputs(7143) <= a;
    layer1_outputs(7144) <= 1'b0;
    layer1_outputs(7145) <= b and not a;
    layer1_outputs(7146) <= not b or a;
    layer1_outputs(7147) <= 1'b0;
    layer1_outputs(7148) <= a and not b;
    layer1_outputs(7149) <= a and not b;
    layer1_outputs(7150) <= not a or b;
    layer1_outputs(7151) <= not (a and b);
    layer1_outputs(7152) <= not a or b;
    layer1_outputs(7153) <= a or b;
    layer1_outputs(7154) <= not b;
    layer1_outputs(7155) <= b and not a;
    layer1_outputs(7156) <= not b;
    layer1_outputs(7157) <= 1'b1;
    layer1_outputs(7158) <= not b;
    layer1_outputs(7159) <= not (a or b);
    layer1_outputs(7160) <= a or b;
    layer1_outputs(7161) <= a and b;
    layer1_outputs(7162) <= not (a and b);
    layer1_outputs(7163) <= b;
    layer1_outputs(7164) <= not (a xor b);
    layer1_outputs(7165) <= 1'b0;
    layer1_outputs(7166) <= not b or a;
    layer1_outputs(7167) <= not (a or b);
    layer1_outputs(7168) <= a xor b;
    layer1_outputs(7169) <= 1'b1;
    layer1_outputs(7170) <= b and not a;
    layer1_outputs(7171) <= not (a or b);
    layer1_outputs(7172) <= a and b;
    layer1_outputs(7173) <= a and not b;
    layer1_outputs(7174) <= a or b;
    layer1_outputs(7175) <= a and b;
    layer1_outputs(7176) <= 1'b0;
    layer1_outputs(7177) <= not (a and b);
    layer1_outputs(7178) <= not b;
    layer1_outputs(7179) <= not (a or b);
    layer1_outputs(7180) <= not b or a;
    layer1_outputs(7181) <= a or b;
    layer1_outputs(7182) <= b and not a;
    layer1_outputs(7183) <= not b or a;
    layer1_outputs(7184) <= not (a xor b);
    layer1_outputs(7185) <= 1'b1;
    layer1_outputs(7186) <= not (a xor b);
    layer1_outputs(7187) <= a;
    layer1_outputs(7188) <= a and b;
    layer1_outputs(7189) <= not (a or b);
    layer1_outputs(7190) <= a xor b;
    layer1_outputs(7191) <= 1'b1;
    layer1_outputs(7192) <= 1'b0;
    layer1_outputs(7193) <= 1'b0;
    layer1_outputs(7194) <= not (a or b);
    layer1_outputs(7195) <= a and not b;
    layer1_outputs(7196) <= not (a and b);
    layer1_outputs(7197) <= not a or b;
    layer1_outputs(7198) <= not a;
    layer1_outputs(7199) <= not (a and b);
    layer1_outputs(7200) <= not b;
    layer1_outputs(7201) <= b;
    layer1_outputs(7202) <= 1'b1;
    layer1_outputs(7203) <= not b;
    layer1_outputs(7204) <= 1'b1;
    layer1_outputs(7205) <= 1'b1;
    layer1_outputs(7206) <= 1'b1;
    layer1_outputs(7207) <= not (a or b);
    layer1_outputs(7208) <= b;
    layer1_outputs(7209) <= b and not a;
    layer1_outputs(7210) <= not (a or b);
    layer1_outputs(7211) <= a or b;
    layer1_outputs(7212) <= a and b;
    layer1_outputs(7213) <= a or b;
    layer1_outputs(7214) <= 1'b0;
    layer1_outputs(7215) <= not b;
    layer1_outputs(7216) <= not b or a;
    layer1_outputs(7217) <= 1'b1;
    layer1_outputs(7218) <= not b or a;
    layer1_outputs(7219) <= a and not b;
    layer1_outputs(7220) <= a or b;
    layer1_outputs(7221) <= 1'b1;
    layer1_outputs(7222) <= b and not a;
    layer1_outputs(7223) <= a and b;
    layer1_outputs(7224) <= not b;
    layer1_outputs(7225) <= a and not b;
    layer1_outputs(7226) <= not (a or b);
    layer1_outputs(7227) <= a and not b;
    layer1_outputs(7228) <= not (a xor b);
    layer1_outputs(7229) <= not (a xor b);
    layer1_outputs(7230) <= not a or b;
    layer1_outputs(7231) <= not b or a;
    layer1_outputs(7232) <= a and not b;
    layer1_outputs(7233) <= 1'b1;
    layer1_outputs(7234) <= a and b;
    layer1_outputs(7235) <= 1'b1;
    layer1_outputs(7236) <= a and b;
    layer1_outputs(7237) <= b and not a;
    layer1_outputs(7238) <= 1'b0;
    layer1_outputs(7239) <= not b or a;
    layer1_outputs(7240) <= b and not a;
    layer1_outputs(7241) <= not a;
    layer1_outputs(7242) <= 1'b1;
    layer1_outputs(7243) <= not b;
    layer1_outputs(7244) <= b and not a;
    layer1_outputs(7245) <= 1'b1;
    layer1_outputs(7246) <= b and not a;
    layer1_outputs(7247) <= not (a or b);
    layer1_outputs(7248) <= not a or b;
    layer1_outputs(7249) <= a and b;
    layer1_outputs(7250) <= not (a or b);
    layer1_outputs(7251) <= b and not a;
    layer1_outputs(7252) <= not (a and b);
    layer1_outputs(7253) <= a and not b;
    layer1_outputs(7254) <= 1'b0;
    layer1_outputs(7255) <= not b;
    layer1_outputs(7256) <= not b;
    layer1_outputs(7257) <= a;
    layer1_outputs(7258) <= not a;
    layer1_outputs(7259) <= b and not a;
    layer1_outputs(7260) <= not (a and b);
    layer1_outputs(7261) <= a and b;
    layer1_outputs(7262) <= not b or a;
    layer1_outputs(7263) <= a xor b;
    layer1_outputs(7264) <= a and b;
    layer1_outputs(7265) <= b and not a;
    layer1_outputs(7266) <= a xor b;
    layer1_outputs(7267) <= not a;
    layer1_outputs(7268) <= b and not a;
    layer1_outputs(7269) <= 1'b1;
    layer1_outputs(7270) <= not (a or b);
    layer1_outputs(7271) <= not b;
    layer1_outputs(7272) <= 1'b1;
    layer1_outputs(7273) <= 1'b1;
    layer1_outputs(7274) <= a and not b;
    layer1_outputs(7275) <= not (a and b);
    layer1_outputs(7276) <= not (a or b);
    layer1_outputs(7277) <= b;
    layer1_outputs(7278) <= 1'b0;
    layer1_outputs(7279) <= not (a or b);
    layer1_outputs(7280) <= 1'b0;
    layer1_outputs(7281) <= a xor b;
    layer1_outputs(7282) <= not (a xor b);
    layer1_outputs(7283) <= a and not b;
    layer1_outputs(7284) <= a;
    layer1_outputs(7285) <= not a or b;
    layer1_outputs(7286) <= 1'b1;
    layer1_outputs(7287) <= not b;
    layer1_outputs(7288) <= 1'b1;
    layer1_outputs(7289) <= b;
    layer1_outputs(7290) <= not a or b;
    layer1_outputs(7291) <= not a;
    layer1_outputs(7292) <= not a;
    layer1_outputs(7293) <= not b or a;
    layer1_outputs(7294) <= not (a or b);
    layer1_outputs(7295) <= a or b;
    layer1_outputs(7296) <= 1'b0;
    layer1_outputs(7297) <= b;
    layer1_outputs(7298) <= b;
    layer1_outputs(7299) <= 1'b0;
    layer1_outputs(7300) <= not (a and b);
    layer1_outputs(7301) <= a xor b;
    layer1_outputs(7302) <= 1'b1;
    layer1_outputs(7303) <= not b;
    layer1_outputs(7304) <= b;
    layer1_outputs(7305) <= not (a or b);
    layer1_outputs(7306) <= a xor b;
    layer1_outputs(7307) <= 1'b0;
    layer1_outputs(7308) <= not (a and b);
    layer1_outputs(7309) <= b;
    layer1_outputs(7310) <= a or b;
    layer1_outputs(7311) <= not a or b;
    layer1_outputs(7312) <= 1'b1;
    layer1_outputs(7313) <= b;
    layer1_outputs(7314) <= not (a or b);
    layer1_outputs(7315) <= not b;
    layer1_outputs(7316) <= a and not b;
    layer1_outputs(7317) <= a and b;
    layer1_outputs(7318) <= not (a or b);
    layer1_outputs(7319) <= not b or a;
    layer1_outputs(7320) <= not (a and b);
    layer1_outputs(7321) <= not (a and b);
    layer1_outputs(7322) <= not (a and b);
    layer1_outputs(7323) <= a and b;
    layer1_outputs(7324) <= b;
    layer1_outputs(7325) <= 1'b1;
    layer1_outputs(7326) <= a or b;
    layer1_outputs(7327) <= b and not a;
    layer1_outputs(7328) <= not (a or b);
    layer1_outputs(7329) <= a;
    layer1_outputs(7330) <= b;
    layer1_outputs(7331) <= a;
    layer1_outputs(7332) <= b;
    layer1_outputs(7333) <= not a or b;
    layer1_outputs(7334) <= b and not a;
    layer1_outputs(7335) <= not a or b;
    layer1_outputs(7336) <= 1'b1;
    layer1_outputs(7337) <= not (a and b);
    layer1_outputs(7338) <= b and not a;
    layer1_outputs(7339) <= not (a xor b);
    layer1_outputs(7340) <= a or b;
    layer1_outputs(7341) <= a;
    layer1_outputs(7342) <= not (a and b);
    layer1_outputs(7343) <= b and not a;
    layer1_outputs(7344) <= b and not a;
    layer1_outputs(7345) <= a;
    layer1_outputs(7346) <= not a or b;
    layer1_outputs(7347) <= b;
    layer1_outputs(7348) <= b;
    layer1_outputs(7349) <= a or b;
    layer1_outputs(7350) <= not (a and b);
    layer1_outputs(7351) <= not (a and b);
    layer1_outputs(7352) <= not (a or b);
    layer1_outputs(7353) <= not (a or b);
    layer1_outputs(7354) <= b;
    layer1_outputs(7355) <= a and not b;
    layer1_outputs(7356) <= a;
    layer1_outputs(7357) <= not (a and b);
    layer1_outputs(7358) <= b and not a;
    layer1_outputs(7359) <= a;
    layer1_outputs(7360) <= 1'b0;
    layer1_outputs(7361) <= 1'b0;
    layer1_outputs(7362) <= not (a and b);
    layer1_outputs(7363) <= not (a or b);
    layer1_outputs(7364) <= not (a and b);
    layer1_outputs(7365) <= a and b;
    layer1_outputs(7366) <= not b or a;
    layer1_outputs(7367) <= not a;
    layer1_outputs(7368) <= a;
    layer1_outputs(7369) <= a;
    layer1_outputs(7370) <= b and not a;
    layer1_outputs(7371) <= not a;
    layer1_outputs(7372) <= not (a or b);
    layer1_outputs(7373) <= not b;
    layer1_outputs(7374) <= not (a or b);
    layer1_outputs(7375) <= b and not a;
    layer1_outputs(7376) <= not (a or b);
    layer1_outputs(7377) <= 1'b1;
    layer1_outputs(7378) <= 1'b0;
    layer1_outputs(7379) <= a;
    layer1_outputs(7380) <= not b;
    layer1_outputs(7381) <= a and not b;
    layer1_outputs(7382) <= not b or a;
    layer1_outputs(7383) <= 1'b1;
    layer1_outputs(7384) <= not (a or b);
    layer1_outputs(7385) <= a and not b;
    layer1_outputs(7386) <= not b or a;
    layer1_outputs(7387) <= not b or a;
    layer1_outputs(7388) <= not b;
    layer1_outputs(7389) <= a;
    layer1_outputs(7390) <= not b;
    layer1_outputs(7391) <= not a or b;
    layer1_outputs(7392) <= 1'b0;
    layer1_outputs(7393) <= not a or b;
    layer1_outputs(7394) <= not (a or b);
    layer1_outputs(7395) <= not (a or b);
    layer1_outputs(7396) <= not b or a;
    layer1_outputs(7397) <= not a;
    layer1_outputs(7398) <= not a;
    layer1_outputs(7399) <= not (a and b);
    layer1_outputs(7400) <= not (a or b);
    layer1_outputs(7401) <= a;
    layer1_outputs(7402) <= 1'b0;
    layer1_outputs(7403) <= a;
    layer1_outputs(7404) <= a;
    layer1_outputs(7405) <= not b;
    layer1_outputs(7406) <= not (a and b);
    layer1_outputs(7407) <= b and not a;
    layer1_outputs(7408) <= a;
    layer1_outputs(7409) <= not (a or b);
    layer1_outputs(7410) <= not b;
    layer1_outputs(7411) <= b and not a;
    layer1_outputs(7412) <= not b or a;
    layer1_outputs(7413) <= not (a or b);
    layer1_outputs(7414) <= a and b;
    layer1_outputs(7415) <= not (a or b);
    layer1_outputs(7416) <= a or b;
    layer1_outputs(7417) <= not b or a;
    layer1_outputs(7418) <= not b or a;
    layer1_outputs(7419) <= a and not b;
    layer1_outputs(7420) <= a;
    layer1_outputs(7421) <= b and not a;
    layer1_outputs(7422) <= not a;
    layer1_outputs(7423) <= a;
    layer1_outputs(7424) <= not a;
    layer1_outputs(7425) <= not b or a;
    layer1_outputs(7426) <= 1'b0;
    layer1_outputs(7427) <= 1'b0;
    layer1_outputs(7428) <= a xor b;
    layer1_outputs(7429) <= not b;
    layer1_outputs(7430) <= a xor b;
    layer1_outputs(7431) <= 1'b0;
    layer1_outputs(7432) <= a and b;
    layer1_outputs(7433) <= a and b;
    layer1_outputs(7434) <= 1'b1;
    layer1_outputs(7435) <= a and not b;
    layer1_outputs(7436) <= a and not b;
    layer1_outputs(7437) <= a or b;
    layer1_outputs(7438) <= not (a xor b);
    layer1_outputs(7439) <= not a;
    layer1_outputs(7440) <= b;
    layer1_outputs(7441) <= a or b;
    layer1_outputs(7442) <= a xor b;
    layer1_outputs(7443) <= 1'b1;
    layer1_outputs(7444) <= b;
    layer1_outputs(7445) <= a xor b;
    layer1_outputs(7446) <= b and not a;
    layer1_outputs(7447) <= b and not a;
    layer1_outputs(7448) <= 1'b1;
    layer1_outputs(7449) <= not a or b;
    layer1_outputs(7450) <= 1'b1;
    layer1_outputs(7451) <= a and not b;
    layer1_outputs(7452) <= a or b;
    layer1_outputs(7453) <= 1'b1;
    layer1_outputs(7454) <= not b;
    layer1_outputs(7455) <= 1'b0;
    layer1_outputs(7456) <= not b;
    layer1_outputs(7457) <= a xor b;
    layer1_outputs(7458) <= a and not b;
    layer1_outputs(7459) <= not (a or b);
    layer1_outputs(7460) <= a and not b;
    layer1_outputs(7461) <= 1'b1;
    layer1_outputs(7462) <= a and not b;
    layer1_outputs(7463) <= a;
    layer1_outputs(7464) <= not b;
    layer1_outputs(7465) <= b and not a;
    layer1_outputs(7466) <= a xor b;
    layer1_outputs(7467) <= 1'b1;
    layer1_outputs(7468) <= a and not b;
    layer1_outputs(7469) <= not b or a;
    layer1_outputs(7470) <= 1'b0;
    layer1_outputs(7471) <= b;
    layer1_outputs(7472) <= a and b;
    layer1_outputs(7473) <= 1'b1;
    layer1_outputs(7474) <= not (a xor b);
    layer1_outputs(7475) <= a and not b;
    layer1_outputs(7476) <= a;
    layer1_outputs(7477) <= 1'b0;
    layer1_outputs(7478) <= b;
    layer1_outputs(7479) <= a and not b;
    layer1_outputs(7480) <= 1'b0;
    layer1_outputs(7481) <= 1'b1;
    layer1_outputs(7482) <= not a;
    layer1_outputs(7483) <= not b;
    layer1_outputs(7484) <= a and b;
    layer1_outputs(7485) <= not a or b;
    layer1_outputs(7486) <= not b;
    layer1_outputs(7487) <= a and b;
    layer1_outputs(7488) <= not (a xor b);
    layer1_outputs(7489) <= a or b;
    layer1_outputs(7490) <= a or b;
    layer1_outputs(7491) <= 1'b1;
    layer1_outputs(7492) <= not a or b;
    layer1_outputs(7493) <= b and not a;
    layer1_outputs(7494) <= not (a and b);
    layer1_outputs(7495) <= not a or b;
    layer1_outputs(7496) <= not (a and b);
    layer1_outputs(7497) <= not (a or b);
    layer1_outputs(7498) <= not a or b;
    layer1_outputs(7499) <= 1'b0;
    layer1_outputs(7500) <= b;
    layer1_outputs(7501) <= b;
    layer1_outputs(7502) <= a or b;
    layer1_outputs(7503) <= a;
    layer1_outputs(7504) <= not (a xor b);
    layer1_outputs(7505) <= b and not a;
    layer1_outputs(7506) <= not (a and b);
    layer1_outputs(7507) <= not (a or b);
    layer1_outputs(7508) <= a or b;
    layer1_outputs(7509) <= not b;
    layer1_outputs(7510) <= a or b;
    layer1_outputs(7511) <= 1'b0;
    layer1_outputs(7512) <= a or b;
    layer1_outputs(7513) <= 1'b1;
    layer1_outputs(7514) <= a and not b;
    layer1_outputs(7515) <= a or b;
    layer1_outputs(7516) <= not a or b;
    layer1_outputs(7517) <= b and not a;
    layer1_outputs(7518) <= b;
    layer1_outputs(7519) <= a or b;
    layer1_outputs(7520) <= 1'b0;
    layer1_outputs(7521) <= a and b;
    layer1_outputs(7522) <= a and not b;
    layer1_outputs(7523) <= not (a or b);
    layer1_outputs(7524) <= 1'b0;
    layer1_outputs(7525) <= b;
    layer1_outputs(7526) <= 1'b1;
    layer1_outputs(7527) <= b;
    layer1_outputs(7528) <= 1'b1;
    layer1_outputs(7529) <= a and not b;
    layer1_outputs(7530) <= 1'b1;
    layer1_outputs(7531) <= a or b;
    layer1_outputs(7532) <= a or b;
    layer1_outputs(7533) <= not (a and b);
    layer1_outputs(7534) <= not (a xor b);
    layer1_outputs(7535) <= not (a and b);
    layer1_outputs(7536) <= a and b;
    layer1_outputs(7537) <= not a or b;
    layer1_outputs(7538) <= 1'b0;
    layer1_outputs(7539) <= not a;
    layer1_outputs(7540) <= b;
    layer1_outputs(7541) <= not a or b;
    layer1_outputs(7542) <= not (a and b);
    layer1_outputs(7543) <= a;
    layer1_outputs(7544) <= not (a and b);
    layer1_outputs(7545) <= not b or a;
    layer1_outputs(7546) <= not b or a;
    layer1_outputs(7547) <= a and not b;
    layer1_outputs(7548) <= a and not b;
    layer1_outputs(7549) <= 1'b0;
    layer1_outputs(7550) <= not b or a;
    layer1_outputs(7551) <= 1'b1;
    layer1_outputs(7552) <= 1'b1;
    layer1_outputs(7553) <= not b or a;
    layer1_outputs(7554) <= not b;
    layer1_outputs(7555) <= a or b;
    layer1_outputs(7556) <= a and not b;
    layer1_outputs(7557) <= a or b;
    layer1_outputs(7558) <= not a or b;
    layer1_outputs(7559) <= 1'b1;
    layer1_outputs(7560) <= a or b;
    layer1_outputs(7561) <= not (a or b);
    layer1_outputs(7562) <= a or b;
    layer1_outputs(7563) <= a and not b;
    layer1_outputs(7564) <= 1'b0;
    layer1_outputs(7565) <= b;
    layer1_outputs(7566) <= not a or b;
    layer1_outputs(7567) <= a and not b;
    layer1_outputs(7568) <= 1'b0;
    layer1_outputs(7569) <= not a or b;
    layer1_outputs(7570) <= 1'b0;
    layer1_outputs(7571) <= a and b;
    layer1_outputs(7572) <= 1'b1;
    layer1_outputs(7573) <= a or b;
    layer1_outputs(7574) <= not a or b;
    layer1_outputs(7575) <= 1'b0;
    layer1_outputs(7576) <= not (a or b);
    layer1_outputs(7577) <= a and b;
    layer1_outputs(7578) <= not (a xor b);
    layer1_outputs(7579) <= a xor b;
    layer1_outputs(7580) <= not b;
    layer1_outputs(7581) <= b;
    layer1_outputs(7582) <= not b or a;
    layer1_outputs(7583) <= a or b;
    layer1_outputs(7584) <= a;
    layer1_outputs(7585) <= not a;
    layer1_outputs(7586) <= not (a and b);
    layer1_outputs(7587) <= b and not a;
    layer1_outputs(7588) <= a or b;
    layer1_outputs(7589) <= not a or b;
    layer1_outputs(7590) <= not a or b;
    layer1_outputs(7591) <= a;
    layer1_outputs(7592) <= 1'b0;
    layer1_outputs(7593) <= b and not a;
    layer1_outputs(7594) <= 1'b0;
    layer1_outputs(7595) <= 1'b1;
    layer1_outputs(7596) <= not (a and b);
    layer1_outputs(7597) <= a and not b;
    layer1_outputs(7598) <= a and b;
    layer1_outputs(7599) <= 1'b1;
    layer1_outputs(7600) <= 1'b0;
    layer1_outputs(7601) <= 1'b1;
    layer1_outputs(7602) <= not b or a;
    layer1_outputs(7603) <= b and not a;
    layer1_outputs(7604) <= b;
    layer1_outputs(7605) <= 1'b1;
    layer1_outputs(7606) <= not (a or b);
    layer1_outputs(7607) <= a;
    layer1_outputs(7608) <= a or b;
    layer1_outputs(7609) <= not a;
    layer1_outputs(7610) <= a;
    layer1_outputs(7611) <= not (a and b);
    layer1_outputs(7612) <= a and b;
    layer1_outputs(7613) <= a and b;
    layer1_outputs(7614) <= 1'b1;
    layer1_outputs(7615) <= b and not a;
    layer1_outputs(7616) <= not a;
    layer1_outputs(7617) <= not b;
    layer1_outputs(7618) <= not (a and b);
    layer1_outputs(7619) <= a and not b;
    layer1_outputs(7620) <= a;
    layer1_outputs(7621) <= not a or b;
    layer1_outputs(7622) <= 1'b1;
    layer1_outputs(7623) <= a and b;
    layer1_outputs(7624) <= b;
    layer1_outputs(7625) <= not (a xor b);
    layer1_outputs(7626) <= b;
    layer1_outputs(7627) <= 1'b0;
    layer1_outputs(7628) <= not b;
    layer1_outputs(7629) <= not (a or b);
    layer1_outputs(7630) <= b and not a;
    layer1_outputs(7631) <= a or b;
    layer1_outputs(7632) <= not b;
    layer1_outputs(7633) <= 1'b1;
    layer1_outputs(7634) <= 1'b1;
    layer1_outputs(7635) <= a;
    layer1_outputs(7636) <= 1'b1;
    layer1_outputs(7637) <= 1'b1;
    layer1_outputs(7638) <= a;
    layer1_outputs(7639) <= a or b;
    layer1_outputs(7640) <= not (a or b);
    layer1_outputs(7641) <= a and b;
    layer1_outputs(7642) <= 1'b1;
    layer1_outputs(7643) <= b and not a;
    layer1_outputs(7644) <= a and not b;
    layer1_outputs(7645) <= not a;
    layer1_outputs(7646) <= b;
    layer1_outputs(7647) <= not a;
    layer1_outputs(7648) <= b;
    layer1_outputs(7649) <= b;
    layer1_outputs(7650) <= b and not a;
    layer1_outputs(7651) <= a and b;
    layer1_outputs(7652) <= a;
    layer1_outputs(7653) <= not a or b;
    layer1_outputs(7654) <= a xor b;
    layer1_outputs(7655) <= 1'b1;
    layer1_outputs(7656) <= not b or a;
    layer1_outputs(7657) <= 1'b1;
    layer1_outputs(7658) <= not a or b;
    layer1_outputs(7659) <= not (a and b);
    layer1_outputs(7660) <= a and b;
    layer1_outputs(7661) <= b and not a;
    layer1_outputs(7662) <= a and b;
    layer1_outputs(7663) <= 1'b0;
    layer1_outputs(7664) <= a;
    layer1_outputs(7665) <= not (a or b);
    layer1_outputs(7666) <= not b;
    layer1_outputs(7667) <= not (a or b);
    layer1_outputs(7668) <= a or b;
    layer1_outputs(7669) <= 1'b1;
    layer1_outputs(7670) <= not b;
    layer1_outputs(7671) <= not a;
    layer1_outputs(7672) <= not (a and b);
    layer1_outputs(7673) <= a;
    layer1_outputs(7674) <= not a or b;
    layer1_outputs(7675) <= 1'b0;
    layer1_outputs(7676) <= not b or a;
    layer1_outputs(7677) <= b;
    layer1_outputs(7678) <= 1'b1;
    layer1_outputs(7679) <= not b or a;
    layer1_outputs(7680) <= not (a and b);
    layer1_outputs(7681) <= not (a and b);
    layer1_outputs(7682) <= 1'b0;
    layer1_outputs(7683) <= not (a and b);
    layer1_outputs(7684) <= b;
    layer1_outputs(7685) <= not (a xor b);
    layer1_outputs(7686) <= not b or a;
    layer1_outputs(7687) <= 1'b1;
    layer1_outputs(7688) <= 1'b1;
    layer1_outputs(7689) <= 1'b0;
    layer1_outputs(7690) <= 1'b0;
    layer1_outputs(7691) <= a and b;
    layer1_outputs(7692) <= not (a and b);
    layer1_outputs(7693) <= b;
    layer1_outputs(7694) <= not b;
    layer1_outputs(7695) <= a and b;
    layer1_outputs(7696) <= b and not a;
    layer1_outputs(7697) <= a;
    layer1_outputs(7698) <= b;
    layer1_outputs(7699) <= 1'b1;
    layer1_outputs(7700) <= not (a and b);
    layer1_outputs(7701) <= 1'b0;
    layer1_outputs(7702) <= not b or a;
    layer1_outputs(7703) <= a and b;
    layer1_outputs(7704) <= a or b;
    layer1_outputs(7705) <= a and not b;
    layer1_outputs(7706) <= b;
    layer1_outputs(7707) <= b;
    layer1_outputs(7708) <= 1'b1;
    layer1_outputs(7709) <= b and not a;
    layer1_outputs(7710) <= not b;
    layer1_outputs(7711) <= b;
    layer1_outputs(7712) <= a and b;
    layer1_outputs(7713) <= a or b;
    layer1_outputs(7714) <= not a or b;
    layer1_outputs(7715) <= a and not b;
    layer1_outputs(7716) <= not a or b;
    layer1_outputs(7717) <= not (a xor b);
    layer1_outputs(7718) <= b;
    layer1_outputs(7719) <= not a or b;
    layer1_outputs(7720) <= 1'b0;
    layer1_outputs(7721) <= a or b;
    layer1_outputs(7722) <= not b or a;
    layer1_outputs(7723) <= not b;
    layer1_outputs(7724) <= 1'b1;
    layer1_outputs(7725) <= not a;
    layer1_outputs(7726) <= not a or b;
    layer1_outputs(7727) <= not (a or b);
    layer1_outputs(7728) <= not (a and b);
    layer1_outputs(7729) <= not a;
    layer1_outputs(7730) <= not a or b;
    layer1_outputs(7731) <= b and not a;
    layer1_outputs(7732) <= a xor b;
    layer1_outputs(7733) <= b and not a;
    layer1_outputs(7734) <= a;
    layer1_outputs(7735) <= a or b;
    layer1_outputs(7736) <= a xor b;
    layer1_outputs(7737) <= b and not a;
    layer1_outputs(7738) <= 1'b1;
    layer1_outputs(7739) <= not a or b;
    layer1_outputs(7740) <= not (a or b);
    layer1_outputs(7741) <= not (a and b);
    layer1_outputs(7742) <= not a or b;
    layer1_outputs(7743) <= b and not a;
    layer1_outputs(7744) <= a or b;
    layer1_outputs(7745) <= not a;
    layer1_outputs(7746) <= a xor b;
    layer1_outputs(7747) <= a or b;
    layer1_outputs(7748) <= not a;
    layer1_outputs(7749) <= b and not a;
    layer1_outputs(7750) <= b;
    layer1_outputs(7751) <= a and not b;
    layer1_outputs(7752) <= b;
    layer1_outputs(7753) <= 1'b1;
    layer1_outputs(7754) <= a or b;
    layer1_outputs(7755) <= not (a or b);
    layer1_outputs(7756) <= b;
    layer1_outputs(7757) <= a and b;
    layer1_outputs(7758) <= b;
    layer1_outputs(7759) <= 1'b1;
    layer1_outputs(7760) <= not a;
    layer1_outputs(7761) <= 1'b1;
    layer1_outputs(7762) <= 1'b0;
    layer1_outputs(7763) <= not (a and b);
    layer1_outputs(7764) <= 1'b1;
    layer1_outputs(7765) <= not (a and b);
    layer1_outputs(7766) <= b and not a;
    layer1_outputs(7767) <= not (a or b);
    layer1_outputs(7768) <= a and b;
    layer1_outputs(7769) <= a and not b;
    layer1_outputs(7770) <= 1'b1;
    layer1_outputs(7771) <= not a;
    layer1_outputs(7772) <= not b;
    layer1_outputs(7773) <= 1'b0;
    layer1_outputs(7774) <= a or b;
    layer1_outputs(7775) <= not a;
    layer1_outputs(7776) <= a and not b;
    layer1_outputs(7777) <= a or b;
    layer1_outputs(7778) <= 1'b1;
    layer1_outputs(7779) <= not (a or b);
    layer1_outputs(7780) <= not (a xor b);
    layer1_outputs(7781) <= 1'b1;
    layer1_outputs(7782) <= not (a and b);
    layer1_outputs(7783) <= 1'b1;
    layer1_outputs(7784) <= b and not a;
    layer1_outputs(7785) <= 1'b1;
    layer1_outputs(7786) <= 1'b0;
    layer1_outputs(7787) <= a;
    layer1_outputs(7788) <= not b or a;
    layer1_outputs(7789) <= b;
    layer1_outputs(7790) <= not a;
    layer1_outputs(7791) <= 1'b1;
    layer1_outputs(7792) <= not a;
    layer1_outputs(7793) <= a and b;
    layer1_outputs(7794) <= not (a xor b);
    layer1_outputs(7795) <= not (a or b);
    layer1_outputs(7796) <= not a;
    layer1_outputs(7797) <= a and not b;
    layer1_outputs(7798) <= a and not b;
    layer1_outputs(7799) <= a and not b;
    layer1_outputs(7800) <= not b;
    layer1_outputs(7801) <= a and b;
    layer1_outputs(7802) <= a and b;
    layer1_outputs(7803) <= 1'b0;
    layer1_outputs(7804) <= 1'b1;
    layer1_outputs(7805) <= 1'b0;
    layer1_outputs(7806) <= a and b;
    layer1_outputs(7807) <= a or b;
    layer1_outputs(7808) <= 1'b1;
    layer1_outputs(7809) <= not (a and b);
    layer1_outputs(7810) <= 1'b0;
    layer1_outputs(7811) <= b;
    layer1_outputs(7812) <= not (a xor b);
    layer1_outputs(7813) <= b and not a;
    layer1_outputs(7814) <= not (a and b);
    layer1_outputs(7815) <= not (a xor b);
    layer1_outputs(7816) <= not b or a;
    layer1_outputs(7817) <= 1'b0;
    layer1_outputs(7818) <= not a;
    layer1_outputs(7819) <= not b or a;
    layer1_outputs(7820) <= not (a or b);
    layer1_outputs(7821) <= not (a and b);
    layer1_outputs(7822) <= a and b;
    layer1_outputs(7823) <= not b;
    layer1_outputs(7824) <= not a or b;
    layer1_outputs(7825) <= a or b;
    layer1_outputs(7826) <= 1'b1;
    layer1_outputs(7827) <= a xor b;
    layer1_outputs(7828) <= 1'b1;
    layer1_outputs(7829) <= 1'b1;
    layer1_outputs(7830) <= a;
    layer1_outputs(7831) <= b and not a;
    layer1_outputs(7832) <= 1'b0;
    layer1_outputs(7833) <= not (a xor b);
    layer1_outputs(7834) <= not a or b;
    layer1_outputs(7835) <= a;
    layer1_outputs(7836) <= not b or a;
    layer1_outputs(7837) <= not (a and b);
    layer1_outputs(7838) <= 1'b0;
    layer1_outputs(7839) <= a or b;
    layer1_outputs(7840) <= not b or a;
    layer1_outputs(7841) <= a and not b;
    layer1_outputs(7842) <= not b or a;
    layer1_outputs(7843) <= not (a and b);
    layer1_outputs(7844) <= a and b;
    layer1_outputs(7845) <= not b or a;
    layer1_outputs(7846) <= not (a and b);
    layer1_outputs(7847) <= 1'b1;
    layer1_outputs(7848) <= b;
    layer1_outputs(7849) <= not (a or b);
    layer1_outputs(7850) <= not a or b;
    layer1_outputs(7851) <= a;
    layer1_outputs(7852) <= 1'b0;
    layer1_outputs(7853) <= 1'b0;
    layer1_outputs(7854) <= b and not a;
    layer1_outputs(7855) <= not b or a;
    layer1_outputs(7856) <= not a;
    layer1_outputs(7857) <= a;
    layer1_outputs(7858) <= a;
    layer1_outputs(7859) <= not b or a;
    layer1_outputs(7860) <= not b;
    layer1_outputs(7861) <= not b;
    layer1_outputs(7862) <= not (a and b);
    layer1_outputs(7863) <= not b or a;
    layer1_outputs(7864) <= a;
    layer1_outputs(7865) <= not (a xor b);
    layer1_outputs(7866) <= a xor b;
    layer1_outputs(7867) <= b;
    layer1_outputs(7868) <= a or b;
    layer1_outputs(7869) <= 1'b1;
    layer1_outputs(7870) <= not a;
    layer1_outputs(7871) <= not (a and b);
    layer1_outputs(7872) <= b;
    layer1_outputs(7873) <= not (a and b);
    layer1_outputs(7874) <= not (a and b);
    layer1_outputs(7875) <= a xor b;
    layer1_outputs(7876) <= a;
    layer1_outputs(7877) <= b and not a;
    layer1_outputs(7878) <= not b;
    layer1_outputs(7879) <= not (a xor b);
    layer1_outputs(7880) <= 1'b0;
    layer1_outputs(7881) <= a and b;
    layer1_outputs(7882) <= not a;
    layer1_outputs(7883) <= not (a or b);
    layer1_outputs(7884) <= not a;
    layer1_outputs(7885) <= not a;
    layer1_outputs(7886) <= not b;
    layer1_outputs(7887) <= not (a or b);
    layer1_outputs(7888) <= not a;
    layer1_outputs(7889) <= not b;
    layer1_outputs(7890) <= a and b;
    layer1_outputs(7891) <= 1'b0;
    layer1_outputs(7892) <= 1'b0;
    layer1_outputs(7893) <= b;
    layer1_outputs(7894) <= not (a and b);
    layer1_outputs(7895) <= a or b;
    layer1_outputs(7896) <= a and b;
    layer1_outputs(7897) <= a or b;
    layer1_outputs(7898) <= a and b;
    layer1_outputs(7899) <= 1'b1;
    layer1_outputs(7900) <= not b or a;
    layer1_outputs(7901) <= b;
    layer1_outputs(7902) <= b and not a;
    layer1_outputs(7903) <= not (a and b);
    layer1_outputs(7904) <= b;
    layer1_outputs(7905) <= not (a and b);
    layer1_outputs(7906) <= a and b;
    layer1_outputs(7907) <= b and not a;
    layer1_outputs(7908) <= not a;
    layer1_outputs(7909) <= 1'b0;
    layer1_outputs(7910) <= 1'b1;
    layer1_outputs(7911) <= a or b;
    layer1_outputs(7912) <= b and not a;
    layer1_outputs(7913) <= b;
    layer1_outputs(7914) <= not (a and b);
    layer1_outputs(7915) <= not a;
    layer1_outputs(7916) <= a and not b;
    layer1_outputs(7917) <= not a;
    layer1_outputs(7918) <= a or b;
    layer1_outputs(7919) <= not (a and b);
    layer1_outputs(7920) <= a;
    layer1_outputs(7921) <= a and not b;
    layer1_outputs(7922) <= not (a or b);
    layer1_outputs(7923) <= a and not b;
    layer1_outputs(7924) <= a;
    layer1_outputs(7925) <= not a or b;
    layer1_outputs(7926) <= not (a or b);
    layer1_outputs(7927) <= 1'b1;
    layer1_outputs(7928) <= a and not b;
    layer1_outputs(7929) <= b and not a;
    layer1_outputs(7930) <= b and not a;
    layer1_outputs(7931) <= not b;
    layer1_outputs(7932) <= not (a and b);
    layer1_outputs(7933) <= a and b;
    layer1_outputs(7934) <= not (a and b);
    layer1_outputs(7935) <= 1'b1;
    layer1_outputs(7936) <= not (a and b);
    layer1_outputs(7937) <= not b or a;
    layer1_outputs(7938) <= 1'b0;
    layer1_outputs(7939) <= a and b;
    layer1_outputs(7940) <= 1'b1;
    layer1_outputs(7941) <= not (a or b);
    layer1_outputs(7942) <= 1'b1;
    layer1_outputs(7943) <= a xor b;
    layer1_outputs(7944) <= not (a or b);
    layer1_outputs(7945) <= a and not b;
    layer1_outputs(7946) <= 1'b1;
    layer1_outputs(7947) <= not a or b;
    layer1_outputs(7948) <= a or b;
    layer1_outputs(7949) <= a or b;
    layer1_outputs(7950) <= a or b;
    layer1_outputs(7951) <= not a;
    layer1_outputs(7952) <= not b;
    layer1_outputs(7953) <= not b or a;
    layer1_outputs(7954) <= not b or a;
    layer1_outputs(7955) <= not (a or b);
    layer1_outputs(7956) <= b;
    layer1_outputs(7957) <= b and not a;
    layer1_outputs(7958) <= a or b;
    layer1_outputs(7959) <= a xor b;
    layer1_outputs(7960) <= b;
    layer1_outputs(7961) <= not (a or b);
    layer1_outputs(7962) <= not b;
    layer1_outputs(7963) <= not b;
    layer1_outputs(7964) <= 1'b0;
    layer1_outputs(7965) <= not a or b;
    layer1_outputs(7966) <= b;
    layer1_outputs(7967) <= not a or b;
    layer1_outputs(7968) <= not b;
    layer1_outputs(7969) <= a;
    layer1_outputs(7970) <= a;
    layer1_outputs(7971) <= 1'b0;
    layer1_outputs(7972) <= 1'b0;
    layer1_outputs(7973) <= 1'b1;
    layer1_outputs(7974) <= not (a and b);
    layer1_outputs(7975) <= a or b;
    layer1_outputs(7976) <= not b or a;
    layer1_outputs(7977) <= not (a xor b);
    layer1_outputs(7978) <= a and b;
    layer1_outputs(7979) <= a xor b;
    layer1_outputs(7980) <= a;
    layer1_outputs(7981) <= not b or a;
    layer1_outputs(7982) <= not a or b;
    layer1_outputs(7983) <= a and b;
    layer1_outputs(7984) <= 1'b0;
    layer1_outputs(7985) <= not (a or b);
    layer1_outputs(7986) <= b and not a;
    layer1_outputs(7987) <= not (a and b);
    layer1_outputs(7988) <= not a or b;
    layer1_outputs(7989) <= a and not b;
    layer1_outputs(7990) <= a and not b;
    layer1_outputs(7991) <= a;
    layer1_outputs(7992) <= not b or a;
    layer1_outputs(7993) <= b;
    layer1_outputs(7994) <= not b;
    layer1_outputs(7995) <= b;
    layer1_outputs(7996) <= a;
    layer1_outputs(7997) <= not b or a;
    layer1_outputs(7998) <= a or b;
    layer1_outputs(7999) <= not (a or b);
    layer1_outputs(8000) <= 1'b0;
    layer1_outputs(8001) <= a or b;
    layer1_outputs(8002) <= not a;
    layer1_outputs(8003) <= a;
    layer1_outputs(8004) <= 1'b1;
    layer1_outputs(8005) <= not (a or b);
    layer1_outputs(8006) <= b and not a;
    layer1_outputs(8007) <= not b or a;
    layer1_outputs(8008) <= a;
    layer1_outputs(8009) <= b and not a;
    layer1_outputs(8010) <= not b or a;
    layer1_outputs(8011) <= a or b;
    layer1_outputs(8012) <= not (a or b);
    layer1_outputs(8013) <= b and not a;
    layer1_outputs(8014) <= a;
    layer1_outputs(8015) <= a and not b;
    layer1_outputs(8016) <= a and b;
    layer1_outputs(8017) <= 1'b0;
    layer1_outputs(8018) <= not b or a;
    layer1_outputs(8019) <= b;
    layer1_outputs(8020) <= not b or a;
    layer1_outputs(8021) <= not (a and b);
    layer1_outputs(8022) <= 1'b0;
    layer1_outputs(8023) <= a;
    layer1_outputs(8024) <= b;
    layer1_outputs(8025) <= a or b;
    layer1_outputs(8026) <= not b;
    layer1_outputs(8027) <= 1'b0;
    layer1_outputs(8028) <= not a or b;
    layer1_outputs(8029) <= not b;
    layer1_outputs(8030) <= b and not a;
    layer1_outputs(8031) <= not (a or b);
    layer1_outputs(8032) <= a and not b;
    layer1_outputs(8033) <= a;
    layer1_outputs(8034) <= a and not b;
    layer1_outputs(8035) <= not a;
    layer1_outputs(8036) <= a and not b;
    layer1_outputs(8037) <= not (a xor b);
    layer1_outputs(8038) <= b and not a;
    layer1_outputs(8039) <= not a;
    layer1_outputs(8040) <= a or b;
    layer1_outputs(8041) <= b and not a;
    layer1_outputs(8042) <= not a or b;
    layer1_outputs(8043) <= 1'b1;
    layer1_outputs(8044) <= a and b;
    layer1_outputs(8045) <= not (a xor b);
    layer1_outputs(8046) <= a and b;
    layer1_outputs(8047) <= a and not b;
    layer1_outputs(8048) <= not a or b;
    layer1_outputs(8049) <= a and b;
    layer1_outputs(8050) <= b and not a;
    layer1_outputs(8051) <= not a or b;
    layer1_outputs(8052) <= not b or a;
    layer1_outputs(8053) <= a;
    layer1_outputs(8054) <= not (a and b);
    layer1_outputs(8055) <= not b or a;
    layer1_outputs(8056) <= b;
    layer1_outputs(8057) <= not b;
    layer1_outputs(8058) <= not a;
    layer1_outputs(8059) <= not (a xor b);
    layer1_outputs(8060) <= a and not b;
    layer1_outputs(8061) <= 1'b0;
    layer1_outputs(8062) <= 1'b0;
    layer1_outputs(8063) <= 1'b1;
    layer1_outputs(8064) <= a or b;
    layer1_outputs(8065) <= a and b;
    layer1_outputs(8066) <= 1'b1;
    layer1_outputs(8067) <= not (a and b);
    layer1_outputs(8068) <= b and not a;
    layer1_outputs(8069) <= not a or b;
    layer1_outputs(8070) <= not a or b;
    layer1_outputs(8071) <= not b or a;
    layer1_outputs(8072) <= not a;
    layer1_outputs(8073) <= a and b;
    layer1_outputs(8074) <= not b;
    layer1_outputs(8075) <= not (a or b);
    layer1_outputs(8076) <= a;
    layer1_outputs(8077) <= a;
    layer1_outputs(8078) <= b and not a;
    layer1_outputs(8079) <= a xor b;
    layer1_outputs(8080) <= not b or a;
    layer1_outputs(8081) <= a or b;
    layer1_outputs(8082) <= a and not b;
    layer1_outputs(8083) <= not b or a;
    layer1_outputs(8084) <= a or b;
    layer1_outputs(8085) <= a and b;
    layer1_outputs(8086) <= a xor b;
    layer1_outputs(8087) <= 1'b0;
    layer1_outputs(8088) <= a or b;
    layer1_outputs(8089) <= not (a or b);
    layer1_outputs(8090) <= b;
    layer1_outputs(8091) <= b and not a;
    layer1_outputs(8092) <= b and not a;
    layer1_outputs(8093) <= not (a and b);
    layer1_outputs(8094) <= b;
    layer1_outputs(8095) <= a or b;
    layer1_outputs(8096) <= 1'b1;
    layer1_outputs(8097) <= not a;
    layer1_outputs(8098) <= not (a and b);
    layer1_outputs(8099) <= not a or b;
    layer1_outputs(8100) <= a or b;
    layer1_outputs(8101) <= a or b;
    layer1_outputs(8102) <= a and b;
    layer1_outputs(8103) <= 1'b0;
    layer1_outputs(8104) <= not a or b;
    layer1_outputs(8105) <= not b or a;
    layer1_outputs(8106) <= a or b;
    layer1_outputs(8107) <= not (a or b);
    layer1_outputs(8108) <= not b;
    layer1_outputs(8109) <= a or b;
    layer1_outputs(8110) <= a;
    layer1_outputs(8111) <= not (a and b);
    layer1_outputs(8112) <= a and b;
    layer1_outputs(8113) <= not b;
    layer1_outputs(8114) <= not b or a;
    layer1_outputs(8115) <= not (a xor b);
    layer1_outputs(8116) <= not b;
    layer1_outputs(8117) <= not a or b;
    layer1_outputs(8118) <= not a or b;
    layer1_outputs(8119) <= not (a and b);
    layer1_outputs(8120) <= a and b;
    layer1_outputs(8121) <= 1'b0;
    layer1_outputs(8122) <= a;
    layer1_outputs(8123) <= a or b;
    layer1_outputs(8124) <= 1'b1;
    layer1_outputs(8125) <= not (a or b);
    layer1_outputs(8126) <= not a;
    layer1_outputs(8127) <= not a or b;
    layer1_outputs(8128) <= not a;
    layer1_outputs(8129) <= a or b;
    layer1_outputs(8130) <= 1'b0;
    layer1_outputs(8131) <= 1'b0;
    layer1_outputs(8132) <= a and b;
    layer1_outputs(8133) <= not a or b;
    layer1_outputs(8134) <= b;
    layer1_outputs(8135) <= not (a or b);
    layer1_outputs(8136) <= not a;
    layer1_outputs(8137) <= 1'b1;
    layer1_outputs(8138) <= not (a and b);
    layer1_outputs(8139) <= not a;
    layer1_outputs(8140) <= 1'b0;
    layer1_outputs(8141) <= a and not b;
    layer1_outputs(8142) <= 1'b1;
    layer1_outputs(8143) <= not b;
    layer1_outputs(8144) <= not (a or b);
    layer1_outputs(8145) <= not (a or b);
    layer1_outputs(8146) <= 1'b1;
    layer1_outputs(8147) <= not b;
    layer1_outputs(8148) <= a and b;
    layer1_outputs(8149) <= 1'b0;
    layer1_outputs(8150) <= 1'b1;
    layer1_outputs(8151) <= b;
    layer1_outputs(8152) <= a;
    layer1_outputs(8153) <= not a or b;
    layer1_outputs(8154) <= a;
    layer1_outputs(8155) <= a and b;
    layer1_outputs(8156) <= not b;
    layer1_outputs(8157) <= a and not b;
    layer1_outputs(8158) <= b and not a;
    layer1_outputs(8159) <= 1'b0;
    layer1_outputs(8160) <= not b;
    layer1_outputs(8161) <= b;
    layer1_outputs(8162) <= a and b;
    layer1_outputs(8163) <= not b;
    layer1_outputs(8164) <= a and b;
    layer1_outputs(8165) <= not (a and b);
    layer1_outputs(8166) <= not (a xor b);
    layer1_outputs(8167) <= not b or a;
    layer1_outputs(8168) <= not a or b;
    layer1_outputs(8169) <= not (a and b);
    layer1_outputs(8170) <= b and not a;
    layer1_outputs(8171) <= a;
    layer1_outputs(8172) <= not b;
    layer1_outputs(8173) <= not b or a;
    layer1_outputs(8174) <= a;
    layer1_outputs(8175) <= a and b;
    layer1_outputs(8176) <= not b or a;
    layer1_outputs(8177) <= not a or b;
    layer1_outputs(8178) <= a;
    layer1_outputs(8179) <= not a or b;
    layer1_outputs(8180) <= not (a xor b);
    layer1_outputs(8181) <= a and b;
    layer1_outputs(8182) <= not a or b;
    layer1_outputs(8183) <= 1'b0;
    layer1_outputs(8184) <= a and not b;
    layer1_outputs(8185) <= not a or b;
    layer1_outputs(8186) <= not a or b;
    layer1_outputs(8187) <= not a;
    layer1_outputs(8188) <= not (a xor b);
    layer1_outputs(8189) <= not a;
    layer1_outputs(8190) <= 1'b0;
    layer1_outputs(8191) <= not a;
    layer1_outputs(8192) <= not (a or b);
    layer1_outputs(8193) <= not (a or b);
    layer1_outputs(8194) <= 1'b1;
    layer1_outputs(8195) <= not a or b;
    layer1_outputs(8196) <= 1'b1;
    layer1_outputs(8197) <= b and not a;
    layer1_outputs(8198) <= not a;
    layer1_outputs(8199) <= b;
    layer1_outputs(8200) <= not a or b;
    layer1_outputs(8201) <= a and not b;
    layer1_outputs(8202) <= not (a and b);
    layer1_outputs(8203) <= a and b;
    layer1_outputs(8204) <= not a or b;
    layer1_outputs(8205) <= not (a and b);
    layer1_outputs(8206) <= not b;
    layer1_outputs(8207) <= not b;
    layer1_outputs(8208) <= not (a and b);
    layer1_outputs(8209) <= 1'b1;
    layer1_outputs(8210) <= not a;
    layer1_outputs(8211) <= not (a and b);
    layer1_outputs(8212) <= not a;
    layer1_outputs(8213) <= a and not b;
    layer1_outputs(8214) <= a;
    layer1_outputs(8215) <= 1'b0;
    layer1_outputs(8216) <= a xor b;
    layer1_outputs(8217) <= not (a and b);
    layer1_outputs(8218) <= a or b;
    layer1_outputs(8219) <= not b or a;
    layer1_outputs(8220) <= not a or b;
    layer1_outputs(8221) <= b and not a;
    layer1_outputs(8222) <= a and b;
    layer1_outputs(8223) <= b and not a;
    layer1_outputs(8224) <= b and not a;
    layer1_outputs(8225) <= not a or b;
    layer1_outputs(8226) <= a and not b;
    layer1_outputs(8227) <= a or b;
    layer1_outputs(8228) <= not (a or b);
    layer1_outputs(8229) <= b;
    layer1_outputs(8230) <= a and not b;
    layer1_outputs(8231) <= a and not b;
    layer1_outputs(8232) <= 1'b1;
    layer1_outputs(8233) <= 1'b0;
    layer1_outputs(8234) <= a and not b;
    layer1_outputs(8235) <= a and b;
    layer1_outputs(8236) <= a;
    layer1_outputs(8237) <= a and b;
    layer1_outputs(8238) <= not (a xor b);
    layer1_outputs(8239) <= not a;
    layer1_outputs(8240) <= a or b;
    layer1_outputs(8241) <= a or b;
    layer1_outputs(8242) <= not (a or b);
    layer1_outputs(8243) <= a or b;
    layer1_outputs(8244) <= not b;
    layer1_outputs(8245) <= not b;
    layer1_outputs(8246) <= not b;
    layer1_outputs(8247) <= 1'b1;
    layer1_outputs(8248) <= 1'b0;
    layer1_outputs(8249) <= not b;
    layer1_outputs(8250) <= a xor b;
    layer1_outputs(8251) <= b and not a;
    layer1_outputs(8252) <= not a or b;
    layer1_outputs(8253) <= 1'b1;
    layer1_outputs(8254) <= 1'b1;
    layer1_outputs(8255) <= not a;
    layer1_outputs(8256) <= b and not a;
    layer1_outputs(8257) <= a and b;
    layer1_outputs(8258) <= not b or a;
    layer1_outputs(8259) <= not a;
    layer1_outputs(8260) <= a or b;
    layer1_outputs(8261) <= a or b;
    layer1_outputs(8262) <= b;
    layer1_outputs(8263) <= 1'b1;
    layer1_outputs(8264) <= not b;
    layer1_outputs(8265) <= a and b;
    layer1_outputs(8266) <= not (a and b);
    layer1_outputs(8267) <= not (a or b);
    layer1_outputs(8268) <= not (a or b);
    layer1_outputs(8269) <= a and not b;
    layer1_outputs(8270) <= a or b;
    layer1_outputs(8271) <= a and not b;
    layer1_outputs(8272) <= a and b;
    layer1_outputs(8273) <= 1'b0;
    layer1_outputs(8274) <= not (a xor b);
    layer1_outputs(8275) <= not (a or b);
    layer1_outputs(8276) <= 1'b0;
    layer1_outputs(8277) <= not (a and b);
    layer1_outputs(8278) <= b and not a;
    layer1_outputs(8279) <= not a;
    layer1_outputs(8280) <= a and b;
    layer1_outputs(8281) <= not (a and b);
    layer1_outputs(8282) <= 1'b1;
    layer1_outputs(8283) <= a xor b;
    layer1_outputs(8284) <= a and not b;
    layer1_outputs(8285) <= not a;
    layer1_outputs(8286) <= b and not a;
    layer1_outputs(8287) <= 1'b1;
    layer1_outputs(8288) <= a and not b;
    layer1_outputs(8289) <= a or b;
    layer1_outputs(8290) <= 1'b0;
    layer1_outputs(8291) <= a and not b;
    layer1_outputs(8292) <= not a or b;
    layer1_outputs(8293) <= 1'b1;
    layer1_outputs(8294) <= not a or b;
    layer1_outputs(8295) <= not (a xor b);
    layer1_outputs(8296) <= b and not a;
    layer1_outputs(8297) <= not (a and b);
    layer1_outputs(8298) <= a or b;
    layer1_outputs(8299) <= not (a or b);
    layer1_outputs(8300) <= not (a or b);
    layer1_outputs(8301) <= not b;
    layer1_outputs(8302) <= not a or b;
    layer1_outputs(8303) <= not (a xor b);
    layer1_outputs(8304) <= b and not a;
    layer1_outputs(8305) <= 1'b1;
    layer1_outputs(8306) <= 1'b0;
    layer1_outputs(8307) <= 1'b1;
    layer1_outputs(8308) <= not a or b;
    layer1_outputs(8309) <= b;
    layer1_outputs(8310) <= a or b;
    layer1_outputs(8311) <= not a or b;
    layer1_outputs(8312) <= b;
    layer1_outputs(8313) <= not (a or b);
    layer1_outputs(8314) <= a or b;
    layer1_outputs(8315) <= not a or b;
    layer1_outputs(8316) <= not a;
    layer1_outputs(8317) <= not b or a;
    layer1_outputs(8318) <= b and not a;
    layer1_outputs(8319) <= a or b;
    layer1_outputs(8320) <= b;
    layer1_outputs(8321) <= not (a or b);
    layer1_outputs(8322) <= 1'b0;
    layer1_outputs(8323) <= 1'b1;
    layer1_outputs(8324) <= not (a or b);
    layer1_outputs(8325) <= a or b;
    layer1_outputs(8326) <= a or b;
    layer1_outputs(8327) <= a;
    layer1_outputs(8328) <= b;
    layer1_outputs(8329) <= not (a and b);
    layer1_outputs(8330) <= not b or a;
    layer1_outputs(8331) <= a;
    layer1_outputs(8332) <= not b or a;
    layer1_outputs(8333) <= a and b;
    layer1_outputs(8334) <= a and b;
    layer1_outputs(8335) <= not a or b;
    layer1_outputs(8336) <= not (a and b);
    layer1_outputs(8337) <= not a or b;
    layer1_outputs(8338) <= a and not b;
    layer1_outputs(8339) <= a and not b;
    layer1_outputs(8340) <= not b or a;
    layer1_outputs(8341) <= a and b;
    layer1_outputs(8342) <= not a;
    layer1_outputs(8343) <= not (a or b);
    layer1_outputs(8344) <= not b;
    layer1_outputs(8345) <= 1'b0;
    layer1_outputs(8346) <= 1'b0;
    layer1_outputs(8347) <= 1'b0;
    layer1_outputs(8348) <= not (a or b);
    layer1_outputs(8349) <= b;
    layer1_outputs(8350) <= a or b;
    layer1_outputs(8351) <= a and not b;
    layer1_outputs(8352) <= not a;
    layer1_outputs(8353) <= 1'b1;
    layer1_outputs(8354) <= a and b;
    layer1_outputs(8355) <= not a;
    layer1_outputs(8356) <= not (a and b);
    layer1_outputs(8357) <= not (a and b);
    layer1_outputs(8358) <= not b;
    layer1_outputs(8359) <= not a or b;
    layer1_outputs(8360) <= b;
    layer1_outputs(8361) <= not a or b;
    layer1_outputs(8362) <= not (a or b);
    layer1_outputs(8363) <= not b or a;
    layer1_outputs(8364) <= not a or b;
    layer1_outputs(8365) <= b;
    layer1_outputs(8366) <= not (a xor b);
    layer1_outputs(8367) <= a xor b;
    layer1_outputs(8368) <= 1'b0;
    layer1_outputs(8369) <= a;
    layer1_outputs(8370) <= b;
    layer1_outputs(8371) <= not b;
    layer1_outputs(8372) <= 1'b0;
    layer1_outputs(8373) <= not b;
    layer1_outputs(8374) <= 1'b0;
    layer1_outputs(8375) <= not (a or b);
    layer1_outputs(8376) <= not (a and b);
    layer1_outputs(8377) <= 1'b0;
    layer1_outputs(8378) <= 1'b0;
    layer1_outputs(8379) <= not b or a;
    layer1_outputs(8380) <= b and not a;
    layer1_outputs(8381) <= not a or b;
    layer1_outputs(8382) <= 1'b1;
    layer1_outputs(8383) <= a;
    layer1_outputs(8384) <= not a or b;
    layer1_outputs(8385) <= a and not b;
    layer1_outputs(8386) <= not b or a;
    layer1_outputs(8387) <= a and b;
    layer1_outputs(8388) <= 1'b0;
    layer1_outputs(8389) <= not a;
    layer1_outputs(8390) <= a and not b;
    layer1_outputs(8391) <= b and not a;
    layer1_outputs(8392) <= a xor b;
    layer1_outputs(8393) <= 1'b0;
    layer1_outputs(8394) <= not b;
    layer1_outputs(8395) <= b and not a;
    layer1_outputs(8396) <= not a;
    layer1_outputs(8397) <= b;
    layer1_outputs(8398) <= a;
    layer1_outputs(8399) <= a;
    layer1_outputs(8400) <= not (a xor b);
    layer1_outputs(8401) <= b and not a;
    layer1_outputs(8402) <= a and b;
    layer1_outputs(8403) <= 1'b0;
    layer1_outputs(8404) <= 1'b1;
    layer1_outputs(8405) <= not (a and b);
    layer1_outputs(8406) <= a xor b;
    layer1_outputs(8407) <= 1'b1;
    layer1_outputs(8408) <= not b;
    layer1_outputs(8409) <= a or b;
    layer1_outputs(8410) <= not a or b;
    layer1_outputs(8411) <= b and not a;
    layer1_outputs(8412) <= not a;
    layer1_outputs(8413) <= a xor b;
    layer1_outputs(8414) <= 1'b1;
    layer1_outputs(8415) <= a and not b;
    layer1_outputs(8416) <= not a or b;
    layer1_outputs(8417) <= not (a and b);
    layer1_outputs(8418) <= b;
    layer1_outputs(8419) <= not b;
    layer1_outputs(8420) <= not (a or b);
    layer1_outputs(8421) <= not (a or b);
    layer1_outputs(8422) <= not (a and b);
    layer1_outputs(8423) <= not (a or b);
    layer1_outputs(8424) <= 1'b1;
    layer1_outputs(8425) <= 1'b0;
    layer1_outputs(8426) <= not b;
    layer1_outputs(8427) <= a and b;
    layer1_outputs(8428) <= not (a or b);
    layer1_outputs(8429) <= not (a or b);
    layer1_outputs(8430) <= not (a and b);
    layer1_outputs(8431) <= b and not a;
    layer1_outputs(8432) <= not (a and b);
    layer1_outputs(8433) <= a or b;
    layer1_outputs(8434) <= 1'b1;
    layer1_outputs(8435) <= not a;
    layer1_outputs(8436) <= b;
    layer1_outputs(8437) <= b;
    layer1_outputs(8438) <= not b;
    layer1_outputs(8439) <= not a;
    layer1_outputs(8440) <= a or b;
    layer1_outputs(8441) <= not (a xor b);
    layer1_outputs(8442) <= not b or a;
    layer1_outputs(8443) <= a xor b;
    layer1_outputs(8444) <= not (a or b);
    layer1_outputs(8445) <= a and b;
    layer1_outputs(8446) <= a and not b;
    layer1_outputs(8447) <= not a;
    layer1_outputs(8448) <= 1'b0;
    layer1_outputs(8449) <= a;
    layer1_outputs(8450) <= 1'b1;
    layer1_outputs(8451) <= not (a and b);
    layer1_outputs(8452) <= not b or a;
    layer1_outputs(8453) <= a and not b;
    layer1_outputs(8454) <= b and not a;
    layer1_outputs(8455) <= not (a and b);
    layer1_outputs(8456) <= a and not b;
    layer1_outputs(8457) <= a and b;
    layer1_outputs(8458) <= a and b;
    layer1_outputs(8459) <= 1'b0;
    layer1_outputs(8460) <= a or b;
    layer1_outputs(8461) <= not b or a;
    layer1_outputs(8462) <= a and b;
    layer1_outputs(8463) <= not (a and b);
    layer1_outputs(8464) <= a;
    layer1_outputs(8465) <= a and b;
    layer1_outputs(8466) <= not a or b;
    layer1_outputs(8467) <= 1'b0;
    layer1_outputs(8468) <= a and not b;
    layer1_outputs(8469) <= b and not a;
    layer1_outputs(8470) <= a and not b;
    layer1_outputs(8471) <= not (a or b);
    layer1_outputs(8472) <= not b or a;
    layer1_outputs(8473) <= a;
    layer1_outputs(8474) <= b and not a;
    layer1_outputs(8475) <= a and b;
    layer1_outputs(8476) <= not (a and b);
    layer1_outputs(8477) <= a or b;
    layer1_outputs(8478) <= 1'b0;
    layer1_outputs(8479) <= a or b;
    layer1_outputs(8480) <= 1'b0;
    layer1_outputs(8481) <= 1'b1;
    layer1_outputs(8482) <= b and not a;
    layer1_outputs(8483) <= a;
    layer1_outputs(8484) <= a xor b;
    layer1_outputs(8485) <= 1'b0;
    layer1_outputs(8486) <= a and not b;
    layer1_outputs(8487) <= not (a or b);
    layer1_outputs(8488) <= 1'b0;
    layer1_outputs(8489) <= not (a or b);
    layer1_outputs(8490) <= b and not a;
    layer1_outputs(8491) <= not (a and b);
    layer1_outputs(8492) <= 1'b0;
    layer1_outputs(8493) <= a and b;
    layer1_outputs(8494) <= a or b;
    layer1_outputs(8495) <= a xor b;
    layer1_outputs(8496) <= b;
    layer1_outputs(8497) <= b;
    layer1_outputs(8498) <= a and b;
    layer1_outputs(8499) <= a and not b;
    layer1_outputs(8500) <= not (a and b);
    layer1_outputs(8501) <= a and not b;
    layer1_outputs(8502) <= not a;
    layer1_outputs(8503) <= a or b;
    layer1_outputs(8504) <= not (a and b);
    layer1_outputs(8505) <= not b;
    layer1_outputs(8506) <= a or b;
    layer1_outputs(8507) <= b;
    layer1_outputs(8508) <= a and b;
    layer1_outputs(8509) <= a;
    layer1_outputs(8510) <= 1'b0;
    layer1_outputs(8511) <= not b or a;
    layer1_outputs(8512) <= b and not a;
    layer1_outputs(8513) <= not (a or b);
    layer1_outputs(8514) <= a;
    layer1_outputs(8515) <= a xor b;
    layer1_outputs(8516) <= a and not b;
    layer1_outputs(8517) <= not (a and b);
    layer1_outputs(8518) <= a or b;
    layer1_outputs(8519) <= 1'b1;
    layer1_outputs(8520) <= not (a and b);
    layer1_outputs(8521) <= not a or b;
    layer1_outputs(8522) <= a and not b;
    layer1_outputs(8523) <= not a or b;
    layer1_outputs(8524) <= b and not a;
    layer1_outputs(8525) <= not (a xor b);
    layer1_outputs(8526) <= not b;
    layer1_outputs(8527) <= not a or b;
    layer1_outputs(8528) <= not (a and b);
    layer1_outputs(8529) <= b and not a;
    layer1_outputs(8530) <= not b;
    layer1_outputs(8531) <= not a;
    layer1_outputs(8532) <= 1'b1;
    layer1_outputs(8533) <= not (a or b);
    layer1_outputs(8534) <= b and not a;
    layer1_outputs(8535) <= not (a xor b);
    layer1_outputs(8536) <= not (a and b);
    layer1_outputs(8537) <= not a or b;
    layer1_outputs(8538) <= b;
    layer1_outputs(8539) <= a;
    layer1_outputs(8540) <= not b or a;
    layer1_outputs(8541) <= 1'b1;
    layer1_outputs(8542) <= 1'b0;
    layer1_outputs(8543) <= not a or b;
    layer1_outputs(8544) <= not (a or b);
    layer1_outputs(8545) <= 1'b1;
    layer1_outputs(8546) <= not (a and b);
    layer1_outputs(8547) <= a and not b;
    layer1_outputs(8548) <= not (a or b);
    layer1_outputs(8549) <= not (a and b);
    layer1_outputs(8550) <= not a;
    layer1_outputs(8551) <= a and b;
    layer1_outputs(8552) <= b and not a;
    layer1_outputs(8553) <= 1'b1;
    layer1_outputs(8554) <= 1'b1;
    layer1_outputs(8555) <= a;
    layer1_outputs(8556) <= not b or a;
    layer1_outputs(8557) <= a or b;
    layer1_outputs(8558) <= a and b;
    layer1_outputs(8559) <= a or b;
    layer1_outputs(8560) <= a;
    layer1_outputs(8561) <= not (a or b);
    layer1_outputs(8562) <= b;
    layer1_outputs(8563) <= a and not b;
    layer1_outputs(8564) <= a xor b;
    layer1_outputs(8565) <= not b or a;
    layer1_outputs(8566) <= b;
    layer1_outputs(8567) <= b;
    layer1_outputs(8568) <= not (a or b);
    layer1_outputs(8569) <= not (a and b);
    layer1_outputs(8570) <= not (a or b);
    layer1_outputs(8571) <= a and not b;
    layer1_outputs(8572) <= not a;
    layer1_outputs(8573) <= b and not a;
    layer1_outputs(8574) <= not (a and b);
    layer1_outputs(8575) <= not a;
    layer1_outputs(8576) <= 1'b0;
    layer1_outputs(8577) <= b and not a;
    layer1_outputs(8578) <= a and not b;
    layer1_outputs(8579) <= a xor b;
    layer1_outputs(8580) <= b and not a;
    layer1_outputs(8581) <= 1'b1;
    layer1_outputs(8582) <= a or b;
    layer1_outputs(8583) <= 1'b0;
    layer1_outputs(8584) <= 1'b1;
    layer1_outputs(8585) <= 1'b0;
    layer1_outputs(8586) <= a or b;
    layer1_outputs(8587) <= not b or a;
    layer1_outputs(8588) <= not a;
    layer1_outputs(8589) <= a and b;
    layer1_outputs(8590) <= a;
    layer1_outputs(8591) <= a and not b;
    layer1_outputs(8592) <= 1'b0;
    layer1_outputs(8593) <= not b;
    layer1_outputs(8594) <= not (a or b);
    layer1_outputs(8595) <= a or b;
    layer1_outputs(8596) <= b and not a;
    layer1_outputs(8597) <= a and not b;
    layer1_outputs(8598) <= not (a and b);
    layer1_outputs(8599) <= not b;
    layer1_outputs(8600) <= b and not a;
    layer1_outputs(8601) <= a and b;
    layer1_outputs(8602) <= not (a and b);
    layer1_outputs(8603) <= not a or b;
    layer1_outputs(8604) <= a;
    layer1_outputs(8605) <= 1'b1;
    layer1_outputs(8606) <= a;
    layer1_outputs(8607) <= not (a and b);
    layer1_outputs(8608) <= a or b;
    layer1_outputs(8609) <= 1'b1;
    layer1_outputs(8610) <= not b;
    layer1_outputs(8611) <= not b;
    layer1_outputs(8612) <= b;
    layer1_outputs(8613) <= not (a xor b);
    layer1_outputs(8614) <= not (a or b);
    layer1_outputs(8615) <= 1'b1;
    layer1_outputs(8616) <= not a or b;
    layer1_outputs(8617) <= a and not b;
    layer1_outputs(8618) <= not a;
    layer1_outputs(8619) <= 1'b1;
    layer1_outputs(8620) <= 1'b1;
    layer1_outputs(8621) <= 1'b0;
    layer1_outputs(8622) <= b and not a;
    layer1_outputs(8623) <= not b or a;
    layer1_outputs(8624) <= not b or a;
    layer1_outputs(8625) <= a and b;
    layer1_outputs(8626) <= a and not b;
    layer1_outputs(8627) <= 1'b0;
    layer1_outputs(8628) <= a and b;
    layer1_outputs(8629) <= b;
    layer1_outputs(8630) <= not b or a;
    layer1_outputs(8631) <= not (a and b);
    layer1_outputs(8632) <= b and not a;
    layer1_outputs(8633) <= a and not b;
    layer1_outputs(8634) <= a and b;
    layer1_outputs(8635) <= a and b;
    layer1_outputs(8636) <= not a;
    layer1_outputs(8637) <= a;
    layer1_outputs(8638) <= not (a or b);
    layer1_outputs(8639) <= a or b;
    layer1_outputs(8640) <= 1'b0;
    layer1_outputs(8641) <= 1'b1;
    layer1_outputs(8642) <= a or b;
    layer1_outputs(8643) <= a or b;
    layer1_outputs(8644) <= a xor b;
    layer1_outputs(8645) <= not (a or b);
    layer1_outputs(8646) <= b and not a;
    layer1_outputs(8647) <= not (a or b);
    layer1_outputs(8648) <= a;
    layer1_outputs(8649) <= not a or b;
    layer1_outputs(8650) <= not (a xor b);
    layer1_outputs(8651) <= 1'b0;
    layer1_outputs(8652) <= not a or b;
    layer1_outputs(8653) <= not b or a;
    layer1_outputs(8654) <= not (a or b);
    layer1_outputs(8655) <= not a or b;
    layer1_outputs(8656) <= 1'b0;
    layer1_outputs(8657) <= b;
    layer1_outputs(8658) <= 1'b0;
    layer1_outputs(8659) <= a or b;
    layer1_outputs(8660) <= not a or b;
    layer1_outputs(8661) <= not (a and b);
    layer1_outputs(8662) <= not b or a;
    layer1_outputs(8663) <= not (a or b);
    layer1_outputs(8664) <= not b;
    layer1_outputs(8665) <= 1'b0;
    layer1_outputs(8666) <= 1'b0;
    layer1_outputs(8667) <= a and not b;
    layer1_outputs(8668) <= 1'b0;
    layer1_outputs(8669) <= 1'b0;
    layer1_outputs(8670) <= 1'b0;
    layer1_outputs(8671) <= b and not a;
    layer1_outputs(8672) <= 1'b0;
    layer1_outputs(8673) <= 1'b1;
    layer1_outputs(8674) <= not (a and b);
    layer1_outputs(8675) <= a or b;
    layer1_outputs(8676) <= 1'b0;
    layer1_outputs(8677) <= a or b;
    layer1_outputs(8678) <= a and b;
    layer1_outputs(8679) <= a or b;
    layer1_outputs(8680) <= 1'b1;
    layer1_outputs(8681) <= not a or b;
    layer1_outputs(8682) <= 1'b1;
    layer1_outputs(8683) <= not b or a;
    layer1_outputs(8684) <= b;
    layer1_outputs(8685) <= a;
    layer1_outputs(8686) <= not a or b;
    layer1_outputs(8687) <= a xor b;
    layer1_outputs(8688) <= not a;
    layer1_outputs(8689) <= b and not a;
    layer1_outputs(8690) <= b;
    layer1_outputs(8691) <= a;
    layer1_outputs(8692) <= not (a and b);
    layer1_outputs(8693) <= a and not b;
    layer1_outputs(8694) <= not (a or b);
    layer1_outputs(8695) <= 1'b0;
    layer1_outputs(8696) <= 1'b0;
    layer1_outputs(8697) <= not b;
    layer1_outputs(8698) <= a and b;
    layer1_outputs(8699) <= a and not b;
    layer1_outputs(8700) <= b and not a;
    layer1_outputs(8701) <= a xor b;
    layer1_outputs(8702) <= not (a or b);
    layer1_outputs(8703) <= a and not b;
    layer1_outputs(8704) <= b and not a;
    layer1_outputs(8705) <= a;
    layer1_outputs(8706) <= not b;
    layer1_outputs(8707) <= not (a or b);
    layer1_outputs(8708) <= not b or a;
    layer1_outputs(8709) <= not b;
    layer1_outputs(8710) <= not b;
    layer1_outputs(8711) <= not (a xor b);
    layer1_outputs(8712) <= not b;
    layer1_outputs(8713) <= a and not b;
    layer1_outputs(8714) <= b;
    layer1_outputs(8715) <= 1'b1;
    layer1_outputs(8716) <= 1'b1;
    layer1_outputs(8717) <= b and not a;
    layer1_outputs(8718) <= a or b;
    layer1_outputs(8719) <= not (a xor b);
    layer1_outputs(8720) <= b;
    layer1_outputs(8721) <= a and not b;
    layer1_outputs(8722) <= not a or b;
    layer1_outputs(8723) <= not b;
    layer1_outputs(8724) <= 1'b0;
    layer1_outputs(8725) <= not (a or b);
    layer1_outputs(8726) <= not b;
    layer1_outputs(8727) <= not (a and b);
    layer1_outputs(8728) <= 1'b1;
    layer1_outputs(8729) <= a and b;
    layer1_outputs(8730) <= a xor b;
    layer1_outputs(8731) <= a and b;
    layer1_outputs(8732) <= not b;
    layer1_outputs(8733) <= 1'b1;
    layer1_outputs(8734) <= a;
    layer1_outputs(8735) <= not a;
    layer1_outputs(8736) <= 1'b1;
    layer1_outputs(8737) <= b;
    layer1_outputs(8738) <= not (a and b);
    layer1_outputs(8739) <= not (a and b);
    layer1_outputs(8740) <= not b;
    layer1_outputs(8741) <= b and not a;
    layer1_outputs(8742) <= not a;
    layer1_outputs(8743) <= 1'b0;
    layer1_outputs(8744) <= a or b;
    layer1_outputs(8745) <= not b or a;
    layer1_outputs(8746) <= a xor b;
    layer1_outputs(8747) <= 1'b0;
    layer1_outputs(8748) <= not (a xor b);
    layer1_outputs(8749) <= not a or b;
    layer1_outputs(8750) <= a;
    layer1_outputs(8751) <= not b or a;
    layer1_outputs(8752) <= 1'b0;
    layer1_outputs(8753) <= not (a or b);
    layer1_outputs(8754) <= not (a and b);
    layer1_outputs(8755) <= a or b;
    layer1_outputs(8756) <= not a;
    layer1_outputs(8757) <= not b;
    layer1_outputs(8758) <= a;
    layer1_outputs(8759) <= a and not b;
    layer1_outputs(8760) <= not b;
    layer1_outputs(8761) <= a or b;
    layer1_outputs(8762) <= not (a and b);
    layer1_outputs(8763) <= a;
    layer1_outputs(8764) <= 1'b0;
    layer1_outputs(8765) <= 1'b0;
    layer1_outputs(8766) <= 1'b1;
    layer1_outputs(8767) <= 1'b1;
    layer1_outputs(8768) <= 1'b0;
    layer1_outputs(8769) <= a;
    layer1_outputs(8770) <= not (a xor b);
    layer1_outputs(8771) <= a or b;
    layer1_outputs(8772) <= 1'b0;
    layer1_outputs(8773) <= a xor b;
    layer1_outputs(8774) <= not b;
    layer1_outputs(8775) <= b and not a;
    layer1_outputs(8776) <= not (a or b);
    layer1_outputs(8777) <= not a or b;
    layer1_outputs(8778) <= a and b;
    layer1_outputs(8779) <= b and not a;
    layer1_outputs(8780) <= a and b;
    layer1_outputs(8781) <= not a;
    layer1_outputs(8782) <= not b or a;
    layer1_outputs(8783) <= not b;
    layer1_outputs(8784) <= not b;
    layer1_outputs(8785) <= not (a or b);
    layer1_outputs(8786) <= a and b;
    layer1_outputs(8787) <= b and not a;
    layer1_outputs(8788) <= a or b;
    layer1_outputs(8789) <= not a or b;
    layer1_outputs(8790) <= 1'b0;
    layer1_outputs(8791) <= not b or a;
    layer1_outputs(8792) <= a;
    layer1_outputs(8793) <= a and not b;
    layer1_outputs(8794) <= a or b;
    layer1_outputs(8795) <= b and not a;
    layer1_outputs(8796) <= not b or a;
    layer1_outputs(8797) <= 1'b0;
    layer1_outputs(8798) <= a or b;
    layer1_outputs(8799) <= a or b;
    layer1_outputs(8800) <= not b;
    layer1_outputs(8801) <= a and b;
    layer1_outputs(8802) <= a;
    layer1_outputs(8803) <= a xor b;
    layer1_outputs(8804) <= not a;
    layer1_outputs(8805) <= a and not b;
    layer1_outputs(8806) <= not (a and b);
    layer1_outputs(8807) <= a and b;
    layer1_outputs(8808) <= not a;
    layer1_outputs(8809) <= a;
    layer1_outputs(8810) <= not b or a;
    layer1_outputs(8811) <= b and not a;
    layer1_outputs(8812) <= not (a xor b);
    layer1_outputs(8813) <= not (a and b);
    layer1_outputs(8814) <= 1'b1;
    layer1_outputs(8815) <= a and b;
    layer1_outputs(8816) <= not b or a;
    layer1_outputs(8817) <= b;
    layer1_outputs(8818) <= not b;
    layer1_outputs(8819) <= a and b;
    layer1_outputs(8820) <= 1'b0;
    layer1_outputs(8821) <= not (a or b);
    layer1_outputs(8822) <= b and not a;
    layer1_outputs(8823) <= b and not a;
    layer1_outputs(8824) <= not (a and b);
    layer1_outputs(8825) <= a or b;
    layer1_outputs(8826) <= a and not b;
    layer1_outputs(8827) <= b and not a;
    layer1_outputs(8828) <= not a;
    layer1_outputs(8829) <= b and not a;
    layer1_outputs(8830) <= a or b;
    layer1_outputs(8831) <= not a;
    layer1_outputs(8832) <= 1'b0;
    layer1_outputs(8833) <= not (a and b);
    layer1_outputs(8834) <= a and not b;
    layer1_outputs(8835) <= not a or b;
    layer1_outputs(8836) <= a and not b;
    layer1_outputs(8837) <= a and b;
    layer1_outputs(8838) <= not b or a;
    layer1_outputs(8839) <= not a or b;
    layer1_outputs(8840) <= not b;
    layer1_outputs(8841) <= not b or a;
    layer1_outputs(8842) <= not b;
    layer1_outputs(8843) <= b;
    layer1_outputs(8844) <= 1'b1;
    layer1_outputs(8845) <= not a;
    layer1_outputs(8846) <= a and b;
    layer1_outputs(8847) <= a or b;
    layer1_outputs(8848) <= b;
    layer1_outputs(8849) <= not (a and b);
    layer1_outputs(8850) <= not (a or b);
    layer1_outputs(8851) <= a and not b;
    layer1_outputs(8852) <= 1'b0;
    layer1_outputs(8853) <= a or b;
    layer1_outputs(8854) <= not a;
    layer1_outputs(8855) <= b;
    layer1_outputs(8856) <= a or b;
    layer1_outputs(8857) <= a or b;
    layer1_outputs(8858) <= b and not a;
    layer1_outputs(8859) <= not (a and b);
    layer1_outputs(8860) <= not a;
    layer1_outputs(8861) <= 1'b0;
    layer1_outputs(8862) <= a and not b;
    layer1_outputs(8863) <= a and b;
    layer1_outputs(8864) <= 1'b1;
    layer1_outputs(8865) <= b;
    layer1_outputs(8866) <= not b;
    layer1_outputs(8867) <= not b or a;
    layer1_outputs(8868) <= not (a and b);
    layer1_outputs(8869) <= not (a and b);
    layer1_outputs(8870) <= a and not b;
    layer1_outputs(8871) <= not (a and b);
    layer1_outputs(8872) <= 1'b0;
    layer1_outputs(8873) <= not a or b;
    layer1_outputs(8874) <= b;
    layer1_outputs(8875) <= 1'b0;
    layer1_outputs(8876) <= b;
    layer1_outputs(8877) <= not (a xor b);
    layer1_outputs(8878) <= a;
    layer1_outputs(8879) <= b and not a;
    layer1_outputs(8880) <= not (a and b);
    layer1_outputs(8881) <= not a;
    layer1_outputs(8882) <= not a or b;
    layer1_outputs(8883) <= a xor b;
    layer1_outputs(8884) <= not (a and b);
    layer1_outputs(8885) <= not (a and b);
    layer1_outputs(8886) <= not b;
    layer1_outputs(8887) <= not (a and b);
    layer1_outputs(8888) <= a or b;
    layer1_outputs(8889) <= b and not a;
    layer1_outputs(8890) <= b;
    layer1_outputs(8891) <= a;
    layer1_outputs(8892) <= a and not b;
    layer1_outputs(8893) <= b and not a;
    layer1_outputs(8894) <= a and not b;
    layer1_outputs(8895) <= not (a and b);
    layer1_outputs(8896) <= a and not b;
    layer1_outputs(8897) <= not (a and b);
    layer1_outputs(8898) <= a;
    layer1_outputs(8899) <= 1'b1;
    layer1_outputs(8900) <= b and not a;
    layer1_outputs(8901) <= not (a or b);
    layer1_outputs(8902) <= b;
    layer1_outputs(8903) <= a;
    layer1_outputs(8904) <= not a;
    layer1_outputs(8905) <= not (a and b);
    layer1_outputs(8906) <= b and not a;
    layer1_outputs(8907) <= b and not a;
    layer1_outputs(8908) <= not b or a;
    layer1_outputs(8909) <= b and not a;
    layer1_outputs(8910) <= not (a or b);
    layer1_outputs(8911) <= a and not b;
    layer1_outputs(8912) <= not (a or b);
    layer1_outputs(8913) <= 1'b1;
    layer1_outputs(8914) <= not a;
    layer1_outputs(8915) <= b;
    layer1_outputs(8916) <= 1'b0;
    layer1_outputs(8917) <= not (a and b);
    layer1_outputs(8918) <= not b or a;
    layer1_outputs(8919) <= a;
    layer1_outputs(8920) <= not b or a;
    layer1_outputs(8921) <= not a;
    layer1_outputs(8922) <= not a;
    layer1_outputs(8923) <= b and not a;
    layer1_outputs(8924) <= not a;
    layer1_outputs(8925) <= b;
    layer1_outputs(8926) <= b and not a;
    layer1_outputs(8927) <= b and not a;
    layer1_outputs(8928) <= not b or a;
    layer1_outputs(8929) <= not (a and b);
    layer1_outputs(8930) <= not a or b;
    layer1_outputs(8931) <= not (a xor b);
    layer1_outputs(8932) <= 1'b0;
    layer1_outputs(8933) <= 1'b0;
    layer1_outputs(8934) <= 1'b1;
    layer1_outputs(8935) <= not a;
    layer1_outputs(8936) <= not b or a;
    layer1_outputs(8937) <= a and not b;
    layer1_outputs(8938) <= not b or a;
    layer1_outputs(8939) <= 1'b0;
    layer1_outputs(8940) <= 1'b1;
    layer1_outputs(8941) <= a;
    layer1_outputs(8942) <= not (a or b);
    layer1_outputs(8943) <= not b;
    layer1_outputs(8944) <= a and not b;
    layer1_outputs(8945) <= a;
    layer1_outputs(8946) <= not b;
    layer1_outputs(8947) <= a and not b;
    layer1_outputs(8948) <= a and not b;
    layer1_outputs(8949) <= b and not a;
    layer1_outputs(8950) <= a or b;
    layer1_outputs(8951) <= a and b;
    layer1_outputs(8952) <= 1'b1;
    layer1_outputs(8953) <= a or b;
    layer1_outputs(8954) <= 1'b0;
    layer1_outputs(8955) <= not a;
    layer1_outputs(8956) <= not b or a;
    layer1_outputs(8957) <= a;
    layer1_outputs(8958) <= not (a xor b);
    layer1_outputs(8959) <= 1'b1;
    layer1_outputs(8960) <= b and not a;
    layer1_outputs(8961) <= not b;
    layer1_outputs(8962) <= not b;
    layer1_outputs(8963) <= a;
    layer1_outputs(8964) <= 1'b0;
    layer1_outputs(8965) <= a and b;
    layer1_outputs(8966) <= not a or b;
    layer1_outputs(8967) <= 1'b1;
    layer1_outputs(8968) <= b;
    layer1_outputs(8969) <= 1'b0;
    layer1_outputs(8970) <= not a;
    layer1_outputs(8971) <= not b or a;
    layer1_outputs(8972) <= not b or a;
    layer1_outputs(8973) <= b;
    layer1_outputs(8974) <= not (a or b);
    layer1_outputs(8975) <= 1'b0;
    layer1_outputs(8976) <= not (a or b);
    layer1_outputs(8977) <= 1'b0;
    layer1_outputs(8978) <= not a or b;
    layer1_outputs(8979) <= not (a and b);
    layer1_outputs(8980) <= b;
    layer1_outputs(8981) <= not b;
    layer1_outputs(8982) <= b and not a;
    layer1_outputs(8983) <= not a;
    layer1_outputs(8984) <= 1'b1;
    layer1_outputs(8985) <= not (a and b);
    layer1_outputs(8986) <= a and not b;
    layer1_outputs(8987) <= a or b;
    layer1_outputs(8988) <= not b or a;
    layer1_outputs(8989) <= 1'b1;
    layer1_outputs(8990) <= 1'b1;
    layer1_outputs(8991) <= not (a xor b);
    layer1_outputs(8992) <= a or b;
    layer1_outputs(8993) <= 1'b0;
    layer1_outputs(8994) <= 1'b1;
    layer1_outputs(8995) <= a;
    layer1_outputs(8996) <= a or b;
    layer1_outputs(8997) <= a and b;
    layer1_outputs(8998) <= a;
    layer1_outputs(8999) <= not (a or b);
    layer1_outputs(9000) <= not (a and b);
    layer1_outputs(9001) <= not b or a;
    layer1_outputs(9002) <= not (a xor b);
    layer1_outputs(9003) <= not a;
    layer1_outputs(9004) <= b;
    layer1_outputs(9005) <= a or b;
    layer1_outputs(9006) <= 1'b1;
    layer1_outputs(9007) <= not (a and b);
    layer1_outputs(9008) <= b and not a;
    layer1_outputs(9009) <= not b;
    layer1_outputs(9010) <= not a or b;
    layer1_outputs(9011) <= not (a xor b);
    layer1_outputs(9012) <= b;
    layer1_outputs(9013) <= b and not a;
    layer1_outputs(9014) <= 1'b1;
    layer1_outputs(9015) <= a or b;
    layer1_outputs(9016) <= not b;
    layer1_outputs(9017) <= not (a and b);
    layer1_outputs(9018) <= a;
    layer1_outputs(9019) <= b and not a;
    layer1_outputs(9020) <= not b or a;
    layer1_outputs(9021) <= b and not a;
    layer1_outputs(9022) <= not (a xor b);
    layer1_outputs(9023) <= 1'b0;
    layer1_outputs(9024) <= a and b;
    layer1_outputs(9025) <= 1'b0;
    layer1_outputs(9026) <= 1'b0;
    layer1_outputs(9027) <= not (a or b);
    layer1_outputs(9028) <= b;
    layer1_outputs(9029) <= not b or a;
    layer1_outputs(9030) <= a and not b;
    layer1_outputs(9031) <= not b;
    layer1_outputs(9032) <= not (a and b);
    layer1_outputs(9033) <= not b;
    layer1_outputs(9034) <= a;
    layer1_outputs(9035) <= not a;
    layer1_outputs(9036) <= a;
    layer1_outputs(9037) <= not a;
    layer1_outputs(9038) <= not (a xor b);
    layer1_outputs(9039) <= b;
    layer1_outputs(9040) <= not a;
    layer1_outputs(9041) <= 1'b0;
    layer1_outputs(9042) <= a;
    layer1_outputs(9043) <= 1'b0;
    layer1_outputs(9044) <= not b;
    layer1_outputs(9045) <= not b;
    layer1_outputs(9046) <= not b or a;
    layer1_outputs(9047) <= not (a or b);
    layer1_outputs(9048) <= not a or b;
    layer1_outputs(9049) <= a and not b;
    layer1_outputs(9050) <= a or b;
    layer1_outputs(9051) <= not b or a;
    layer1_outputs(9052) <= 1'b1;
    layer1_outputs(9053) <= not a;
    layer1_outputs(9054) <= not b or a;
    layer1_outputs(9055) <= not (a or b);
    layer1_outputs(9056) <= not (a and b);
    layer1_outputs(9057) <= not (a xor b);
    layer1_outputs(9058) <= a and b;
    layer1_outputs(9059) <= a and b;
    layer1_outputs(9060) <= not a;
    layer1_outputs(9061) <= 1'b1;
    layer1_outputs(9062) <= not a;
    layer1_outputs(9063) <= a and b;
    layer1_outputs(9064) <= a and not b;
    layer1_outputs(9065) <= b and not a;
    layer1_outputs(9066) <= a xor b;
    layer1_outputs(9067) <= a;
    layer1_outputs(9068) <= b;
    layer1_outputs(9069) <= not b;
    layer1_outputs(9070) <= a and b;
    layer1_outputs(9071) <= b;
    layer1_outputs(9072) <= not b or a;
    layer1_outputs(9073) <= not a;
    layer1_outputs(9074) <= not b or a;
    layer1_outputs(9075) <= not b or a;
    layer1_outputs(9076) <= not b or a;
    layer1_outputs(9077) <= 1'b1;
    layer1_outputs(9078) <= not a;
    layer1_outputs(9079) <= 1'b1;
    layer1_outputs(9080) <= b and not a;
    layer1_outputs(9081) <= b;
    layer1_outputs(9082) <= 1'b1;
    layer1_outputs(9083) <= 1'b1;
    layer1_outputs(9084) <= not b or a;
    layer1_outputs(9085) <= not a;
    layer1_outputs(9086) <= b;
    layer1_outputs(9087) <= not (a and b);
    layer1_outputs(9088) <= a xor b;
    layer1_outputs(9089) <= 1'b1;
    layer1_outputs(9090) <= a xor b;
    layer1_outputs(9091) <= 1'b0;
    layer1_outputs(9092) <= 1'b0;
    layer1_outputs(9093) <= a and not b;
    layer1_outputs(9094) <= b and not a;
    layer1_outputs(9095) <= b and not a;
    layer1_outputs(9096) <= 1'b1;
    layer1_outputs(9097) <= a and not b;
    layer1_outputs(9098) <= a;
    layer1_outputs(9099) <= not a or b;
    layer1_outputs(9100) <= a and b;
    layer1_outputs(9101) <= not b;
    layer1_outputs(9102) <= a or b;
    layer1_outputs(9103) <= b and not a;
    layer1_outputs(9104) <= 1'b0;
    layer1_outputs(9105) <= not a or b;
    layer1_outputs(9106) <= a or b;
    layer1_outputs(9107) <= not b;
    layer1_outputs(9108) <= not (a or b);
    layer1_outputs(9109) <= a;
    layer1_outputs(9110) <= a xor b;
    layer1_outputs(9111) <= a xor b;
    layer1_outputs(9112) <= not (a and b);
    layer1_outputs(9113) <= not a;
    layer1_outputs(9114) <= not (a xor b);
    layer1_outputs(9115) <= 1'b1;
    layer1_outputs(9116) <= a;
    layer1_outputs(9117) <= b;
    layer1_outputs(9118) <= not b;
    layer1_outputs(9119) <= a;
    layer1_outputs(9120) <= not b or a;
    layer1_outputs(9121) <= not b or a;
    layer1_outputs(9122) <= not (a or b);
    layer1_outputs(9123) <= 1'b0;
    layer1_outputs(9124) <= a xor b;
    layer1_outputs(9125) <= b and not a;
    layer1_outputs(9126) <= not a or b;
    layer1_outputs(9127) <= b and not a;
    layer1_outputs(9128) <= b;
    layer1_outputs(9129) <= a or b;
    layer1_outputs(9130) <= b and not a;
    layer1_outputs(9131) <= not a;
    layer1_outputs(9132) <= a and not b;
    layer1_outputs(9133) <= b;
    layer1_outputs(9134) <= a and b;
    layer1_outputs(9135) <= a and b;
    layer1_outputs(9136) <= b and not a;
    layer1_outputs(9137) <= 1'b0;
    layer1_outputs(9138) <= b;
    layer1_outputs(9139) <= not b;
    layer1_outputs(9140) <= not (a or b);
    layer1_outputs(9141) <= not b or a;
    layer1_outputs(9142) <= not b;
    layer1_outputs(9143) <= 1'b1;
    layer1_outputs(9144) <= a or b;
    layer1_outputs(9145) <= 1'b1;
    layer1_outputs(9146) <= 1'b1;
    layer1_outputs(9147) <= not (a xor b);
    layer1_outputs(9148) <= a or b;
    layer1_outputs(9149) <= a or b;
    layer1_outputs(9150) <= a and b;
    layer1_outputs(9151) <= a and b;
    layer1_outputs(9152) <= a;
    layer1_outputs(9153) <= not a or b;
    layer1_outputs(9154) <= not (a xor b);
    layer1_outputs(9155) <= not (a and b);
    layer1_outputs(9156) <= a and not b;
    layer1_outputs(9157) <= a and b;
    layer1_outputs(9158) <= not a;
    layer1_outputs(9159) <= a and b;
    layer1_outputs(9160) <= not b;
    layer1_outputs(9161) <= a or b;
    layer1_outputs(9162) <= not (a or b);
    layer1_outputs(9163) <= not a or b;
    layer1_outputs(9164) <= a and not b;
    layer1_outputs(9165) <= not b or a;
    layer1_outputs(9166) <= a and not b;
    layer1_outputs(9167) <= not b;
    layer1_outputs(9168) <= not a;
    layer1_outputs(9169) <= a and not b;
    layer1_outputs(9170) <= a;
    layer1_outputs(9171) <= b;
    layer1_outputs(9172) <= not a or b;
    layer1_outputs(9173) <= a;
    layer1_outputs(9174) <= not (a and b);
    layer1_outputs(9175) <= a and b;
    layer1_outputs(9176) <= not (a xor b);
    layer1_outputs(9177) <= not b or a;
    layer1_outputs(9178) <= not (a or b);
    layer1_outputs(9179) <= not a;
    layer1_outputs(9180) <= 1'b0;
    layer1_outputs(9181) <= not (a and b);
    layer1_outputs(9182) <= not (a or b);
    layer1_outputs(9183) <= a or b;
    layer1_outputs(9184) <= 1'b1;
    layer1_outputs(9185) <= not a or b;
    layer1_outputs(9186) <= not (a and b);
    layer1_outputs(9187) <= not (a and b);
    layer1_outputs(9188) <= 1'b0;
    layer1_outputs(9189) <= a and b;
    layer1_outputs(9190) <= a and b;
    layer1_outputs(9191) <= a;
    layer1_outputs(9192) <= not b;
    layer1_outputs(9193) <= a or b;
    layer1_outputs(9194) <= 1'b0;
    layer1_outputs(9195) <= a or b;
    layer1_outputs(9196) <= not a or b;
    layer1_outputs(9197) <= 1'b1;
    layer1_outputs(9198) <= 1'b1;
    layer1_outputs(9199) <= 1'b1;
    layer1_outputs(9200) <= not (a and b);
    layer1_outputs(9201) <= not b or a;
    layer1_outputs(9202) <= not (a xor b);
    layer1_outputs(9203) <= not b or a;
    layer1_outputs(9204) <= not b;
    layer1_outputs(9205) <= a;
    layer1_outputs(9206) <= a and not b;
    layer1_outputs(9207) <= not a or b;
    layer1_outputs(9208) <= 1'b1;
    layer1_outputs(9209) <= not b;
    layer1_outputs(9210) <= not (a and b);
    layer1_outputs(9211) <= not b;
    layer1_outputs(9212) <= a and not b;
    layer1_outputs(9213) <= a and not b;
    layer1_outputs(9214) <= a or b;
    layer1_outputs(9215) <= not (a and b);
    layer1_outputs(9216) <= 1'b0;
    layer1_outputs(9217) <= b;
    layer1_outputs(9218) <= b;
    layer1_outputs(9219) <= a and not b;
    layer1_outputs(9220) <= not (a xor b);
    layer1_outputs(9221) <= b;
    layer1_outputs(9222) <= 1'b0;
    layer1_outputs(9223) <= a or b;
    layer1_outputs(9224) <= a or b;
    layer1_outputs(9225) <= a or b;
    layer1_outputs(9226) <= not a or b;
    layer1_outputs(9227) <= b and not a;
    layer1_outputs(9228) <= not a or b;
    layer1_outputs(9229) <= not b or a;
    layer1_outputs(9230) <= 1'b0;
    layer1_outputs(9231) <= a or b;
    layer1_outputs(9232) <= a;
    layer1_outputs(9233) <= a and b;
    layer1_outputs(9234) <= not b;
    layer1_outputs(9235) <= 1'b0;
    layer1_outputs(9236) <= b and not a;
    layer1_outputs(9237) <= b;
    layer1_outputs(9238) <= not a or b;
    layer1_outputs(9239) <= 1'b1;
    layer1_outputs(9240) <= 1'b0;
    layer1_outputs(9241) <= 1'b1;
    layer1_outputs(9242) <= a or b;
    layer1_outputs(9243) <= not (a or b);
    layer1_outputs(9244) <= not b or a;
    layer1_outputs(9245) <= not (a xor b);
    layer1_outputs(9246) <= 1'b1;
    layer1_outputs(9247) <= not a or b;
    layer1_outputs(9248) <= b and not a;
    layer1_outputs(9249) <= not b;
    layer1_outputs(9250) <= a or b;
    layer1_outputs(9251) <= not b;
    layer1_outputs(9252) <= not (a xor b);
    layer1_outputs(9253) <= not a;
    layer1_outputs(9254) <= b and not a;
    layer1_outputs(9255) <= b;
    layer1_outputs(9256) <= a;
    layer1_outputs(9257) <= a;
    layer1_outputs(9258) <= not a or b;
    layer1_outputs(9259) <= a and not b;
    layer1_outputs(9260) <= not (a and b);
    layer1_outputs(9261) <= not (a or b);
    layer1_outputs(9262) <= not a or b;
    layer1_outputs(9263) <= not b;
    layer1_outputs(9264) <= not a or b;
    layer1_outputs(9265) <= b and not a;
    layer1_outputs(9266) <= a and b;
    layer1_outputs(9267) <= 1'b1;
    layer1_outputs(9268) <= 1'b0;
    layer1_outputs(9269) <= a and b;
    layer1_outputs(9270) <= not b or a;
    layer1_outputs(9271) <= not (a or b);
    layer1_outputs(9272) <= b;
    layer1_outputs(9273) <= not b or a;
    layer1_outputs(9274) <= not b or a;
    layer1_outputs(9275) <= a or b;
    layer1_outputs(9276) <= not a or b;
    layer1_outputs(9277) <= a or b;
    layer1_outputs(9278) <= not (a or b);
    layer1_outputs(9279) <= 1'b0;
    layer1_outputs(9280) <= a and not b;
    layer1_outputs(9281) <= a xor b;
    layer1_outputs(9282) <= a;
    layer1_outputs(9283) <= not a or b;
    layer1_outputs(9284) <= a;
    layer1_outputs(9285) <= not b or a;
    layer1_outputs(9286) <= not (a or b);
    layer1_outputs(9287) <= not b or a;
    layer1_outputs(9288) <= not (a and b);
    layer1_outputs(9289) <= b and not a;
    layer1_outputs(9290) <= a and b;
    layer1_outputs(9291) <= not b;
    layer1_outputs(9292) <= 1'b0;
    layer1_outputs(9293) <= b;
    layer1_outputs(9294) <= not a or b;
    layer1_outputs(9295) <= 1'b1;
    layer1_outputs(9296) <= a;
    layer1_outputs(9297) <= b and not a;
    layer1_outputs(9298) <= not (a and b);
    layer1_outputs(9299) <= not a;
    layer1_outputs(9300) <= b;
    layer1_outputs(9301) <= a;
    layer1_outputs(9302) <= a or b;
    layer1_outputs(9303) <= a and not b;
    layer1_outputs(9304) <= not (a xor b);
    layer1_outputs(9305) <= 1'b0;
    layer1_outputs(9306) <= 1'b0;
    layer1_outputs(9307) <= not a;
    layer1_outputs(9308) <= b and not a;
    layer1_outputs(9309) <= not a or b;
    layer1_outputs(9310) <= 1'b0;
    layer1_outputs(9311) <= b;
    layer1_outputs(9312) <= not b or a;
    layer1_outputs(9313) <= not b;
    layer1_outputs(9314) <= a and not b;
    layer1_outputs(9315) <= b and not a;
    layer1_outputs(9316) <= b and not a;
    layer1_outputs(9317) <= b;
    layer1_outputs(9318) <= not b or a;
    layer1_outputs(9319) <= a or b;
    layer1_outputs(9320) <= b and not a;
    layer1_outputs(9321) <= a or b;
    layer1_outputs(9322) <= b;
    layer1_outputs(9323) <= not b;
    layer1_outputs(9324) <= 1'b1;
    layer1_outputs(9325) <= a and not b;
    layer1_outputs(9326) <= a and b;
    layer1_outputs(9327) <= not b or a;
    layer1_outputs(9328) <= 1'b1;
    layer1_outputs(9329) <= a and not b;
    layer1_outputs(9330) <= not b or a;
    layer1_outputs(9331) <= a and b;
    layer1_outputs(9332) <= 1'b1;
    layer1_outputs(9333) <= not b or a;
    layer1_outputs(9334) <= not (a or b);
    layer1_outputs(9335) <= not (a and b);
    layer1_outputs(9336) <= a and b;
    layer1_outputs(9337) <= not (a or b);
    layer1_outputs(9338) <= not (a and b);
    layer1_outputs(9339) <= b and not a;
    layer1_outputs(9340) <= a or b;
    layer1_outputs(9341) <= not (a and b);
    layer1_outputs(9342) <= not (a or b);
    layer1_outputs(9343) <= not a or b;
    layer1_outputs(9344) <= not (a xor b);
    layer1_outputs(9345) <= not a or b;
    layer1_outputs(9346) <= not b;
    layer1_outputs(9347) <= a xor b;
    layer1_outputs(9348) <= a and b;
    layer1_outputs(9349) <= not a;
    layer1_outputs(9350) <= b and not a;
    layer1_outputs(9351) <= 1'b1;
    layer1_outputs(9352) <= a and b;
    layer1_outputs(9353) <= not a or b;
    layer1_outputs(9354) <= not b or a;
    layer1_outputs(9355) <= a or b;
    layer1_outputs(9356) <= not (a and b);
    layer1_outputs(9357) <= a;
    layer1_outputs(9358) <= not b;
    layer1_outputs(9359) <= b;
    layer1_outputs(9360) <= 1'b1;
    layer1_outputs(9361) <= not b;
    layer1_outputs(9362) <= a;
    layer1_outputs(9363) <= a or b;
    layer1_outputs(9364) <= not (a or b);
    layer1_outputs(9365) <= b;
    layer1_outputs(9366) <= not b;
    layer1_outputs(9367) <= 1'b0;
    layer1_outputs(9368) <= a;
    layer1_outputs(9369) <= b;
    layer1_outputs(9370) <= b;
    layer1_outputs(9371) <= 1'b0;
    layer1_outputs(9372) <= not b or a;
    layer1_outputs(9373) <= a;
    layer1_outputs(9374) <= not a;
    layer1_outputs(9375) <= 1'b0;
    layer1_outputs(9376) <= a or b;
    layer1_outputs(9377) <= 1'b0;
    layer1_outputs(9378) <= not b;
    layer1_outputs(9379) <= a or b;
    layer1_outputs(9380) <= 1'b0;
    layer1_outputs(9381) <= not a;
    layer1_outputs(9382) <= not b;
    layer1_outputs(9383) <= 1'b0;
    layer1_outputs(9384) <= not (a xor b);
    layer1_outputs(9385) <= not (a or b);
    layer1_outputs(9386) <= a and not b;
    layer1_outputs(9387) <= a and not b;
    layer1_outputs(9388) <= not b or a;
    layer1_outputs(9389) <= 1'b0;
    layer1_outputs(9390) <= b and not a;
    layer1_outputs(9391) <= not (a and b);
    layer1_outputs(9392) <= not (a and b);
    layer1_outputs(9393) <= not (a or b);
    layer1_outputs(9394) <= not b;
    layer1_outputs(9395) <= b and not a;
    layer1_outputs(9396) <= 1'b1;
    layer1_outputs(9397) <= 1'b1;
    layer1_outputs(9398) <= not a or b;
    layer1_outputs(9399) <= a and not b;
    layer1_outputs(9400) <= not a;
    layer1_outputs(9401) <= a;
    layer1_outputs(9402) <= not (a xor b);
    layer1_outputs(9403) <= b and not a;
    layer1_outputs(9404) <= not b or a;
    layer1_outputs(9405) <= 1'b0;
    layer1_outputs(9406) <= a;
    layer1_outputs(9407) <= not a or b;
    layer1_outputs(9408) <= not b or a;
    layer1_outputs(9409) <= b;
    layer1_outputs(9410) <= b and not a;
    layer1_outputs(9411) <= not (a and b);
    layer1_outputs(9412) <= a;
    layer1_outputs(9413) <= b;
    layer1_outputs(9414) <= b and not a;
    layer1_outputs(9415) <= a and not b;
    layer1_outputs(9416) <= 1'b0;
    layer1_outputs(9417) <= not a or b;
    layer1_outputs(9418) <= 1'b0;
    layer1_outputs(9419) <= not (a and b);
    layer1_outputs(9420) <= not (a or b);
    layer1_outputs(9421) <= a and b;
    layer1_outputs(9422) <= not b;
    layer1_outputs(9423) <= b;
    layer1_outputs(9424) <= not (a or b);
    layer1_outputs(9425) <= not b or a;
    layer1_outputs(9426) <= a or b;
    layer1_outputs(9427) <= not b;
    layer1_outputs(9428) <= not a or b;
    layer1_outputs(9429) <= not a;
    layer1_outputs(9430) <= not (a or b);
    layer1_outputs(9431) <= a and b;
    layer1_outputs(9432) <= a and not b;
    layer1_outputs(9433) <= b and not a;
    layer1_outputs(9434) <= 1'b0;
    layer1_outputs(9435) <= not b;
    layer1_outputs(9436) <= not b;
    layer1_outputs(9437) <= 1'b0;
    layer1_outputs(9438) <= a and not b;
    layer1_outputs(9439) <= a and b;
    layer1_outputs(9440) <= not (a or b);
    layer1_outputs(9441) <= 1'b0;
    layer1_outputs(9442) <= 1'b1;
    layer1_outputs(9443) <= a or b;
    layer1_outputs(9444) <= not b;
    layer1_outputs(9445) <= not (a or b);
    layer1_outputs(9446) <= a and not b;
    layer1_outputs(9447) <= 1'b0;
    layer1_outputs(9448) <= a;
    layer1_outputs(9449) <= 1'b0;
    layer1_outputs(9450) <= b;
    layer1_outputs(9451) <= 1'b0;
    layer1_outputs(9452) <= 1'b1;
    layer1_outputs(9453) <= b and not a;
    layer1_outputs(9454) <= a and b;
    layer1_outputs(9455) <= a and not b;
    layer1_outputs(9456) <= a or b;
    layer1_outputs(9457) <= a or b;
    layer1_outputs(9458) <= a and b;
    layer1_outputs(9459) <= a;
    layer1_outputs(9460) <= not (a and b);
    layer1_outputs(9461) <= a and b;
    layer1_outputs(9462) <= 1'b0;
    layer1_outputs(9463) <= b;
    layer1_outputs(9464) <= not b or a;
    layer1_outputs(9465) <= 1'b0;
    layer1_outputs(9466) <= not (a xor b);
    layer1_outputs(9467) <= b and not a;
    layer1_outputs(9468) <= a and not b;
    layer1_outputs(9469) <= not (a and b);
    layer1_outputs(9470) <= a and b;
    layer1_outputs(9471) <= not a;
    layer1_outputs(9472) <= 1'b0;
    layer1_outputs(9473) <= not (a or b);
    layer1_outputs(9474) <= 1'b1;
    layer1_outputs(9475) <= not (a and b);
    layer1_outputs(9476) <= 1'b1;
    layer1_outputs(9477) <= a and b;
    layer1_outputs(9478) <= a and not b;
    layer1_outputs(9479) <= b and not a;
    layer1_outputs(9480) <= not (a and b);
    layer1_outputs(9481) <= 1'b0;
    layer1_outputs(9482) <= a;
    layer1_outputs(9483) <= a;
    layer1_outputs(9484) <= a and not b;
    layer1_outputs(9485) <= a;
    layer1_outputs(9486) <= not (a and b);
    layer1_outputs(9487) <= not a or b;
    layer1_outputs(9488) <= a;
    layer1_outputs(9489) <= a;
    layer1_outputs(9490) <= b;
    layer1_outputs(9491) <= not a or b;
    layer1_outputs(9492) <= not b or a;
    layer1_outputs(9493) <= not a or b;
    layer1_outputs(9494) <= not (a or b);
    layer1_outputs(9495) <= not a or b;
    layer1_outputs(9496) <= 1'b1;
    layer1_outputs(9497) <= a;
    layer1_outputs(9498) <= a and not b;
    layer1_outputs(9499) <= a;
    layer1_outputs(9500) <= not b;
    layer1_outputs(9501) <= a or b;
    layer1_outputs(9502) <= 1'b1;
    layer1_outputs(9503) <= 1'b1;
    layer1_outputs(9504) <= not b;
    layer1_outputs(9505) <= a and not b;
    layer1_outputs(9506) <= a;
    layer1_outputs(9507) <= not (a and b);
    layer1_outputs(9508) <= not (a and b);
    layer1_outputs(9509) <= not a or b;
    layer1_outputs(9510) <= not a;
    layer1_outputs(9511) <= a;
    layer1_outputs(9512) <= not (a or b);
    layer1_outputs(9513) <= not (a and b);
    layer1_outputs(9514) <= not b or a;
    layer1_outputs(9515) <= not a;
    layer1_outputs(9516) <= a xor b;
    layer1_outputs(9517) <= not (a and b);
    layer1_outputs(9518) <= a or b;
    layer1_outputs(9519) <= not a;
    layer1_outputs(9520) <= 1'b0;
    layer1_outputs(9521) <= b and not a;
    layer1_outputs(9522) <= a;
    layer1_outputs(9523) <= not a;
    layer1_outputs(9524) <= not (a or b);
    layer1_outputs(9525) <= not a or b;
    layer1_outputs(9526) <= 1'b1;
    layer1_outputs(9527) <= not a;
    layer1_outputs(9528) <= not (a or b);
    layer1_outputs(9529) <= not a or b;
    layer1_outputs(9530) <= not a;
    layer1_outputs(9531) <= b and not a;
    layer1_outputs(9532) <= a and not b;
    layer1_outputs(9533) <= not b or a;
    layer1_outputs(9534) <= a;
    layer1_outputs(9535) <= b and not a;
    layer1_outputs(9536) <= not (a and b);
    layer1_outputs(9537) <= not (a or b);
    layer1_outputs(9538) <= 1'b0;
    layer1_outputs(9539) <= not a or b;
    layer1_outputs(9540) <= a and not b;
    layer1_outputs(9541) <= not (a and b);
    layer1_outputs(9542) <= a;
    layer1_outputs(9543) <= a or b;
    layer1_outputs(9544) <= a and b;
    layer1_outputs(9545) <= a and b;
    layer1_outputs(9546) <= a or b;
    layer1_outputs(9547) <= a xor b;
    layer1_outputs(9548) <= 1'b0;
    layer1_outputs(9549) <= not b or a;
    layer1_outputs(9550) <= not b;
    layer1_outputs(9551) <= not b;
    layer1_outputs(9552) <= not b;
    layer1_outputs(9553) <= a xor b;
    layer1_outputs(9554) <= not (a or b);
    layer1_outputs(9555) <= not (a and b);
    layer1_outputs(9556) <= a or b;
    layer1_outputs(9557) <= 1'b1;
    layer1_outputs(9558) <= not (a or b);
    layer1_outputs(9559) <= b;
    layer1_outputs(9560) <= not b;
    layer1_outputs(9561) <= a or b;
    layer1_outputs(9562) <= not a;
    layer1_outputs(9563) <= not (a and b);
    layer1_outputs(9564) <= a or b;
    layer1_outputs(9565) <= a and not b;
    layer1_outputs(9566) <= a;
    layer1_outputs(9567) <= not b or a;
    layer1_outputs(9568) <= 1'b0;
    layer1_outputs(9569) <= b and not a;
    layer1_outputs(9570) <= not a or b;
    layer1_outputs(9571) <= not a or b;
    layer1_outputs(9572) <= not b;
    layer1_outputs(9573) <= not (a or b);
    layer1_outputs(9574) <= a and not b;
    layer1_outputs(9575) <= a and not b;
    layer1_outputs(9576) <= not a or b;
    layer1_outputs(9577) <= a and b;
    layer1_outputs(9578) <= not (a and b);
    layer1_outputs(9579) <= a;
    layer1_outputs(9580) <= 1'b1;
    layer1_outputs(9581) <= not b or a;
    layer1_outputs(9582) <= not a or b;
    layer1_outputs(9583) <= not a or b;
    layer1_outputs(9584) <= a xor b;
    layer1_outputs(9585) <= b;
    layer1_outputs(9586) <= a;
    layer1_outputs(9587) <= a and not b;
    layer1_outputs(9588) <= not a;
    layer1_outputs(9589) <= not a or b;
    layer1_outputs(9590) <= not a or b;
    layer1_outputs(9591) <= not (a xor b);
    layer1_outputs(9592) <= 1'b0;
    layer1_outputs(9593) <= a and b;
    layer1_outputs(9594) <= a and b;
    layer1_outputs(9595) <= not b or a;
    layer1_outputs(9596) <= not (a or b);
    layer1_outputs(9597) <= not a or b;
    layer1_outputs(9598) <= not (a or b);
    layer1_outputs(9599) <= a and not b;
    layer1_outputs(9600) <= not a;
    layer1_outputs(9601) <= not (a or b);
    layer1_outputs(9602) <= a and not b;
    layer1_outputs(9603) <= not a;
    layer1_outputs(9604) <= a and b;
    layer1_outputs(9605) <= not a;
    layer1_outputs(9606) <= 1'b1;
    layer1_outputs(9607) <= not b or a;
    layer1_outputs(9608) <= not a or b;
    layer1_outputs(9609) <= a and not b;
    layer1_outputs(9610) <= a and b;
    layer1_outputs(9611) <= not (a or b);
    layer1_outputs(9612) <= b and not a;
    layer1_outputs(9613) <= not a or b;
    layer1_outputs(9614) <= not a or b;
    layer1_outputs(9615) <= a;
    layer1_outputs(9616) <= a and b;
    layer1_outputs(9617) <= not (a or b);
    layer1_outputs(9618) <= not (a and b);
    layer1_outputs(9619) <= a;
    layer1_outputs(9620) <= b and not a;
    layer1_outputs(9621) <= not a or b;
    layer1_outputs(9622) <= not a;
    layer1_outputs(9623) <= a;
    layer1_outputs(9624) <= a and not b;
    layer1_outputs(9625) <= a or b;
    layer1_outputs(9626) <= 1'b0;
    layer1_outputs(9627) <= not a or b;
    layer1_outputs(9628) <= 1'b1;
    layer1_outputs(9629) <= not b or a;
    layer1_outputs(9630) <= not a;
    layer1_outputs(9631) <= not (a or b);
    layer1_outputs(9632) <= not a;
    layer1_outputs(9633) <= not b;
    layer1_outputs(9634) <= b and not a;
    layer1_outputs(9635) <= not b;
    layer1_outputs(9636) <= b;
    layer1_outputs(9637) <= a or b;
    layer1_outputs(9638) <= not b;
    layer1_outputs(9639) <= a or b;
    layer1_outputs(9640) <= b and not a;
    layer1_outputs(9641) <= not a or b;
    layer1_outputs(9642) <= b;
    layer1_outputs(9643) <= b and not a;
    layer1_outputs(9644) <= 1'b1;
    layer1_outputs(9645) <= a or b;
    layer1_outputs(9646) <= b;
    layer1_outputs(9647) <= 1'b1;
    layer1_outputs(9648) <= not b;
    layer1_outputs(9649) <= a and not b;
    layer1_outputs(9650) <= a and b;
    layer1_outputs(9651) <= b and not a;
    layer1_outputs(9652) <= not (a or b);
    layer1_outputs(9653) <= b;
    layer1_outputs(9654) <= not b;
    layer1_outputs(9655) <= not a or b;
    layer1_outputs(9656) <= not (a xor b);
    layer1_outputs(9657) <= a;
    layer1_outputs(9658) <= not a or b;
    layer1_outputs(9659) <= a and b;
    layer1_outputs(9660) <= not b;
    layer1_outputs(9661) <= not a;
    layer1_outputs(9662) <= not (a and b);
    layer1_outputs(9663) <= a and not b;
    layer1_outputs(9664) <= a and b;
    layer1_outputs(9665) <= not b;
    layer1_outputs(9666) <= b and not a;
    layer1_outputs(9667) <= 1'b1;
    layer1_outputs(9668) <= not a;
    layer1_outputs(9669) <= not b or a;
    layer1_outputs(9670) <= b and not a;
    layer1_outputs(9671) <= not b;
    layer1_outputs(9672) <= a and not b;
    layer1_outputs(9673) <= not a or b;
    layer1_outputs(9674) <= b and not a;
    layer1_outputs(9675) <= not a or b;
    layer1_outputs(9676) <= not a;
    layer1_outputs(9677) <= not (a and b);
    layer1_outputs(9678) <= b and not a;
    layer1_outputs(9679) <= not a or b;
    layer1_outputs(9680) <= a and b;
    layer1_outputs(9681) <= 1'b0;
    layer1_outputs(9682) <= not (a or b);
    layer1_outputs(9683) <= not (a and b);
    layer1_outputs(9684) <= 1'b1;
    layer1_outputs(9685) <= 1'b1;
    layer1_outputs(9686) <= not (a and b);
    layer1_outputs(9687) <= 1'b1;
    layer1_outputs(9688) <= not b or a;
    layer1_outputs(9689) <= not a or b;
    layer1_outputs(9690) <= not b;
    layer1_outputs(9691) <= 1'b0;
    layer1_outputs(9692) <= 1'b0;
    layer1_outputs(9693) <= a and b;
    layer1_outputs(9694) <= not a or b;
    layer1_outputs(9695) <= not b;
    layer1_outputs(9696) <= b and not a;
    layer1_outputs(9697) <= 1'b0;
    layer1_outputs(9698) <= a and not b;
    layer1_outputs(9699) <= not (a xor b);
    layer1_outputs(9700) <= 1'b0;
    layer1_outputs(9701) <= not (a or b);
    layer1_outputs(9702) <= 1'b0;
    layer1_outputs(9703) <= not a or b;
    layer1_outputs(9704) <= a and not b;
    layer1_outputs(9705) <= b;
    layer1_outputs(9706) <= a and not b;
    layer1_outputs(9707) <= not b or a;
    layer1_outputs(9708) <= not a or b;
    layer1_outputs(9709) <= b;
    layer1_outputs(9710) <= a and b;
    layer1_outputs(9711) <= b;
    layer1_outputs(9712) <= not a;
    layer1_outputs(9713) <= a or b;
    layer1_outputs(9714) <= not (a and b);
    layer1_outputs(9715) <= a and not b;
    layer1_outputs(9716) <= not a;
    layer1_outputs(9717) <= b and not a;
    layer1_outputs(9718) <= 1'b1;
    layer1_outputs(9719) <= a;
    layer1_outputs(9720) <= not (a and b);
    layer1_outputs(9721) <= 1'b1;
    layer1_outputs(9722) <= a;
    layer1_outputs(9723) <= not (a or b);
    layer1_outputs(9724) <= a or b;
    layer1_outputs(9725) <= a;
    layer1_outputs(9726) <= not b or a;
    layer1_outputs(9727) <= not (a or b);
    layer1_outputs(9728) <= 1'b0;
    layer1_outputs(9729) <= 1'b0;
    layer1_outputs(9730) <= not (a xor b);
    layer1_outputs(9731) <= b and not a;
    layer1_outputs(9732) <= not b;
    layer1_outputs(9733) <= not b;
    layer1_outputs(9734) <= a;
    layer1_outputs(9735) <= a and not b;
    layer1_outputs(9736) <= a and b;
    layer1_outputs(9737) <= a;
    layer1_outputs(9738) <= not a or b;
    layer1_outputs(9739) <= a;
    layer1_outputs(9740) <= not b;
    layer1_outputs(9741) <= not a or b;
    layer1_outputs(9742) <= a and not b;
    layer1_outputs(9743) <= a or b;
    layer1_outputs(9744) <= 1'b0;
    layer1_outputs(9745) <= not a or b;
    layer1_outputs(9746) <= a;
    layer1_outputs(9747) <= not a;
    layer1_outputs(9748) <= a and not b;
    layer1_outputs(9749) <= not a or b;
    layer1_outputs(9750) <= a;
    layer1_outputs(9751) <= 1'b1;
    layer1_outputs(9752) <= b and not a;
    layer1_outputs(9753) <= 1'b0;
    layer1_outputs(9754) <= not (a and b);
    layer1_outputs(9755) <= 1'b0;
    layer1_outputs(9756) <= a or b;
    layer1_outputs(9757) <= a and not b;
    layer1_outputs(9758) <= b and not a;
    layer1_outputs(9759) <= b;
    layer1_outputs(9760) <= not b;
    layer1_outputs(9761) <= a or b;
    layer1_outputs(9762) <= 1'b0;
    layer1_outputs(9763) <= a and b;
    layer1_outputs(9764) <= not b or a;
    layer1_outputs(9765) <= not (a xor b);
    layer1_outputs(9766) <= a xor b;
    layer1_outputs(9767) <= not b or a;
    layer1_outputs(9768) <= b and not a;
    layer1_outputs(9769) <= not b or a;
    layer1_outputs(9770) <= not (a xor b);
    layer1_outputs(9771) <= not b or a;
    layer1_outputs(9772) <= b and not a;
    layer1_outputs(9773) <= 1'b1;
    layer1_outputs(9774) <= not a or b;
    layer1_outputs(9775) <= 1'b1;
    layer1_outputs(9776) <= a and b;
    layer1_outputs(9777) <= not (a and b);
    layer1_outputs(9778) <= a xor b;
    layer1_outputs(9779) <= not a;
    layer1_outputs(9780) <= 1'b0;
    layer1_outputs(9781) <= not a or b;
    layer1_outputs(9782) <= 1'b1;
    layer1_outputs(9783) <= not (a and b);
    layer1_outputs(9784) <= 1'b1;
    layer1_outputs(9785) <= a or b;
    layer1_outputs(9786) <= not b or a;
    layer1_outputs(9787) <= a or b;
    layer1_outputs(9788) <= not b or a;
    layer1_outputs(9789) <= not b or a;
    layer1_outputs(9790) <= not b or a;
    layer1_outputs(9791) <= not b;
    layer1_outputs(9792) <= 1'b0;
    layer1_outputs(9793) <= not a or b;
    layer1_outputs(9794) <= 1'b1;
    layer1_outputs(9795) <= not a or b;
    layer1_outputs(9796) <= not a;
    layer1_outputs(9797) <= not b or a;
    layer1_outputs(9798) <= not b;
    layer1_outputs(9799) <= 1'b0;
    layer1_outputs(9800) <= not a or b;
    layer1_outputs(9801) <= b;
    layer1_outputs(9802) <= not (a xor b);
    layer1_outputs(9803) <= a and not b;
    layer1_outputs(9804) <= not (a and b);
    layer1_outputs(9805) <= not b or a;
    layer1_outputs(9806) <= b and not a;
    layer1_outputs(9807) <= not b;
    layer1_outputs(9808) <= a or b;
    layer1_outputs(9809) <= not a or b;
    layer1_outputs(9810) <= 1'b0;
    layer1_outputs(9811) <= a and not b;
    layer1_outputs(9812) <= 1'b0;
    layer1_outputs(9813) <= 1'b0;
    layer1_outputs(9814) <= a and b;
    layer1_outputs(9815) <= b;
    layer1_outputs(9816) <= 1'b0;
    layer1_outputs(9817) <= not a;
    layer1_outputs(9818) <= 1'b0;
    layer1_outputs(9819) <= 1'b1;
    layer1_outputs(9820) <= b;
    layer1_outputs(9821) <= not (a or b);
    layer1_outputs(9822) <= b;
    layer1_outputs(9823) <= 1'b1;
    layer1_outputs(9824) <= 1'b1;
    layer1_outputs(9825) <= not a or b;
    layer1_outputs(9826) <= not a or b;
    layer1_outputs(9827) <= not a;
    layer1_outputs(9828) <= a and b;
    layer1_outputs(9829) <= a and b;
    layer1_outputs(9830) <= not a or b;
    layer1_outputs(9831) <= a or b;
    layer1_outputs(9832) <= a and b;
    layer1_outputs(9833) <= a and b;
    layer1_outputs(9834) <= not a;
    layer1_outputs(9835) <= not a;
    layer1_outputs(9836) <= a;
    layer1_outputs(9837) <= b;
    layer1_outputs(9838) <= a and not b;
    layer1_outputs(9839) <= not (a xor b);
    layer1_outputs(9840) <= 1'b1;
    layer1_outputs(9841) <= not a or b;
    layer1_outputs(9842) <= not (a and b);
    layer1_outputs(9843) <= not (a or b);
    layer1_outputs(9844) <= not b;
    layer1_outputs(9845) <= not (a xor b);
    layer1_outputs(9846) <= 1'b0;
    layer1_outputs(9847) <= not b;
    layer1_outputs(9848) <= a;
    layer1_outputs(9849) <= a;
    layer1_outputs(9850) <= 1'b0;
    layer1_outputs(9851) <= a;
    layer1_outputs(9852) <= not b or a;
    layer1_outputs(9853) <= not a or b;
    layer1_outputs(9854) <= 1'b1;
    layer1_outputs(9855) <= not b or a;
    layer1_outputs(9856) <= not a or b;
    layer1_outputs(9857) <= not a or b;
    layer1_outputs(9858) <= a or b;
    layer1_outputs(9859) <= 1'b1;
    layer1_outputs(9860) <= 1'b1;
    layer1_outputs(9861) <= not b or a;
    layer1_outputs(9862) <= not b or a;
    layer1_outputs(9863) <= not (a and b);
    layer1_outputs(9864) <= not (a or b);
    layer1_outputs(9865) <= a or b;
    layer1_outputs(9866) <= a and not b;
    layer1_outputs(9867) <= not a;
    layer1_outputs(9868) <= a and b;
    layer1_outputs(9869) <= b;
    layer1_outputs(9870) <= 1'b1;
    layer1_outputs(9871) <= a or b;
    layer1_outputs(9872) <= a and b;
    layer1_outputs(9873) <= 1'b0;
    layer1_outputs(9874) <= not b;
    layer1_outputs(9875) <= not a or b;
    layer1_outputs(9876) <= not a;
    layer1_outputs(9877) <= not a;
    layer1_outputs(9878) <= a or b;
    layer1_outputs(9879) <= a and b;
    layer1_outputs(9880) <= not b;
    layer1_outputs(9881) <= b and not a;
    layer1_outputs(9882) <= 1'b0;
    layer1_outputs(9883) <= 1'b0;
    layer1_outputs(9884) <= not (a and b);
    layer1_outputs(9885) <= 1'b0;
    layer1_outputs(9886) <= 1'b0;
    layer1_outputs(9887) <= 1'b0;
    layer1_outputs(9888) <= not a;
    layer1_outputs(9889) <= not a;
    layer1_outputs(9890) <= not a;
    layer1_outputs(9891) <= a or b;
    layer1_outputs(9892) <= not b or a;
    layer1_outputs(9893) <= a or b;
    layer1_outputs(9894) <= not (a or b);
    layer1_outputs(9895) <= a and not b;
    layer1_outputs(9896) <= 1'b1;
    layer1_outputs(9897) <= a;
    layer1_outputs(9898) <= not b or a;
    layer1_outputs(9899) <= a or b;
    layer1_outputs(9900) <= not b;
    layer1_outputs(9901) <= not (a or b);
    layer1_outputs(9902) <= not b or a;
    layer1_outputs(9903) <= not (a xor b);
    layer1_outputs(9904) <= 1'b0;
    layer1_outputs(9905) <= a and b;
    layer1_outputs(9906) <= not a or b;
    layer1_outputs(9907) <= a and not b;
    layer1_outputs(9908) <= 1'b1;
    layer1_outputs(9909) <= b and not a;
    layer1_outputs(9910) <= not (a and b);
    layer1_outputs(9911) <= not (a or b);
    layer1_outputs(9912) <= a xor b;
    layer1_outputs(9913) <= not a;
    layer1_outputs(9914) <= 1'b1;
    layer1_outputs(9915) <= not b;
    layer1_outputs(9916) <= a;
    layer1_outputs(9917) <= not (a or b);
    layer1_outputs(9918) <= a or b;
    layer1_outputs(9919) <= not a;
    layer1_outputs(9920) <= not (a and b);
    layer1_outputs(9921) <= 1'b0;
    layer1_outputs(9922) <= b and not a;
    layer1_outputs(9923) <= a;
    layer1_outputs(9924) <= a and b;
    layer1_outputs(9925) <= not (a and b);
    layer1_outputs(9926) <= not b;
    layer1_outputs(9927) <= not a or b;
    layer1_outputs(9928) <= not a or b;
    layer1_outputs(9929) <= b and not a;
    layer1_outputs(9930) <= not (a and b);
    layer1_outputs(9931) <= not b;
    layer1_outputs(9932) <= not b;
    layer1_outputs(9933) <= not a;
    layer1_outputs(9934) <= 1'b1;
    layer1_outputs(9935) <= a and b;
    layer1_outputs(9936) <= a and b;
    layer1_outputs(9937) <= a and not b;
    layer1_outputs(9938) <= not (a and b);
    layer1_outputs(9939) <= a;
    layer1_outputs(9940) <= not a or b;
    layer1_outputs(9941) <= 1'b0;
    layer1_outputs(9942) <= not b;
    layer1_outputs(9943) <= a and not b;
    layer1_outputs(9944) <= a and b;
    layer1_outputs(9945) <= not (a and b);
    layer1_outputs(9946) <= b;
    layer1_outputs(9947) <= not a;
    layer1_outputs(9948) <= a or b;
    layer1_outputs(9949) <= a and not b;
    layer1_outputs(9950) <= not a or b;
    layer1_outputs(9951) <= not b or a;
    layer1_outputs(9952) <= 1'b0;
    layer1_outputs(9953) <= 1'b0;
    layer1_outputs(9954) <= 1'b1;
    layer1_outputs(9955) <= not a or b;
    layer1_outputs(9956) <= not a or b;
    layer1_outputs(9957) <= not b;
    layer1_outputs(9958) <= a and not b;
    layer1_outputs(9959) <= 1'b1;
    layer1_outputs(9960) <= a and b;
    layer1_outputs(9961) <= not (a and b);
    layer1_outputs(9962) <= 1'b1;
    layer1_outputs(9963) <= a and not b;
    layer1_outputs(9964) <= not (a xor b);
    layer1_outputs(9965) <= a and b;
    layer1_outputs(9966) <= not (a xor b);
    layer1_outputs(9967) <= a;
    layer1_outputs(9968) <= a and not b;
    layer1_outputs(9969) <= not a;
    layer1_outputs(9970) <= b;
    layer1_outputs(9971) <= not b;
    layer1_outputs(9972) <= a;
    layer1_outputs(9973) <= 1'b1;
    layer1_outputs(9974) <= not b or a;
    layer1_outputs(9975) <= a xor b;
    layer1_outputs(9976) <= not a;
    layer1_outputs(9977) <= not (a or b);
    layer1_outputs(9978) <= not (a and b);
    layer1_outputs(9979) <= not (a or b);
    layer1_outputs(9980) <= not b;
    layer1_outputs(9981) <= b;
    layer1_outputs(9982) <= b and not a;
    layer1_outputs(9983) <= 1'b0;
    layer1_outputs(9984) <= b;
    layer1_outputs(9985) <= not (a and b);
    layer1_outputs(9986) <= b and not a;
    layer1_outputs(9987) <= not (a or b);
    layer1_outputs(9988) <= a and not b;
    layer1_outputs(9989) <= 1'b0;
    layer1_outputs(9990) <= not b;
    layer1_outputs(9991) <= a and b;
    layer1_outputs(9992) <= 1'b0;
    layer1_outputs(9993) <= b;
    layer1_outputs(9994) <= a and b;
    layer1_outputs(9995) <= a or b;
    layer1_outputs(9996) <= not a;
    layer1_outputs(9997) <= a or b;
    layer1_outputs(9998) <= not a or b;
    layer1_outputs(9999) <= a and b;
    layer1_outputs(10000) <= a and b;
    layer1_outputs(10001) <= not b or a;
    layer1_outputs(10002) <= b and not a;
    layer1_outputs(10003) <= not (a and b);
    layer1_outputs(10004) <= b and not a;
    layer1_outputs(10005) <= not a or b;
    layer1_outputs(10006) <= a;
    layer1_outputs(10007) <= a and not b;
    layer1_outputs(10008) <= not (a or b);
    layer1_outputs(10009) <= b and not a;
    layer1_outputs(10010) <= a or b;
    layer1_outputs(10011) <= a xor b;
    layer1_outputs(10012) <= not a;
    layer1_outputs(10013) <= not b;
    layer1_outputs(10014) <= not a;
    layer1_outputs(10015) <= a and b;
    layer1_outputs(10016) <= a;
    layer1_outputs(10017) <= a and b;
    layer1_outputs(10018) <= 1'b1;
    layer1_outputs(10019) <= not (a and b);
    layer1_outputs(10020) <= not a;
    layer1_outputs(10021) <= 1'b1;
    layer1_outputs(10022) <= not (a and b);
    layer1_outputs(10023) <= not (a xor b);
    layer1_outputs(10024) <= not a or b;
    layer1_outputs(10025) <= a and not b;
    layer1_outputs(10026) <= not (a or b);
    layer1_outputs(10027) <= not b;
    layer1_outputs(10028) <= not b or a;
    layer1_outputs(10029) <= b;
    layer1_outputs(10030) <= a or b;
    layer1_outputs(10031) <= b and not a;
    layer1_outputs(10032) <= 1'b1;
    layer1_outputs(10033) <= a and not b;
    layer1_outputs(10034) <= not (a and b);
    layer1_outputs(10035) <= b;
    layer1_outputs(10036) <= not b or a;
    layer1_outputs(10037) <= not b or a;
    layer1_outputs(10038) <= not (a and b);
    layer1_outputs(10039) <= not (a and b);
    layer1_outputs(10040) <= 1'b1;
    layer1_outputs(10041) <= not b or a;
    layer1_outputs(10042) <= b;
    layer1_outputs(10043) <= not b or a;
    layer1_outputs(10044) <= not b or a;
    layer1_outputs(10045) <= not a;
    layer1_outputs(10046) <= a and b;
    layer1_outputs(10047) <= 1'b0;
    layer1_outputs(10048) <= a or b;
    layer1_outputs(10049) <= a;
    layer1_outputs(10050) <= not a or b;
    layer1_outputs(10051) <= 1'b1;
    layer1_outputs(10052) <= b;
    layer1_outputs(10053) <= 1'b0;
    layer1_outputs(10054) <= not a or b;
    layer1_outputs(10055) <= not b or a;
    layer1_outputs(10056) <= not b or a;
    layer1_outputs(10057) <= not (a and b);
    layer1_outputs(10058) <= a and not b;
    layer1_outputs(10059) <= 1'b0;
    layer1_outputs(10060) <= not (a or b);
    layer1_outputs(10061) <= a xor b;
    layer1_outputs(10062) <= not (a or b);
    layer1_outputs(10063) <= b and not a;
    layer1_outputs(10064) <= not a;
    layer1_outputs(10065) <= not a;
    layer1_outputs(10066) <= b and not a;
    layer1_outputs(10067) <= a xor b;
    layer1_outputs(10068) <= 1'b1;
    layer1_outputs(10069) <= b;
    layer1_outputs(10070) <= 1'b0;
    layer1_outputs(10071) <= a;
    layer1_outputs(10072) <= not a or b;
    layer1_outputs(10073) <= a and not b;
    layer1_outputs(10074) <= not (a or b);
    layer1_outputs(10075) <= 1'b1;
    layer1_outputs(10076) <= not b;
    layer1_outputs(10077) <= a or b;
    layer1_outputs(10078) <= a and b;
    layer1_outputs(10079) <= not a or b;
    layer1_outputs(10080) <= not (a and b);
    layer1_outputs(10081) <= not (a and b);
    layer1_outputs(10082) <= not a;
    layer1_outputs(10083) <= a xor b;
    layer1_outputs(10084) <= a;
    layer1_outputs(10085) <= a;
    layer1_outputs(10086) <= b;
    layer1_outputs(10087) <= b and not a;
    layer1_outputs(10088) <= b and not a;
    layer1_outputs(10089) <= a or b;
    layer1_outputs(10090) <= not b;
    layer1_outputs(10091) <= a or b;
    layer1_outputs(10092) <= b;
    layer1_outputs(10093) <= not a;
    layer1_outputs(10094) <= a;
    layer1_outputs(10095) <= b;
    layer1_outputs(10096) <= a and not b;
    layer1_outputs(10097) <= a or b;
    layer1_outputs(10098) <= a and not b;
    layer1_outputs(10099) <= a or b;
    layer1_outputs(10100) <= 1'b1;
    layer1_outputs(10101) <= not (a or b);
    layer1_outputs(10102) <= 1'b1;
    layer1_outputs(10103) <= not b or a;
    layer1_outputs(10104) <= not a or b;
    layer1_outputs(10105) <= not (a xor b);
    layer1_outputs(10106) <= not a or b;
    layer1_outputs(10107) <= not (a or b);
    layer1_outputs(10108) <= not a or b;
    layer1_outputs(10109) <= a;
    layer1_outputs(10110) <= not (a and b);
    layer1_outputs(10111) <= not a or b;
    layer1_outputs(10112) <= a and b;
    layer1_outputs(10113) <= not b;
    layer1_outputs(10114) <= not (a and b);
    layer1_outputs(10115) <= a;
    layer1_outputs(10116) <= a and not b;
    layer1_outputs(10117) <= not b;
    layer1_outputs(10118) <= 1'b1;
    layer1_outputs(10119) <= not a;
    layer1_outputs(10120) <= not (a and b);
    layer1_outputs(10121) <= a and b;
    layer1_outputs(10122) <= a and b;
    layer1_outputs(10123) <= a;
    layer1_outputs(10124) <= b and not a;
    layer1_outputs(10125) <= not b;
    layer1_outputs(10126) <= not b;
    layer1_outputs(10127) <= not a;
    layer1_outputs(10128) <= not (a xor b);
    layer1_outputs(10129) <= a xor b;
    layer1_outputs(10130) <= 1'b0;
    layer1_outputs(10131) <= not a;
    layer1_outputs(10132) <= b and not a;
    layer1_outputs(10133) <= a xor b;
    layer1_outputs(10134) <= not (a xor b);
    layer1_outputs(10135) <= not a;
    layer1_outputs(10136) <= not (a xor b);
    layer1_outputs(10137) <= b;
    layer1_outputs(10138) <= b;
    layer1_outputs(10139) <= not a;
    layer1_outputs(10140) <= a and b;
    layer1_outputs(10141) <= a;
    layer1_outputs(10142) <= 1'b1;
    layer1_outputs(10143) <= b;
    layer1_outputs(10144) <= b and not a;
    layer1_outputs(10145) <= not (a xor b);
    layer1_outputs(10146) <= not a;
    layer1_outputs(10147) <= a;
    layer1_outputs(10148) <= 1'b1;
    layer1_outputs(10149) <= 1'b1;
    layer1_outputs(10150) <= not b;
    layer1_outputs(10151) <= b and not a;
    layer1_outputs(10152) <= not b or a;
    layer1_outputs(10153) <= not a or b;
    layer1_outputs(10154) <= b and not a;
    layer1_outputs(10155) <= a or b;
    layer1_outputs(10156) <= not a or b;
    layer1_outputs(10157) <= not b or a;
    layer1_outputs(10158) <= not b;
    layer1_outputs(10159) <= not (a and b);
    layer1_outputs(10160) <= not (a xor b);
    layer1_outputs(10161) <= a or b;
    layer1_outputs(10162) <= a xor b;
    layer1_outputs(10163) <= not a;
    layer1_outputs(10164) <= not a or b;
    layer1_outputs(10165) <= not (a or b);
    layer1_outputs(10166) <= 1'b1;
    layer1_outputs(10167) <= not b or a;
    layer1_outputs(10168) <= a and b;
    layer1_outputs(10169) <= 1'b0;
    layer1_outputs(10170) <= b and not a;
    layer1_outputs(10171) <= a;
    layer1_outputs(10172) <= a xor b;
    layer1_outputs(10173) <= a and not b;
    layer1_outputs(10174) <= b;
    layer1_outputs(10175) <= not a;
    layer1_outputs(10176) <= 1'b0;
    layer1_outputs(10177) <= 1'b1;
    layer1_outputs(10178) <= 1'b1;
    layer1_outputs(10179) <= not (a or b);
    layer1_outputs(10180) <= not (a or b);
    layer1_outputs(10181) <= not a or b;
    layer1_outputs(10182) <= 1'b1;
    layer1_outputs(10183) <= b;
    layer1_outputs(10184) <= not b;
    layer1_outputs(10185) <= a or b;
    layer1_outputs(10186) <= not a or b;
    layer1_outputs(10187) <= 1'b1;
    layer1_outputs(10188) <= not (a or b);
    layer1_outputs(10189) <= not b or a;
    layer1_outputs(10190) <= not b;
    layer1_outputs(10191) <= a;
    layer1_outputs(10192) <= b and not a;
    layer1_outputs(10193) <= not b or a;
    layer1_outputs(10194) <= not a or b;
    layer1_outputs(10195) <= 1'b0;
    layer1_outputs(10196) <= not a or b;
    layer1_outputs(10197) <= a and b;
    layer1_outputs(10198) <= not b or a;
    layer1_outputs(10199) <= not (a and b);
    layer1_outputs(10200) <= not a;
    layer1_outputs(10201) <= not (a xor b);
    layer1_outputs(10202) <= a and not b;
    layer1_outputs(10203) <= not (a or b);
    layer1_outputs(10204) <= 1'b1;
    layer1_outputs(10205) <= not a or b;
    layer1_outputs(10206) <= a;
    layer1_outputs(10207) <= 1'b0;
    layer1_outputs(10208) <= 1'b0;
    layer1_outputs(10209) <= not (a or b);
    layer1_outputs(10210) <= not a;
    layer1_outputs(10211) <= 1'b0;
    layer1_outputs(10212) <= a or b;
    layer1_outputs(10213) <= a or b;
    layer1_outputs(10214) <= a;
    layer1_outputs(10215) <= a;
    layer1_outputs(10216) <= not (a or b);
    layer1_outputs(10217) <= b;
    layer1_outputs(10218) <= not b;
    layer1_outputs(10219) <= b and not a;
    layer1_outputs(10220) <= not a;
    layer1_outputs(10221) <= not (a xor b);
    layer1_outputs(10222) <= b and not a;
    layer1_outputs(10223) <= not a or b;
    layer1_outputs(10224) <= 1'b1;
    layer1_outputs(10225) <= not b or a;
    layer1_outputs(10226) <= b and not a;
    layer1_outputs(10227) <= a xor b;
    layer1_outputs(10228) <= 1'b0;
    layer1_outputs(10229) <= a or b;
    layer1_outputs(10230) <= not b;
    layer1_outputs(10231) <= b and not a;
    layer1_outputs(10232) <= not (a or b);
    layer1_outputs(10233) <= 1'b1;
    layer1_outputs(10234) <= a and not b;
    layer1_outputs(10235) <= not a;
    layer1_outputs(10236) <= 1'b0;
    layer1_outputs(10237) <= 1'b1;
    layer1_outputs(10238) <= not (a xor b);
    layer1_outputs(10239) <= a and b;
    layer2_outputs(0) <= 1'b0;
    layer2_outputs(1) <= b and not a;
    layer2_outputs(2) <= not a or b;
    layer2_outputs(3) <= a and not b;
    layer2_outputs(4) <= not b;
    layer2_outputs(5) <= not (a and b);
    layer2_outputs(6) <= 1'b0;
    layer2_outputs(7) <= a xor b;
    layer2_outputs(8) <= a;
    layer2_outputs(9) <= a or b;
    layer2_outputs(10) <= not a or b;
    layer2_outputs(11) <= not (a and b);
    layer2_outputs(12) <= a;
    layer2_outputs(13) <= not (a and b);
    layer2_outputs(14) <= not (a or b);
    layer2_outputs(15) <= b;
    layer2_outputs(16) <= not (a and b);
    layer2_outputs(17) <= not (a or b);
    layer2_outputs(18) <= not a or b;
    layer2_outputs(19) <= a or b;
    layer2_outputs(20) <= not (a and b);
    layer2_outputs(21) <= not b or a;
    layer2_outputs(22) <= a;
    layer2_outputs(23) <= a or b;
    layer2_outputs(24) <= not (a or b);
    layer2_outputs(25) <= not (a or b);
    layer2_outputs(26) <= a and b;
    layer2_outputs(27) <= a or b;
    layer2_outputs(28) <= not a or b;
    layer2_outputs(29) <= not a;
    layer2_outputs(30) <= a xor b;
    layer2_outputs(31) <= not b or a;
    layer2_outputs(32) <= not b;
    layer2_outputs(33) <= 1'b1;
    layer2_outputs(34) <= not a or b;
    layer2_outputs(35) <= b;
    layer2_outputs(36) <= a or b;
    layer2_outputs(37) <= 1'b1;
    layer2_outputs(38) <= not (a xor b);
    layer2_outputs(39) <= 1'b0;
    layer2_outputs(40) <= a;
    layer2_outputs(41) <= b and not a;
    layer2_outputs(42) <= not (a and b);
    layer2_outputs(43) <= a and not b;
    layer2_outputs(44) <= not a;
    layer2_outputs(45) <= 1'b1;
    layer2_outputs(46) <= not a;
    layer2_outputs(47) <= 1'b0;
    layer2_outputs(48) <= 1'b0;
    layer2_outputs(49) <= a xor b;
    layer2_outputs(50) <= 1'b1;
    layer2_outputs(51) <= b and not a;
    layer2_outputs(52) <= a and not b;
    layer2_outputs(53) <= not (a xor b);
    layer2_outputs(54) <= b;
    layer2_outputs(55) <= a and b;
    layer2_outputs(56) <= not b;
    layer2_outputs(57) <= b;
    layer2_outputs(58) <= a and b;
    layer2_outputs(59) <= not (a or b);
    layer2_outputs(60) <= not b or a;
    layer2_outputs(61) <= a and b;
    layer2_outputs(62) <= a;
    layer2_outputs(63) <= a and b;
    layer2_outputs(64) <= 1'b0;
    layer2_outputs(65) <= 1'b0;
    layer2_outputs(66) <= a and not b;
    layer2_outputs(67) <= not (a or b);
    layer2_outputs(68) <= 1'b1;
    layer2_outputs(69) <= a;
    layer2_outputs(70) <= a and b;
    layer2_outputs(71) <= b and not a;
    layer2_outputs(72) <= a or b;
    layer2_outputs(73) <= a;
    layer2_outputs(74) <= 1'b0;
    layer2_outputs(75) <= b;
    layer2_outputs(76) <= b;
    layer2_outputs(77) <= b and not a;
    layer2_outputs(78) <= 1'b0;
    layer2_outputs(79) <= not (a or b);
    layer2_outputs(80) <= not a;
    layer2_outputs(81) <= a or b;
    layer2_outputs(82) <= b;
    layer2_outputs(83) <= a and not b;
    layer2_outputs(84) <= b and not a;
    layer2_outputs(85) <= not (a or b);
    layer2_outputs(86) <= 1'b0;
    layer2_outputs(87) <= not b;
    layer2_outputs(88) <= b and not a;
    layer2_outputs(89) <= b;
    layer2_outputs(90) <= a and b;
    layer2_outputs(91) <= not b;
    layer2_outputs(92) <= not a;
    layer2_outputs(93) <= not (a and b);
    layer2_outputs(94) <= 1'b1;
    layer2_outputs(95) <= a;
    layer2_outputs(96) <= 1'b0;
    layer2_outputs(97) <= a xor b;
    layer2_outputs(98) <= a and b;
    layer2_outputs(99) <= not a or b;
    layer2_outputs(100) <= 1'b1;
    layer2_outputs(101) <= not (a and b);
    layer2_outputs(102) <= not b or a;
    layer2_outputs(103) <= not b;
    layer2_outputs(104) <= not (a and b);
    layer2_outputs(105) <= 1'b0;
    layer2_outputs(106) <= not b or a;
    layer2_outputs(107) <= not (a xor b);
    layer2_outputs(108) <= 1'b1;
    layer2_outputs(109) <= 1'b1;
    layer2_outputs(110) <= 1'b1;
    layer2_outputs(111) <= a and not b;
    layer2_outputs(112) <= not (a xor b);
    layer2_outputs(113) <= not (a and b);
    layer2_outputs(114) <= not a or b;
    layer2_outputs(115) <= not (a and b);
    layer2_outputs(116) <= not (a xor b);
    layer2_outputs(117) <= a xor b;
    layer2_outputs(118) <= 1'b0;
    layer2_outputs(119) <= a xor b;
    layer2_outputs(120) <= not (a or b);
    layer2_outputs(121) <= b and not a;
    layer2_outputs(122) <= a and b;
    layer2_outputs(123) <= a;
    layer2_outputs(124) <= b;
    layer2_outputs(125) <= a;
    layer2_outputs(126) <= a or b;
    layer2_outputs(127) <= a and not b;
    layer2_outputs(128) <= 1'b1;
    layer2_outputs(129) <= not b;
    layer2_outputs(130) <= a;
    layer2_outputs(131) <= not b;
    layer2_outputs(132) <= b;
    layer2_outputs(133) <= not a;
    layer2_outputs(134) <= b;
    layer2_outputs(135) <= not (a or b);
    layer2_outputs(136) <= b and not a;
    layer2_outputs(137) <= not b;
    layer2_outputs(138) <= not (a and b);
    layer2_outputs(139) <= b and not a;
    layer2_outputs(140) <= not b;
    layer2_outputs(141) <= not (a or b);
    layer2_outputs(142) <= 1'b1;
    layer2_outputs(143) <= not (a and b);
    layer2_outputs(144) <= 1'b1;
    layer2_outputs(145) <= 1'b0;
    layer2_outputs(146) <= not (a xor b);
    layer2_outputs(147) <= 1'b1;
    layer2_outputs(148) <= a and b;
    layer2_outputs(149) <= a and not b;
    layer2_outputs(150) <= not (a or b);
    layer2_outputs(151) <= 1'b1;
    layer2_outputs(152) <= b;
    layer2_outputs(153) <= 1'b1;
    layer2_outputs(154) <= 1'b1;
    layer2_outputs(155) <= 1'b0;
    layer2_outputs(156) <= not (a and b);
    layer2_outputs(157) <= 1'b0;
    layer2_outputs(158) <= a and b;
    layer2_outputs(159) <= 1'b0;
    layer2_outputs(160) <= not a;
    layer2_outputs(161) <= not a or b;
    layer2_outputs(162) <= b and not a;
    layer2_outputs(163) <= 1'b0;
    layer2_outputs(164) <= not (a and b);
    layer2_outputs(165) <= a xor b;
    layer2_outputs(166) <= not (a or b);
    layer2_outputs(167) <= not (a or b);
    layer2_outputs(168) <= 1'b0;
    layer2_outputs(169) <= b and not a;
    layer2_outputs(170) <= not a or b;
    layer2_outputs(171) <= not a;
    layer2_outputs(172) <= not (a and b);
    layer2_outputs(173) <= 1'b1;
    layer2_outputs(174) <= a and not b;
    layer2_outputs(175) <= not b or a;
    layer2_outputs(176) <= a and b;
    layer2_outputs(177) <= b and not a;
    layer2_outputs(178) <= a and b;
    layer2_outputs(179) <= not (a and b);
    layer2_outputs(180) <= a or b;
    layer2_outputs(181) <= not b or a;
    layer2_outputs(182) <= not a or b;
    layer2_outputs(183) <= 1'b1;
    layer2_outputs(184) <= 1'b1;
    layer2_outputs(185) <= not (a xor b);
    layer2_outputs(186) <= 1'b0;
    layer2_outputs(187) <= not b or a;
    layer2_outputs(188) <= a and not b;
    layer2_outputs(189) <= 1'b0;
    layer2_outputs(190) <= 1'b1;
    layer2_outputs(191) <= a or b;
    layer2_outputs(192) <= not (a or b);
    layer2_outputs(193) <= b;
    layer2_outputs(194) <= not a;
    layer2_outputs(195) <= a and not b;
    layer2_outputs(196) <= not (a and b);
    layer2_outputs(197) <= a and not b;
    layer2_outputs(198) <= b;
    layer2_outputs(199) <= 1'b0;
    layer2_outputs(200) <= a and b;
    layer2_outputs(201) <= a and b;
    layer2_outputs(202) <= b;
    layer2_outputs(203) <= a and not b;
    layer2_outputs(204) <= b and not a;
    layer2_outputs(205) <= a and b;
    layer2_outputs(206) <= not (a and b);
    layer2_outputs(207) <= not b;
    layer2_outputs(208) <= a and b;
    layer2_outputs(209) <= a and not b;
    layer2_outputs(210) <= 1'b1;
    layer2_outputs(211) <= a or b;
    layer2_outputs(212) <= 1'b1;
    layer2_outputs(213) <= a and not b;
    layer2_outputs(214) <= a and not b;
    layer2_outputs(215) <= not b;
    layer2_outputs(216) <= a;
    layer2_outputs(217) <= not b or a;
    layer2_outputs(218) <= 1'b1;
    layer2_outputs(219) <= 1'b1;
    layer2_outputs(220) <= not (a or b);
    layer2_outputs(221) <= not a or b;
    layer2_outputs(222) <= b and not a;
    layer2_outputs(223) <= not (a or b);
    layer2_outputs(224) <= not (a xor b);
    layer2_outputs(225) <= a;
    layer2_outputs(226) <= not (a or b);
    layer2_outputs(227) <= not a or b;
    layer2_outputs(228) <= not (a or b);
    layer2_outputs(229) <= a and not b;
    layer2_outputs(230) <= not b;
    layer2_outputs(231) <= 1'b1;
    layer2_outputs(232) <= a and b;
    layer2_outputs(233) <= a and b;
    layer2_outputs(234) <= b and not a;
    layer2_outputs(235) <= a;
    layer2_outputs(236) <= a or b;
    layer2_outputs(237) <= not b or a;
    layer2_outputs(238) <= a xor b;
    layer2_outputs(239) <= a and b;
    layer2_outputs(240) <= a;
    layer2_outputs(241) <= 1'b0;
    layer2_outputs(242) <= a and not b;
    layer2_outputs(243) <= not (a xor b);
    layer2_outputs(244) <= not b;
    layer2_outputs(245) <= b and not a;
    layer2_outputs(246) <= b;
    layer2_outputs(247) <= not a;
    layer2_outputs(248) <= 1'b1;
    layer2_outputs(249) <= a or b;
    layer2_outputs(250) <= not b;
    layer2_outputs(251) <= b;
    layer2_outputs(252) <= not b;
    layer2_outputs(253) <= a or b;
    layer2_outputs(254) <= not b or a;
    layer2_outputs(255) <= not (a and b);
    layer2_outputs(256) <= a;
    layer2_outputs(257) <= a and not b;
    layer2_outputs(258) <= not b or a;
    layer2_outputs(259) <= 1'b1;
    layer2_outputs(260) <= b;
    layer2_outputs(261) <= a and b;
    layer2_outputs(262) <= b;
    layer2_outputs(263) <= b and not a;
    layer2_outputs(264) <= 1'b0;
    layer2_outputs(265) <= not b or a;
    layer2_outputs(266) <= a;
    layer2_outputs(267) <= a;
    layer2_outputs(268) <= not a;
    layer2_outputs(269) <= b;
    layer2_outputs(270) <= 1'b0;
    layer2_outputs(271) <= a and b;
    layer2_outputs(272) <= not (a and b);
    layer2_outputs(273) <= b;
    layer2_outputs(274) <= not (a xor b);
    layer2_outputs(275) <= 1'b0;
    layer2_outputs(276) <= a and not b;
    layer2_outputs(277) <= not b;
    layer2_outputs(278) <= a and not b;
    layer2_outputs(279) <= not (a or b);
    layer2_outputs(280) <= a;
    layer2_outputs(281) <= a and b;
    layer2_outputs(282) <= b and not a;
    layer2_outputs(283) <= a and not b;
    layer2_outputs(284) <= not a;
    layer2_outputs(285) <= b and not a;
    layer2_outputs(286) <= a or b;
    layer2_outputs(287) <= a and b;
    layer2_outputs(288) <= a and b;
    layer2_outputs(289) <= b;
    layer2_outputs(290) <= 1'b1;
    layer2_outputs(291) <= a xor b;
    layer2_outputs(292) <= a;
    layer2_outputs(293) <= a and not b;
    layer2_outputs(294) <= not (a and b);
    layer2_outputs(295) <= b and not a;
    layer2_outputs(296) <= a;
    layer2_outputs(297) <= not (a or b);
    layer2_outputs(298) <= not (a xor b);
    layer2_outputs(299) <= a and not b;
    layer2_outputs(300) <= 1'b0;
    layer2_outputs(301) <= not b;
    layer2_outputs(302) <= a;
    layer2_outputs(303) <= 1'b0;
    layer2_outputs(304) <= b and not a;
    layer2_outputs(305) <= not a or b;
    layer2_outputs(306) <= not a or b;
    layer2_outputs(307) <= 1'b0;
    layer2_outputs(308) <= b;
    layer2_outputs(309) <= not b;
    layer2_outputs(310) <= not b or a;
    layer2_outputs(311) <= not (a and b);
    layer2_outputs(312) <= not (a xor b);
    layer2_outputs(313) <= not a or b;
    layer2_outputs(314) <= not b;
    layer2_outputs(315) <= 1'b0;
    layer2_outputs(316) <= a and not b;
    layer2_outputs(317) <= a and b;
    layer2_outputs(318) <= 1'b1;
    layer2_outputs(319) <= a and b;
    layer2_outputs(320) <= not a or b;
    layer2_outputs(321) <= not a;
    layer2_outputs(322) <= a or b;
    layer2_outputs(323) <= a and b;
    layer2_outputs(324) <= not a or b;
    layer2_outputs(325) <= not a;
    layer2_outputs(326) <= a and b;
    layer2_outputs(327) <= not (a and b);
    layer2_outputs(328) <= a;
    layer2_outputs(329) <= not (a and b);
    layer2_outputs(330) <= a;
    layer2_outputs(331) <= a xor b;
    layer2_outputs(332) <= not b or a;
    layer2_outputs(333) <= not (a or b);
    layer2_outputs(334) <= not (a or b);
    layer2_outputs(335) <= not a or b;
    layer2_outputs(336) <= not (a or b);
    layer2_outputs(337) <= a or b;
    layer2_outputs(338) <= not (a xor b);
    layer2_outputs(339) <= not (a and b);
    layer2_outputs(340) <= not a;
    layer2_outputs(341) <= not a;
    layer2_outputs(342) <= 1'b1;
    layer2_outputs(343) <= 1'b0;
    layer2_outputs(344) <= 1'b1;
    layer2_outputs(345) <= 1'b1;
    layer2_outputs(346) <= a and b;
    layer2_outputs(347) <= 1'b0;
    layer2_outputs(348) <= not (a xor b);
    layer2_outputs(349) <= b;
    layer2_outputs(350) <= 1'b0;
    layer2_outputs(351) <= b and not a;
    layer2_outputs(352) <= a xor b;
    layer2_outputs(353) <= a;
    layer2_outputs(354) <= not b;
    layer2_outputs(355) <= not a or b;
    layer2_outputs(356) <= not a;
    layer2_outputs(357) <= b and not a;
    layer2_outputs(358) <= not b;
    layer2_outputs(359) <= 1'b0;
    layer2_outputs(360) <= 1'b0;
    layer2_outputs(361) <= not a;
    layer2_outputs(362) <= not (a and b);
    layer2_outputs(363) <= not (a or b);
    layer2_outputs(364) <= b;
    layer2_outputs(365) <= not b or a;
    layer2_outputs(366) <= not a;
    layer2_outputs(367) <= 1'b0;
    layer2_outputs(368) <= not (a and b);
    layer2_outputs(369) <= not (a or b);
    layer2_outputs(370) <= not b or a;
    layer2_outputs(371) <= a and b;
    layer2_outputs(372) <= not a or b;
    layer2_outputs(373) <= a and b;
    layer2_outputs(374) <= a and not b;
    layer2_outputs(375) <= 1'b1;
    layer2_outputs(376) <= a;
    layer2_outputs(377) <= not (a and b);
    layer2_outputs(378) <= not (a and b);
    layer2_outputs(379) <= a and b;
    layer2_outputs(380) <= not a;
    layer2_outputs(381) <= not b;
    layer2_outputs(382) <= 1'b1;
    layer2_outputs(383) <= a and b;
    layer2_outputs(384) <= not (a and b);
    layer2_outputs(385) <= a or b;
    layer2_outputs(386) <= not (a and b);
    layer2_outputs(387) <= not a;
    layer2_outputs(388) <= b and not a;
    layer2_outputs(389) <= not b or a;
    layer2_outputs(390) <= a and not b;
    layer2_outputs(391) <= a xor b;
    layer2_outputs(392) <= not a or b;
    layer2_outputs(393) <= not (a and b);
    layer2_outputs(394) <= not (a or b);
    layer2_outputs(395) <= not b or a;
    layer2_outputs(396) <= not a or b;
    layer2_outputs(397) <= not (a and b);
    layer2_outputs(398) <= not (a and b);
    layer2_outputs(399) <= not (a and b);
    layer2_outputs(400) <= 1'b1;
    layer2_outputs(401) <= a or b;
    layer2_outputs(402) <= a;
    layer2_outputs(403) <= b;
    layer2_outputs(404) <= b and not a;
    layer2_outputs(405) <= not a or b;
    layer2_outputs(406) <= not a;
    layer2_outputs(407) <= not b;
    layer2_outputs(408) <= 1'b1;
    layer2_outputs(409) <= not a or b;
    layer2_outputs(410) <= a or b;
    layer2_outputs(411) <= a and b;
    layer2_outputs(412) <= a and not b;
    layer2_outputs(413) <= 1'b0;
    layer2_outputs(414) <= not a;
    layer2_outputs(415) <= not (a or b);
    layer2_outputs(416) <= a;
    layer2_outputs(417) <= a or b;
    layer2_outputs(418) <= 1'b0;
    layer2_outputs(419) <= not (a and b);
    layer2_outputs(420) <= not b or a;
    layer2_outputs(421) <= not a;
    layer2_outputs(422) <= not a or b;
    layer2_outputs(423) <= a or b;
    layer2_outputs(424) <= 1'b1;
    layer2_outputs(425) <= not (a or b);
    layer2_outputs(426) <= 1'b0;
    layer2_outputs(427) <= not (a and b);
    layer2_outputs(428) <= not (a and b);
    layer2_outputs(429) <= not b;
    layer2_outputs(430) <= not a or b;
    layer2_outputs(431) <= not b;
    layer2_outputs(432) <= a and not b;
    layer2_outputs(433) <= a and not b;
    layer2_outputs(434) <= a;
    layer2_outputs(435) <= a xor b;
    layer2_outputs(436) <= not a or b;
    layer2_outputs(437) <= not (a and b);
    layer2_outputs(438) <= a;
    layer2_outputs(439) <= b and not a;
    layer2_outputs(440) <= not (a xor b);
    layer2_outputs(441) <= b;
    layer2_outputs(442) <= not a or b;
    layer2_outputs(443) <= not b or a;
    layer2_outputs(444) <= a or b;
    layer2_outputs(445) <= 1'b0;
    layer2_outputs(446) <= not (a or b);
    layer2_outputs(447) <= a;
    layer2_outputs(448) <= not (a xor b);
    layer2_outputs(449) <= 1'b1;
    layer2_outputs(450) <= not (a or b);
    layer2_outputs(451) <= a;
    layer2_outputs(452) <= not (a or b);
    layer2_outputs(453) <= not b or a;
    layer2_outputs(454) <= not b or a;
    layer2_outputs(455) <= 1'b0;
    layer2_outputs(456) <= a and b;
    layer2_outputs(457) <= not (a and b);
    layer2_outputs(458) <= a;
    layer2_outputs(459) <= not b;
    layer2_outputs(460) <= b;
    layer2_outputs(461) <= a and not b;
    layer2_outputs(462) <= 1'b0;
    layer2_outputs(463) <= 1'b0;
    layer2_outputs(464) <= a and b;
    layer2_outputs(465) <= not (a or b);
    layer2_outputs(466) <= not b;
    layer2_outputs(467) <= not (a or b);
    layer2_outputs(468) <= a and not b;
    layer2_outputs(469) <= b and not a;
    layer2_outputs(470) <= a;
    layer2_outputs(471) <= 1'b1;
    layer2_outputs(472) <= a;
    layer2_outputs(473) <= b and not a;
    layer2_outputs(474) <= not (a or b);
    layer2_outputs(475) <= a and not b;
    layer2_outputs(476) <= b and not a;
    layer2_outputs(477) <= a xor b;
    layer2_outputs(478) <= not (a or b);
    layer2_outputs(479) <= not (a and b);
    layer2_outputs(480) <= 1'b1;
    layer2_outputs(481) <= not b or a;
    layer2_outputs(482) <= b;
    layer2_outputs(483) <= 1'b1;
    layer2_outputs(484) <= b;
    layer2_outputs(485) <= a;
    layer2_outputs(486) <= b;
    layer2_outputs(487) <= not (a or b);
    layer2_outputs(488) <= a and b;
    layer2_outputs(489) <= 1'b1;
    layer2_outputs(490) <= not (a or b);
    layer2_outputs(491) <= 1'b0;
    layer2_outputs(492) <= b and not a;
    layer2_outputs(493) <= not b;
    layer2_outputs(494) <= not a or b;
    layer2_outputs(495) <= not a or b;
    layer2_outputs(496) <= a and not b;
    layer2_outputs(497) <= 1'b0;
    layer2_outputs(498) <= a;
    layer2_outputs(499) <= 1'b1;
    layer2_outputs(500) <= not (a xor b);
    layer2_outputs(501) <= a;
    layer2_outputs(502) <= a or b;
    layer2_outputs(503) <= 1'b0;
    layer2_outputs(504) <= a and not b;
    layer2_outputs(505) <= a or b;
    layer2_outputs(506) <= a or b;
    layer2_outputs(507) <= 1'b1;
    layer2_outputs(508) <= a and not b;
    layer2_outputs(509) <= not (a and b);
    layer2_outputs(510) <= not b or a;
    layer2_outputs(511) <= b and not a;
    layer2_outputs(512) <= not b or a;
    layer2_outputs(513) <= not (a and b);
    layer2_outputs(514) <= 1'b0;
    layer2_outputs(515) <= 1'b0;
    layer2_outputs(516) <= 1'b0;
    layer2_outputs(517) <= b and not a;
    layer2_outputs(518) <= not b or a;
    layer2_outputs(519) <= not a or b;
    layer2_outputs(520) <= not a or b;
    layer2_outputs(521) <= 1'b1;
    layer2_outputs(522) <= not a;
    layer2_outputs(523) <= a;
    layer2_outputs(524) <= b;
    layer2_outputs(525) <= a and not b;
    layer2_outputs(526) <= not (a or b);
    layer2_outputs(527) <= a or b;
    layer2_outputs(528) <= a;
    layer2_outputs(529) <= not (a or b);
    layer2_outputs(530) <= a;
    layer2_outputs(531) <= 1'b1;
    layer2_outputs(532) <= not b or a;
    layer2_outputs(533) <= not a or b;
    layer2_outputs(534) <= 1'b0;
    layer2_outputs(535) <= not (a or b);
    layer2_outputs(536) <= 1'b1;
    layer2_outputs(537) <= a or b;
    layer2_outputs(538) <= not b;
    layer2_outputs(539) <= 1'b0;
    layer2_outputs(540) <= b;
    layer2_outputs(541) <= 1'b1;
    layer2_outputs(542) <= not b;
    layer2_outputs(543) <= a and not b;
    layer2_outputs(544) <= b and not a;
    layer2_outputs(545) <= not a or b;
    layer2_outputs(546) <= a and not b;
    layer2_outputs(547) <= a and not b;
    layer2_outputs(548) <= 1'b1;
    layer2_outputs(549) <= not a or b;
    layer2_outputs(550) <= a xor b;
    layer2_outputs(551) <= a and not b;
    layer2_outputs(552) <= 1'b0;
    layer2_outputs(553) <= a and not b;
    layer2_outputs(554) <= a or b;
    layer2_outputs(555) <= not b or a;
    layer2_outputs(556) <= not a or b;
    layer2_outputs(557) <= a and b;
    layer2_outputs(558) <= b;
    layer2_outputs(559) <= b and not a;
    layer2_outputs(560) <= a;
    layer2_outputs(561) <= 1'b1;
    layer2_outputs(562) <= b;
    layer2_outputs(563) <= not a;
    layer2_outputs(564) <= a or b;
    layer2_outputs(565) <= not a or b;
    layer2_outputs(566) <= not a or b;
    layer2_outputs(567) <= not a or b;
    layer2_outputs(568) <= a and not b;
    layer2_outputs(569) <= 1'b1;
    layer2_outputs(570) <= not (a and b);
    layer2_outputs(571) <= a and not b;
    layer2_outputs(572) <= b;
    layer2_outputs(573) <= a;
    layer2_outputs(574) <= not b;
    layer2_outputs(575) <= a or b;
    layer2_outputs(576) <= b;
    layer2_outputs(577) <= 1'b1;
    layer2_outputs(578) <= a xor b;
    layer2_outputs(579) <= 1'b0;
    layer2_outputs(580) <= not (a or b);
    layer2_outputs(581) <= not b or a;
    layer2_outputs(582) <= not a;
    layer2_outputs(583) <= not a;
    layer2_outputs(584) <= not (a or b);
    layer2_outputs(585) <= not a or b;
    layer2_outputs(586) <= not b;
    layer2_outputs(587) <= a and b;
    layer2_outputs(588) <= 1'b0;
    layer2_outputs(589) <= a and b;
    layer2_outputs(590) <= not a or b;
    layer2_outputs(591) <= 1'b0;
    layer2_outputs(592) <= 1'b0;
    layer2_outputs(593) <= a;
    layer2_outputs(594) <= a and b;
    layer2_outputs(595) <= b;
    layer2_outputs(596) <= b;
    layer2_outputs(597) <= a and not b;
    layer2_outputs(598) <= a;
    layer2_outputs(599) <= a and b;
    layer2_outputs(600) <= a and b;
    layer2_outputs(601) <= not b;
    layer2_outputs(602) <= not (a xor b);
    layer2_outputs(603) <= not b;
    layer2_outputs(604) <= not b or a;
    layer2_outputs(605) <= not (a xor b);
    layer2_outputs(606) <= not (a xor b);
    layer2_outputs(607) <= 1'b1;
    layer2_outputs(608) <= 1'b0;
    layer2_outputs(609) <= 1'b0;
    layer2_outputs(610) <= not a or b;
    layer2_outputs(611) <= b;
    layer2_outputs(612) <= not (a and b);
    layer2_outputs(613) <= a and not b;
    layer2_outputs(614) <= 1'b1;
    layer2_outputs(615) <= 1'b0;
    layer2_outputs(616) <= 1'b0;
    layer2_outputs(617) <= not (a and b);
    layer2_outputs(618) <= a;
    layer2_outputs(619) <= b and not a;
    layer2_outputs(620) <= not a or b;
    layer2_outputs(621) <= 1'b0;
    layer2_outputs(622) <= not b or a;
    layer2_outputs(623) <= not a or b;
    layer2_outputs(624) <= not a or b;
    layer2_outputs(625) <= 1'b0;
    layer2_outputs(626) <= not a or b;
    layer2_outputs(627) <= a and b;
    layer2_outputs(628) <= not b or a;
    layer2_outputs(629) <= a xor b;
    layer2_outputs(630) <= 1'b0;
    layer2_outputs(631) <= not (a or b);
    layer2_outputs(632) <= not b or a;
    layer2_outputs(633) <= b;
    layer2_outputs(634) <= a and b;
    layer2_outputs(635) <= not a or b;
    layer2_outputs(636) <= a and not b;
    layer2_outputs(637) <= not a or b;
    layer2_outputs(638) <= b and not a;
    layer2_outputs(639) <= not b or a;
    layer2_outputs(640) <= not (a or b);
    layer2_outputs(641) <= a or b;
    layer2_outputs(642) <= not (a xor b);
    layer2_outputs(643) <= b;
    layer2_outputs(644) <= not a;
    layer2_outputs(645) <= 1'b0;
    layer2_outputs(646) <= not a or b;
    layer2_outputs(647) <= not a;
    layer2_outputs(648) <= not b or a;
    layer2_outputs(649) <= not a or b;
    layer2_outputs(650) <= a and b;
    layer2_outputs(651) <= b and not a;
    layer2_outputs(652) <= not (a and b);
    layer2_outputs(653) <= a and b;
    layer2_outputs(654) <= b and not a;
    layer2_outputs(655) <= not (a or b);
    layer2_outputs(656) <= not a or b;
    layer2_outputs(657) <= b and not a;
    layer2_outputs(658) <= a and b;
    layer2_outputs(659) <= a;
    layer2_outputs(660) <= not a or b;
    layer2_outputs(661) <= not b;
    layer2_outputs(662) <= 1'b1;
    layer2_outputs(663) <= a and not b;
    layer2_outputs(664) <= 1'b1;
    layer2_outputs(665) <= b and not a;
    layer2_outputs(666) <= a and b;
    layer2_outputs(667) <= not (a and b);
    layer2_outputs(668) <= a;
    layer2_outputs(669) <= a and not b;
    layer2_outputs(670) <= a and b;
    layer2_outputs(671) <= 1'b1;
    layer2_outputs(672) <= b and not a;
    layer2_outputs(673) <= 1'b1;
    layer2_outputs(674) <= a;
    layer2_outputs(675) <= a;
    layer2_outputs(676) <= not (a or b);
    layer2_outputs(677) <= a or b;
    layer2_outputs(678) <= 1'b0;
    layer2_outputs(679) <= not (a or b);
    layer2_outputs(680) <= not b or a;
    layer2_outputs(681) <= not a or b;
    layer2_outputs(682) <= 1'b1;
    layer2_outputs(683) <= b and not a;
    layer2_outputs(684) <= a or b;
    layer2_outputs(685) <= not b or a;
    layer2_outputs(686) <= not a;
    layer2_outputs(687) <= not a;
    layer2_outputs(688) <= 1'b1;
    layer2_outputs(689) <= not (a xor b);
    layer2_outputs(690) <= not a;
    layer2_outputs(691) <= 1'b1;
    layer2_outputs(692) <= not a or b;
    layer2_outputs(693) <= b and not a;
    layer2_outputs(694) <= a;
    layer2_outputs(695) <= not a or b;
    layer2_outputs(696) <= not (a or b);
    layer2_outputs(697) <= not a or b;
    layer2_outputs(698) <= a and not b;
    layer2_outputs(699) <= a xor b;
    layer2_outputs(700) <= 1'b0;
    layer2_outputs(701) <= not b;
    layer2_outputs(702) <= not (a or b);
    layer2_outputs(703) <= 1'b1;
    layer2_outputs(704) <= not (a or b);
    layer2_outputs(705) <= a xor b;
    layer2_outputs(706) <= a and not b;
    layer2_outputs(707) <= a xor b;
    layer2_outputs(708) <= 1'b1;
    layer2_outputs(709) <= a and b;
    layer2_outputs(710) <= a and b;
    layer2_outputs(711) <= not a;
    layer2_outputs(712) <= a or b;
    layer2_outputs(713) <= a and not b;
    layer2_outputs(714) <= 1'b0;
    layer2_outputs(715) <= 1'b1;
    layer2_outputs(716) <= b;
    layer2_outputs(717) <= not (a xor b);
    layer2_outputs(718) <= not a or b;
    layer2_outputs(719) <= not (a and b);
    layer2_outputs(720) <= b;
    layer2_outputs(721) <= not a;
    layer2_outputs(722) <= not (a or b);
    layer2_outputs(723) <= not b or a;
    layer2_outputs(724) <= b;
    layer2_outputs(725) <= a and not b;
    layer2_outputs(726) <= a;
    layer2_outputs(727) <= 1'b0;
    layer2_outputs(728) <= b and not a;
    layer2_outputs(729) <= a or b;
    layer2_outputs(730) <= not b or a;
    layer2_outputs(731) <= a or b;
    layer2_outputs(732) <= a;
    layer2_outputs(733) <= a;
    layer2_outputs(734) <= not b or a;
    layer2_outputs(735) <= not b or a;
    layer2_outputs(736) <= 1'b0;
    layer2_outputs(737) <= b;
    layer2_outputs(738) <= a or b;
    layer2_outputs(739) <= not b;
    layer2_outputs(740) <= b;
    layer2_outputs(741) <= not (a or b);
    layer2_outputs(742) <= not (a or b);
    layer2_outputs(743) <= not (a and b);
    layer2_outputs(744) <= not (a and b);
    layer2_outputs(745) <= b and not a;
    layer2_outputs(746) <= 1'b1;
    layer2_outputs(747) <= 1'b1;
    layer2_outputs(748) <= b;
    layer2_outputs(749) <= a;
    layer2_outputs(750) <= a and not b;
    layer2_outputs(751) <= not (a or b);
    layer2_outputs(752) <= b and not a;
    layer2_outputs(753) <= a and not b;
    layer2_outputs(754) <= a and not b;
    layer2_outputs(755) <= not b;
    layer2_outputs(756) <= not b or a;
    layer2_outputs(757) <= a and b;
    layer2_outputs(758) <= a and not b;
    layer2_outputs(759) <= a;
    layer2_outputs(760) <= a xor b;
    layer2_outputs(761) <= not b;
    layer2_outputs(762) <= not (a or b);
    layer2_outputs(763) <= not (a and b);
    layer2_outputs(764) <= not a or b;
    layer2_outputs(765) <= not (a and b);
    layer2_outputs(766) <= a and not b;
    layer2_outputs(767) <= 1'b1;
    layer2_outputs(768) <= b;
    layer2_outputs(769) <= not b;
    layer2_outputs(770) <= b and not a;
    layer2_outputs(771) <= b and not a;
    layer2_outputs(772) <= a and not b;
    layer2_outputs(773) <= not (a and b);
    layer2_outputs(774) <= 1'b1;
    layer2_outputs(775) <= not b or a;
    layer2_outputs(776) <= not (a or b);
    layer2_outputs(777) <= b and not a;
    layer2_outputs(778) <= 1'b1;
    layer2_outputs(779) <= not a;
    layer2_outputs(780) <= not b or a;
    layer2_outputs(781) <= 1'b0;
    layer2_outputs(782) <= 1'b1;
    layer2_outputs(783) <= 1'b1;
    layer2_outputs(784) <= a;
    layer2_outputs(785) <= a;
    layer2_outputs(786) <= a and not b;
    layer2_outputs(787) <= not b or a;
    layer2_outputs(788) <= not (a and b);
    layer2_outputs(789) <= not b;
    layer2_outputs(790) <= a and not b;
    layer2_outputs(791) <= a or b;
    layer2_outputs(792) <= not (a and b);
    layer2_outputs(793) <= a xor b;
    layer2_outputs(794) <= not (a or b);
    layer2_outputs(795) <= a xor b;
    layer2_outputs(796) <= not (a and b);
    layer2_outputs(797) <= a and not b;
    layer2_outputs(798) <= a and not b;
    layer2_outputs(799) <= not b or a;
    layer2_outputs(800) <= a and not b;
    layer2_outputs(801) <= not (a or b);
    layer2_outputs(802) <= not b or a;
    layer2_outputs(803) <= 1'b1;
    layer2_outputs(804) <= 1'b0;
    layer2_outputs(805) <= not (a or b);
    layer2_outputs(806) <= a and not b;
    layer2_outputs(807) <= not (a or b);
    layer2_outputs(808) <= b;
    layer2_outputs(809) <= a and not b;
    layer2_outputs(810) <= a or b;
    layer2_outputs(811) <= 1'b0;
    layer2_outputs(812) <= 1'b1;
    layer2_outputs(813) <= b and not a;
    layer2_outputs(814) <= b;
    layer2_outputs(815) <= a and b;
    layer2_outputs(816) <= a and not b;
    layer2_outputs(817) <= b and not a;
    layer2_outputs(818) <= a and b;
    layer2_outputs(819) <= a and b;
    layer2_outputs(820) <= a and not b;
    layer2_outputs(821) <= not b or a;
    layer2_outputs(822) <= b and not a;
    layer2_outputs(823) <= not (a or b);
    layer2_outputs(824) <= 1'b0;
    layer2_outputs(825) <= a and b;
    layer2_outputs(826) <= a and b;
    layer2_outputs(827) <= a and b;
    layer2_outputs(828) <= a and not b;
    layer2_outputs(829) <= a and b;
    layer2_outputs(830) <= a and b;
    layer2_outputs(831) <= a and not b;
    layer2_outputs(832) <= not (a or b);
    layer2_outputs(833) <= a and b;
    layer2_outputs(834) <= not a or b;
    layer2_outputs(835) <= 1'b0;
    layer2_outputs(836) <= not b;
    layer2_outputs(837) <= not a;
    layer2_outputs(838) <= 1'b0;
    layer2_outputs(839) <= a or b;
    layer2_outputs(840) <= not (a or b);
    layer2_outputs(841) <= not (a or b);
    layer2_outputs(842) <= a and not b;
    layer2_outputs(843) <= 1'b1;
    layer2_outputs(844) <= not a or b;
    layer2_outputs(845) <= 1'b1;
    layer2_outputs(846) <= a and not b;
    layer2_outputs(847) <= b and not a;
    layer2_outputs(848) <= 1'b1;
    layer2_outputs(849) <= a;
    layer2_outputs(850) <= not a or b;
    layer2_outputs(851) <= not (a and b);
    layer2_outputs(852) <= b;
    layer2_outputs(853) <= not a or b;
    layer2_outputs(854) <= b and not a;
    layer2_outputs(855) <= not a;
    layer2_outputs(856) <= not a or b;
    layer2_outputs(857) <= not b;
    layer2_outputs(858) <= not b;
    layer2_outputs(859) <= b;
    layer2_outputs(860) <= not (a or b);
    layer2_outputs(861) <= a and b;
    layer2_outputs(862) <= not a;
    layer2_outputs(863) <= 1'b1;
    layer2_outputs(864) <= 1'b1;
    layer2_outputs(865) <= 1'b0;
    layer2_outputs(866) <= b and not a;
    layer2_outputs(867) <= 1'b1;
    layer2_outputs(868) <= not b or a;
    layer2_outputs(869) <= not a;
    layer2_outputs(870) <= 1'b1;
    layer2_outputs(871) <= 1'b0;
    layer2_outputs(872) <= not a or b;
    layer2_outputs(873) <= a and not b;
    layer2_outputs(874) <= not (a and b);
    layer2_outputs(875) <= 1'b1;
    layer2_outputs(876) <= a or b;
    layer2_outputs(877) <= a and not b;
    layer2_outputs(878) <= not (a xor b);
    layer2_outputs(879) <= not b;
    layer2_outputs(880) <= 1'b1;
    layer2_outputs(881) <= not (a and b);
    layer2_outputs(882) <= a and not b;
    layer2_outputs(883) <= a or b;
    layer2_outputs(884) <= not (a or b);
    layer2_outputs(885) <= not b or a;
    layer2_outputs(886) <= not b;
    layer2_outputs(887) <= a or b;
    layer2_outputs(888) <= a and not b;
    layer2_outputs(889) <= b;
    layer2_outputs(890) <= a;
    layer2_outputs(891) <= not a or b;
    layer2_outputs(892) <= 1'b1;
    layer2_outputs(893) <= b;
    layer2_outputs(894) <= a xor b;
    layer2_outputs(895) <= not b or a;
    layer2_outputs(896) <= not a or b;
    layer2_outputs(897) <= not (a or b);
    layer2_outputs(898) <= not (a or b);
    layer2_outputs(899) <= b and not a;
    layer2_outputs(900) <= not b;
    layer2_outputs(901) <= a and b;
    layer2_outputs(902) <= not a or b;
    layer2_outputs(903) <= b and not a;
    layer2_outputs(904) <= not a or b;
    layer2_outputs(905) <= b and not a;
    layer2_outputs(906) <= not (a or b);
    layer2_outputs(907) <= not a or b;
    layer2_outputs(908) <= not a or b;
    layer2_outputs(909) <= not b or a;
    layer2_outputs(910) <= 1'b0;
    layer2_outputs(911) <= 1'b1;
    layer2_outputs(912) <= not a or b;
    layer2_outputs(913) <= a and b;
    layer2_outputs(914) <= a and not b;
    layer2_outputs(915) <= a;
    layer2_outputs(916) <= not b;
    layer2_outputs(917) <= a and b;
    layer2_outputs(918) <= a and not b;
    layer2_outputs(919) <= a and not b;
    layer2_outputs(920) <= not b;
    layer2_outputs(921) <= a or b;
    layer2_outputs(922) <= not b or a;
    layer2_outputs(923) <= a xor b;
    layer2_outputs(924) <= a xor b;
    layer2_outputs(925) <= 1'b0;
    layer2_outputs(926) <= not (a xor b);
    layer2_outputs(927) <= not (a and b);
    layer2_outputs(928) <= not b;
    layer2_outputs(929) <= not (a and b);
    layer2_outputs(930) <= b;
    layer2_outputs(931) <= not a or b;
    layer2_outputs(932) <= 1'b0;
    layer2_outputs(933) <= a and not b;
    layer2_outputs(934) <= not a;
    layer2_outputs(935) <= b and not a;
    layer2_outputs(936) <= 1'b0;
    layer2_outputs(937) <= a and b;
    layer2_outputs(938) <= not b;
    layer2_outputs(939) <= a and not b;
    layer2_outputs(940) <= a or b;
    layer2_outputs(941) <= not a;
    layer2_outputs(942) <= not b or a;
    layer2_outputs(943) <= a and b;
    layer2_outputs(944) <= not (a or b);
    layer2_outputs(945) <= b;
    layer2_outputs(946) <= b and not a;
    layer2_outputs(947) <= b;
    layer2_outputs(948) <= not a or b;
    layer2_outputs(949) <= not (a and b);
    layer2_outputs(950) <= 1'b0;
    layer2_outputs(951) <= a;
    layer2_outputs(952) <= not a or b;
    layer2_outputs(953) <= a;
    layer2_outputs(954) <= a;
    layer2_outputs(955) <= a;
    layer2_outputs(956) <= not (a xor b);
    layer2_outputs(957) <= not a or b;
    layer2_outputs(958) <= 1'b1;
    layer2_outputs(959) <= b;
    layer2_outputs(960) <= not (a xor b);
    layer2_outputs(961) <= a or b;
    layer2_outputs(962) <= 1'b0;
    layer2_outputs(963) <= 1'b1;
    layer2_outputs(964) <= a xor b;
    layer2_outputs(965) <= a or b;
    layer2_outputs(966) <= a or b;
    layer2_outputs(967) <= not (a or b);
    layer2_outputs(968) <= a and not b;
    layer2_outputs(969) <= 1'b1;
    layer2_outputs(970) <= b and not a;
    layer2_outputs(971) <= not a or b;
    layer2_outputs(972) <= not (a or b);
    layer2_outputs(973) <= 1'b0;
    layer2_outputs(974) <= a;
    layer2_outputs(975) <= not (a and b);
    layer2_outputs(976) <= 1'b0;
    layer2_outputs(977) <= a or b;
    layer2_outputs(978) <= not (a or b);
    layer2_outputs(979) <= not a;
    layer2_outputs(980) <= not b;
    layer2_outputs(981) <= a and not b;
    layer2_outputs(982) <= a and b;
    layer2_outputs(983) <= 1'b0;
    layer2_outputs(984) <= a;
    layer2_outputs(985) <= a or b;
    layer2_outputs(986) <= not b or a;
    layer2_outputs(987) <= b;
    layer2_outputs(988) <= not b;
    layer2_outputs(989) <= a xor b;
    layer2_outputs(990) <= not b or a;
    layer2_outputs(991) <= not (a and b);
    layer2_outputs(992) <= not a or b;
    layer2_outputs(993) <= not (a and b);
    layer2_outputs(994) <= not b;
    layer2_outputs(995) <= not a;
    layer2_outputs(996) <= not (a and b);
    layer2_outputs(997) <= a and b;
    layer2_outputs(998) <= b and not a;
    layer2_outputs(999) <= b and not a;
    layer2_outputs(1000) <= not (a or b);
    layer2_outputs(1001) <= not b or a;
    layer2_outputs(1002) <= a;
    layer2_outputs(1003) <= not (a and b);
    layer2_outputs(1004) <= b;
    layer2_outputs(1005) <= not b;
    layer2_outputs(1006) <= a;
    layer2_outputs(1007) <= a or b;
    layer2_outputs(1008) <= a;
    layer2_outputs(1009) <= not a or b;
    layer2_outputs(1010) <= 1'b1;
    layer2_outputs(1011) <= 1'b1;
    layer2_outputs(1012) <= b;
    layer2_outputs(1013) <= a and not b;
    layer2_outputs(1014) <= a and not b;
    layer2_outputs(1015) <= b;
    layer2_outputs(1016) <= a xor b;
    layer2_outputs(1017) <= not (a xor b);
    layer2_outputs(1018) <= 1'b0;
    layer2_outputs(1019) <= 1'b0;
    layer2_outputs(1020) <= not b;
    layer2_outputs(1021) <= a;
    layer2_outputs(1022) <= b;
    layer2_outputs(1023) <= 1'b1;
    layer2_outputs(1024) <= 1'b0;
    layer2_outputs(1025) <= 1'b1;
    layer2_outputs(1026) <= a and b;
    layer2_outputs(1027) <= a and not b;
    layer2_outputs(1028) <= not a;
    layer2_outputs(1029) <= not (a xor b);
    layer2_outputs(1030) <= a and b;
    layer2_outputs(1031) <= not b;
    layer2_outputs(1032) <= 1'b1;
    layer2_outputs(1033) <= 1'b0;
    layer2_outputs(1034) <= not (a and b);
    layer2_outputs(1035) <= not b;
    layer2_outputs(1036) <= not b or a;
    layer2_outputs(1037) <= 1'b0;
    layer2_outputs(1038) <= 1'b0;
    layer2_outputs(1039) <= not b;
    layer2_outputs(1040) <= b and not a;
    layer2_outputs(1041) <= a;
    layer2_outputs(1042) <= not (a xor b);
    layer2_outputs(1043) <= a and not b;
    layer2_outputs(1044) <= a and not b;
    layer2_outputs(1045) <= 1'b0;
    layer2_outputs(1046) <= b and not a;
    layer2_outputs(1047) <= b and not a;
    layer2_outputs(1048) <= b;
    layer2_outputs(1049) <= a and b;
    layer2_outputs(1050) <= not (a or b);
    layer2_outputs(1051) <= 1'b1;
    layer2_outputs(1052) <= not b or a;
    layer2_outputs(1053) <= not a;
    layer2_outputs(1054) <= not a or b;
    layer2_outputs(1055) <= not (a xor b);
    layer2_outputs(1056) <= not (a and b);
    layer2_outputs(1057) <= a and not b;
    layer2_outputs(1058) <= not (a or b);
    layer2_outputs(1059) <= a and b;
    layer2_outputs(1060) <= not (a xor b);
    layer2_outputs(1061) <= not a or b;
    layer2_outputs(1062) <= not (a xor b);
    layer2_outputs(1063) <= not (a xor b);
    layer2_outputs(1064) <= b;
    layer2_outputs(1065) <= 1'b0;
    layer2_outputs(1066) <= a or b;
    layer2_outputs(1067) <= a or b;
    layer2_outputs(1068) <= not (a and b);
    layer2_outputs(1069) <= a and not b;
    layer2_outputs(1070) <= not (a or b);
    layer2_outputs(1071) <= b and not a;
    layer2_outputs(1072) <= not b;
    layer2_outputs(1073) <= not (a and b);
    layer2_outputs(1074) <= not (a xor b);
    layer2_outputs(1075) <= a;
    layer2_outputs(1076) <= 1'b1;
    layer2_outputs(1077) <= 1'b0;
    layer2_outputs(1078) <= a;
    layer2_outputs(1079) <= not a or b;
    layer2_outputs(1080) <= a and not b;
    layer2_outputs(1081) <= a;
    layer2_outputs(1082) <= 1'b1;
    layer2_outputs(1083) <= 1'b0;
    layer2_outputs(1084) <= a or b;
    layer2_outputs(1085) <= a and b;
    layer2_outputs(1086) <= not a or b;
    layer2_outputs(1087) <= 1'b1;
    layer2_outputs(1088) <= a and not b;
    layer2_outputs(1089) <= not b;
    layer2_outputs(1090) <= not (a and b);
    layer2_outputs(1091) <= not a;
    layer2_outputs(1092) <= a;
    layer2_outputs(1093) <= not b or a;
    layer2_outputs(1094) <= a or b;
    layer2_outputs(1095) <= not (a and b);
    layer2_outputs(1096) <= not (a or b);
    layer2_outputs(1097) <= b and not a;
    layer2_outputs(1098) <= not b;
    layer2_outputs(1099) <= b;
    layer2_outputs(1100) <= 1'b0;
    layer2_outputs(1101) <= 1'b1;
    layer2_outputs(1102) <= a;
    layer2_outputs(1103) <= b and not a;
    layer2_outputs(1104) <= not a or b;
    layer2_outputs(1105) <= a or b;
    layer2_outputs(1106) <= a or b;
    layer2_outputs(1107) <= not (a or b);
    layer2_outputs(1108) <= a;
    layer2_outputs(1109) <= not b or a;
    layer2_outputs(1110) <= not a or b;
    layer2_outputs(1111) <= not a or b;
    layer2_outputs(1112) <= a or b;
    layer2_outputs(1113) <= not b;
    layer2_outputs(1114) <= not (a and b);
    layer2_outputs(1115) <= b and not a;
    layer2_outputs(1116) <= b and not a;
    layer2_outputs(1117) <= not a;
    layer2_outputs(1118) <= a;
    layer2_outputs(1119) <= b;
    layer2_outputs(1120) <= a or b;
    layer2_outputs(1121) <= not b or a;
    layer2_outputs(1122) <= 1'b1;
    layer2_outputs(1123) <= a or b;
    layer2_outputs(1124) <= 1'b0;
    layer2_outputs(1125) <= not b or a;
    layer2_outputs(1126) <= b and not a;
    layer2_outputs(1127) <= not b;
    layer2_outputs(1128) <= not (a or b);
    layer2_outputs(1129) <= b;
    layer2_outputs(1130) <= a and b;
    layer2_outputs(1131) <= b and not a;
    layer2_outputs(1132) <= b and not a;
    layer2_outputs(1133) <= a;
    layer2_outputs(1134) <= 1'b0;
    layer2_outputs(1135) <= b and not a;
    layer2_outputs(1136) <= not (a or b);
    layer2_outputs(1137) <= a and b;
    layer2_outputs(1138) <= 1'b1;
    layer2_outputs(1139) <= not b;
    layer2_outputs(1140) <= a and not b;
    layer2_outputs(1141) <= not b;
    layer2_outputs(1142) <= a and b;
    layer2_outputs(1143) <= not b;
    layer2_outputs(1144) <= not (a and b);
    layer2_outputs(1145) <= not (a or b);
    layer2_outputs(1146) <= 1'b1;
    layer2_outputs(1147) <= a or b;
    layer2_outputs(1148) <= not (a and b);
    layer2_outputs(1149) <= a or b;
    layer2_outputs(1150) <= not a;
    layer2_outputs(1151) <= not (a or b);
    layer2_outputs(1152) <= 1'b0;
    layer2_outputs(1153) <= b and not a;
    layer2_outputs(1154) <= a;
    layer2_outputs(1155) <= a and not b;
    layer2_outputs(1156) <= not b;
    layer2_outputs(1157) <= b and not a;
    layer2_outputs(1158) <= a;
    layer2_outputs(1159) <= a or b;
    layer2_outputs(1160) <= not b or a;
    layer2_outputs(1161) <= a;
    layer2_outputs(1162) <= not a;
    layer2_outputs(1163) <= 1'b1;
    layer2_outputs(1164) <= a and b;
    layer2_outputs(1165) <= not (a and b);
    layer2_outputs(1166) <= a and not b;
    layer2_outputs(1167) <= not a;
    layer2_outputs(1168) <= 1'b1;
    layer2_outputs(1169) <= 1'b1;
    layer2_outputs(1170) <= a and b;
    layer2_outputs(1171) <= a;
    layer2_outputs(1172) <= 1'b0;
    layer2_outputs(1173) <= b and not a;
    layer2_outputs(1174) <= not (a and b);
    layer2_outputs(1175) <= not a;
    layer2_outputs(1176) <= a;
    layer2_outputs(1177) <= a and not b;
    layer2_outputs(1178) <= not b or a;
    layer2_outputs(1179) <= a and b;
    layer2_outputs(1180) <= a and not b;
    layer2_outputs(1181) <= a and b;
    layer2_outputs(1182) <= a and b;
    layer2_outputs(1183) <= a and b;
    layer2_outputs(1184) <= 1'b1;
    layer2_outputs(1185) <= not b or a;
    layer2_outputs(1186) <= 1'b1;
    layer2_outputs(1187) <= a or b;
    layer2_outputs(1188) <= 1'b0;
    layer2_outputs(1189) <= a and b;
    layer2_outputs(1190) <= not (a or b);
    layer2_outputs(1191) <= 1'b1;
    layer2_outputs(1192) <= a;
    layer2_outputs(1193) <= not b or a;
    layer2_outputs(1194) <= not (a and b);
    layer2_outputs(1195) <= not a or b;
    layer2_outputs(1196) <= a and b;
    layer2_outputs(1197) <= not a or b;
    layer2_outputs(1198) <= a;
    layer2_outputs(1199) <= a;
    layer2_outputs(1200) <= a and b;
    layer2_outputs(1201) <= 1'b1;
    layer2_outputs(1202) <= not b or a;
    layer2_outputs(1203) <= a and b;
    layer2_outputs(1204) <= not a;
    layer2_outputs(1205) <= 1'b0;
    layer2_outputs(1206) <= a and not b;
    layer2_outputs(1207) <= 1'b1;
    layer2_outputs(1208) <= not b or a;
    layer2_outputs(1209) <= a and not b;
    layer2_outputs(1210) <= not a or b;
    layer2_outputs(1211) <= not b or a;
    layer2_outputs(1212) <= a or b;
    layer2_outputs(1213) <= a;
    layer2_outputs(1214) <= not b;
    layer2_outputs(1215) <= not b;
    layer2_outputs(1216) <= 1'b0;
    layer2_outputs(1217) <= not (a or b);
    layer2_outputs(1218) <= a and not b;
    layer2_outputs(1219) <= 1'b0;
    layer2_outputs(1220) <= not b;
    layer2_outputs(1221) <= 1'b1;
    layer2_outputs(1222) <= b and not a;
    layer2_outputs(1223) <= not b or a;
    layer2_outputs(1224) <= a;
    layer2_outputs(1225) <= not a;
    layer2_outputs(1226) <= 1'b1;
    layer2_outputs(1227) <= b;
    layer2_outputs(1228) <= a and not b;
    layer2_outputs(1229) <= b and not a;
    layer2_outputs(1230) <= not a;
    layer2_outputs(1231) <= not b;
    layer2_outputs(1232) <= a;
    layer2_outputs(1233) <= a or b;
    layer2_outputs(1234) <= not b or a;
    layer2_outputs(1235) <= b;
    layer2_outputs(1236) <= 1'b1;
    layer2_outputs(1237) <= a;
    layer2_outputs(1238) <= b;
    layer2_outputs(1239) <= b;
    layer2_outputs(1240) <= not b;
    layer2_outputs(1241) <= 1'b0;
    layer2_outputs(1242) <= b;
    layer2_outputs(1243) <= 1'b0;
    layer2_outputs(1244) <= not (a or b);
    layer2_outputs(1245) <= 1'b1;
    layer2_outputs(1246) <= a;
    layer2_outputs(1247) <= not a or b;
    layer2_outputs(1248) <= not (a and b);
    layer2_outputs(1249) <= not b or a;
    layer2_outputs(1250) <= not a;
    layer2_outputs(1251) <= not (a and b);
    layer2_outputs(1252) <= not a or b;
    layer2_outputs(1253) <= not (a or b);
    layer2_outputs(1254) <= not (a or b);
    layer2_outputs(1255) <= 1'b0;
    layer2_outputs(1256) <= 1'b1;
    layer2_outputs(1257) <= a;
    layer2_outputs(1258) <= b and not a;
    layer2_outputs(1259) <= b;
    layer2_outputs(1260) <= 1'b1;
    layer2_outputs(1261) <= 1'b0;
    layer2_outputs(1262) <= not b or a;
    layer2_outputs(1263) <= not a;
    layer2_outputs(1264) <= not a or b;
    layer2_outputs(1265) <= a or b;
    layer2_outputs(1266) <= b;
    layer2_outputs(1267) <= b;
    layer2_outputs(1268) <= not a or b;
    layer2_outputs(1269) <= a and b;
    layer2_outputs(1270) <= b;
    layer2_outputs(1271) <= not a;
    layer2_outputs(1272) <= not (a or b);
    layer2_outputs(1273) <= b and not a;
    layer2_outputs(1274) <= 1'b0;
    layer2_outputs(1275) <= not b;
    layer2_outputs(1276) <= a or b;
    layer2_outputs(1277) <= 1'b1;
    layer2_outputs(1278) <= not (a or b);
    layer2_outputs(1279) <= a and not b;
    layer2_outputs(1280) <= b;
    layer2_outputs(1281) <= a;
    layer2_outputs(1282) <= not (a and b);
    layer2_outputs(1283) <= 1'b0;
    layer2_outputs(1284) <= 1'b0;
    layer2_outputs(1285) <= a;
    layer2_outputs(1286) <= 1'b1;
    layer2_outputs(1287) <= a and not b;
    layer2_outputs(1288) <= b;
    layer2_outputs(1289) <= not b or a;
    layer2_outputs(1290) <= b;
    layer2_outputs(1291) <= b and not a;
    layer2_outputs(1292) <= not b or a;
    layer2_outputs(1293) <= a or b;
    layer2_outputs(1294) <= not b;
    layer2_outputs(1295) <= not a;
    layer2_outputs(1296) <= not (a or b);
    layer2_outputs(1297) <= b and not a;
    layer2_outputs(1298) <= not b;
    layer2_outputs(1299) <= b and not a;
    layer2_outputs(1300) <= 1'b0;
    layer2_outputs(1301) <= not (a or b);
    layer2_outputs(1302) <= b;
    layer2_outputs(1303) <= not (a and b);
    layer2_outputs(1304) <= a or b;
    layer2_outputs(1305) <= not a;
    layer2_outputs(1306) <= not (a and b);
    layer2_outputs(1307) <= 1'b0;
    layer2_outputs(1308) <= b and not a;
    layer2_outputs(1309) <= not b or a;
    layer2_outputs(1310) <= 1'b0;
    layer2_outputs(1311) <= 1'b1;
    layer2_outputs(1312) <= 1'b0;
    layer2_outputs(1313) <= not a or b;
    layer2_outputs(1314) <= a and b;
    layer2_outputs(1315) <= a and b;
    layer2_outputs(1316) <= a or b;
    layer2_outputs(1317) <= not a;
    layer2_outputs(1318) <= 1'b0;
    layer2_outputs(1319) <= not a or b;
    layer2_outputs(1320) <= a or b;
    layer2_outputs(1321) <= not a or b;
    layer2_outputs(1322) <= 1'b1;
    layer2_outputs(1323) <= 1'b0;
    layer2_outputs(1324) <= a;
    layer2_outputs(1325) <= not (a and b);
    layer2_outputs(1326) <= 1'b1;
    layer2_outputs(1327) <= b;
    layer2_outputs(1328) <= a or b;
    layer2_outputs(1329) <= not (a and b);
    layer2_outputs(1330) <= not b;
    layer2_outputs(1331) <= not b or a;
    layer2_outputs(1332) <= not (a xor b);
    layer2_outputs(1333) <= a or b;
    layer2_outputs(1334) <= a;
    layer2_outputs(1335) <= not a;
    layer2_outputs(1336) <= not a;
    layer2_outputs(1337) <= a and not b;
    layer2_outputs(1338) <= not (a and b);
    layer2_outputs(1339) <= a and b;
    layer2_outputs(1340) <= not (a xor b);
    layer2_outputs(1341) <= 1'b0;
    layer2_outputs(1342) <= a;
    layer2_outputs(1343) <= not b or a;
    layer2_outputs(1344) <= not (a and b);
    layer2_outputs(1345) <= 1'b1;
    layer2_outputs(1346) <= a;
    layer2_outputs(1347) <= not (a and b);
    layer2_outputs(1348) <= b and not a;
    layer2_outputs(1349) <= not (a xor b);
    layer2_outputs(1350) <= 1'b0;
    layer2_outputs(1351) <= not b or a;
    layer2_outputs(1352) <= a;
    layer2_outputs(1353) <= a or b;
    layer2_outputs(1354) <= 1'b1;
    layer2_outputs(1355) <= not (a or b);
    layer2_outputs(1356) <= 1'b1;
    layer2_outputs(1357) <= 1'b0;
    layer2_outputs(1358) <= b;
    layer2_outputs(1359) <= a and not b;
    layer2_outputs(1360) <= b;
    layer2_outputs(1361) <= 1'b1;
    layer2_outputs(1362) <= a or b;
    layer2_outputs(1363) <= not a or b;
    layer2_outputs(1364) <= b and not a;
    layer2_outputs(1365) <= not (a and b);
    layer2_outputs(1366) <= not b;
    layer2_outputs(1367) <= a or b;
    layer2_outputs(1368) <= not b;
    layer2_outputs(1369) <= not (a and b);
    layer2_outputs(1370) <= b and not a;
    layer2_outputs(1371) <= not a;
    layer2_outputs(1372) <= a or b;
    layer2_outputs(1373) <= a;
    layer2_outputs(1374) <= b;
    layer2_outputs(1375) <= not a or b;
    layer2_outputs(1376) <= 1'b0;
    layer2_outputs(1377) <= a;
    layer2_outputs(1378) <= not a or b;
    layer2_outputs(1379) <= a and b;
    layer2_outputs(1380) <= not b;
    layer2_outputs(1381) <= not a;
    layer2_outputs(1382) <= b;
    layer2_outputs(1383) <= 1'b1;
    layer2_outputs(1384) <= a and not b;
    layer2_outputs(1385) <= 1'b0;
    layer2_outputs(1386) <= 1'b1;
    layer2_outputs(1387) <= 1'b1;
    layer2_outputs(1388) <= b and not a;
    layer2_outputs(1389) <= b;
    layer2_outputs(1390) <= not (a and b);
    layer2_outputs(1391) <= b;
    layer2_outputs(1392) <= not b or a;
    layer2_outputs(1393) <= b;
    layer2_outputs(1394) <= a and not b;
    layer2_outputs(1395) <= b and not a;
    layer2_outputs(1396) <= a;
    layer2_outputs(1397) <= not (a and b);
    layer2_outputs(1398) <= not (a and b);
    layer2_outputs(1399) <= a and not b;
    layer2_outputs(1400) <= 1'b1;
    layer2_outputs(1401) <= not a or b;
    layer2_outputs(1402) <= a;
    layer2_outputs(1403) <= a and not b;
    layer2_outputs(1404) <= not (a xor b);
    layer2_outputs(1405) <= 1'b0;
    layer2_outputs(1406) <= not (a or b);
    layer2_outputs(1407) <= not a;
    layer2_outputs(1408) <= a;
    layer2_outputs(1409) <= b and not a;
    layer2_outputs(1410) <= a;
    layer2_outputs(1411) <= b and not a;
    layer2_outputs(1412) <= not (a and b);
    layer2_outputs(1413) <= not a;
    layer2_outputs(1414) <= not (a or b);
    layer2_outputs(1415) <= 1'b1;
    layer2_outputs(1416) <= 1'b0;
    layer2_outputs(1417) <= not (a xor b);
    layer2_outputs(1418) <= not a or b;
    layer2_outputs(1419) <= a;
    layer2_outputs(1420) <= not b or a;
    layer2_outputs(1421) <= a or b;
    layer2_outputs(1422) <= not (a and b);
    layer2_outputs(1423) <= not a;
    layer2_outputs(1424) <= not b or a;
    layer2_outputs(1425) <= b;
    layer2_outputs(1426) <= not a;
    layer2_outputs(1427) <= not b;
    layer2_outputs(1428) <= not (a or b);
    layer2_outputs(1429) <= a or b;
    layer2_outputs(1430) <= a;
    layer2_outputs(1431) <= a or b;
    layer2_outputs(1432) <= b;
    layer2_outputs(1433) <= a;
    layer2_outputs(1434) <= not b or a;
    layer2_outputs(1435) <= b and not a;
    layer2_outputs(1436) <= not b or a;
    layer2_outputs(1437) <= a;
    layer2_outputs(1438) <= not (a and b);
    layer2_outputs(1439) <= a or b;
    layer2_outputs(1440) <= a or b;
    layer2_outputs(1441) <= not (a or b);
    layer2_outputs(1442) <= a and not b;
    layer2_outputs(1443) <= not a or b;
    layer2_outputs(1444) <= b;
    layer2_outputs(1445) <= not b or a;
    layer2_outputs(1446) <= b;
    layer2_outputs(1447) <= not (a or b);
    layer2_outputs(1448) <= 1'b1;
    layer2_outputs(1449) <= a and b;
    layer2_outputs(1450) <= a or b;
    layer2_outputs(1451) <= not a;
    layer2_outputs(1452) <= 1'b1;
    layer2_outputs(1453) <= b;
    layer2_outputs(1454) <= not (a and b);
    layer2_outputs(1455) <= 1'b0;
    layer2_outputs(1456) <= 1'b1;
    layer2_outputs(1457) <= not (a or b);
    layer2_outputs(1458) <= 1'b0;
    layer2_outputs(1459) <= 1'b0;
    layer2_outputs(1460) <= not b;
    layer2_outputs(1461) <= not b or a;
    layer2_outputs(1462) <= not (a or b);
    layer2_outputs(1463) <= not a;
    layer2_outputs(1464) <= not (a or b);
    layer2_outputs(1465) <= b and not a;
    layer2_outputs(1466) <= not a;
    layer2_outputs(1467) <= not a;
    layer2_outputs(1468) <= not b;
    layer2_outputs(1469) <= not a or b;
    layer2_outputs(1470) <= not a or b;
    layer2_outputs(1471) <= b and not a;
    layer2_outputs(1472) <= a xor b;
    layer2_outputs(1473) <= not a;
    layer2_outputs(1474) <= not (a or b);
    layer2_outputs(1475) <= a and b;
    layer2_outputs(1476) <= not a;
    layer2_outputs(1477) <= 1'b0;
    layer2_outputs(1478) <= not b or a;
    layer2_outputs(1479) <= 1'b0;
    layer2_outputs(1480) <= not b or a;
    layer2_outputs(1481) <= not (a or b);
    layer2_outputs(1482) <= not b;
    layer2_outputs(1483) <= 1'b1;
    layer2_outputs(1484) <= not b or a;
    layer2_outputs(1485) <= a xor b;
    layer2_outputs(1486) <= b;
    layer2_outputs(1487) <= not a;
    layer2_outputs(1488) <= a and b;
    layer2_outputs(1489) <= not a;
    layer2_outputs(1490) <= not b or a;
    layer2_outputs(1491) <= not (a and b);
    layer2_outputs(1492) <= 1'b0;
    layer2_outputs(1493) <= 1'b0;
    layer2_outputs(1494) <= a and not b;
    layer2_outputs(1495) <= a xor b;
    layer2_outputs(1496) <= a or b;
    layer2_outputs(1497) <= a and b;
    layer2_outputs(1498) <= b and not a;
    layer2_outputs(1499) <= b;
    layer2_outputs(1500) <= not a or b;
    layer2_outputs(1501) <= a;
    layer2_outputs(1502) <= not b;
    layer2_outputs(1503) <= not a or b;
    layer2_outputs(1504) <= a and not b;
    layer2_outputs(1505) <= not a;
    layer2_outputs(1506) <= a or b;
    layer2_outputs(1507) <= b;
    layer2_outputs(1508) <= not a or b;
    layer2_outputs(1509) <= not (a and b);
    layer2_outputs(1510) <= a;
    layer2_outputs(1511) <= a;
    layer2_outputs(1512) <= not (a xor b);
    layer2_outputs(1513) <= not a or b;
    layer2_outputs(1514) <= 1'b1;
    layer2_outputs(1515) <= not a;
    layer2_outputs(1516) <= b and not a;
    layer2_outputs(1517) <= b and not a;
    layer2_outputs(1518) <= not b;
    layer2_outputs(1519) <= not (a or b);
    layer2_outputs(1520) <= b;
    layer2_outputs(1521) <= not b or a;
    layer2_outputs(1522) <= a;
    layer2_outputs(1523) <= not a;
    layer2_outputs(1524) <= not (a or b);
    layer2_outputs(1525) <= 1'b0;
    layer2_outputs(1526) <= b and not a;
    layer2_outputs(1527) <= b;
    layer2_outputs(1528) <= a;
    layer2_outputs(1529) <= a;
    layer2_outputs(1530) <= a or b;
    layer2_outputs(1531) <= a or b;
    layer2_outputs(1532) <= a and not b;
    layer2_outputs(1533) <= not (a xor b);
    layer2_outputs(1534) <= a and not b;
    layer2_outputs(1535) <= a;
    layer2_outputs(1536) <= b;
    layer2_outputs(1537) <= not (a and b);
    layer2_outputs(1538) <= b;
    layer2_outputs(1539) <= b and not a;
    layer2_outputs(1540) <= b;
    layer2_outputs(1541) <= a or b;
    layer2_outputs(1542) <= 1'b0;
    layer2_outputs(1543) <= 1'b1;
    layer2_outputs(1544) <= not a;
    layer2_outputs(1545) <= 1'b0;
    layer2_outputs(1546) <= 1'b1;
    layer2_outputs(1547) <= not a;
    layer2_outputs(1548) <= a and not b;
    layer2_outputs(1549) <= not (a and b);
    layer2_outputs(1550) <= not (a and b);
    layer2_outputs(1551) <= 1'b0;
    layer2_outputs(1552) <= 1'b1;
    layer2_outputs(1553) <= a and b;
    layer2_outputs(1554) <= not (a or b);
    layer2_outputs(1555) <= a or b;
    layer2_outputs(1556) <= a;
    layer2_outputs(1557) <= not (a xor b);
    layer2_outputs(1558) <= 1'b0;
    layer2_outputs(1559) <= a or b;
    layer2_outputs(1560) <= 1'b0;
    layer2_outputs(1561) <= a or b;
    layer2_outputs(1562) <= not a;
    layer2_outputs(1563) <= not b;
    layer2_outputs(1564) <= not (a xor b);
    layer2_outputs(1565) <= not a;
    layer2_outputs(1566) <= 1'b1;
    layer2_outputs(1567) <= b and not a;
    layer2_outputs(1568) <= a;
    layer2_outputs(1569) <= not b or a;
    layer2_outputs(1570) <= not (a and b);
    layer2_outputs(1571) <= not (a and b);
    layer2_outputs(1572) <= a;
    layer2_outputs(1573) <= not b or a;
    layer2_outputs(1574) <= a and b;
    layer2_outputs(1575) <= not (a or b);
    layer2_outputs(1576) <= 1'b1;
    layer2_outputs(1577) <= not b or a;
    layer2_outputs(1578) <= not (a or b);
    layer2_outputs(1579) <= a or b;
    layer2_outputs(1580) <= not b or a;
    layer2_outputs(1581) <= not b or a;
    layer2_outputs(1582) <= a or b;
    layer2_outputs(1583) <= not b or a;
    layer2_outputs(1584) <= a;
    layer2_outputs(1585) <= a and b;
    layer2_outputs(1586) <= not (a xor b);
    layer2_outputs(1587) <= a and not b;
    layer2_outputs(1588) <= not b or a;
    layer2_outputs(1589) <= not a or b;
    layer2_outputs(1590) <= 1'b1;
    layer2_outputs(1591) <= not a;
    layer2_outputs(1592) <= a;
    layer2_outputs(1593) <= b and not a;
    layer2_outputs(1594) <= a or b;
    layer2_outputs(1595) <= 1'b1;
    layer2_outputs(1596) <= not b;
    layer2_outputs(1597) <= b and not a;
    layer2_outputs(1598) <= not a or b;
    layer2_outputs(1599) <= 1'b0;
    layer2_outputs(1600) <= a and not b;
    layer2_outputs(1601) <= not b;
    layer2_outputs(1602) <= 1'b0;
    layer2_outputs(1603) <= not a or b;
    layer2_outputs(1604) <= a or b;
    layer2_outputs(1605) <= a and b;
    layer2_outputs(1606) <= not a or b;
    layer2_outputs(1607) <= not (a and b);
    layer2_outputs(1608) <= not a;
    layer2_outputs(1609) <= not a or b;
    layer2_outputs(1610) <= not b;
    layer2_outputs(1611) <= not b;
    layer2_outputs(1612) <= not (a and b);
    layer2_outputs(1613) <= 1'b0;
    layer2_outputs(1614) <= not (a or b);
    layer2_outputs(1615) <= b and not a;
    layer2_outputs(1616) <= 1'b0;
    layer2_outputs(1617) <= a or b;
    layer2_outputs(1618) <= 1'b1;
    layer2_outputs(1619) <= not a or b;
    layer2_outputs(1620) <= a or b;
    layer2_outputs(1621) <= not (a or b);
    layer2_outputs(1622) <= a and not b;
    layer2_outputs(1623) <= a or b;
    layer2_outputs(1624) <= a and not b;
    layer2_outputs(1625) <= 1'b0;
    layer2_outputs(1626) <= 1'b1;
    layer2_outputs(1627) <= not b or a;
    layer2_outputs(1628) <= a or b;
    layer2_outputs(1629) <= not a;
    layer2_outputs(1630) <= not b or a;
    layer2_outputs(1631) <= not (a or b);
    layer2_outputs(1632) <= 1'b0;
    layer2_outputs(1633) <= not (a and b);
    layer2_outputs(1634) <= 1'b0;
    layer2_outputs(1635) <= not b or a;
    layer2_outputs(1636) <= 1'b0;
    layer2_outputs(1637) <= not (a or b);
    layer2_outputs(1638) <= a and b;
    layer2_outputs(1639) <= not a;
    layer2_outputs(1640) <= not (a or b);
    layer2_outputs(1641) <= not a;
    layer2_outputs(1642) <= a xor b;
    layer2_outputs(1643) <= a xor b;
    layer2_outputs(1644) <= 1'b1;
    layer2_outputs(1645) <= a and not b;
    layer2_outputs(1646) <= a or b;
    layer2_outputs(1647) <= not a or b;
    layer2_outputs(1648) <= b and not a;
    layer2_outputs(1649) <= b and not a;
    layer2_outputs(1650) <= not b or a;
    layer2_outputs(1651) <= 1'b0;
    layer2_outputs(1652) <= not a;
    layer2_outputs(1653) <= not (a or b);
    layer2_outputs(1654) <= a and not b;
    layer2_outputs(1655) <= not b or a;
    layer2_outputs(1656) <= 1'b0;
    layer2_outputs(1657) <= b;
    layer2_outputs(1658) <= b;
    layer2_outputs(1659) <= not a or b;
    layer2_outputs(1660) <= not b or a;
    layer2_outputs(1661) <= b;
    layer2_outputs(1662) <= not (a and b);
    layer2_outputs(1663) <= b;
    layer2_outputs(1664) <= b and not a;
    layer2_outputs(1665) <= b and not a;
    layer2_outputs(1666) <= b and not a;
    layer2_outputs(1667) <= not a;
    layer2_outputs(1668) <= not a or b;
    layer2_outputs(1669) <= a and b;
    layer2_outputs(1670) <= 1'b1;
    layer2_outputs(1671) <= a or b;
    layer2_outputs(1672) <= not (a and b);
    layer2_outputs(1673) <= a and b;
    layer2_outputs(1674) <= not b or a;
    layer2_outputs(1675) <= 1'b0;
    layer2_outputs(1676) <= a or b;
    layer2_outputs(1677) <= not a or b;
    layer2_outputs(1678) <= not (a xor b);
    layer2_outputs(1679) <= 1'b1;
    layer2_outputs(1680) <= not (a xor b);
    layer2_outputs(1681) <= 1'b0;
    layer2_outputs(1682) <= 1'b0;
    layer2_outputs(1683) <= not (a or b);
    layer2_outputs(1684) <= b and not a;
    layer2_outputs(1685) <= b;
    layer2_outputs(1686) <= a or b;
    layer2_outputs(1687) <= a;
    layer2_outputs(1688) <= not a or b;
    layer2_outputs(1689) <= a or b;
    layer2_outputs(1690) <= not (a or b);
    layer2_outputs(1691) <= 1'b1;
    layer2_outputs(1692) <= a and not b;
    layer2_outputs(1693) <= not a;
    layer2_outputs(1694) <= 1'b0;
    layer2_outputs(1695) <= 1'b0;
    layer2_outputs(1696) <= a and b;
    layer2_outputs(1697) <= a;
    layer2_outputs(1698) <= a;
    layer2_outputs(1699) <= a xor b;
    layer2_outputs(1700) <= not b;
    layer2_outputs(1701) <= b;
    layer2_outputs(1702) <= a;
    layer2_outputs(1703) <= b and not a;
    layer2_outputs(1704) <= b and not a;
    layer2_outputs(1705) <= not b;
    layer2_outputs(1706) <= not (a and b);
    layer2_outputs(1707) <= not a or b;
    layer2_outputs(1708) <= 1'b0;
    layer2_outputs(1709) <= a and not b;
    layer2_outputs(1710) <= b and not a;
    layer2_outputs(1711) <= 1'b0;
    layer2_outputs(1712) <= not b or a;
    layer2_outputs(1713) <= not a or b;
    layer2_outputs(1714) <= not b;
    layer2_outputs(1715) <= b and not a;
    layer2_outputs(1716) <= b and not a;
    layer2_outputs(1717) <= b and not a;
    layer2_outputs(1718) <= not a or b;
    layer2_outputs(1719) <= b and not a;
    layer2_outputs(1720) <= not (a and b);
    layer2_outputs(1721) <= a;
    layer2_outputs(1722) <= not (a and b);
    layer2_outputs(1723) <= a xor b;
    layer2_outputs(1724) <= not b;
    layer2_outputs(1725) <= a and not b;
    layer2_outputs(1726) <= b and not a;
    layer2_outputs(1727) <= a and b;
    layer2_outputs(1728) <= not (a and b);
    layer2_outputs(1729) <= not a;
    layer2_outputs(1730) <= a and b;
    layer2_outputs(1731) <= 1'b0;
    layer2_outputs(1732) <= a xor b;
    layer2_outputs(1733) <= a and b;
    layer2_outputs(1734) <= not b;
    layer2_outputs(1735) <= not a or b;
    layer2_outputs(1736) <= not a;
    layer2_outputs(1737) <= b;
    layer2_outputs(1738) <= a or b;
    layer2_outputs(1739) <= b and not a;
    layer2_outputs(1740) <= not (a and b);
    layer2_outputs(1741) <= not a or b;
    layer2_outputs(1742) <= not a or b;
    layer2_outputs(1743) <= not b;
    layer2_outputs(1744) <= 1'b1;
    layer2_outputs(1745) <= 1'b0;
    layer2_outputs(1746) <= not a or b;
    layer2_outputs(1747) <= not b;
    layer2_outputs(1748) <= 1'b1;
    layer2_outputs(1749) <= a or b;
    layer2_outputs(1750) <= 1'b1;
    layer2_outputs(1751) <= not a or b;
    layer2_outputs(1752) <= 1'b1;
    layer2_outputs(1753) <= b and not a;
    layer2_outputs(1754) <= b;
    layer2_outputs(1755) <= b and not a;
    layer2_outputs(1756) <= not (a or b);
    layer2_outputs(1757) <= a or b;
    layer2_outputs(1758) <= not b;
    layer2_outputs(1759) <= a xor b;
    layer2_outputs(1760) <= b and not a;
    layer2_outputs(1761) <= a and not b;
    layer2_outputs(1762) <= b and not a;
    layer2_outputs(1763) <= a or b;
    layer2_outputs(1764) <= not (a and b);
    layer2_outputs(1765) <= not (a or b);
    layer2_outputs(1766) <= a;
    layer2_outputs(1767) <= not b or a;
    layer2_outputs(1768) <= a;
    layer2_outputs(1769) <= a and b;
    layer2_outputs(1770) <= 1'b1;
    layer2_outputs(1771) <= not a or b;
    layer2_outputs(1772) <= a;
    layer2_outputs(1773) <= 1'b1;
    layer2_outputs(1774) <= b and not a;
    layer2_outputs(1775) <= not a;
    layer2_outputs(1776) <= not b or a;
    layer2_outputs(1777) <= not a;
    layer2_outputs(1778) <= a and b;
    layer2_outputs(1779) <= a xor b;
    layer2_outputs(1780) <= a or b;
    layer2_outputs(1781) <= a xor b;
    layer2_outputs(1782) <= 1'b0;
    layer2_outputs(1783) <= a;
    layer2_outputs(1784) <= b;
    layer2_outputs(1785) <= not b;
    layer2_outputs(1786) <= not a;
    layer2_outputs(1787) <= a and not b;
    layer2_outputs(1788) <= b;
    layer2_outputs(1789) <= a;
    layer2_outputs(1790) <= a and b;
    layer2_outputs(1791) <= b and not a;
    layer2_outputs(1792) <= a or b;
    layer2_outputs(1793) <= a or b;
    layer2_outputs(1794) <= b and not a;
    layer2_outputs(1795) <= 1'b1;
    layer2_outputs(1796) <= not (a xor b);
    layer2_outputs(1797) <= not b;
    layer2_outputs(1798) <= b;
    layer2_outputs(1799) <= not a or b;
    layer2_outputs(1800) <= not a;
    layer2_outputs(1801) <= a;
    layer2_outputs(1802) <= b;
    layer2_outputs(1803) <= a and b;
    layer2_outputs(1804) <= not (a xor b);
    layer2_outputs(1805) <= b;
    layer2_outputs(1806) <= not (a xor b);
    layer2_outputs(1807) <= a;
    layer2_outputs(1808) <= a or b;
    layer2_outputs(1809) <= a or b;
    layer2_outputs(1810) <= a and not b;
    layer2_outputs(1811) <= not (a and b);
    layer2_outputs(1812) <= a and b;
    layer2_outputs(1813) <= not b or a;
    layer2_outputs(1814) <= not (a xor b);
    layer2_outputs(1815) <= not a or b;
    layer2_outputs(1816) <= a and b;
    layer2_outputs(1817) <= b and not a;
    layer2_outputs(1818) <= a and b;
    layer2_outputs(1819) <= b and not a;
    layer2_outputs(1820) <= 1'b0;
    layer2_outputs(1821) <= not b;
    layer2_outputs(1822) <= a and not b;
    layer2_outputs(1823) <= a and not b;
    layer2_outputs(1824) <= not b;
    layer2_outputs(1825) <= b;
    layer2_outputs(1826) <= not b or a;
    layer2_outputs(1827) <= b;
    layer2_outputs(1828) <= not b or a;
    layer2_outputs(1829) <= a and b;
    layer2_outputs(1830) <= 1'b0;
    layer2_outputs(1831) <= a and b;
    layer2_outputs(1832) <= a or b;
    layer2_outputs(1833) <= not a;
    layer2_outputs(1834) <= b;
    layer2_outputs(1835) <= not (a or b);
    layer2_outputs(1836) <= not a or b;
    layer2_outputs(1837) <= not a or b;
    layer2_outputs(1838) <= 1'b1;
    layer2_outputs(1839) <= 1'b1;
    layer2_outputs(1840) <= a and b;
    layer2_outputs(1841) <= a and not b;
    layer2_outputs(1842) <= 1'b1;
    layer2_outputs(1843) <= not (a xor b);
    layer2_outputs(1844) <= not a or b;
    layer2_outputs(1845) <= not b or a;
    layer2_outputs(1846) <= not (a or b);
    layer2_outputs(1847) <= not (a and b);
    layer2_outputs(1848) <= b;
    layer2_outputs(1849) <= a or b;
    layer2_outputs(1850) <= 1'b0;
    layer2_outputs(1851) <= not (a or b);
    layer2_outputs(1852) <= 1'b1;
    layer2_outputs(1853) <= not a;
    layer2_outputs(1854) <= not b;
    layer2_outputs(1855) <= not b or a;
    layer2_outputs(1856) <= not a or b;
    layer2_outputs(1857) <= not (a or b);
    layer2_outputs(1858) <= a and b;
    layer2_outputs(1859) <= not a or b;
    layer2_outputs(1860) <= a or b;
    layer2_outputs(1861) <= not b or a;
    layer2_outputs(1862) <= not (a and b);
    layer2_outputs(1863) <= a and b;
    layer2_outputs(1864) <= not a;
    layer2_outputs(1865) <= not (a or b);
    layer2_outputs(1866) <= not (a xor b);
    layer2_outputs(1867) <= not (a xor b);
    layer2_outputs(1868) <= not b or a;
    layer2_outputs(1869) <= 1'b0;
    layer2_outputs(1870) <= 1'b1;
    layer2_outputs(1871) <= not a;
    layer2_outputs(1872) <= b and not a;
    layer2_outputs(1873) <= a and not b;
    layer2_outputs(1874) <= not b;
    layer2_outputs(1875) <= not (a and b);
    layer2_outputs(1876) <= a and b;
    layer2_outputs(1877) <= a and b;
    layer2_outputs(1878) <= b;
    layer2_outputs(1879) <= b;
    layer2_outputs(1880) <= b;
    layer2_outputs(1881) <= 1'b1;
    layer2_outputs(1882) <= a and b;
    layer2_outputs(1883) <= not b or a;
    layer2_outputs(1884) <= b and not a;
    layer2_outputs(1885) <= a and not b;
    layer2_outputs(1886) <= 1'b0;
    layer2_outputs(1887) <= not a;
    layer2_outputs(1888) <= not a or b;
    layer2_outputs(1889) <= 1'b1;
    layer2_outputs(1890) <= not b;
    layer2_outputs(1891) <= not a;
    layer2_outputs(1892) <= not b;
    layer2_outputs(1893) <= a;
    layer2_outputs(1894) <= b;
    layer2_outputs(1895) <= a xor b;
    layer2_outputs(1896) <= not a;
    layer2_outputs(1897) <= b and not a;
    layer2_outputs(1898) <= a xor b;
    layer2_outputs(1899) <= b and not a;
    layer2_outputs(1900) <= not b or a;
    layer2_outputs(1901) <= a;
    layer2_outputs(1902) <= not a;
    layer2_outputs(1903) <= not b or a;
    layer2_outputs(1904) <= 1'b1;
    layer2_outputs(1905) <= not (a and b);
    layer2_outputs(1906) <= b;
    layer2_outputs(1907) <= not (a or b);
    layer2_outputs(1908) <= a and b;
    layer2_outputs(1909) <= not (a xor b);
    layer2_outputs(1910) <= 1'b0;
    layer2_outputs(1911) <= a;
    layer2_outputs(1912) <= a and not b;
    layer2_outputs(1913) <= not b;
    layer2_outputs(1914) <= a and b;
    layer2_outputs(1915) <= not a or b;
    layer2_outputs(1916) <= 1'b1;
    layer2_outputs(1917) <= b and not a;
    layer2_outputs(1918) <= not a;
    layer2_outputs(1919) <= not (a or b);
    layer2_outputs(1920) <= not (a and b);
    layer2_outputs(1921) <= not a;
    layer2_outputs(1922) <= not a;
    layer2_outputs(1923) <= a or b;
    layer2_outputs(1924) <= b;
    layer2_outputs(1925) <= 1'b1;
    layer2_outputs(1926) <= not b;
    layer2_outputs(1927) <= b;
    layer2_outputs(1928) <= a;
    layer2_outputs(1929) <= a or b;
    layer2_outputs(1930) <= 1'b1;
    layer2_outputs(1931) <= not a;
    layer2_outputs(1932) <= a and b;
    layer2_outputs(1933) <= not a;
    layer2_outputs(1934) <= a or b;
    layer2_outputs(1935) <= 1'b0;
    layer2_outputs(1936) <= 1'b0;
    layer2_outputs(1937) <= not (a xor b);
    layer2_outputs(1938) <= a and not b;
    layer2_outputs(1939) <= not (a or b);
    layer2_outputs(1940) <= a;
    layer2_outputs(1941) <= a and b;
    layer2_outputs(1942) <= not (a or b);
    layer2_outputs(1943) <= a and not b;
    layer2_outputs(1944) <= b and not a;
    layer2_outputs(1945) <= 1'b1;
    layer2_outputs(1946) <= not (a and b);
    layer2_outputs(1947) <= not b;
    layer2_outputs(1948) <= not (a or b);
    layer2_outputs(1949) <= not (a or b);
    layer2_outputs(1950) <= a;
    layer2_outputs(1951) <= b;
    layer2_outputs(1952) <= 1'b1;
    layer2_outputs(1953) <= not (a and b);
    layer2_outputs(1954) <= a or b;
    layer2_outputs(1955) <= not b or a;
    layer2_outputs(1956) <= not b or a;
    layer2_outputs(1957) <= b;
    layer2_outputs(1958) <= not a or b;
    layer2_outputs(1959) <= a xor b;
    layer2_outputs(1960) <= b and not a;
    layer2_outputs(1961) <= 1'b1;
    layer2_outputs(1962) <= a or b;
    layer2_outputs(1963) <= 1'b1;
    layer2_outputs(1964) <= a and b;
    layer2_outputs(1965) <= not b or a;
    layer2_outputs(1966) <= not (a or b);
    layer2_outputs(1967) <= not b or a;
    layer2_outputs(1968) <= not a or b;
    layer2_outputs(1969) <= not a;
    layer2_outputs(1970) <= 1'b1;
    layer2_outputs(1971) <= not a;
    layer2_outputs(1972) <= 1'b1;
    layer2_outputs(1973) <= not (a or b);
    layer2_outputs(1974) <= a or b;
    layer2_outputs(1975) <= not b or a;
    layer2_outputs(1976) <= 1'b1;
    layer2_outputs(1977) <= 1'b1;
    layer2_outputs(1978) <= not b;
    layer2_outputs(1979) <= not (a or b);
    layer2_outputs(1980) <= not a or b;
    layer2_outputs(1981) <= a or b;
    layer2_outputs(1982) <= a and not b;
    layer2_outputs(1983) <= not a;
    layer2_outputs(1984) <= not b or a;
    layer2_outputs(1985) <= not b or a;
    layer2_outputs(1986) <= not b;
    layer2_outputs(1987) <= not (a or b);
    layer2_outputs(1988) <= a and b;
    layer2_outputs(1989) <= b;
    layer2_outputs(1990) <= not a or b;
    layer2_outputs(1991) <= b and not a;
    layer2_outputs(1992) <= 1'b0;
    layer2_outputs(1993) <= a or b;
    layer2_outputs(1994) <= not b or a;
    layer2_outputs(1995) <= not b or a;
    layer2_outputs(1996) <= not (a xor b);
    layer2_outputs(1997) <= not a;
    layer2_outputs(1998) <= b;
    layer2_outputs(1999) <= not a;
    layer2_outputs(2000) <= 1'b0;
    layer2_outputs(2001) <= not a;
    layer2_outputs(2002) <= 1'b0;
    layer2_outputs(2003) <= not a;
    layer2_outputs(2004) <= a;
    layer2_outputs(2005) <= a and b;
    layer2_outputs(2006) <= 1'b1;
    layer2_outputs(2007) <= not b;
    layer2_outputs(2008) <= not (a or b);
    layer2_outputs(2009) <= not (a xor b);
    layer2_outputs(2010) <= a or b;
    layer2_outputs(2011) <= not b or a;
    layer2_outputs(2012) <= a xor b;
    layer2_outputs(2013) <= a and not b;
    layer2_outputs(2014) <= 1'b0;
    layer2_outputs(2015) <= 1'b1;
    layer2_outputs(2016) <= not b or a;
    layer2_outputs(2017) <= not b or a;
    layer2_outputs(2018) <= a and not b;
    layer2_outputs(2019) <= not b or a;
    layer2_outputs(2020) <= a and b;
    layer2_outputs(2021) <= 1'b0;
    layer2_outputs(2022) <= not a;
    layer2_outputs(2023) <= a xor b;
    layer2_outputs(2024) <= 1'b1;
    layer2_outputs(2025) <= 1'b0;
    layer2_outputs(2026) <= not (a xor b);
    layer2_outputs(2027) <= b and not a;
    layer2_outputs(2028) <= 1'b1;
    layer2_outputs(2029) <= not (a or b);
    layer2_outputs(2030) <= not b;
    layer2_outputs(2031) <= b and not a;
    layer2_outputs(2032) <= not (a and b);
    layer2_outputs(2033) <= a;
    layer2_outputs(2034) <= not a or b;
    layer2_outputs(2035) <= not b or a;
    layer2_outputs(2036) <= a and not b;
    layer2_outputs(2037) <= a and b;
    layer2_outputs(2038) <= not a;
    layer2_outputs(2039) <= a and b;
    layer2_outputs(2040) <= not b or a;
    layer2_outputs(2041) <= not (a or b);
    layer2_outputs(2042) <= not b or a;
    layer2_outputs(2043) <= 1'b1;
    layer2_outputs(2044) <= a;
    layer2_outputs(2045) <= a;
    layer2_outputs(2046) <= b;
    layer2_outputs(2047) <= a or b;
    layer2_outputs(2048) <= not (a xor b);
    layer2_outputs(2049) <= 1'b1;
    layer2_outputs(2050) <= a and not b;
    layer2_outputs(2051) <= not (a or b);
    layer2_outputs(2052) <= not a or b;
    layer2_outputs(2053) <= a and b;
    layer2_outputs(2054) <= b;
    layer2_outputs(2055) <= b;
    layer2_outputs(2056) <= not (a or b);
    layer2_outputs(2057) <= 1'b1;
    layer2_outputs(2058) <= 1'b0;
    layer2_outputs(2059) <= not a or b;
    layer2_outputs(2060) <= b;
    layer2_outputs(2061) <= not (a xor b);
    layer2_outputs(2062) <= b and not a;
    layer2_outputs(2063) <= b and not a;
    layer2_outputs(2064) <= a or b;
    layer2_outputs(2065) <= not b or a;
    layer2_outputs(2066) <= not a;
    layer2_outputs(2067) <= not a or b;
    layer2_outputs(2068) <= a and b;
    layer2_outputs(2069) <= not a or b;
    layer2_outputs(2070) <= 1'b1;
    layer2_outputs(2071) <= b and not a;
    layer2_outputs(2072) <= a and b;
    layer2_outputs(2073) <= b;
    layer2_outputs(2074) <= not (a and b);
    layer2_outputs(2075) <= 1'b1;
    layer2_outputs(2076) <= not b;
    layer2_outputs(2077) <= a or b;
    layer2_outputs(2078) <= not (a xor b);
    layer2_outputs(2079) <= a and b;
    layer2_outputs(2080) <= 1'b0;
    layer2_outputs(2081) <= 1'b0;
    layer2_outputs(2082) <= not b;
    layer2_outputs(2083) <= not (a and b);
    layer2_outputs(2084) <= a;
    layer2_outputs(2085) <= 1'b0;
    layer2_outputs(2086) <= 1'b0;
    layer2_outputs(2087) <= 1'b0;
    layer2_outputs(2088) <= b and not a;
    layer2_outputs(2089) <= a or b;
    layer2_outputs(2090) <= a or b;
    layer2_outputs(2091) <= not b;
    layer2_outputs(2092) <= a or b;
    layer2_outputs(2093) <= not a;
    layer2_outputs(2094) <= not (a and b);
    layer2_outputs(2095) <= not a or b;
    layer2_outputs(2096) <= not a;
    layer2_outputs(2097) <= not b;
    layer2_outputs(2098) <= a and not b;
    layer2_outputs(2099) <= a and b;
    layer2_outputs(2100) <= a and not b;
    layer2_outputs(2101) <= not b or a;
    layer2_outputs(2102) <= b and not a;
    layer2_outputs(2103) <= a and b;
    layer2_outputs(2104) <= not a;
    layer2_outputs(2105) <= b;
    layer2_outputs(2106) <= a and b;
    layer2_outputs(2107) <= 1'b1;
    layer2_outputs(2108) <= not a or b;
    layer2_outputs(2109) <= b and not a;
    layer2_outputs(2110) <= b and not a;
    layer2_outputs(2111) <= not b or a;
    layer2_outputs(2112) <= not b or a;
    layer2_outputs(2113) <= not b;
    layer2_outputs(2114) <= b;
    layer2_outputs(2115) <= not b;
    layer2_outputs(2116) <= a and b;
    layer2_outputs(2117) <= a and not b;
    layer2_outputs(2118) <= not b;
    layer2_outputs(2119) <= 1'b1;
    layer2_outputs(2120) <= b;
    layer2_outputs(2121) <= a;
    layer2_outputs(2122) <= not (a and b);
    layer2_outputs(2123) <= not (a or b);
    layer2_outputs(2124) <= 1'b0;
    layer2_outputs(2125) <= not a;
    layer2_outputs(2126) <= a or b;
    layer2_outputs(2127) <= not (a or b);
    layer2_outputs(2128) <= not b or a;
    layer2_outputs(2129) <= not (a and b);
    layer2_outputs(2130) <= a or b;
    layer2_outputs(2131) <= a or b;
    layer2_outputs(2132) <= not (a xor b);
    layer2_outputs(2133) <= a and not b;
    layer2_outputs(2134) <= 1'b0;
    layer2_outputs(2135) <= not (a or b);
    layer2_outputs(2136) <= not a;
    layer2_outputs(2137) <= b;
    layer2_outputs(2138) <= 1'b0;
    layer2_outputs(2139) <= 1'b0;
    layer2_outputs(2140) <= a;
    layer2_outputs(2141) <= b;
    layer2_outputs(2142) <= not a;
    layer2_outputs(2143) <= not a;
    layer2_outputs(2144) <= 1'b0;
    layer2_outputs(2145) <= 1'b0;
    layer2_outputs(2146) <= not (a and b);
    layer2_outputs(2147) <= a;
    layer2_outputs(2148) <= not b or a;
    layer2_outputs(2149) <= a or b;
    layer2_outputs(2150) <= not b;
    layer2_outputs(2151) <= not (a and b);
    layer2_outputs(2152) <= not b or a;
    layer2_outputs(2153) <= 1'b1;
    layer2_outputs(2154) <= not a or b;
    layer2_outputs(2155) <= not (a or b);
    layer2_outputs(2156) <= a and b;
    layer2_outputs(2157) <= a or b;
    layer2_outputs(2158) <= b;
    layer2_outputs(2159) <= not b;
    layer2_outputs(2160) <= a and not b;
    layer2_outputs(2161) <= a and not b;
    layer2_outputs(2162) <= not (a xor b);
    layer2_outputs(2163) <= 1'b0;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= not a or b;
    layer2_outputs(2166) <= 1'b0;
    layer2_outputs(2167) <= not a;
    layer2_outputs(2168) <= not (a and b);
    layer2_outputs(2169) <= not (a or b);
    layer2_outputs(2170) <= a and b;
    layer2_outputs(2171) <= b;
    layer2_outputs(2172) <= a and not b;
    layer2_outputs(2173) <= b;
    layer2_outputs(2174) <= not a or b;
    layer2_outputs(2175) <= not (a or b);
    layer2_outputs(2176) <= not b or a;
    layer2_outputs(2177) <= not b or a;
    layer2_outputs(2178) <= not (a or b);
    layer2_outputs(2179) <= b and not a;
    layer2_outputs(2180) <= b;
    layer2_outputs(2181) <= not a;
    layer2_outputs(2182) <= not b;
    layer2_outputs(2183) <= not (a and b);
    layer2_outputs(2184) <= not (a and b);
    layer2_outputs(2185) <= a and not b;
    layer2_outputs(2186) <= b and not a;
    layer2_outputs(2187) <= a and b;
    layer2_outputs(2188) <= b and not a;
    layer2_outputs(2189) <= a and b;
    layer2_outputs(2190) <= not (a or b);
    layer2_outputs(2191) <= 1'b0;
    layer2_outputs(2192) <= not (a or b);
    layer2_outputs(2193) <= not (a or b);
    layer2_outputs(2194) <= 1'b0;
    layer2_outputs(2195) <= a;
    layer2_outputs(2196) <= b;
    layer2_outputs(2197) <= not a or b;
    layer2_outputs(2198) <= not b or a;
    layer2_outputs(2199) <= b and not a;
    layer2_outputs(2200) <= not a;
    layer2_outputs(2201) <= not b or a;
    layer2_outputs(2202) <= not b;
    layer2_outputs(2203) <= a and not b;
    layer2_outputs(2204) <= not (a or b);
    layer2_outputs(2205) <= 1'b0;
    layer2_outputs(2206) <= not (a and b);
    layer2_outputs(2207) <= not a or b;
    layer2_outputs(2208) <= b;
    layer2_outputs(2209) <= a and b;
    layer2_outputs(2210) <= 1'b1;
    layer2_outputs(2211) <= a and b;
    layer2_outputs(2212) <= 1'b1;
    layer2_outputs(2213) <= not b;
    layer2_outputs(2214) <= not (a and b);
    layer2_outputs(2215) <= 1'b1;
    layer2_outputs(2216) <= a;
    layer2_outputs(2217) <= not (a or b);
    layer2_outputs(2218) <= a and b;
    layer2_outputs(2219) <= a or b;
    layer2_outputs(2220) <= b and not a;
    layer2_outputs(2221) <= not (a and b);
    layer2_outputs(2222) <= not a;
    layer2_outputs(2223) <= a and b;
    layer2_outputs(2224) <= 1'b0;
    layer2_outputs(2225) <= not (a or b);
    layer2_outputs(2226) <= not b or a;
    layer2_outputs(2227) <= not a;
    layer2_outputs(2228) <= not b or a;
    layer2_outputs(2229) <= a and not b;
    layer2_outputs(2230) <= not a;
    layer2_outputs(2231) <= not a or b;
    layer2_outputs(2232) <= not b or a;
    layer2_outputs(2233) <= not (a or b);
    layer2_outputs(2234) <= 1'b0;
    layer2_outputs(2235) <= not a or b;
    layer2_outputs(2236) <= not (a or b);
    layer2_outputs(2237) <= 1'b0;
    layer2_outputs(2238) <= a or b;
    layer2_outputs(2239) <= not (a and b);
    layer2_outputs(2240) <= not (a or b);
    layer2_outputs(2241) <= not b;
    layer2_outputs(2242) <= b and not a;
    layer2_outputs(2243) <= a or b;
    layer2_outputs(2244) <= not a;
    layer2_outputs(2245) <= 1'b1;
    layer2_outputs(2246) <= 1'b0;
    layer2_outputs(2247) <= a;
    layer2_outputs(2248) <= b;
    layer2_outputs(2249) <= not b or a;
    layer2_outputs(2250) <= not (a and b);
    layer2_outputs(2251) <= 1'b1;
    layer2_outputs(2252) <= not (a and b);
    layer2_outputs(2253) <= b;
    layer2_outputs(2254) <= b;
    layer2_outputs(2255) <= not a;
    layer2_outputs(2256) <= not b;
    layer2_outputs(2257) <= b and not a;
    layer2_outputs(2258) <= a and b;
    layer2_outputs(2259) <= 1'b0;
    layer2_outputs(2260) <= b;
    layer2_outputs(2261) <= a and not b;
    layer2_outputs(2262) <= a or b;
    layer2_outputs(2263) <= not a;
    layer2_outputs(2264) <= a and not b;
    layer2_outputs(2265) <= a and not b;
    layer2_outputs(2266) <= a and b;
    layer2_outputs(2267) <= b and not a;
    layer2_outputs(2268) <= not a;
    layer2_outputs(2269) <= a and b;
    layer2_outputs(2270) <= a and b;
    layer2_outputs(2271) <= a xor b;
    layer2_outputs(2272) <= not (a and b);
    layer2_outputs(2273) <= a and b;
    layer2_outputs(2274) <= not (a xor b);
    layer2_outputs(2275) <= not b;
    layer2_outputs(2276) <= not (a xor b);
    layer2_outputs(2277) <= not b;
    layer2_outputs(2278) <= not (a xor b);
    layer2_outputs(2279) <= 1'b0;
    layer2_outputs(2280) <= not b or a;
    layer2_outputs(2281) <= not b or a;
    layer2_outputs(2282) <= 1'b1;
    layer2_outputs(2283) <= not b;
    layer2_outputs(2284) <= not b;
    layer2_outputs(2285) <= not b or a;
    layer2_outputs(2286) <= not (a and b);
    layer2_outputs(2287) <= a or b;
    layer2_outputs(2288) <= 1'b1;
    layer2_outputs(2289) <= 1'b0;
    layer2_outputs(2290) <= a;
    layer2_outputs(2291) <= not (a or b);
    layer2_outputs(2292) <= a and b;
    layer2_outputs(2293) <= not (a xor b);
    layer2_outputs(2294) <= not (a and b);
    layer2_outputs(2295) <= b;
    layer2_outputs(2296) <= a;
    layer2_outputs(2297) <= not b or a;
    layer2_outputs(2298) <= 1'b1;
    layer2_outputs(2299) <= b and not a;
    layer2_outputs(2300) <= not b or a;
    layer2_outputs(2301) <= not (a or b);
    layer2_outputs(2302) <= not (a or b);
    layer2_outputs(2303) <= not a;
    layer2_outputs(2304) <= 1'b1;
    layer2_outputs(2305) <= a;
    layer2_outputs(2306) <= b;
    layer2_outputs(2307) <= not b or a;
    layer2_outputs(2308) <= a xor b;
    layer2_outputs(2309) <= a and not b;
    layer2_outputs(2310) <= not (a or b);
    layer2_outputs(2311) <= not a or b;
    layer2_outputs(2312) <= a and not b;
    layer2_outputs(2313) <= not (a and b);
    layer2_outputs(2314) <= a and b;
    layer2_outputs(2315) <= not (a or b);
    layer2_outputs(2316) <= not a or b;
    layer2_outputs(2317) <= a and not b;
    layer2_outputs(2318) <= not a or b;
    layer2_outputs(2319) <= not a or b;
    layer2_outputs(2320) <= b and not a;
    layer2_outputs(2321) <= not a or b;
    layer2_outputs(2322) <= not b or a;
    layer2_outputs(2323) <= a;
    layer2_outputs(2324) <= a;
    layer2_outputs(2325) <= a xor b;
    layer2_outputs(2326) <= not b or a;
    layer2_outputs(2327) <= b and not a;
    layer2_outputs(2328) <= not b;
    layer2_outputs(2329) <= a or b;
    layer2_outputs(2330) <= not (a and b);
    layer2_outputs(2331) <= 1'b1;
    layer2_outputs(2332) <= 1'b0;
    layer2_outputs(2333) <= 1'b1;
    layer2_outputs(2334) <= not b or a;
    layer2_outputs(2335) <= not b;
    layer2_outputs(2336) <= not (a xor b);
    layer2_outputs(2337) <= a and not b;
    layer2_outputs(2338) <= not a or b;
    layer2_outputs(2339) <= not b or a;
    layer2_outputs(2340) <= 1'b1;
    layer2_outputs(2341) <= a and b;
    layer2_outputs(2342) <= not a or b;
    layer2_outputs(2343) <= b;
    layer2_outputs(2344) <= 1'b1;
    layer2_outputs(2345) <= a;
    layer2_outputs(2346) <= not a or b;
    layer2_outputs(2347) <= b;
    layer2_outputs(2348) <= a and b;
    layer2_outputs(2349) <= a and b;
    layer2_outputs(2350) <= b;
    layer2_outputs(2351) <= not a;
    layer2_outputs(2352) <= 1'b1;
    layer2_outputs(2353) <= a and not b;
    layer2_outputs(2354) <= not (a and b);
    layer2_outputs(2355) <= a or b;
    layer2_outputs(2356) <= not a;
    layer2_outputs(2357) <= b;
    layer2_outputs(2358) <= 1'b1;
    layer2_outputs(2359) <= not b or a;
    layer2_outputs(2360) <= not (a xor b);
    layer2_outputs(2361) <= not a;
    layer2_outputs(2362) <= b and not a;
    layer2_outputs(2363) <= not (a or b);
    layer2_outputs(2364) <= b;
    layer2_outputs(2365) <= 1'b0;
    layer2_outputs(2366) <= 1'b1;
    layer2_outputs(2367) <= not (a or b);
    layer2_outputs(2368) <= a;
    layer2_outputs(2369) <= a or b;
    layer2_outputs(2370) <= 1'b0;
    layer2_outputs(2371) <= a;
    layer2_outputs(2372) <= 1'b0;
    layer2_outputs(2373) <= a or b;
    layer2_outputs(2374) <= a xor b;
    layer2_outputs(2375) <= not b;
    layer2_outputs(2376) <= a and b;
    layer2_outputs(2377) <= a;
    layer2_outputs(2378) <= 1'b1;
    layer2_outputs(2379) <= not b;
    layer2_outputs(2380) <= b and not a;
    layer2_outputs(2381) <= b and not a;
    layer2_outputs(2382) <= a and b;
    layer2_outputs(2383) <= not (a and b);
    layer2_outputs(2384) <= b and not a;
    layer2_outputs(2385) <= a or b;
    layer2_outputs(2386) <= a;
    layer2_outputs(2387) <= not a or b;
    layer2_outputs(2388) <= b;
    layer2_outputs(2389) <= not (a xor b);
    layer2_outputs(2390) <= 1'b0;
    layer2_outputs(2391) <= a xor b;
    layer2_outputs(2392) <= a or b;
    layer2_outputs(2393) <= 1'b1;
    layer2_outputs(2394) <= a or b;
    layer2_outputs(2395) <= b and not a;
    layer2_outputs(2396) <= not (a or b);
    layer2_outputs(2397) <= not (a or b);
    layer2_outputs(2398) <= b;
    layer2_outputs(2399) <= not b;
    layer2_outputs(2400) <= 1'b1;
    layer2_outputs(2401) <= not (a and b);
    layer2_outputs(2402) <= not b or a;
    layer2_outputs(2403) <= not (a and b);
    layer2_outputs(2404) <= not (a or b);
    layer2_outputs(2405) <= not b or a;
    layer2_outputs(2406) <= 1'b0;
    layer2_outputs(2407) <= a and not b;
    layer2_outputs(2408) <= 1'b1;
    layer2_outputs(2409) <= b and not a;
    layer2_outputs(2410) <= a or b;
    layer2_outputs(2411) <= a and not b;
    layer2_outputs(2412) <= not a;
    layer2_outputs(2413) <= 1'b1;
    layer2_outputs(2414) <= a xor b;
    layer2_outputs(2415) <= not (a or b);
    layer2_outputs(2416) <= not (a or b);
    layer2_outputs(2417) <= not a;
    layer2_outputs(2418) <= a and not b;
    layer2_outputs(2419) <= b and not a;
    layer2_outputs(2420) <= 1'b0;
    layer2_outputs(2421) <= not b or a;
    layer2_outputs(2422) <= b and not a;
    layer2_outputs(2423) <= 1'b1;
    layer2_outputs(2424) <= a and b;
    layer2_outputs(2425) <= not a;
    layer2_outputs(2426) <= a and b;
    layer2_outputs(2427) <= b;
    layer2_outputs(2428) <= 1'b1;
    layer2_outputs(2429) <= not b or a;
    layer2_outputs(2430) <= a and not b;
    layer2_outputs(2431) <= a;
    layer2_outputs(2432) <= not (a xor b);
    layer2_outputs(2433) <= not b or a;
    layer2_outputs(2434) <= not a;
    layer2_outputs(2435) <= 1'b1;
    layer2_outputs(2436) <= 1'b0;
    layer2_outputs(2437) <= not a or b;
    layer2_outputs(2438) <= not a or b;
    layer2_outputs(2439) <= not (a or b);
    layer2_outputs(2440) <= a and b;
    layer2_outputs(2441) <= 1'b0;
    layer2_outputs(2442) <= b;
    layer2_outputs(2443) <= a and b;
    layer2_outputs(2444) <= a and not b;
    layer2_outputs(2445) <= not b or a;
    layer2_outputs(2446) <= b;
    layer2_outputs(2447) <= 1'b0;
    layer2_outputs(2448) <= not (a and b);
    layer2_outputs(2449) <= b and not a;
    layer2_outputs(2450) <= a or b;
    layer2_outputs(2451) <= b;
    layer2_outputs(2452) <= not b or a;
    layer2_outputs(2453) <= 1'b1;
    layer2_outputs(2454) <= b and not a;
    layer2_outputs(2455) <= not a or b;
    layer2_outputs(2456) <= not b;
    layer2_outputs(2457) <= not a or b;
    layer2_outputs(2458) <= not (a or b);
    layer2_outputs(2459) <= b;
    layer2_outputs(2460) <= not a or b;
    layer2_outputs(2461) <= not a or b;
    layer2_outputs(2462) <= a and not b;
    layer2_outputs(2463) <= not (a and b);
    layer2_outputs(2464) <= a or b;
    layer2_outputs(2465) <= a or b;
    layer2_outputs(2466) <= not a or b;
    layer2_outputs(2467) <= b and not a;
    layer2_outputs(2468) <= a;
    layer2_outputs(2469) <= a xor b;
    layer2_outputs(2470) <= a and b;
    layer2_outputs(2471) <= not (a or b);
    layer2_outputs(2472) <= a;
    layer2_outputs(2473) <= not (a and b);
    layer2_outputs(2474) <= 1'b1;
    layer2_outputs(2475) <= not b or a;
    layer2_outputs(2476) <= a xor b;
    layer2_outputs(2477) <= b and not a;
    layer2_outputs(2478) <= a;
    layer2_outputs(2479) <= 1'b0;
    layer2_outputs(2480) <= 1'b0;
    layer2_outputs(2481) <= not a or b;
    layer2_outputs(2482) <= a or b;
    layer2_outputs(2483) <= not a;
    layer2_outputs(2484) <= 1'b1;
    layer2_outputs(2485) <= not (a or b);
    layer2_outputs(2486) <= a;
    layer2_outputs(2487) <= 1'b1;
    layer2_outputs(2488) <= not (a or b);
    layer2_outputs(2489) <= not a or b;
    layer2_outputs(2490) <= a or b;
    layer2_outputs(2491) <= b and not a;
    layer2_outputs(2492) <= a and not b;
    layer2_outputs(2493) <= a and b;
    layer2_outputs(2494) <= a;
    layer2_outputs(2495) <= not (a or b);
    layer2_outputs(2496) <= not (a or b);
    layer2_outputs(2497) <= 1'b1;
    layer2_outputs(2498) <= a and not b;
    layer2_outputs(2499) <= b and not a;
    layer2_outputs(2500) <= not b;
    layer2_outputs(2501) <= 1'b0;
    layer2_outputs(2502) <= b;
    layer2_outputs(2503) <= not a;
    layer2_outputs(2504) <= 1'b0;
    layer2_outputs(2505) <= not b or a;
    layer2_outputs(2506) <= a or b;
    layer2_outputs(2507) <= not (a xor b);
    layer2_outputs(2508) <= not (a xor b);
    layer2_outputs(2509) <= a xor b;
    layer2_outputs(2510) <= not a;
    layer2_outputs(2511) <= 1'b1;
    layer2_outputs(2512) <= not b or a;
    layer2_outputs(2513) <= 1'b0;
    layer2_outputs(2514) <= a or b;
    layer2_outputs(2515) <= 1'b0;
    layer2_outputs(2516) <= not b;
    layer2_outputs(2517) <= not a;
    layer2_outputs(2518) <= 1'b0;
    layer2_outputs(2519) <= a and b;
    layer2_outputs(2520) <= 1'b1;
    layer2_outputs(2521) <= b and not a;
    layer2_outputs(2522) <= not (a or b);
    layer2_outputs(2523) <= not (a or b);
    layer2_outputs(2524) <= a and b;
    layer2_outputs(2525) <= not (a and b);
    layer2_outputs(2526) <= not (a or b);
    layer2_outputs(2527) <= not a;
    layer2_outputs(2528) <= not b;
    layer2_outputs(2529) <= not (a xor b);
    layer2_outputs(2530) <= a;
    layer2_outputs(2531) <= b;
    layer2_outputs(2532) <= not (a and b);
    layer2_outputs(2533) <= not b or a;
    layer2_outputs(2534) <= b;
    layer2_outputs(2535) <= not b;
    layer2_outputs(2536) <= not b or a;
    layer2_outputs(2537) <= a and b;
    layer2_outputs(2538) <= b;
    layer2_outputs(2539) <= not (a and b);
    layer2_outputs(2540) <= a;
    layer2_outputs(2541) <= a and not b;
    layer2_outputs(2542) <= a or b;
    layer2_outputs(2543) <= a;
    layer2_outputs(2544) <= not b or a;
    layer2_outputs(2545) <= not b or a;
    layer2_outputs(2546) <= not a or b;
    layer2_outputs(2547) <= not a;
    layer2_outputs(2548) <= not b;
    layer2_outputs(2549) <= a or b;
    layer2_outputs(2550) <= not (a and b);
    layer2_outputs(2551) <= a or b;
    layer2_outputs(2552) <= a and not b;
    layer2_outputs(2553) <= not a or b;
    layer2_outputs(2554) <= not b or a;
    layer2_outputs(2555) <= a or b;
    layer2_outputs(2556) <= a and not b;
    layer2_outputs(2557) <= not b or a;
    layer2_outputs(2558) <= not (a xor b);
    layer2_outputs(2559) <= not (a or b);
    layer2_outputs(2560) <= not a;
    layer2_outputs(2561) <= not (a xor b);
    layer2_outputs(2562) <= b and not a;
    layer2_outputs(2563) <= not b or a;
    layer2_outputs(2564) <= a and b;
    layer2_outputs(2565) <= b and not a;
    layer2_outputs(2566) <= not (a or b);
    layer2_outputs(2567) <= 1'b0;
    layer2_outputs(2568) <= a;
    layer2_outputs(2569) <= 1'b1;
    layer2_outputs(2570) <= not (a and b);
    layer2_outputs(2571) <= a and b;
    layer2_outputs(2572) <= 1'b0;
    layer2_outputs(2573) <= 1'b1;
    layer2_outputs(2574) <= not a;
    layer2_outputs(2575) <= 1'b0;
    layer2_outputs(2576) <= b and not a;
    layer2_outputs(2577) <= not (a and b);
    layer2_outputs(2578) <= not a or b;
    layer2_outputs(2579) <= not b;
    layer2_outputs(2580) <= not a or b;
    layer2_outputs(2581) <= a xor b;
    layer2_outputs(2582) <= not a or b;
    layer2_outputs(2583) <= a and b;
    layer2_outputs(2584) <= not a;
    layer2_outputs(2585) <= not b;
    layer2_outputs(2586) <= a xor b;
    layer2_outputs(2587) <= not a;
    layer2_outputs(2588) <= not (a and b);
    layer2_outputs(2589) <= 1'b1;
    layer2_outputs(2590) <= 1'b1;
    layer2_outputs(2591) <= a or b;
    layer2_outputs(2592) <= a or b;
    layer2_outputs(2593) <= not b;
    layer2_outputs(2594) <= not (a or b);
    layer2_outputs(2595) <= a or b;
    layer2_outputs(2596) <= not b or a;
    layer2_outputs(2597) <= not a or b;
    layer2_outputs(2598) <= not a;
    layer2_outputs(2599) <= b and not a;
    layer2_outputs(2600) <= a;
    layer2_outputs(2601) <= b and not a;
    layer2_outputs(2602) <= a or b;
    layer2_outputs(2603) <= a and b;
    layer2_outputs(2604) <= b;
    layer2_outputs(2605) <= not b;
    layer2_outputs(2606) <= not (a and b);
    layer2_outputs(2607) <= not a;
    layer2_outputs(2608) <= 1'b0;
    layer2_outputs(2609) <= b;
    layer2_outputs(2610) <= not a;
    layer2_outputs(2611) <= not (a or b);
    layer2_outputs(2612) <= not a or b;
    layer2_outputs(2613) <= a and not b;
    layer2_outputs(2614) <= a and b;
    layer2_outputs(2615) <= a and not b;
    layer2_outputs(2616) <= a and b;
    layer2_outputs(2617) <= b and not a;
    layer2_outputs(2618) <= not a;
    layer2_outputs(2619) <= a;
    layer2_outputs(2620) <= a or b;
    layer2_outputs(2621) <= a and not b;
    layer2_outputs(2622) <= not b or a;
    layer2_outputs(2623) <= not b;
    layer2_outputs(2624) <= 1'b1;
    layer2_outputs(2625) <= not a;
    layer2_outputs(2626) <= not b;
    layer2_outputs(2627) <= not (a or b);
    layer2_outputs(2628) <= a;
    layer2_outputs(2629) <= not (a xor b);
    layer2_outputs(2630) <= not b or a;
    layer2_outputs(2631) <= b and not a;
    layer2_outputs(2632) <= 1'b1;
    layer2_outputs(2633) <= a and not b;
    layer2_outputs(2634) <= a and b;
    layer2_outputs(2635) <= not (a and b);
    layer2_outputs(2636) <= b and not a;
    layer2_outputs(2637) <= a and b;
    layer2_outputs(2638) <= b;
    layer2_outputs(2639) <= 1'b1;
    layer2_outputs(2640) <= 1'b1;
    layer2_outputs(2641) <= a xor b;
    layer2_outputs(2642) <= not b;
    layer2_outputs(2643) <= a;
    layer2_outputs(2644) <= 1'b1;
    layer2_outputs(2645) <= a or b;
    layer2_outputs(2646) <= a and not b;
    layer2_outputs(2647) <= a;
    layer2_outputs(2648) <= not b;
    layer2_outputs(2649) <= not (a and b);
    layer2_outputs(2650) <= not (a and b);
    layer2_outputs(2651) <= a and b;
    layer2_outputs(2652) <= 1'b1;
    layer2_outputs(2653) <= a or b;
    layer2_outputs(2654) <= b and not a;
    layer2_outputs(2655) <= a or b;
    layer2_outputs(2656) <= not (a or b);
    layer2_outputs(2657) <= a and b;
    layer2_outputs(2658) <= 1'b1;
    layer2_outputs(2659) <= not b or a;
    layer2_outputs(2660) <= a or b;
    layer2_outputs(2661) <= not (a and b);
    layer2_outputs(2662) <= a;
    layer2_outputs(2663) <= not a or b;
    layer2_outputs(2664) <= not (a and b);
    layer2_outputs(2665) <= 1'b0;
    layer2_outputs(2666) <= not (a or b);
    layer2_outputs(2667) <= b;
    layer2_outputs(2668) <= b;
    layer2_outputs(2669) <= not (a xor b);
    layer2_outputs(2670) <= a;
    layer2_outputs(2671) <= not b or a;
    layer2_outputs(2672) <= a and b;
    layer2_outputs(2673) <= not a;
    layer2_outputs(2674) <= a;
    layer2_outputs(2675) <= a and not b;
    layer2_outputs(2676) <= a;
    layer2_outputs(2677) <= not b or a;
    layer2_outputs(2678) <= 1'b0;
    layer2_outputs(2679) <= a or b;
    layer2_outputs(2680) <= not b;
    layer2_outputs(2681) <= b;
    layer2_outputs(2682) <= not a or b;
    layer2_outputs(2683) <= 1'b0;
    layer2_outputs(2684) <= b;
    layer2_outputs(2685) <= 1'b1;
    layer2_outputs(2686) <= not b or a;
    layer2_outputs(2687) <= not (a or b);
    layer2_outputs(2688) <= a;
    layer2_outputs(2689) <= b;
    layer2_outputs(2690) <= 1'b1;
    layer2_outputs(2691) <= 1'b0;
    layer2_outputs(2692) <= not b or a;
    layer2_outputs(2693) <= 1'b0;
    layer2_outputs(2694) <= not a or b;
    layer2_outputs(2695) <= not (a or b);
    layer2_outputs(2696) <= not a or b;
    layer2_outputs(2697) <= not a or b;
    layer2_outputs(2698) <= not a;
    layer2_outputs(2699) <= a and b;
    layer2_outputs(2700) <= a or b;
    layer2_outputs(2701) <= a and b;
    layer2_outputs(2702) <= a and not b;
    layer2_outputs(2703) <= 1'b1;
    layer2_outputs(2704) <= a and b;
    layer2_outputs(2705) <= 1'b1;
    layer2_outputs(2706) <= 1'b1;
    layer2_outputs(2707) <= not a or b;
    layer2_outputs(2708) <= a;
    layer2_outputs(2709) <= 1'b1;
    layer2_outputs(2710) <= a or b;
    layer2_outputs(2711) <= not b or a;
    layer2_outputs(2712) <= b;
    layer2_outputs(2713) <= not a;
    layer2_outputs(2714) <= 1'b1;
    layer2_outputs(2715) <= not a;
    layer2_outputs(2716) <= 1'b1;
    layer2_outputs(2717) <= not b;
    layer2_outputs(2718) <= 1'b1;
    layer2_outputs(2719) <= not (a or b);
    layer2_outputs(2720) <= 1'b0;
    layer2_outputs(2721) <= not (a and b);
    layer2_outputs(2722) <= 1'b1;
    layer2_outputs(2723) <= not b;
    layer2_outputs(2724) <= a and b;
    layer2_outputs(2725) <= a and b;
    layer2_outputs(2726) <= 1'b1;
    layer2_outputs(2727) <= a and b;
    layer2_outputs(2728) <= not (a or b);
    layer2_outputs(2729) <= a;
    layer2_outputs(2730) <= not (a or b);
    layer2_outputs(2731) <= not (a or b);
    layer2_outputs(2732) <= a xor b;
    layer2_outputs(2733) <= a and not b;
    layer2_outputs(2734) <= a xor b;
    layer2_outputs(2735) <= b and not a;
    layer2_outputs(2736) <= 1'b0;
    layer2_outputs(2737) <= 1'b0;
    layer2_outputs(2738) <= not b or a;
    layer2_outputs(2739) <= a;
    layer2_outputs(2740) <= b and not a;
    layer2_outputs(2741) <= not b or a;
    layer2_outputs(2742) <= a;
    layer2_outputs(2743) <= not b or a;
    layer2_outputs(2744) <= b and not a;
    layer2_outputs(2745) <= 1'b0;
    layer2_outputs(2746) <= not a or b;
    layer2_outputs(2747) <= a or b;
    layer2_outputs(2748) <= a and b;
    layer2_outputs(2749) <= not (a or b);
    layer2_outputs(2750) <= not (a and b);
    layer2_outputs(2751) <= not b;
    layer2_outputs(2752) <= not b;
    layer2_outputs(2753) <= not b or a;
    layer2_outputs(2754) <= a xor b;
    layer2_outputs(2755) <= not b;
    layer2_outputs(2756) <= b;
    layer2_outputs(2757) <= not b;
    layer2_outputs(2758) <= not (a or b);
    layer2_outputs(2759) <= not (a or b);
    layer2_outputs(2760) <= not a;
    layer2_outputs(2761) <= a and not b;
    layer2_outputs(2762) <= a;
    layer2_outputs(2763) <= 1'b1;
    layer2_outputs(2764) <= not a;
    layer2_outputs(2765) <= b;
    layer2_outputs(2766) <= a or b;
    layer2_outputs(2767) <= a and not b;
    layer2_outputs(2768) <= a and not b;
    layer2_outputs(2769) <= 1'b1;
    layer2_outputs(2770) <= a;
    layer2_outputs(2771) <= a or b;
    layer2_outputs(2772) <= 1'b1;
    layer2_outputs(2773) <= not a or b;
    layer2_outputs(2774) <= not b or a;
    layer2_outputs(2775) <= not a;
    layer2_outputs(2776) <= not a;
    layer2_outputs(2777) <= not a or b;
    layer2_outputs(2778) <= a or b;
    layer2_outputs(2779) <= not a or b;
    layer2_outputs(2780) <= not (a or b);
    layer2_outputs(2781) <= not (a or b);
    layer2_outputs(2782) <= not (a and b);
    layer2_outputs(2783) <= not a;
    layer2_outputs(2784) <= not (a or b);
    layer2_outputs(2785) <= b and not a;
    layer2_outputs(2786) <= a and not b;
    layer2_outputs(2787) <= not b;
    layer2_outputs(2788) <= 1'b1;
    layer2_outputs(2789) <= not a;
    layer2_outputs(2790) <= b and not a;
    layer2_outputs(2791) <= b and not a;
    layer2_outputs(2792) <= not a;
    layer2_outputs(2793) <= 1'b0;
    layer2_outputs(2794) <= 1'b0;
    layer2_outputs(2795) <= not b or a;
    layer2_outputs(2796) <= b and not a;
    layer2_outputs(2797) <= not (a xor b);
    layer2_outputs(2798) <= not b or a;
    layer2_outputs(2799) <= b;
    layer2_outputs(2800) <= a and b;
    layer2_outputs(2801) <= not (a or b);
    layer2_outputs(2802) <= a and not b;
    layer2_outputs(2803) <= not (a and b);
    layer2_outputs(2804) <= 1'b0;
    layer2_outputs(2805) <= 1'b1;
    layer2_outputs(2806) <= a and b;
    layer2_outputs(2807) <= 1'b0;
    layer2_outputs(2808) <= a or b;
    layer2_outputs(2809) <= 1'b1;
    layer2_outputs(2810) <= not (a or b);
    layer2_outputs(2811) <= b;
    layer2_outputs(2812) <= not b;
    layer2_outputs(2813) <= b;
    layer2_outputs(2814) <= b and not a;
    layer2_outputs(2815) <= a;
    layer2_outputs(2816) <= b and not a;
    layer2_outputs(2817) <= not b or a;
    layer2_outputs(2818) <= not a or b;
    layer2_outputs(2819) <= not (a or b);
    layer2_outputs(2820) <= not a;
    layer2_outputs(2821) <= not b or a;
    layer2_outputs(2822) <= not (a or b);
    layer2_outputs(2823) <= 1'b0;
    layer2_outputs(2824) <= b and not a;
    layer2_outputs(2825) <= b and not a;
    layer2_outputs(2826) <= not b or a;
    layer2_outputs(2827) <= not a or b;
    layer2_outputs(2828) <= not b or a;
    layer2_outputs(2829) <= a or b;
    layer2_outputs(2830) <= a and not b;
    layer2_outputs(2831) <= 1'b1;
    layer2_outputs(2832) <= a and not b;
    layer2_outputs(2833) <= not (a or b);
    layer2_outputs(2834) <= not (a and b);
    layer2_outputs(2835) <= a and not b;
    layer2_outputs(2836) <= 1'b0;
    layer2_outputs(2837) <= a and not b;
    layer2_outputs(2838) <= not b;
    layer2_outputs(2839) <= a or b;
    layer2_outputs(2840) <= 1'b1;
    layer2_outputs(2841) <= not b;
    layer2_outputs(2842) <= 1'b1;
    layer2_outputs(2843) <= 1'b0;
    layer2_outputs(2844) <= a and not b;
    layer2_outputs(2845) <= a and b;
    layer2_outputs(2846) <= a xor b;
    layer2_outputs(2847) <= 1'b1;
    layer2_outputs(2848) <= a;
    layer2_outputs(2849) <= a and not b;
    layer2_outputs(2850) <= a and not b;
    layer2_outputs(2851) <= 1'b0;
    layer2_outputs(2852) <= not b or a;
    layer2_outputs(2853) <= not (a and b);
    layer2_outputs(2854) <= not b;
    layer2_outputs(2855) <= a;
    layer2_outputs(2856) <= a;
    layer2_outputs(2857) <= 1'b0;
    layer2_outputs(2858) <= not b;
    layer2_outputs(2859) <= not a;
    layer2_outputs(2860) <= not b or a;
    layer2_outputs(2861) <= 1'b0;
    layer2_outputs(2862) <= a;
    layer2_outputs(2863) <= not (a and b);
    layer2_outputs(2864) <= not (a and b);
    layer2_outputs(2865) <= b and not a;
    layer2_outputs(2866) <= not (a or b);
    layer2_outputs(2867) <= not (a and b);
    layer2_outputs(2868) <= a and b;
    layer2_outputs(2869) <= a and b;
    layer2_outputs(2870) <= 1'b0;
    layer2_outputs(2871) <= b and not a;
    layer2_outputs(2872) <= a xor b;
    layer2_outputs(2873) <= not (a or b);
    layer2_outputs(2874) <= not a;
    layer2_outputs(2875) <= 1'b1;
    layer2_outputs(2876) <= a and not b;
    layer2_outputs(2877) <= a and b;
    layer2_outputs(2878) <= a or b;
    layer2_outputs(2879) <= b and not a;
    layer2_outputs(2880) <= 1'b1;
    layer2_outputs(2881) <= a and b;
    layer2_outputs(2882) <= a or b;
    layer2_outputs(2883) <= a xor b;
    layer2_outputs(2884) <= a and b;
    layer2_outputs(2885) <= a and not b;
    layer2_outputs(2886) <= not a or b;
    layer2_outputs(2887) <= 1'b0;
    layer2_outputs(2888) <= not (a and b);
    layer2_outputs(2889) <= not (a or b);
    layer2_outputs(2890) <= not a;
    layer2_outputs(2891) <= not b or a;
    layer2_outputs(2892) <= not (a xor b);
    layer2_outputs(2893) <= a and not b;
    layer2_outputs(2894) <= b and not a;
    layer2_outputs(2895) <= a;
    layer2_outputs(2896) <= a and not b;
    layer2_outputs(2897) <= not b or a;
    layer2_outputs(2898) <= 1'b1;
    layer2_outputs(2899) <= not b;
    layer2_outputs(2900) <= b;
    layer2_outputs(2901) <= not b;
    layer2_outputs(2902) <= 1'b0;
    layer2_outputs(2903) <= 1'b0;
    layer2_outputs(2904) <= not (a or b);
    layer2_outputs(2905) <= b;
    layer2_outputs(2906) <= a or b;
    layer2_outputs(2907) <= 1'b1;
    layer2_outputs(2908) <= b;
    layer2_outputs(2909) <= 1'b0;
    layer2_outputs(2910) <= not a or b;
    layer2_outputs(2911) <= not a or b;
    layer2_outputs(2912) <= a or b;
    layer2_outputs(2913) <= not a;
    layer2_outputs(2914) <= a and b;
    layer2_outputs(2915) <= a and b;
    layer2_outputs(2916) <= 1'b0;
    layer2_outputs(2917) <= a and not b;
    layer2_outputs(2918) <= a;
    layer2_outputs(2919) <= a and b;
    layer2_outputs(2920) <= a and not b;
    layer2_outputs(2921) <= a or b;
    layer2_outputs(2922) <= 1'b1;
    layer2_outputs(2923) <= 1'b1;
    layer2_outputs(2924) <= not (a and b);
    layer2_outputs(2925) <= not b or a;
    layer2_outputs(2926) <= not (a and b);
    layer2_outputs(2927) <= a or b;
    layer2_outputs(2928) <= b;
    layer2_outputs(2929) <= not b or a;
    layer2_outputs(2930) <= not b;
    layer2_outputs(2931) <= a and not b;
    layer2_outputs(2932) <= 1'b0;
    layer2_outputs(2933) <= 1'b0;
    layer2_outputs(2934) <= b and not a;
    layer2_outputs(2935) <= not (a xor b);
    layer2_outputs(2936) <= not a or b;
    layer2_outputs(2937) <= not b or a;
    layer2_outputs(2938) <= not (a and b);
    layer2_outputs(2939) <= b and not a;
    layer2_outputs(2940) <= 1'b1;
    layer2_outputs(2941) <= a and not b;
    layer2_outputs(2942) <= not a or b;
    layer2_outputs(2943) <= 1'b1;
    layer2_outputs(2944) <= 1'b1;
    layer2_outputs(2945) <= not b;
    layer2_outputs(2946) <= a or b;
    layer2_outputs(2947) <= a or b;
    layer2_outputs(2948) <= not b;
    layer2_outputs(2949) <= a and b;
    layer2_outputs(2950) <= a and b;
    layer2_outputs(2951) <= a and not b;
    layer2_outputs(2952) <= a and not b;
    layer2_outputs(2953) <= not (a or b);
    layer2_outputs(2954) <= 1'b1;
    layer2_outputs(2955) <= a and b;
    layer2_outputs(2956) <= a and not b;
    layer2_outputs(2957) <= a or b;
    layer2_outputs(2958) <= not a;
    layer2_outputs(2959) <= b;
    layer2_outputs(2960) <= not b or a;
    layer2_outputs(2961) <= not (a and b);
    layer2_outputs(2962) <= a;
    layer2_outputs(2963) <= a or b;
    layer2_outputs(2964) <= 1'b1;
    layer2_outputs(2965) <= not (a or b);
    layer2_outputs(2966) <= not (a xor b);
    layer2_outputs(2967) <= b and not a;
    layer2_outputs(2968) <= not (a or b);
    layer2_outputs(2969) <= b;
    layer2_outputs(2970) <= a or b;
    layer2_outputs(2971) <= not (a xor b);
    layer2_outputs(2972) <= not a;
    layer2_outputs(2973) <= not (a and b);
    layer2_outputs(2974) <= a and not b;
    layer2_outputs(2975) <= 1'b1;
    layer2_outputs(2976) <= 1'b0;
    layer2_outputs(2977) <= not a;
    layer2_outputs(2978) <= 1'b1;
    layer2_outputs(2979) <= a and not b;
    layer2_outputs(2980) <= not b or a;
    layer2_outputs(2981) <= a and b;
    layer2_outputs(2982) <= not a or b;
    layer2_outputs(2983) <= a;
    layer2_outputs(2984) <= not (a xor b);
    layer2_outputs(2985) <= a or b;
    layer2_outputs(2986) <= not b or a;
    layer2_outputs(2987) <= a and not b;
    layer2_outputs(2988) <= a;
    layer2_outputs(2989) <= not a;
    layer2_outputs(2990) <= not a;
    layer2_outputs(2991) <= a and not b;
    layer2_outputs(2992) <= not a;
    layer2_outputs(2993) <= b and not a;
    layer2_outputs(2994) <= not b or a;
    layer2_outputs(2995) <= a or b;
    layer2_outputs(2996) <= not (a and b);
    layer2_outputs(2997) <= not a;
    layer2_outputs(2998) <= a or b;
    layer2_outputs(2999) <= a and b;
    layer2_outputs(3000) <= a or b;
    layer2_outputs(3001) <= not (a or b);
    layer2_outputs(3002) <= not (a and b);
    layer2_outputs(3003) <= a or b;
    layer2_outputs(3004) <= a and b;
    layer2_outputs(3005) <= b and not a;
    layer2_outputs(3006) <= not (a and b);
    layer2_outputs(3007) <= not b;
    layer2_outputs(3008) <= not (a and b);
    layer2_outputs(3009) <= not b;
    layer2_outputs(3010) <= not b;
    layer2_outputs(3011) <= not (a or b);
    layer2_outputs(3012) <= not a;
    layer2_outputs(3013) <= not a or b;
    layer2_outputs(3014) <= not a or b;
    layer2_outputs(3015) <= b and not a;
    layer2_outputs(3016) <= not a;
    layer2_outputs(3017) <= not (a or b);
    layer2_outputs(3018) <= b;
    layer2_outputs(3019) <= 1'b0;
    layer2_outputs(3020) <= b and not a;
    layer2_outputs(3021) <= not b;
    layer2_outputs(3022) <= 1'b1;
    layer2_outputs(3023) <= not a;
    layer2_outputs(3024) <= not b;
    layer2_outputs(3025) <= 1'b0;
    layer2_outputs(3026) <= not b;
    layer2_outputs(3027) <= not a or b;
    layer2_outputs(3028) <= 1'b1;
    layer2_outputs(3029) <= not (a and b);
    layer2_outputs(3030) <= 1'b0;
    layer2_outputs(3031) <= not (a and b);
    layer2_outputs(3032) <= not (a or b);
    layer2_outputs(3033) <= a or b;
    layer2_outputs(3034) <= not (a or b);
    layer2_outputs(3035) <= not a;
    layer2_outputs(3036) <= a;
    layer2_outputs(3037) <= not (a or b);
    layer2_outputs(3038) <= not a or b;
    layer2_outputs(3039) <= a and not b;
    layer2_outputs(3040) <= not b or a;
    layer2_outputs(3041) <= a or b;
    layer2_outputs(3042) <= 1'b0;
    layer2_outputs(3043) <= 1'b0;
    layer2_outputs(3044) <= a xor b;
    layer2_outputs(3045) <= b and not a;
    layer2_outputs(3046) <= not b or a;
    layer2_outputs(3047) <= not b or a;
    layer2_outputs(3048) <= not (a or b);
    layer2_outputs(3049) <= a;
    layer2_outputs(3050) <= a or b;
    layer2_outputs(3051) <= a or b;
    layer2_outputs(3052) <= a xor b;
    layer2_outputs(3053) <= 1'b1;
    layer2_outputs(3054) <= b;
    layer2_outputs(3055) <= not b or a;
    layer2_outputs(3056) <= not (a and b);
    layer2_outputs(3057) <= a and not b;
    layer2_outputs(3058) <= a and b;
    layer2_outputs(3059) <= not b;
    layer2_outputs(3060) <= not a;
    layer2_outputs(3061) <= 1'b1;
    layer2_outputs(3062) <= 1'b0;
    layer2_outputs(3063) <= a and not b;
    layer2_outputs(3064) <= a;
    layer2_outputs(3065) <= 1'b0;
    layer2_outputs(3066) <= not (a xor b);
    layer2_outputs(3067) <= not a;
    layer2_outputs(3068) <= a;
    layer2_outputs(3069) <= a or b;
    layer2_outputs(3070) <= 1'b0;
    layer2_outputs(3071) <= a and b;
    layer2_outputs(3072) <= 1'b1;
    layer2_outputs(3073) <= not b;
    layer2_outputs(3074) <= not b or a;
    layer2_outputs(3075) <= b;
    layer2_outputs(3076) <= not b;
    layer2_outputs(3077) <= not a;
    layer2_outputs(3078) <= a or b;
    layer2_outputs(3079) <= not (a and b);
    layer2_outputs(3080) <= not (a or b);
    layer2_outputs(3081) <= b and not a;
    layer2_outputs(3082) <= a xor b;
    layer2_outputs(3083) <= not a;
    layer2_outputs(3084) <= a and not b;
    layer2_outputs(3085) <= not b or a;
    layer2_outputs(3086) <= a;
    layer2_outputs(3087) <= not (a and b);
    layer2_outputs(3088) <= a;
    layer2_outputs(3089) <= b and not a;
    layer2_outputs(3090) <= not b;
    layer2_outputs(3091) <= not a;
    layer2_outputs(3092) <= not (a and b);
    layer2_outputs(3093) <= a;
    layer2_outputs(3094) <= not b;
    layer2_outputs(3095) <= a;
    layer2_outputs(3096) <= b and not a;
    layer2_outputs(3097) <= not a or b;
    layer2_outputs(3098) <= a or b;
    layer2_outputs(3099) <= a xor b;
    layer2_outputs(3100) <= not a or b;
    layer2_outputs(3101) <= a xor b;
    layer2_outputs(3102) <= not a;
    layer2_outputs(3103) <= a;
    layer2_outputs(3104) <= a and b;
    layer2_outputs(3105) <= not a or b;
    layer2_outputs(3106) <= a;
    layer2_outputs(3107) <= not a or b;
    layer2_outputs(3108) <= not a or b;
    layer2_outputs(3109) <= a and b;
    layer2_outputs(3110) <= not (a xor b);
    layer2_outputs(3111) <= a xor b;
    layer2_outputs(3112) <= not a or b;
    layer2_outputs(3113) <= not b or a;
    layer2_outputs(3114) <= a or b;
    layer2_outputs(3115) <= not (a or b);
    layer2_outputs(3116) <= not (a or b);
    layer2_outputs(3117) <= not a or b;
    layer2_outputs(3118) <= not b;
    layer2_outputs(3119) <= b and not a;
    layer2_outputs(3120) <= a and b;
    layer2_outputs(3121) <= 1'b0;
    layer2_outputs(3122) <= not b;
    layer2_outputs(3123) <= not (a and b);
    layer2_outputs(3124) <= not a or b;
    layer2_outputs(3125) <= a xor b;
    layer2_outputs(3126) <= b;
    layer2_outputs(3127) <= a;
    layer2_outputs(3128) <= not (a and b);
    layer2_outputs(3129) <= not (a and b);
    layer2_outputs(3130) <= 1'b0;
    layer2_outputs(3131) <= not a or b;
    layer2_outputs(3132) <= 1'b0;
    layer2_outputs(3133) <= not a;
    layer2_outputs(3134) <= a and b;
    layer2_outputs(3135) <= not b;
    layer2_outputs(3136) <= not (a or b);
    layer2_outputs(3137) <= a and b;
    layer2_outputs(3138) <= b and not a;
    layer2_outputs(3139) <= a and not b;
    layer2_outputs(3140) <= not (a and b);
    layer2_outputs(3141) <= not b or a;
    layer2_outputs(3142) <= b;
    layer2_outputs(3143) <= 1'b1;
    layer2_outputs(3144) <= not b or a;
    layer2_outputs(3145) <= not (a xor b);
    layer2_outputs(3146) <= 1'b0;
    layer2_outputs(3147) <= 1'b0;
    layer2_outputs(3148) <= not a;
    layer2_outputs(3149) <= a;
    layer2_outputs(3150) <= not (a and b);
    layer2_outputs(3151) <= not b;
    layer2_outputs(3152) <= a xor b;
    layer2_outputs(3153) <= not (a and b);
    layer2_outputs(3154) <= not a;
    layer2_outputs(3155) <= not (a xor b);
    layer2_outputs(3156) <= 1'b1;
    layer2_outputs(3157) <= 1'b0;
    layer2_outputs(3158) <= not b or a;
    layer2_outputs(3159) <= a xor b;
    layer2_outputs(3160) <= not (a or b);
    layer2_outputs(3161) <= not a;
    layer2_outputs(3162) <= b;
    layer2_outputs(3163) <= a and not b;
    layer2_outputs(3164) <= not a;
    layer2_outputs(3165) <= a or b;
    layer2_outputs(3166) <= not (a and b);
    layer2_outputs(3167) <= not a or b;
    layer2_outputs(3168) <= not b or a;
    layer2_outputs(3169) <= not (a and b);
    layer2_outputs(3170) <= not (a or b);
    layer2_outputs(3171) <= b;
    layer2_outputs(3172) <= a or b;
    layer2_outputs(3173) <= b and not a;
    layer2_outputs(3174) <= a or b;
    layer2_outputs(3175) <= a xor b;
    layer2_outputs(3176) <= not (a or b);
    layer2_outputs(3177) <= not (a or b);
    layer2_outputs(3178) <= a and b;
    layer2_outputs(3179) <= not (a or b);
    layer2_outputs(3180) <= not a;
    layer2_outputs(3181) <= not b;
    layer2_outputs(3182) <= not a;
    layer2_outputs(3183) <= 1'b0;
    layer2_outputs(3184) <= 1'b1;
    layer2_outputs(3185) <= not b or a;
    layer2_outputs(3186) <= a or b;
    layer2_outputs(3187) <= b and not a;
    layer2_outputs(3188) <= b and not a;
    layer2_outputs(3189) <= a xor b;
    layer2_outputs(3190) <= a and not b;
    layer2_outputs(3191) <= not b or a;
    layer2_outputs(3192) <= a and not b;
    layer2_outputs(3193) <= a;
    layer2_outputs(3194) <= a and not b;
    layer2_outputs(3195) <= not a;
    layer2_outputs(3196) <= a;
    layer2_outputs(3197) <= not b or a;
    layer2_outputs(3198) <= a and b;
    layer2_outputs(3199) <= not a or b;
    layer2_outputs(3200) <= a or b;
    layer2_outputs(3201) <= a;
    layer2_outputs(3202) <= not a;
    layer2_outputs(3203) <= a or b;
    layer2_outputs(3204) <= a and not b;
    layer2_outputs(3205) <= a;
    layer2_outputs(3206) <= a;
    layer2_outputs(3207) <= a and not b;
    layer2_outputs(3208) <= not (a or b);
    layer2_outputs(3209) <= not (a and b);
    layer2_outputs(3210) <= not (a and b);
    layer2_outputs(3211) <= b and not a;
    layer2_outputs(3212) <= a or b;
    layer2_outputs(3213) <= 1'b0;
    layer2_outputs(3214) <= a and not b;
    layer2_outputs(3215) <= not b or a;
    layer2_outputs(3216) <= a or b;
    layer2_outputs(3217) <= 1'b1;
    layer2_outputs(3218) <= not (a and b);
    layer2_outputs(3219) <= not a;
    layer2_outputs(3220) <= a and not b;
    layer2_outputs(3221) <= 1'b1;
    layer2_outputs(3222) <= 1'b0;
    layer2_outputs(3223) <= not b or a;
    layer2_outputs(3224) <= not b or a;
    layer2_outputs(3225) <= b and not a;
    layer2_outputs(3226) <= not (a xor b);
    layer2_outputs(3227) <= not a or b;
    layer2_outputs(3228) <= not (a or b);
    layer2_outputs(3229) <= 1'b1;
    layer2_outputs(3230) <= a;
    layer2_outputs(3231) <= b;
    layer2_outputs(3232) <= not (a and b);
    layer2_outputs(3233) <= 1'b1;
    layer2_outputs(3234) <= a and not b;
    layer2_outputs(3235) <= a and b;
    layer2_outputs(3236) <= not b;
    layer2_outputs(3237) <= not (a or b);
    layer2_outputs(3238) <= 1'b1;
    layer2_outputs(3239) <= not a;
    layer2_outputs(3240) <= not b or a;
    layer2_outputs(3241) <= not a;
    layer2_outputs(3242) <= 1'b0;
    layer2_outputs(3243) <= b;
    layer2_outputs(3244) <= not b;
    layer2_outputs(3245) <= 1'b0;
    layer2_outputs(3246) <= a;
    layer2_outputs(3247) <= 1'b0;
    layer2_outputs(3248) <= not (a or b);
    layer2_outputs(3249) <= not (a or b);
    layer2_outputs(3250) <= b and not a;
    layer2_outputs(3251) <= 1'b0;
    layer2_outputs(3252) <= not b or a;
    layer2_outputs(3253) <= a and b;
    layer2_outputs(3254) <= b;
    layer2_outputs(3255) <= a and not b;
    layer2_outputs(3256) <= 1'b1;
    layer2_outputs(3257) <= a or b;
    layer2_outputs(3258) <= 1'b0;
    layer2_outputs(3259) <= a and b;
    layer2_outputs(3260) <= not b;
    layer2_outputs(3261) <= a or b;
    layer2_outputs(3262) <= not b or a;
    layer2_outputs(3263) <= not (a xor b);
    layer2_outputs(3264) <= 1'b0;
    layer2_outputs(3265) <= not (a or b);
    layer2_outputs(3266) <= not (a and b);
    layer2_outputs(3267) <= 1'b0;
    layer2_outputs(3268) <= not b;
    layer2_outputs(3269) <= a;
    layer2_outputs(3270) <= a or b;
    layer2_outputs(3271) <= a and b;
    layer2_outputs(3272) <= not a;
    layer2_outputs(3273) <= 1'b1;
    layer2_outputs(3274) <= not b or a;
    layer2_outputs(3275) <= a and b;
    layer2_outputs(3276) <= not (a xor b);
    layer2_outputs(3277) <= b and not a;
    layer2_outputs(3278) <= not b;
    layer2_outputs(3279) <= a and b;
    layer2_outputs(3280) <= 1'b0;
    layer2_outputs(3281) <= not a or b;
    layer2_outputs(3282) <= a;
    layer2_outputs(3283) <= 1'b0;
    layer2_outputs(3284) <= 1'b0;
    layer2_outputs(3285) <= a and not b;
    layer2_outputs(3286) <= b;
    layer2_outputs(3287) <= not a;
    layer2_outputs(3288) <= a or b;
    layer2_outputs(3289) <= a or b;
    layer2_outputs(3290) <= not a;
    layer2_outputs(3291) <= not a or b;
    layer2_outputs(3292) <= not a;
    layer2_outputs(3293) <= a;
    layer2_outputs(3294) <= a and b;
    layer2_outputs(3295) <= not a or b;
    layer2_outputs(3296) <= not b;
    layer2_outputs(3297) <= not (a and b);
    layer2_outputs(3298) <= not (a or b);
    layer2_outputs(3299) <= 1'b1;
    layer2_outputs(3300) <= a or b;
    layer2_outputs(3301) <= not b;
    layer2_outputs(3302) <= a or b;
    layer2_outputs(3303) <= a and not b;
    layer2_outputs(3304) <= not (a and b);
    layer2_outputs(3305) <= b;
    layer2_outputs(3306) <= not (a and b);
    layer2_outputs(3307) <= a;
    layer2_outputs(3308) <= a and not b;
    layer2_outputs(3309) <= b;
    layer2_outputs(3310) <= not a;
    layer2_outputs(3311) <= a and not b;
    layer2_outputs(3312) <= 1'b1;
    layer2_outputs(3313) <= a;
    layer2_outputs(3314) <= a and b;
    layer2_outputs(3315) <= not (a xor b);
    layer2_outputs(3316) <= a and b;
    layer2_outputs(3317) <= not a;
    layer2_outputs(3318) <= not (a and b);
    layer2_outputs(3319) <= b;
    layer2_outputs(3320) <= a xor b;
    layer2_outputs(3321) <= not b or a;
    layer2_outputs(3322) <= not (a or b);
    layer2_outputs(3323) <= a and not b;
    layer2_outputs(3324) <= 1'b1;
    layer2_outputs(3325) <= a and not b;
    layer2_outputs(3326) <= not b;
    layer2_outputs(3327) <= not b;
    layer2_outputs(3328) <= a and not b;
    layer2_outputs(3329) <= not a or b;
    layer2_outputs(3330) <= not b or a;
    layer2_outputs(3331) <= 1'b0;
    layer2_outputs(3332) <= 1'b0;
    layer2_outputs(3333) <= not a or b;
    layer2_outputs(3334) <= b;
    layer2_outputs(3335) <= not b or a;
    layer2_outputs(3336) <= not b or a;
    layer2_outputs(3337) <= not a;
    layer2_outputs(3338) <= 1'b1;
    layer2_outputs(3339) <= b and not a;
    layer2_outputs(3340) <= not a or b;
    layer2_outputs(3341) <= a or b;
    layer2_outputs(3342) <= not b or a;
    layer2_outputs(3343) <= 1'b0;
    layer2_outputs(3344) <= not (a or b);
    layer2_outputs(3345) <= not a;
    layer2_outputs(3346) <= a and b;
    layer2_outputs(3347) <= not b or a;
    layer2_outputs(3348) <= a and b;
    layer2_outputs(3349) <= not a or b;
    layer2_outputs(3350) <= not (a and b);
    layer2_outputs(3351) <= a;
    layer2_outputs(3352) <= 1'b0;
    layer2_outputs(3353) <= not (a or b);
    layer2_outputs(3354) <= a and not b;
    layer2_outputs(3355) <= a xor b;
    layer2_outputs(3356) <= not (a or b);
    layer2_outputs(3357) <= not a or b;
    layer2_outputs(3358) <= not (a or b);
    layer2_outputs(3359) <= a and b;
    layer2_outputs(3360) <= 1'b0;
    layer2_outputs(3361) <= not a or b;
    layer2_outputs(3362) <= a or b;
    layer2_outputs(3363) <= not b or a;
    layer2_outputs(3364) <= 1'b1;
    layer2_outputs(3365) <= not (a or b);
    layer2_outputs(3366) <= not a or b;
    layer2_outputs(3367) <= 1'b0;
    layer2_outputs(3368) <= 1'b1;
    layer2_outputs(3369) <= not (a and b);
    layer2_outputs(3370) <= a or b;
    layer2_outputs(3371) <= 1'b0;
    layer2_outputs(3372) <= b;
    layer2_outputs(3373) <= 1'b1;
    layer2_outputs(3374) <= a;
    layer2_outputs(3375) <= not b;
    layer2_outputs(3376) <= a or b;
    layer2_outputs(3377) <= not b or a;
    layer2_outputs(3378) <= a and b;
    layer2_outputs(3379) <= not a;
    layer2_outputs(3380) <= not a;
    layer2_outputs(3381) <= b and not a;
    layer2_outputs(3382) <= a and b;
    layer2_outputs(3383) <= not a or b;
    layer2_outputs(3384) <= not b or a;
    layer2_outputs(3385) <= not b or a;
    layer2_outputs(3386) <= not (a or b);
    layer2_outputs(3387) <= not b or a;
    layer2_outputs(3388) <= a and b;
    layer2_outputs(3389) <= a or b;
    layer2_outputs(3390) <= not a or b;
    layer2_outputs(3391) <= not a;
    layer2_outputs(3392) <= not a or b;
    layer2_outputs(3393) <= b;
    layer2_outputs(3394) <= a;
    layer2_outputs(3395) <= a and not b;
    layer2_outputs(3396) <= a and b;
    layer2_outputs(3397) <= 1'b0;
    layer2_outputs(3398) <= not b or a;
    layer2_outputs(3399) <= not (a and b);
    layer2_outputs(3400) <= b and not a;
    layer2_outputs(3401) <= b;
    layer2_outputs(3402) <= 1'b0;
    layer2_outputs(3403) <= not b;
    layer2_outputs(3404) <= 1'b0;
    layer2_outputs(3405) <= a;
    layer2_outputs(3406) <= not (a or b);
    layer2_outputs(3407) <= not b or a;
    layer2_outputs(3408) <= not (a and b);
    layer2_outputs(3409) <= not a or b;
    layer2_outputs(3410) <= a;
    layer2_outputs(3411) <= not a or b;
    layer2_outputs(3412) <= not b;
    layer2_outputs(3413) <= not (a or b);
    layer2_outputs(3414) <= a and not b;
    layer2_outputs(3415) <= b and not a;
    layer2_outputs(3416) <= not a;
    layer2_outputs(3417) <= not b;
    layer2_outputs(3418) <= not (a or b);
    layer2_outputs(3419) <= 1'b0;
    layer2_outputs(3420) <= 1'b0;
    layer2_outputs(3421) <= 1'b0;
    layer2_outputs(3422) <= not b;
    layer2_outputs(3423) <= not a or b;
    layer2_outputs(3424) <= not (a and b);
    layer2_outputs(3425) <= not (a and b);
    layer2_outputs(3426) <= not b or a;
    layer2_outputs(3427) <= not b or a;
    layer2_outputs(3428) <= not (a and b);
    layer2_outputs(3429) <= not a or b;
    layer2_outputs(3430) <= 1'b0;
    layer2_outputs(3431) <= 1'b1;
    layer2_outputs(3432) <= a or b;
    layer2_outputs(3433) <= b and not a;
    layer2_outputs(3434) <= a xor b;
    layer2_outputs(3435) <= a xor b;
    layer2_outputs(3436) <= b;
    layer2_outputs(3437) <= not a;
    layer2_outputs(3438) <= 1'b1;
    layer2_outputs(3439) <= not a or b;
    layer2_outputs(3440) <= 1'b1;
    layer2_outputs(3441) <= not (a or b);
    layer2_outputs(3442) <= a or b;
    layer2_outputs(3443) <= not b;
    layer2_outputs(3444) <= 1'b0;
    layer2_outputs(3445) <= a and b;
    layer2_outputs(3446) <= not b or a;
    layer2_outputs(3447) <= 1'b1;
    layer2_outputs(3448) <= a and not b;
    layer2_outputs(3449) <= not b or a;
    layer2_outputs(3450) <= b and not a;
    layer2_outputs(3451) <= not (a or b);
    layer2_outputs(3452) <= not a or b;
    layer2_outputs(3453) <= b and not a;
    layer2_outputs(3454) <= b;
    layer2_outputs(3455) <= a;
    layer2_outputs(3456) <= not b or a;
    layer2_outputs(3457) <= a;
    layer2_outputs(3458) <= not (a and b);
    layer2_outputs(3459) <= not b or a;
    layer2_outputs(3460) <= not (a or b);
    layer2_outputs(3461) <= b and not a;
    layer2_outputs(3462) <= 1'b0;
    layer2_outputs(3463) <= not b or a;
    layer2_outputs(3464) <= a or b;
    layer2_outputs(3465) <= not a;
    layer2_outputs(3466) <= not (a and b);
    layer2_outputs(3467) <= b;
    layer2_outputs(3468) <= a or b;
    layer2_outputs(3469) <= not (a or b);
    layer2_outputs(3470) <= a and b;
    layer2_outputs(3471) <= not (a or b);
    layer2_outputs(3472) <= not (a or b);
    layer2_outputs(3473) <= a or b;
    layer2_outputs(3474) <= not b;
    layer2_outputs(3475) <= not (a and b);
    layer2_outputs(3476) <= 1'b0;
    layer2_outputs(3477) <= not b or a;
    layer2_outputs(3478) <= 1'b1;
    layer2_outputs(3479) <= not (a or b);
    layer2_outputs(3480) <= b;
    layer2_outputs(3481) <= not a or b;
    layer2_outputs(3482) <= a or b;
    layer2_outputs(3483) <= 1'b1;
    layer2_outputs(3484) <= a and b;
    layer2_outputs(3485) <= b;
    layer2_outputs(3486) <= a and b;
    layer2_outputs(3487) <= 1'b0;
    layer2_outputs(3488) <= not (a or b);
    layer2_outputs(3489) <= a and b;
    layer2_outputs(3490) <= a xor b;
    layer2_outputs(3491) <= b and not a;
    layer2_outputs(3492) <= not a;
    layer2_outputs(3493) <= a and not b;
    layer2_outputs(3494) <= a and not b;
    layer2_outputs(3495) <= not b or a;
    layer2_outputs(3496) <= b;
    layer2_outputs(3497) <= not (a or b);
    layer2_outputs(3498) <= not b or a;
    layer2_outputs(3499) <= 1'b1;
    layer2_outputs(3500) <= not a;
    layer2_outputs(3501) <= not b or a;
    layer2_outputs(3502) <= not (a or b);
    layer2_outputs(3503) <= b and not a;
    layer2_outputs(3504) <= not a;
    layer2_outputs(3505) <= a and b;
    layer2_outputs(3506) <= 1'b1;
    layer2_outputs(3507) <= not b;
    layer2_outputs(3508) <= 1'b0;
    layer2_outputs(3509) <= a and b;
    layer2_outputs(3510) <= b;
    layer2_outputs(3511) <= b;
    layer2_outputs(3512) <= not a;
    layer2_outputs(3513) <= 1'b1;
    layer2_outputs(3514) <= a and not b;
    layer2_outputs(3515) <= 1'b1;
    layer2_outputs(3516) <= 1'b1;
    layer2_outputs(3517) <= a and not b;
    layer2_outputs(3518) <= 1'b1;
    layer2_outputs(3519) <= 1'b0;
    layer2_outputs(3520) <= 1'b1;
    layer2_outputs(3521) <= not (a or b);
    layer2_outputs(3522) <= not (a xor b);
    layer2_outputs(3523) <= 1'b0;
    layer2_outputs(3524) <= not b;
    layer2_outputs(3525) <= 1'b0;
    layer2_outputs(3526) <= 1'b1;
    layer2_outputs(3527) <= not b;
    layer2_outputs(3528) <= not (a or b);
    layer2_outputs(3529) <= b;
    layer2_outputs(3530) <= a xor b;
    layer2_outputs(3531) <= not a or b;
    layer2_outputs(3532) <= not b;
    layer2_outputs(3533) <= b and not a;
    layer2_outputs(3534) <= a or b;
    layer2_outputs(3535) <= 1'b0;
    layer2_outputs(3536) <= a and b;
    layer2_outputs(3537) <= a or b;
    layer2_outputs(3538) <= not a;
    layer2_outputs(3539) <= a xor b;
    layer2_outputs(3540) <= not b;
    layer2_outputs(3541) <= not a;
    layer2_outputs(3542) <= 1'b1;
    layer2_outputs(3543) <= not b or a;
    layer2_outputs(3544) <= 1'b0;
    layer2_outputs(3545) <= b and not a;
    layer2_outputs(3546) <= b;
    layer2_outputs(3547) <= 1'b0;
    layer2_outputs(3548) <= not a or b;
    layer2_outputs(3549) <= not b or a;
    layer2_outputs(3550) <= a or b;
    layer2_outputs(3551) <= b and not a;
    layer2_outputs(3552) <= a and b;
    layer2_outputs(3553) <= a and not b;
    layer2_outputs(3554) <= not b or a;
    layer2_outputs(3555) <= 1'b0;
    layer2_outputs(3556) <= 1'b1;
    layer2_outputs(3557) <= 1'b0;
    layer2_outputs(3558) <= not b or a;
    layer2_outputs(3559) <= not b;
    layer2_outputs(3560) <= a and b;
    layer2_outputs(3561) <= not (a or b);
    layer2_outputs(3562) <= not a;
    layer2_outputs(3563) <= b and not a;
    layer2_outputs(3564) <= not b or a;
    layer2_outputs(3565) <= not b;
    layer2_outputs(3566) <= not (a or b);
    layer2_outputs(3567) <= b;
    layer2_outputs(3568) <= b and not a;
    layer2_outputs(3569) <= 1'b1;
    layer2_outputs(3570) <= 1'b0;
    layer2_outputs(3571) <= not a or b;
    layer2_outputs(3572) <= a and not b;
    layer2_outputs(3573) <= a and b;
    layer2_outputs(3574) <= not b or a;
    layer2_outputs(3575) <= b;
    layer2_outputs(3576) <= 1'b1;
    layer2_outputs(3577) <= not b;
    layer2_outputs(3578) <= not (a and b);
    layer2_outputs(3579) <= a and not b;
    layer2_outputs(3580) <= not b;
    layer2_outputs(3581) <= not (a and b);
    layer2_outputs(3582) <= a;
    layer2_outputs(3583) <= b;
    layer2_outputs(3584) <= 1'b0;
    layer2_outputs(3585) <= 1'b0;
    layer2_outputs(3586) <= a and not b;
    layer2_outputs(3587) <= a or b;
    layer2_outputs(3588) <= b and not a;
    layer2_outputs(3589) <= not a or b;
    layer2_outputs(3590) <= 1'b0;
    layer2_outputs(3591) <= a;
    layer2_outputs(3592) <= not a;
    layer2_outputs(3593) <= 1'b1;
    layer2_outputs(3594) <= 1'b1;
    layer2_outputs(3595) <= 1'b0;
    layer2_outputs(3596) <= b;
    layer2_outputs(3597) <= a xor b;
    layer2_outputs(3598) <= not a or b;
    layer2_outputs(3599) <= a;
    layer2_outputs(3600) <= a and not b;
    layer2_outputs(3601) <= b and not a;
    layer2_outputs(3602) <= not (a and b);
    layer2_outputs(3603) <= a and b;
    layer2_outputs(3604) <= not a;
    layer2_outputs(3605) <= not b;
    layer2_outputs(3606) <= a and b;
    layer2_outputs(3607) <= 1'b0;
    layer2_outputs(3608) <= a and not b;
    layer2_outputs(3609) <= not (a and b);
    layer2_outputs(3610) <= not a or b;
    layer2_outputs(3611) <= 1'b0;
    layer2_outputs(3612) <= 1'b1;
    layer2_outputs(3613) <= a and not b;
    layer2_outputs(3614) <= a and not b;
    layer2_outputs(3615) <= not a;
    layer2_outputs(3616) <= 1'b1;
    layer2_outputs(3617) <= a and b;
    layer2_outputs(3618) <= not b or a;
    layer2_outputs(3619) <= not a;
    layer2_outputs(3620) <= not (a and b);
    layer2_outputs(3621) <= not a or b;
    layer2_outputs(3622) <= not (a or b);
    layer2_outputs(3623) <= not a or b;
    layer2_outputs(3624) <= 1'b0;
    layer2_outputs(3625) <= a xor b;
    layer2_outputs(3626) <= not b;
    layer2_outputs(3627) <= 1'b1;
    layer2_outputs(3628) <= 1'b1;
    layer2_outputs(3629) <= b;
    layer2_outputs(3630) <= a and b;
    layer2_outputs(3631) <= a;
    layer2_outputs(3632) <= 1'b0;
    layer2_outputs(3633) <= a and b;
    layer2_outputs(3634) <= not a or b;
    layer2_outputs(3635) <= not b or a;
    layer2_outputs(3636) <= not a or b;
    layer2_outputs(3637) <= b;
    layer2_outputs(3638) <= 1'b0;
    layer2_outputs(3639) <= b and not a;
    layer2_outputs(3640) <= not a or b;
    layer2_outputs(3641) <= not b;
    layer2_outputs(3642) <= not a or b;
    layer2_outputs(3643) <= a;
    layer2_outputs(3644) <= a and b;
    layer2_outputs(3645) <= not b;
    layer2_outputs(3646) <= not (a and b);
    layer2_outputs(3647) <= not a or b;
    layer2_outputs(3648) <= a and not b;
    layer2_outputs(3649) <= b and not a;
    layer2_outputs(3650) <= b and not a;
    layer2_outputs(3651) <= 1'b1;
    layer2_outputs(3652) <= b and not a;
    layer2_outputs(3653) <= a xor b;
    layer2_outputs(3654) <= b and not a;
    layer2_outputs(3655) <= a;
    layer2_outputs(3656) <= not a;
    layer2_outputs(3657) <= not a;
    layer2_outputs(3658) <= 1'b1;
    layer2_outputs(3659) <= not (a and b);
    layer2_outputs(3660) <= a;
    layer2_outputs(3661) <= a and not b;
    layer2_outputs(3662) <= a;
    layer2_outputs(3663) <= not a or b;
    layer2_outputs(3664) <= not (a xor b);
    layer2_outputs(3665) <= not a;
    layer2_outputs(3666) <= not b or a;
    layer2_outputs(3667) <= 1'b1;
    layer2_outputs(3668) <= a and b;
    layer2_outputs(3669) <= not a or b;
    layer2_outputs(3670) <= not (a or b);
    layer2_outputs(3671) <= not (a xor b);
    layer2_outputs(3672) <= not b;
    layer2_outputs(3673) <= not a;
    layer2_outputs(3674) <= b and not a;
    layer2_outputs(3675) <= not (a xor b);
    layer2_outputs(3676) <= not a or b;
    layer2_outputs(3677) <= not (a or b);
    layer2_outputs(3678) <= a xor b;
    layer2_outputs(3679) <= not b or a;
    layer2_outputs(3680) <= a;
    layer2_outputs(3681) <= not a;
    layer2_outputs(3682) <= b;
    layer2_outputs(3683) <= b;
    layer2_outputs(3684) <= a and not b;
    layer2_outputs(3685) <= a and b;
    layer2_outputs(3686) <= not (a and b);
    layer2_outputs(3687) <= a and not b;
    layer2_outputs(3688) <= a;
    layer2_outputs(3689) <= 1'b0;
    layer2_outputs(3690) <= 1'b0;
    layer2_outputs(3691) <= b;
    layer2_outputs(3692) <= 1'b0;
    layer2_outputs(3693) <= b;
    layer2_outputs(3694) <= b and not a;
    layer2_outputs(3695) <= a and not b;
    layer2_outputs(3696) <= not b;
    layer2_outputs(3697) <= 1'b0;
    layer2_outputs(3698) <= not b;
    layer2_outputs(3699) <= 1'b1;
    layer2_outputs(3700) <= 1'b0;
    layer2_outputs(3701) <= not a or b;
    layer2_outputs(3702) <= b and not a;
    layer2_outputs(3703) <= a and b;
    layer2_outputs(3704) <= 1'b0;
    layer2_outputs(3705) <= 1'b0;
    layer2_outputs(3706) <= not (a or b);
    layer2_outputs(3707) <= b;
    layer2_outputs(3708) <= b and not a;
    layer2_outputs(3709) <= 1'b0;
    layer2_outputs(3710) <= 1'b0;
    layer2_outputs(3711) <= b;
    layer2_outputs(3712) <= not (a and b);
    layer2_outputs(3713) <= a and not b;
    layer2_outputs(3714) <= 1'b0;
    layer2_outputs(3715) <= 1'b0;
    layer2_outputs(3716) <= a and not b;
    layer2_outputs(3717) <= 1'b0;
    layer2_outputs(3718) <= not a;
    layer2_outputs(3719) <= 1'b0;
    layer2_outputs(3720) <= b and not a;
    layer2_outputs(3721) <= b;
    layer2_outputs(3722) <= a and not b;
    layer2_outputs(3723) <= a and not b;
    layer2_outputs(3724) <= not (a or b);
    layer2_outputs(3725) <= not a;
    layer2_outputs(3726) <= b and not a;
    layer2_outputs(3727) <= not (a and b);
    layer2_outputs(3728) <= not (a and b);
    layer2_outputs(3729) <= a and b;
    layer2_outputs(3730) <= b;
    layer2_outputs(3731) <= a;
    layer2_outputs(3732) <= 1'b1;
    layer2_outputs(3733) <= a and b;
    layer2_outputs(3734) <= a and not b;
    layer2_outputs(3735) <= b;
    layer2_outputs(3736) <= not (a and b);
    layer2_outputs(3737) <= a and b;
    layer2_outputs(3738) <= not (a or b);
    layer2_outputs(3739) <= 1'b1;
    layer2_outputs(3740) <= b;
    layer2_outputs(3741) <= not a;
    layer2_outputs(3742) <= a and b;
    layer2_outputs(3743) <= a or b;
    layer2_outputs(3744) <= 1'b1;
    layer2_outputs(3745) <= not a;
    layer2_outputs(3746) <= 1'b0;
    layer2_outputs(3747) <= not a;
    layer2_outputs(3748) <= not (a and b);
    layer2_outputs(3749) <= not a or b;
    layer2_outputs(3750) <= a and not b;
    layer2_outputs(3751) <= not b or a;
    layer2_outputs(3752) <= not (a or b);
    layer2_outputs(3753) <= a and b;
    layer2_outputs(3754) <= a and b;
    layer2_outputs(3755) <= a;
    layer2_outputs(3756) <= a;
    layer2_outputs(3757) <= not b or a;
    layer2_outputs(3758) <= b;
    layer2_outputs(3759) <= b and not a;
    layer2_outputs(3760) <= 1'b1;
    layer2_outputs(3761) <= a and not b;
    layer2_outputs(3762) <= 1'b1;
    layer2_outputs(3763) <= not b;
    layer2_outputs(3764) <= b;
    layer2_outputs(3765) <= b and not a;
    layer2_outputs(3766) <= not (a or b);
    layer2_outputs(3767) <= a and b;
    layer2_outputs(3768) <= b and not a;
    layer2_outputs(3769) <= a and not b;
    layer2_outputs(3770) <= a;
    layer2_outputs(3771) <= not b or a;
    layer2_outputs(3772) <= not a or b;
    layer2_outputs(3773) <= 1'b1;
    layer2_outputs(3774) <= 1'b0;
    layer2_outputs(3775) <= a or b;
    layer2_outputs(3776) <= 1'b1;
    layer2_outputs(3777) <= not (a and b);
    layer2_outputs(3778) <= a and not b;
    layer2_outputs(3779) <= a or b;
    layer2_outputs(3780) <= b and not a;
    layer2_outputs(3781) <= b;
    layer2_outputs(3782) <= not (a or b);
    layer2_outputs(3783) <= not (a and b);
    layer2_outputs(3784) <= not a or b;
    layer2_outputs(3785) <= a and b;
    layer2_outputs(3786) <= not b;
    layer2_outputs(3787) <= a and not b;
    layer2_outputs(3788) <= b and not a;
    layer2_outputs(3789) <= not (a and b);
    layer2_outputs(3790) <= not b or a;
    layer2_outputs(3791) <= 1'b0;
    layer2_outputs(3792) <= not b or a;
    layer2_outputs(3793) <= b and not a;
    layer2_outputs(3794) <= a;
    layer2_outputs(3795) <= not b or a;
    layer2_outputs(3796) <= not a or b;
    layer2_outputs(3797) <= 1'b0;
    layer2_outputs(3798) <= not b;
    layer2_outputs(3799) <= a xor b;
    layer2_outputs(3800) <= 1'b0;
    layer2_outputs(3801) <= not a;
    layer2_outputs(3802) <= a xor b;
    layer2_outputs(3803) <= not b or a;
    layer2_outputs(3804) <= not b or a;
    layer2_outputs(3805) <= not b;
    layer2_outputs(3806) <= not a or b;
    layer2_outputs(3807) <= a;
    layer2_outputs(3808) <= not a or b;
    layer2_outputs(3809) <= a and b;
    layer2_outputs(3810) <= b and not a;
    layer2_outputs(3811) <= not (a and b);
    layer2_outputs(3812) <= not a or b;
    layer2_outputs(3813) <= 1'b0;
    layer2_outputs(3814) <= 1'b1;
    layer2_outputs(3815) <= 1'b0;
    layer2_outputs(3816) <= not (a and b);
    layer2_outputs(3817) <= not b or a;
    layer2_outputs(3818) <= a or b;
    layer2_outputs(3819) <= a;
    layer2_outputs(3820) <= b and not a;
    layer2_outputs(3821) <= a xor b;
    layer2_outputs(3822) <= b and not a;
    layer2_outputs(3823) <= not a or b;
    layer2_outputs(3824) <= 1'b0;
    layer2_outputs(3825) <= 1'b0;
    layer2_outputs(3826) <= not (a and b);
    layer2_outputs(3827) <= not b or a;
    layer2_outputs(3828) <= not (a xor b);
    layer2_outputs(3829) <= 1'b1;
    layer2_outputs(3830) <= a and not b;
    layer2_outputs(3831) <= not (a and b);
    layer2_outputs(3832) <= 1'b0;
    layer2_outputs(3833) <= a and not b;
    layer2_outputs(3834) <= 1'b1;
    layer2_outputs(3835) <= not (a and b);
    layer2_outputs(3836) <= not a;
    layer2_outputs(3837) <= not b or a;
    layer2_outputs(3838) <= not a or b;
    layer2_outputs(3839) <= not b or a;
    layer2_outputs(3840) <= 1'b1;
    layer2_outputs(3841) <= 1'b0;
    layer2_outputs(3842) <= a or b;
    layer2_outputs(3843) <= not b or a;
    layer2_outputs(3844) <= not (a and b);
    layer2_outputs(3845) <= 1'b1;
    layer2_outputs(3846) <= 1'b0;
    layer2_outputs(3847) <= not a;
    layer2_outputs(3848) <= a and b;
    layer2_outputs(3849) <= a and b;
    layer2_outputs(3850) <= a and not b;
    layer2_outputs(3851) <= a xor b;
    layer2_outputs(3852) <= a and not b;
    layer2_outputs(3853) <= b and not a;
    layer2_outputs(3854) <= not a or b;
    layer2_outputs(3855) <= b and not a;
    layer2_outputs(3856) <= a or b;
    layer2_outputs(3857) <= a xor b;
    layer2_outputs(3858) <= a;
    layer2_outputs(3859) <= b and not a;
    layer2_outputs(3860) <= not (a and b);
    layer2_outputs(3861) <= not (a and b);
    layer2_outputs(3862) <= not b or a;
    layer2_outputs(3863) <= b;
    layer2_outputs(3864) <= 1'b0;
    layer2_outputs(3865) <= not (a or b);
    layer2_outputs(3866) <= not a;
    layer2_outputs(3867) <= b;
    layer2_outputs(3868) <= b and not a;
    layer2_outputs(3869) <= not (a and b);
    layer2_outputs(3870) <= a xor b;
    layer2_outputs(3871) <= a;
    layer2_outputs(3872) <= a and not b;
    layer2_outputs(3873) <= 1'b1;
    layer2_outputs(3874) <= b and not a;
    layer2_outputs(3875) <= not (a or b);
    layer2_outputs(3876) <= b;
    layer2_outputs(3877) <= a and not b;
    layer2_outputs(3878) <= a or b;
    layer2_outputs(3879) <= b;
    layer2_outputs(3880) <= a;
    layer2_outputs(3881) <= a and b;
    layer2_outputs(3882) <= b and not a;
    layer2_outputs(3883) <= 1'b0;
    layer2_outputs(3884) <= not (a and b);
    layer2_outputs(3885) <= a or b;
    layer2_outputs(3886) <= a and b;
    layer2_outputs(3887) <= a;
    layer2_outputs(3888) <= not a or b;
    layer2_outputs(3889) <= not b or a;
    layer2_outputs(3890) <= a or b;
    layer2_outputs(3891) <= 1'b0;
    layer2_outputs(3892) <= b;
    layer2_outputs(3893) <= a;
    layer2_outputs(3894) <= not a;
    layer2_outputs(3895) <= b;
    layer2_outputs(3896) <= not b or a;
    layer2_outputs(3897) <= not a;
    layer2_outputs(3898) <= 1'b1;
    layer2_outputs(3899) <= a and b;
    layer2_outputs(3900) <= a and not b;
    layer2_outputs(3901) <= 1'b1;
    layer2_outputs(3902) <= b;
    layer2_outputs(3903) <= 1'b1;
    layer2_outputs(3904) <= not b;
    layer2_outputs(3905) <= not a or b;
    layer2_outputs(3906) <= 1'b1;
    layer2_outputs(3907) <= 1'b1;
    layer2_outputs(3908) <= 1'b1;
    layer2_outputs(3909) <= not (a and b);
    layer2_outputs(3910) <= 1'b1;
    layer2_outputs(3911) <= 1'b1;
    layer2_outputs(3912) <= 1'b0;
    layer2_outputs(3913) <= a and not b;
    layer2_outputs(3914) <= a or b;
    layer2_outputs(3915) <= not b;
    layer2_outputs(3916) <= 1'b0;
    layer2_outputs(3917) <= b and not a;
    layer2_outputs(3918) <= b;
    layer2_outputs(3919) <= a;
    layer2_outputs(3920) <= not b or a;
    layer2_outputs(3921) <= 1'b1;
    layer2_outputs(3922) <= 1'b1;
    layer2_outputs(3923) <= 1'b1;
    layer2_outputs(3924) <= not a or b;
    layer2_outputs(3925) <= 1'b0;
    layer2_outputs(3926) <= not (a or b);
    layer2_outputs(3927) <= not (a and b);
    layer2_outputs(3928) <= 1'b0;
    layer2_outputs(3929) <= 1'b0;
    layer2_outputs(3930) <= not (a or b);
    layer2_outputs(3931) <= not b;
    layer2_outputs(3932) <= 1'b0;
    layer2_outputs(3933) <= not a or b;
    layer2_outputs(3934) <= not b or a;
    layer2_outputs(3935) <= a and b;
    layer2_outputs(3936) <= 1'b1;
    layer2_outputs(3937) <= not (a and b);
    layer2_outputs(3938) <= not b or a;
    layer2_outputs(3939) <= a and b;
    layer2_outputs(3940) <= 1'b1;
    layer2_outputs(3941) <= not a or b;
    layer2_outputs(3942) <= not a or b;
    layer2_outputs(3943) <= not b;
    layer2_outputs(3944) <= b;
    layer2_outputs(3945) <= a and not b;
    layer2_outputs(3946) <= a;
    layer2_outputs(3947) <= not (a and b);
    layer2_outputs(3948) <= not (a and b);
    layer2_outputs(3949) <= b and not a;
    layer2_outputs(3950) <= 1'b1;
    layer2_outputs(3951) <= a;
    layer2_outputs(3952) <= not a;
    layer2_outputs(3953) <= a or b;
    layer2_outputs(3954) <= not (a or b);
    layer2_outputs(3955) <= a and not b;
    layer2_outputs(3956) <= not b or a;
    layer2_outputs(3957) <= a and not b;
    layer2_outputs(3958) <= 1'b1;
    layer2_outputs(3959) <= not (a or b);
    layer2_outputs(3960) <= a or b;
    layer2_outputs(3961) <= a or b;
    layer2_outputs(3962) <= a and not b;
    layer2_outputs(3963) <= not (a and b);
    layer2_outputs(3964) <= not (a and b);
    layer2_outputs(3965) <= not a;
    layer2_outputs(3966) <= not b or a;
    layer2_outputs(3967) <= 1'b0;
    layer2_outputs(3968) <= a or b;
    layer2_outputs(3969) <= b;
    layer2_outputs(3970) <= not (a and b);
    layer2_outputs(3971) <= not a;
    layer2_outputs(3972) <= a;
    layer2_outputs(3973) <= b;
    layer2_outputs(3974) <= not (a xor b);
    layer2_outputs(3975) <= b and not a;
    layer2_outputs(3976) <= a;
    layer2_outputs(3977) <= 1'b1;
    layer2_outputs(3978) <= 1'b1;
    layer2_outputs(3979) <= not (a or b);
    layer2_outputs(3980) <= not a;
    layer2_outputs(3981) <= a or b;
    layer2_outputs(3982) <= not (a or b);
    layer2_outputs(3983) <= not a or b;
    layer2_outputs(3984) <= 1'b1;
    layer2_outputs(3985) <= not a or b;
    layer2_outputs(3986) <= a xor b;
    layer2_outputs(3987) <= not a or b;
    layer2_outputs(3988) <= a or b;
    layer2_outputs(3989) <= 1'b1;
    layer2_outputs(3990) <= a and not b;
    layer2_outputs(3991) <= 1'b0;
    layer2_outputs(3992) <= a and not b;
    layer2_outputs(3993) <= 1'b1;
    layer2_outputs(3994) <= a and not b;
    layer2_outputs(3995) <= a and not b;
    layer2_outputs(3996) <= a and b;
    layer2_outputs(3997) <= a and not b;
    layer2_outputs(3998) <= not b;
    layer2_outputs(3999) <= a xor b;
    layer2_outputs(4000) <= 1'b1;
    layer2_outputs(4001) <= b and not a;
    layer2_outputs(4002) <= 1'b0;
    layer2_outputs(4003) <= a;
    layer2_outputs(4004) <= not a;
    layer2_outputs(4005) <= b and not a;
    layer2_outputs(4006) <= a and b;
    layer2_outputs(4007) <= a or b;
    layer2_outputs(4008) <= not b;
    layer2_outputs(4009) <= not b;
    layer2_outputs(4010) <= not (a or b);
    layer2_outputs(4011) <= 1'b0;
    layer2_outputs(4012) <= a or b;
    layer2_outputs(4013) <= 1'b1;
    layer2_outputs(4014) <= 1'b0;
    layer2_outputs(4015) <= a or b;
    layer2_outputs(4016) <= not (a xor b);
    layer2_outputs(4017) <= not (a or b);
    layer2_outputs(4018) <= a and not b;
    layer2_outputs(4019) <= not (a and b);
    layer2_outputs(4020) <= not b or a;
    layer2_outputs(4021) <= a;
    layer2_outputs(4022) <= a or b;
    layer2_outputs(4023) <= not (a and b);
    layer2_outputs(4024) <= a or b;
    layer2_outputs(4025) <= a and not b;
    layer2_outputs(4026) <= not (a xor b);
    layer2_outputs(4027) <= a and b;
    layer2_outputs(4028) <= b;
    layer2_outputs(4029) <= 1'b0;
    layer2_outputs(4030) <= 1'b1;
    layer2_outputs(4031) <= a xor b;
    layer2_outputs(4032) <= not a;
    layer2_outputs(4033) <= not (a and b);
    layer2_outputs(4034) <= not b or a;
    layer2_outputs(4035) <= not b;
    layer2_outputs(4036) <= 1'b0;
    layer2_outputs(4037) <= b and not a;
    layer2_outputs(4038) <= a;
    layer2_outputs(4039) <= a and b;
    layer2_outputs(4040) <= 1'b1;
    layer2_outputs(4041) <= a xor b;
    layer2_outputs(4042) <= 1'b1;
    layer2_outputs(4043) <= a;
    layer2_outputs(4044) <= a or b;
    layer2_outputs(4045) <= 1'b1;
    layer2_outputs(4046) <= 1'b1;
    layer2_outputs(4047) <= 1'b0;
    layer2_outputs(4048) <= a;
    layer2_outputs(4049) <= a and b;
    layer2_outputs(4050) <= 1'b1;
    layer2_outputs(4051) <= not a;
    layer2_outputs(4052) <= not (a or b);
    layer2_outputs(4053) <= not a;
    layer2_outputs(4054) <= not (a or b);
    layer2_outputs(4055) <= b and not a;
    layer2_outputs(4056) <= a and not b;
    layer2_outputs(4057) <= a and not b;
    layer2_outputs(4058) <= a xor b;
    layer2_outputs(4059) <= not a;
    layer2_outputs(4060) <= not b;
    layer2_outputs(4061) <= not (a and b);
    layer2_outputs(4062) <= not (a or b);
    layer2_outputs(4063) <= not b or a;
    layer2_outputs(4064) <= not a or b;
    layer2_outputs(4065) <= a and not b;
    layer2_outputs(4066) <= a;
    layer2_outputs(4067) <= a xor b;
    layer2_outputs(4068) <= a and not b;
    layer2_outputs(4069) <= a or b;
    layer2_outputs(4070) <= a and not b;
    layer2_outputs(4071) <= 1'b1;
    layer2_outputs(4072) <= b;
    layer2_outputs(4073) <= not (a or b);
    layer2_outputs(4074) <= a or b;
    layer2_outputs(4075) <= not b or a;
    layer2_outputs(4076) <= not (a xor b);
    layer2_outputs(4077) <= not b;
    layer2_outputs(4078) <= not b or a;
    layer2_outputs(4079) <= not a or b;
    layer2_outputs(4080) <= b and not a;
    layer2_outputs(4081) <= 1'b0;
    layer2_outputs(4082) <= 1'b0;
    layer2_outputs(4083) <= a;
    layer2_outputs(4084) <= 1'b1;
    layer2_outputs(4085) <= b;
    layer2_outputs(4086) <= 1'b0;
    layer2_outputs(4087) <= 1'b1;
    layer2_outputs(4088) <= b and not a;
    layer2_outputs(4089) <= a xor b;
    layer2_outputs(4090) <= not b;
    layer2_outputs(4091) <= 1'b0;
    layer2_outputs(4092) <= 1'b0;
    layer2_outputs(4093) <= 1'b0;
    layer2_outputs(4094) <= not a or b;
    layer2_outputs(4095) <= b;
    layer2_outputs(4096) <= 1'b1;
    layer2_outputs(4097) <= not (a and b);
    layer2_outputs(4098) <= not (a and b);
    layer2_outputs(4099) <= b and not a;
    layer2_outputs(4100) <= a and b;
    layer2_outputs(4101) <= not a or b;
    layer2_outputs(4102) <= 1'b0;
    layer2_outputs(4103) <= 1'b1;
    layer2_outputs(4104) <= not a or b;
    layer2_outputs(4105) <= not b or a;
    layer2_outputs(4106) <= a or b;
    layer2_outputs(4107) <= not (a xor b);
    layer2_outputs(4108) <= not b or a;
    layer2_outputs(4109) <= not a;
    layer2_outputs(4110) <= not (a xor b);
    layer2_outputs(4111) <= a;
    layer2_outputs(4112) <= a or b;
    layer2_outputs(4113) <= not a or b;
    layer2_outputs(4114) <= b;
    layer2_outputs(4115) <= 1'b1;
    layer2_outputs(4116) <= not (a and b);
    layer2_outputs(4117) <= not (a and b);
    layer2_outputs(4118) <= not (a or b);
    layer2_outputs(4119) <= a and b;
    layer2_outputs(4120) <= not (a and b);
    layer2_outputs(4121) <= not b;
    layer2_outputs(4122) <= b and not a;
    layer2_outputs(4123) <= a and not b;
    layer2_outputs(4124) <= b and not a;
    layer2_outputs(4125) <= 1'b0;
    layer2_outputs(4126) <= a;
    layer2_outputs(4127) <= not a;
    layer2_outputs(4128) <= not a;
    layer2_outputs(4129) <= not (a xor b);
    layer2_outputs(4130) <= not (a or b);
    layer2_outputs(4131) <= 1'b1;
    layer2_outputs(4132) <= a or b;
    layer2_outputs(4133) <= not a or b;
    layer2_outputs(4134) <= 1'b0;
    layer2_outputs(4135) <= not b;
    layer2_outputs(4136) <= not a or b;
    layer2_outputs(4137) <= a or b;
    layer2_outputs(4138) <= not (a or b);
    layer2_outputs(4139) <= 1'b0;
    layer2_outputs(4140) <= not a;
    layer2_outputs(4141) <= not a or b;
    layer2_outputs(4142) <= 1'b1;
    layer2_outputs(4143) <= 1'b0;
    layer2_outputs(4144) <= not (a or b);
    layer2_outputs(4145) <= not b or a;
    layer2_outputs(4146) <= 1'b1;
    layer2_outputs(4147) <= not b;
    layer2_outputs(4148) <= a and b;
    layer2_outputs(4149) <= a and b;
    layer2_outputs(4150) <= a;
    layer2_outputs(4151) <= not a or b;
    layer2_outputs(4152) <= not (a or b);
    layer2_outputs(4153) <= a;
    layer2_outputs(4154) <= a;
    layer2_outputs(4155) <= not b or a;
    layer2_outputs(4156) <= a and not b;
    layer2_outputs(4157) <= not (a or b);
    layer2_outputs(4158) <= not (a or b);
    layer2_outputs(4159) <= 1'b1;
    layer2_outputs(4160) <= 1'b1;
    layer2_outputs(4161) <= a and b;
    layer2_outputs(4162) <= not (a and b);
    layer2_outputs(4163) <= not a or b;
    layer2_outputs(4164) <= not (a and b);
    layer2_outputs(4165) <= not (a xor b);
    layer2_outputs(4166) <= not (a or b);
    layer2_outputs(4167) <= b;
    layer2_outputs(4168) <= a and not b;
    layer2_outputs(4169) <= a or b;
    layer2_outputs(4170) <= not (a xor b);
    layer2_outputs(4171) <= a and not b;
    layer2_outputs(4172) <= not (a xor b);
    layer2_outputs(4173) <= not a;
    layer2_outputs(4174) <= a and not b;
    layer2_outputs(4175) <= not (a xor b);
    layer2_outputs(4176) <= a and b;
    layer2_outputs(4177) <= a xor b;
    layer2_outputs(4178) <= not (a and b);
    layer2_outputs(4179) <= a and b;
    layer2_outputs(4180) <= a and b;
    layer2_outputs(4181) <= not b or a;
    layer2_outputs(4182) <= a;
    layer2_outputs(4183) <= a and b;
    layer2_outputs(4184) <= not b or a;
    layer2_outputs(4185) <= 1'b0;
    layer2_outputs(4186) <= a;
    layer2_outputs(4187) <= a;
    layer2_outputs(4188) <= a and not b;
    layer2_outputs(4189) <= 1'b0;
    layer2_outputs(4190) <= not (a and b);
    layer2_outputs(4191) <= 1'b1;
    layer2_outputs(4192) <= 1'b1;
    layer2_outputs(4193) <= not (a and b);
    layer2_outputs(4194) <= a or b;
    layer2_outputs(4195) <= a and b;
    layer2_outputs(4196) <= not b or a;
    layer2_outputs(4197) <= not (a and b);
    layer2_outputs(4198) <= a or b;
    layer2_outputs(4199) <= a and b;
    layer2_outputs(4200) <= not a;
    layer2_outputs(4201) <= not a;
    layer2_outputs(4202) <= a or b;
    layer2_outputs(4203) <= not a or b;
    layer2_outputs(4204) <= a and not b;
    layer2_outputs(4205) <= a xor b;
    layer2_outputs(4206) <= a xor b;
    layer2_outputs(4207) <= a and b;
    layer2_outputs(4208) <= 1'b0;
    layer2_outputs(4209) <= not b or a;
    layer2_outputs(4210) <= b;
    layer2_outputs(4211) <= a or b;
    layer2_outputs(4212) <= a or b;
    layer2_outputs(4213) <= 1'b0;
    layer2_outputs(4214) <= a;
    layer2_outputs(4215) <= not a or b;
    layer2_outputs(4216) <= 1'b1;
    layer2_outputs(4217) <= not a;
    layer2_outputs(4218) <= not b;
    layer2_outputs(4219) <= a or b;
    layer2_outputs(4220) <= not a;
    layer2_outputs(4221) <= a or b;
    layer2_outputs(4222) <= a and b;
    layer2_outputs(4223) <= b and not a;
    layer2_outputs(4224) <= not a or b;
    layer2_outputs(4225) <= 1'b0;
    layer2_outputs(4226) <= not (a xor b);
    layer2_outputs(4227) <= not a;
    layer2_outputs(4228) <= a or b;
    layer2_outputs(4229) <= 1'b0;
    layer2_outputs(4230) <= b and not a;
    layer2_outputs(4231) <= 1'b1;
    layer2_outputs(4232) <= a and not b;
    layer2_outputs(4233) <= not (a or b);
    layer2_outputs(4234) <= a and b;
    layer2_outputs(4235) <= a or b;
    layer2_outputs(4236) <= b and not a;
    layer2_outputs(4237) <= a;
    layer2_outputs(4238) <= 1'b0;
    layer2_outputs(4239) <= b and not a;
    layer2_outputs(4240) <= b and not a;
    layer2_outputs(4241) <= not a;
    layer2_outputs(4242) <= a and not b;
    layer2_outputs(4243) <= b;
    layer2_outputs(4244) <= not a;
    layer2_outputs(4245) <= b;
    layer2_outputs(4246) <= not (a xor b);
    layer2_outputs(4247) <= a or b;
    layer2_outputs(4248) <= 1'b1;
    layer2_outputs(4249) <= 1'b0;
    layer2_outputs(4250) <= not a or b;
    layer2_outputs(4251) <= b and not a;
    layer2_outputs(4252) <= a or b;
    layer2_outputs(4253) <= not (a xor b);
    layer2_outputs(4254) <= a and b;
    layer2_outputs(4255) <= 1'b1;
    layer2_outputs(4256) <= a;
    layer2_outputs(4257) <= not (a and b);
    layer2_outputs(4258) <= not b;
    layer2_outputs(4259) <= not b or a;
    layer2_outputs(4260) <= a and b;
    layer2_outputs(4261) <= a;
    layer2_outputs(4262) <= 1'b0;
    layer2_outputs(4263) <= not b;
    layer2_outputs(4264) <= 1'b1;
    layer2_outputs(4265) <= a and b;
    layer2_outputs(4266) <= not b;
    layer2_outputs(4267) <= not a or b;
    layer2_outputs(4268) <= 1'b1;
    layer2_outputs(4269) <= not b;
    layer2_outputs(4270) <= not (a or b);
    layer2_outputs(4271) <= a;
    layer2_outputs(4272) <= not a;
    layer2_outputs(4273) <= a xor b;
    layer2_outputs(4274) <= a or b;
    layer2_outputs(4275) <= b;
    layer2_outputs(4276) <= a and not b;
    layer2_outputs(4277) <= 1'b1;
    layer2_outputs(4278) <= not a;
    layer2_outputs(4279) <= 1'b0;
    layer2_outputs(4280) <= a or b;
    layer2_outputs(4281) <= not (a or b);
    layer2_outputs(4282) <= a xor b;
    layer2_outputs(4283) <= 1'b1;
    layer2_outputs(4284) <= not (a or b);
    layer2_outputs(4285) <= 1'b1;
    layer2_outputs(4286) <= not (a and b);
    layer2_outputs(4287) <= a and b;
    layer2_outputs(4288) <= not a;
    layer2_outputs(4289) <= 1'b0;
    layer2_outputs(4290) <= not b or a;
    layer2_outputs(4291) <= not b or a;
    layer2_outputs(4292) <= b;
    layer2_outputs(4293) <= not (a or b);
    layer2_outputs(4294) <= a and not b;
    layer2_outputs(4295) <= 1'b1;
    layer2_outputs(4296) <= not b or a;
    layer2_outputs(4297) <= not a;
    layer2_outputs(4298) <= not (a or b);
    layer2_outputs(4299) <= a and not b;
    layer2_outputs(4300) <= a and not b;
    layer2_outputs(4301) <= a and not b;
    layer2_outputs(4302) <= 1'b1;
    layer2_outputs(4303) <= not (a and b);
    layer2_outputs(4304) <= not a;
    layer2_outputs(4305) <= not a or b;
    layer2_outputs(4306) <= not (a and b);
    layer2_outputs(4307) <= not a or b;
    layer2_outputs(4308) <= a and b;
    layer2_outputs(4309) <= b and not a;
    layer2_outputs(4310) <= 1'b0;
    layer2_outputs(4311) <= b;
    layer2_outputs(4312) <= 1'b0;
    layer2_outputs(4313) <= not (a and b);
    layer2_outputs(4314) <= a and not b;
    layer2_outputs(4315) <= b and not a;
    layer2_outputs(4316) <= not a;
    layer2_outputs(4317) <= not a;
    layer2_outputs(4318) <= a and b;
    layer2_outputs(4319) <= a or b;
    layer2_outputs(4320) <= 1'b0;
    layer2_outputs(4321) <= not b or a;
    layer2_outputs(4322) <= b;
    layer2_outputs(4323) <= b;
    layer2_outputs(4324) <= 1'b0;
    layer2_outputs(4325) <= not a;
    layer2_outputs(4326) <= not a;
    layer2_outputs(4327) <= not (a or b);
    layer2_outputs(4328) <= a and not b;
    layer2_outputs(4329) <= not a;
    layer2_outputs(4330) <= not b;
    layer2_outputs(4331) <= not a;
    layer2_outputs(4332) <= not b or a;
    layer2_outputs(4333) <= 1'b1;
    layer2_outputs(4334) <= not b;
    layer2_outputs(4335) <= 1'b1;
    layer2_outputs(4336) <= not b;
    layer2_outputs(4337) <= a and not b;
    layer2_outputs(4338) <= a and not b;
    layer2_outputs(4339) <= b;
    layer2_outputs(4340) <= not (a or b);
    layer2_outputs(4341) <= not b or a;
    layer2_outputs(4342) <= a;
    layer2_outputs(4343) <= not a or b;
    layer2_outputs(4344) <= not b;
    layer2_outputs(4345) <= b and not a;
    layer2_outputs(4346) <= a and not b;
    layer2_outputs(4347) <= 1'b0;
    layer2_outputs(4348) <= a or b;
    layer2_outputs(4349) <= a;
    layer2_outputs(4350) <= not a;
    layer2_outputs(4351) <= not (a xor b);
    layer2_outputs(4352) <= a or b;
    layer2_outputs(4353) <= not (a and b);
    layer2_outputs(4354) <= a and b;
    layer2_outputs(4355) <= a and b;
    layer2_outputs(4356) <= a xor b;
    layer2_outputs(4357) <= a and not b;
    layer2_outputs(4358) <= a and not b;
    layer2_outputs(4359) <= not (a or b);
    layer2_outputs(4360) <= not (a xor b);
    layer2_outputs(4361) <= not (a or b);
    layer2_outputs(4362) <= a or b;
    layer2_outputs(4363) <= a and b;
    layer2_outputs(4364) <= a and not b;
    layer2_outputs(4365) <= not (a and b);
    layer2_outputs(4366) <= a and not b;
    layer2_outputs(4367) <= a;
    layer2_outputs(4368) <= a and b;
    layer2_outputs(4369) <= a and not b;
    layer2_outputs(4370) <= a;
    layer2_outputs(4371) <= not b;
    layer2_outputs(4372) <= not (a and b);
    layer2_outputs(4373) <= not b;
    layer2_outputs(4374) <= not a or b;
    layer2_outputs(4375) <= not a;
    layer2_outputs(4376) <= a and b;
    layer2_outputs(4377) <= not (a or b);
    layer2_outputs(4378) <= not (a and b);
    layer2_outputs(4379) <= not b or a;
    layer2_outputs(4380) <= 1'b1;
    layer2_outputs(4381) <= not a;
    layer2_outputs(4382) <= 1'b0;
    layer2_outputs(4383) <= 1'b1;
    layer2_outputs(4384) <= not (a and b);
    layer2_outputs(4385) <= a and b;
    layer2_outputs(4386) <= b;
    layer2_outputs(4387) <= not a;
    layer2_outputs(4388) <= not b;
    layer2_outputs(4389) <= not b or a;
    layer2_outputs(4390) <= not b or a;
    layer2_outputs(4391) <= b and not a;
    layer2_outputs(4392) <= a or b;
    layer2_outputs(4393) <= 1'b0;
    layer2_outputs(4394) <= not (a or b);
    layer2_outputs(4395) <= not (a or b);
    layer2_outputs(4396) <= not a;
    layer2_outputs(4397) <= not b or a;
    layer2_outputs(4398) <= not b;
    layer2_outputs(4399) <= a and not b;
    layer2_outputs(4400) <= 1'b1;
    layer2_outputs(4401) <= a;
    layer2_outputs(4402) <= 1'b1;
    layer2_outputs(4403) <= a and not b;
    layer2_outputs(4404) <= a;
    layer2_outputs(4405) <= a and not b;
    layer2_outputs(4406) <= not b or a;
    layer2_outputs(4407) <= not (a and b);
    layer2_outputs(4408) <= not a or b;
    layer2_outputs(4409) <= not a or b;
    layer2_outputs(4410) <= b and not a;
    layer2_outputs(4411) <= not a or b;
    layer2_outputs(4412) <= not a;
    layer2_outputs(4413) <= not b;
    layer2_outputs(4414) <= 1'b0;
    layer2_outputs(4415) <= not a or b;
    layer2_outputs(4416) <= 1'b0;
    layer2_outputs(4417) <= not b;
    layer2_outputs(4418) <= a or b;
    layer2_outputs(4419) <= a;
    layer2_outputs(4420) <= a or b;
    layer2_outputs(4421) <= b;
    layer2_outputs(4422) <= a and b;
    layer2_outputs(4423) <= a and b;
    layer2_outputs(4424) <= not a;
    layer2_outputs(4425) <= not (a and b);
    layer2_outputs(4426) <= 1'b0;
    layer2_outputs(4427) <= a and b;
    layer2_outputs(4428) <= 1'b0;
    layer2_outputs(4429) <= b and not a;
    layer2_outputs(4430) <= a or b;
    layer2_outputs(4431) <= 1'b0;
    layer2_outputs(4432) <= a and not b;
    layer2_outputs(4433) <= a and b;
    layer2_outputs(4434) <= not a;
    layer2_outputs(4435) <= not (a or b);
    layer2_outputs(4436) <= not (a and b);
    layer2_outputs(4437) <= a or b;
    layer2_outputs(4438) <= a and not b;
    layer2_outputs(4439) <= 1'b1;
    layer2_outputs(4440) <= not (a xor b);
    layer2_outputs(4441) <= a and not b;
    layer2_outputs(4442) <= not b;
    layer2_outputs(4443) <= not a;
    layer2_outputs(4444) <= b and not a;
    layer2_outputs(4445) <= 1'b0;
    layer2_outputs(4446) <= a and not b;
    layer2_outputs(4447) <= 1'b0;
    layer2_outputs(4448) <= not a or b;
    layer2_outputs(4449) <= not (a and b);
    layer2_outputs(4450) <= a or b;
    layer2_outputs(4451) <= not (a or b);
    layer2_outputs(4452) <= not b or a;
    layer2_outputs(4453) <= not (a or b);
    layer2_outputs(4454) <= b and not a;
    layer2_outputs(4455) <= 1'b1;
    layer2_outputs(4456) <= not (a or b);
    layer2_outputs(4457) <= not b;
    layer2_outputs(4458) <= not b or a;
    layer2_outputs(4459) <= 1'b1;
    layer2_outputs(4460) <= not (a or b);
    layer2_outputs(4461) <= not b or a;
    layer2_outputs(4462) <= a and b;
    layer2_outputs(4463) <= 1'b0;
    layer2_outputs(4464) <= a or b;
    layer2_outputs(4465) <= not b;
    layer2_outputs(4466) <= b and not a;
    layer2_outputs(4467) <= a and b;
    layer2_outputs(4468) <= a and not b;
    layer2_outputs(4469) <= not a or b;
    layer2_outputs(4470) <= 1'b1;
    layer2_outputs(4471) <= not (a and b);
    layer2_outputs(4472) <= not b or a;
    layer2_outputs(4473) <= a or b;
    layer2_outputs(4474) <= not a or b;
    layer2_outputs(4475) <= a and b;
    layer2_outputs(4476) <= not (a or b);
    layer2_outputs(4477) <= not b or a;
    layer2_outputs(4478) <= 1'b1;
    layer2_outputs(4479) <= a or b;
    layer2_outputs(4480) <= not (a or b);
    layer2_outputs(4481) <= not b or a;
    layer2_outputs(4482) <= a and not b;
    layer2_outputs(4483) <= a;
    layer2_outputs(4484) <= a and b;
    layer2_outputs(4485) <= not b or a;
    layer2_outputs(4486) <= not a or b;
    layer2_outputs(4487) <= b and not a;
    layer2_outputs(4488) <= not a or b;
    layer2_outputs(4489) <= a;
    layer2_outputs(4490) <= a and b;
    layer2_outputs(4491) <= not (a or b);
    layer2_outputs(4492) <= a or b;
    layer2_outputs(4493) <= not a;
    layer2_outputs(4494) <= not (a and b);
    layer2_outputs(4495) <= a and b;
    layer2_outputs(4496) <= b;
    layer2_outputs(4497) <= a;
    layer2_outputs(4498) <= a or b;
    layer2_outputs(4499) <= a xor b;
    layer2_outputs(4500) <= a or b;
    layer2_outputs(4501) <= a;
    layer2_outputs(4502) <= a or b;
    layer2_outputs(4503) <= not a;
    layer2_outputs(4504) <= 1'b1;
    layer2_outputs(4505) <= 1'b1;
    layer2_outputs(4506) <= 1'b0;
    layer2_outputs(4507) <= not b or a;
    layer2_outputs(4508) <= b and not a;
    layer2_outputs(4509) <= b;
    layer2_outputs(4510) <= not a or b;
    layer2_outputs(4511) <= a and not b;
    layer2_outputs(4512) <= not b or a;
    layer2_outputs(4513) <= 1'b0;
    layer2_outputs(4514) <= 1'b0;
    layer2_outputs(4515) <= 1'b0;
    layer2_outputs(4516) <= 1'b1;
    layer2_outputs(4517) <= 1'b0;
    layer2_outputs(4518) <= a and b;
    layer2_outputs(4519) <= 1'b0;
    layer2_outputs(4520) <= 1'b0;
    layer2_outputs(4521) <= a;
    layer2_outputs(4522) <= not b;
    layer2_outputs(4523) <= b;
    layer2_outputs(4524) <= not a;
    layer2_outputs(4525) <= a;
    layer2_outputs(4526) <= not (a or b);
    layer2_outputs(4527) <= not (a and b);
    layer2_outputs(4528) <= not b or a;
    layer2_outputs(4529) <= a and not b;
    layer2_outputs(4530) <= a or b;
    layer2_outputs(4531) <= not b;
    layer2_outputs(4532) <= b;
    layer2_outputs(4533) <= b and not a;
    layer2_outputs(4534) <= a and b;
    layer2_outputs(4535) <= not b;
    layer2_outputs(4536) <= not (a xor b);
    layer2_outputs(4537) <= not (a or b);
    layer2_outputs(4538) <= not (a or b);
    layer2_outputs(4539) <= a;
    layer2_outputs(4540) <= not b;
    layer2_outputs(4541) <= a;
    layer2_outputs(4542) <= b;
    layer2_outputs(4543) <= b;
    layer2_outputs(4544) <= b;
    layer2_outputs(4545) <= 1'b0;
    layer2_outputs(4546) <= a and not b;
    layer2_outputs(4547) <= a and not b;
    layer2_outputs(4548) <= b and not a;
    layer2_outputs(4549) <= a xor b;
    layer2_outputs(4550) <= not b;
    layer2_outputs(4551) <= not (a and b);
    layer2_outputs(4552) <= 1'b1;
    layer2_outputs(4553) <= 1'b0;
    layer2_outputs(4554) <= not (a and b);
    layer2_outputs(4555) <= a and b;
    layer2_outputs(4556) <= a or b;
    layer2_outputs(4557) <= a and b;
    layer2_outputs(4558) <= a;
    layer2_outputs(4559) <= 1'b0;
    layer2_outputs(4560) <= 1'b1;
    layer2_outputs(4561) <= not a;
    layer2_outputs(4562) <= a and b;
    layer2_outputs(4563) <= a or b;
    layer2_outputs(4564) <= a and b;
    layer2_outputs(4565) <= a and b;
    layer2_outputs(4566) <= not a or b;
    layer2_outputs(4567) <= 1'b1;
    layer2_outputs(4568) <= not b;
    layer2_outputs(4569) <= 1'b1;
    layer2_outputs(4570) <= a and b;
    layer2_outputs(4571) <= a and b;
    layer2_outputs(4572) <= not (a and b);
    layer2_outputs(4573) <= a;
    layer2_outputs(4574) <= 1'b0;
    layer2_outputs(4575) <= b;
    layer2_outputs(4576) <= b and not a;
    layer2_outputs(4577) <= a or b;
    layer2_outputs(4578) <= not a;
    layer2_outputs(4579) <= b and not a;
    layer2_outputs(4580) <= 1'b0;
    layer2_outputs(4581) <= 1'b1;
    layer2_outputs(4582) <= a and not b;
    layer2_outputs(4583) <= a and not b;
    layer2_outputs(4584) <= not (a and b);
    layer2_outputs(4585) <= not (a and b);
    layer2_outputs(4586) <= b and not a;
    layer2_outputs(4587) <= a and not b;
    layer2_outputs(4588) <= not b;
    layer2_outputs(4589) <= b and not a;
    layer2_outputs(4590) <= not (a and b);
    layer2_outputs(4591) <= not a;
    layer2_outputs(4592) <= a and not b;
    layer2_outputs(4593) <= not (a or b);
    layer2_outputs(4594) <= not (a and b);
    layer2_outputs(4595) <= not a or b;
    layer2_outputs(4596) <= b and not a;
    layer2_outputs(4597) <= b and not a;
    layer2_outputs(4598) <= a and not b;
    layer2_outputs(4599) <= a xor b;
    layer2_outputs(4600) <= not b;
    layer2_outputs(4601) <= 1'b0;
    layer2_outputs(4602) <= 1'b0;
    layer2_outputs(4603) <= a and b;
    layer2_outputs(4604) <= not (a and b);
    layer2_outputs(4605) <= not (a and b);
    layer2_outputs(4606) <= 1'b1;
    layer2_outputs(4607) <= 1'b1;
    layer2_outputs(4608) <= not b or a;
    layer2_outputs(4609) <= 1'b1;
    layer2_outputs(4610) <= a or b;
    layer2_outputs(4611) <= not a;
    layer2_outputs(4612) <= 1'b1;
    layer2_outputs(4613) <= not (a or b);
    layer2_outputs(4614) <= not b or a;
    layer2_outputs(4615) <= a and not b;
    layer2_outputs(4616) <= not b;
    layer2_outputs(4617) <= a or b;
    layer2_outputs(4618) <= not (a or b);
    layer2_outputs(4619) <= not b;
    layer2_outputs(4620) <= b and not a;
    layer2_outputs(4621) <= a and b;
    layer2_outputs(4622) <= a;
    layer2_outputs(4623) <= a;
    layer2_outputs(4624) <= not a or b;
    layer2_outputs(4625) <= not (a xor b);
    layer2_outputs(4626) <= not (a xor b);
    layer2_outputs(4627) <= not b;
    layer2_outputs(4628) <= a and not b;
    layer2_outputs(4629) <= not b or a;
    layer2_outputs(4630) <= not (a xor b);
    layer2_outputs(4631) <= not b;
    layer2_outputs(4632) <= not (a xor b);
    layer2_outputs(4633) <= not a or b;
    layer2_outputs(4634) <= not a or b;
    layer2_outputs(4635) <= not (a xor b);
    layer2_outputs(4636) <= not (a xor b);
    layer2_outputs(4637) <= 1'b1;
    layer2_outputs(4638) <= a or b;
    layer2_outputs(4639) <= not b or a;
    layer2_outputs(4640) <= not b or a;
    layer2_outputs(4641) <= 1'b0;
    layer2_outputs(4642) <= not b;
    layer2_outputs(4643) <= b and not a;
    layer2_outputs(4644) <= b;
    layer2_outputs(4645) <= not (a or b);
    layer2_outputs(4646) <= b;
    layer2_outputs(4647) <= not (a and b);
    layer2_outputs(4648) <= a and b;
    layer2_outputs(4649) <= not (a or b);
    layer2_outputs(4650) <= not a or b;
    layer2_outputs(4651) <= b and not a;
    layer2_outputs(4652) <= a or b;
    layer2_outputs(4653) <= not (a and b);
    layer2_outputs(4654) <= not b or a;
    layer2_outputs(4655) <= not (a or b);
    layer2_outputs(4656) <= b and not a;
    layer2_outputs(4657) <= 1'b0;
    layer2_outputs(4658) <= not a;
    layer2_outputs(4659) <= 1'b1;
    layer2_outputs(4660) <= not a or b;
    layer2_outputs(4661) <= a xor b;
    layer2_outputs(4662) <= 1'b0;
    layer2_outputs(4663) <= b;
    layer2_outputs(4664) <= b and not a;
    layer2_outputs(4665) <= not b;
    layer2_outputs(4666) <= not a or b;
    layer2_outputs(4667) <= not (a or b);
    layer2_outputs(4668) <= not (a and b);
    layer2_outputs(4669) <= a xor b;
    layer2_outputs(4670) <= a or b;
    layer2_outputs(4671) <= b;
    layer2_outputs(4672) <= not (a and b);
    layer2_outputs(4673) <= 1'b1;
    layer2_outputs(4674) <= a and not b;
    layer2_outputs(4675) <= not a or b;
    layer2_outputs(4676) <= 1'b0;
    layer2_outputs(4677) <= 1'b1;
    layer2_outputs(4678) <= 1'b1;
    layer2_outputs(4679) <= 1'b0;
    layer2_outputs(4680) <= 1'b0;
    layer2_outputs(4681) <= not (a xor b);
    layer2_outputs(4682) <= not (a xor b);
    layer2_outputs(4683) <= a;
    layer2_outputs(4684) <= b and not a;
    layer2_outputs(4685) <= not (a or b);
    layer2_outputs(4686) <= a and b;
    layer2_outputs(4687) <= not b;
    layer2_outputs(4688) <= b and not a;
    layer2_outputs(4689) <= not a or b;
    layer2_outputs(4690) <= not (a or b);
    layer2_outputs(4691) <= a or b;
    layer2_outputs(4692) <= a or b;
    layer2_outputs(4693) <= not b;
    layer2_outputs(4694) <= 1'b1;
    layer2_outputs(4695) <= not (a and b);
    layer2_outputs(4696) <= b and not a;
    layer2_outputs(4697) <= b;
    layer2_outputs(4698) <= not (a and b);
    layer2_outputs(4699) <= not a or b;
    layer2_outputs(4700) <= b and not a;
    layer2_outputs(4701) <= not a or b;
    layer2_outputs(4702) <= not (a xor b);
    layer2_outputs(4703) <= not (a or b);
    layer2_outputs(4704) <= not a;
    layer2_outputs(4705) <= b;
    layer2_outputs(4706) <= a or b;
    layer2_outputs(4707) <= a or b;
    layer2_outputs(4708) <= a and not b;
    layer2_outputs(4709) <= a and b;
    layer2_outputs(4710) <= a and not b;
    layer2_outputs(4711) <= not (a xor b);
    layer2_outputs(4712) <= a or b;
    layer2_outputs(4713) <= a and b;
    layer2_outputs(4714) <= not (a and b);
    layer2_outputs(4715) <= a and not b;
    layer2_outputs(4716) <= not (a or b);
    layer2_outputs(4717) <= not (a or b);
    layer2_outputs(4718) <= a and not b;
    layer2_outputs(4719) <= b;
    layer2_outputs(4720) <= not a or b;
    layer2_outputs(4721) <= a and b;
    layer2_outputs(4722) <= not (a xor b);
    layer2_outputs(4723) <= not a;
    layer2_outputs(4724) <= 1'b1;
    layer2_outputs(4725) <= not b;
    layer2_outputs(4726) <= 1'b0;
    layer2_outputs(4727) <= 1'b1;
    layer2_outputs(4728) <= not (a and b);
    layer2_outputs(4729) <= a or b;
    layer2_outputs(4730) <= 1'b1;
    layer2_outputs(4731) <= a;
    layer2_outputs(4732) <= 1'b1;
    layer2_outputs(4733) <= not (a or b);
    layer2_outputs(4734) <= not (a and b);
    layer2_outputs(4735) <= not (a or b);
    layer2_outputs(4736) <= not (a or b);
    layer2_outputs(4737) <= b;
    layer2_outputs(4738) <= not b or a;
    layer2_outputs(4739) <= a and not b;
    layer2_outputs(4740) <= a or b;
    layer2_outputs(4741) <= b;
    layer2_outputs(4742) <= a or b;
    layer2_outputs(4743) <= not b;
    layer2_outputs(4744) <= not b or a;
    layer2_outputs(4745) <= not a or b;
    layer2_outputs(4746) <= not a or b;
    layer2_outputs(4747) <= not a;
    layer2_outputs(4748) <= not b;
    layer2_outputs(4749) <= not b or a;
    layer2_outputs(4750) <= not b;
    layer2_outputs(4751) <= 1'b0;
    layer2_outputs(4752) <= not (a and b);
    layer2_outputs(4753) <= b;
    layer2_outputs(4754) <= not (a and b);
    layer2_outputs(4755) <= a or b;
    layer2_outputs(4756) <= a and b;
    layer2_outputs(4757) <= not (a and b);
    layer2_outputs(4758) <= not a;
    layer2_outputs(4759) <= 1'b1;
    layer2_outputs(4760) <= not (a or b);
    layer2_outputs(4761) <= not a or b;
    layer2_outputs(4762) <= not b or a;
    layer2_outputs(4763) <= a and not b;
    layer2_outputs(4764) <= b and not a;
    layer2_outputs(4765) <= not a or b;
    layer2_outputs(4766) <= 1'b0;
    layer2_outputs(4767) <= b;
    layer2_outputs(4768) <= not b;
    layer2_outputs(4769) <= b;
    layer2_outputs(4770) <= a;
    layer2_outputs(4771) <= 1'b1;
    layer2_outputs(4772) <= not (a and b);
    layer2_outputs(4773) <= a and not b;
    layer2_outputs(4774) <= b and not a;
    layer2_outputs(4775) <= 1'b0;
    layer2_outputs(4776) <= a and not b;
    layer2_outputs(4777) <= a and not b;
    layer2_outputs(4778) <= a or b;
    layer2_outputs(4779) <= not b or a;
    layer2_outputs(4780) <= b;
    layer2_outputs(4781) <= b;
    layer2_outputs(4782) <= a and not b;
    layer2_outputs(4783) <= a and not b;
    layer2_outputs(4784) <= not b or a;
    layer2_outputs(4785) <= not b;
    layer2_outputs(4786) <= 1'b0;
    layer2_outputs(4787) <= not a;
    layer2_outputs(4788) <= 1'b1;
    layer2_outputs(4789) <= not a or b;
    layer2_outputs(4790) <= a or b;
    layer2_outputs(4791) <= a and b;
    layer2_outputs(4792) <= not b or a;
    layer2_outputs(4793) <= b;
    layer2_outputs(4794) <= a or b;
    layer2_outputs(4795) <= not a;
    layer2_outputs(4796) <= 1'b1;
    layer2_outputs(4797) <= a or b;
    layer2_outputs(4798) <= a and not b;
    layer2_outputs(4799) <= a xor b;
    layer2_outputs(4800) <= 1'b1;
    layer2_outputs(4801) <= not a or b;
    layer2_outputs(4802) <= not (a or b);
    layer2_outputs(4803) <= 1'b0;
    layer2_outputs(4804) <= b and not a;
    layer2_outputs(4805) <= 1'b0;
    layer2_outputs(4806) <= not (a and b);
    layer2_outputs(4807) <= not b or a;
    layer2_outputs(4808) <= b;
    layer2_outputs(4809) <= not b;
    layer2_outputs(4810) <= 1'b1;
    layer2_outputs(4811) <= 1'b1;
    layer2_outputs(4812) <= 1'b1;
    layer2_outputs(4813) <= not (a and b);
    layer2_outputs(4814) <= not a;
    layer2_outputs(4815) <= 1'b0;
    layer2_outputs(4816) <= 1'b1;
    layer2_outputs(4817) <= 1'b1;
    layer2_outputs(4818) <= a and not b;
    layer2_outputs(4819) <= not a or b;
    layer2_outputs(4820) <= 1'b1;
    layer2_outputs(4821) <= a or b;
    layer2_outputs(4822) <= 1'b1;
    layer2_outputs(4823) <= not b or a;
    layer2_outputs(4824) <= not a or b;
    layer2_outputs(4825) <= a and not b;
    layer2_outputs(4826) <= a and not b;
    layer2_outputs(4827) <= not (a or b);
    layer2_outputs(4828) <= not b or a;
    layer2_outputs(4829) <= 1'b0;
    layer2_outputs(4830) <= not b;
    layer2_outputs(4831) <= b;
    layer2_outputs(4832) <= not (a or b);
    layer2_outputs(4833) <= not b or a;
    layer2_outputs(4834) <= not a;
    layer2_outputs(4835) <= b and not a;
    layer2_outputs(4836) <= not (a xor b);
    layer2_outputs(4837) <= b and not a;
    layer2_outputs(4838) <= a and b;
    layer2_outputs(4839) <= 1'b0;
    layer2_outputs(4840) <= a and not b;
    layer2_outputs(4841) <= b and not a;
    layer2_outputs(4842) <= not b or a;
    layer2_outputs(4843) <= 1'b1;
    layer2_outputs(4844) <= not (a and b);
    layer2_outputs(4845) <= a or b;
    layer2_outputs(4846) <= a and b;
    layer2_outputs(4847) <= not b;
    layer2_outputs(4848) <= not a or b;
    layer2_outputs(4849) <= 1'b1;
    layer2_outputs(4850) <= a and not b;
    layer2_outputs(4851) <= a or b;
    layer2_outputs(4852) <= not a or b;
    layer2_outputs(4853) <= not b or a;
    layer2_outputs(4854) <= a and not b;
    layer2_outputs(4855) <= 1'b1;
    layer2_outputs(4856) <= 1'b0;
    layer2_outputs(4857) <= 1'b1;
    layer2_outputs(4858) <= not (a xor b);
    layer2_outputs(4859) <= a or b;
    layer2_outputs(4860) <= b;
    layer2_outputs(4861) <= not (a and b);
    layer2_outputs(4862) <= b and not a;
    layer2_outputs(4863) <= 1'b1;
    layer2_outputs(4864) <= not a or b;
    layer2_outputs(4865) <= a xor b;
    layer2_outputs(4866) <= a and not b;
    layer2_outputs(4867) <= a or b;
    layer2_outputs(4868) <= a or b;
    layer2_outputs(4869) <= not a or b;
    layer2_outputs(4870) <= 1'b0;
    layer2_outputs(4871) <= a and b;
    layer2_outputs(4872) <= not a;
    layer2_outputs(4873) <= 1'b1;
    layer2_outputs(4874) <= a and b;
    layer2_outputs(4875) <= not b;
    layer2_outputs(4876) <= not a or b;
    layer2_outputs(4877) <= a or b;
    layer2_outputs(4878) <= not (a or b);
    layer2_outputs(4879) <= not (a xor b);
    layer2_outputs(4880) <= 1'b0;
    layer2_outputs(4881) <= a or b;
    layer2_outputs(4882) <= not (a or b);
    layer2_outputs(4883) <= a and not b;
    layer2_outputs(4884) <= a;
    layer2_outputs(4885) <= not (a and b);
    layer2_outputs(4886) <= not a;
    layer2_outputs(4887) <= a or b;
    layer2_outputs(4888) <= not (a and b);
    layer2_outputs(4889) <= b and not a;
    layer2_outputs(4890) <= not (a xor b);
    layer2_outputs(4891) <= a or b;
    layer2_outputs(4892) <= not b;
    layer2_outputs(4893) <= 1'b0;
    layer2_outputs(4894) <= 1'b1;
    layer2_outputs(4895) <= not (a and b);
    layer2_outputs(4896) <= a or b;
    layer2_outputs(4897) <= not b;
    layer2_outputs(4898) <= a and b;
    layer2_outputs(4899) <= b;
    layer2_outputs(4900) <= 1'b1;
    layer2_outputs(4901) <= a and b;
    layer2_outputs(4902) <= a xor b;
    layer2_outputs(4903) <= 1'b0;
    layer2_outputs(4904) <= 1'b0;
    layer2_outputs(4905) <= 1'b0;
    layer2_outputs(4906) <= 1'b1;
    layer2_outputs(4907) <= not (a or b);
    layer2_outputs(4908) <= not a;
    layer2_outputs(4909) <= not (a or b);
    layer2_outputs(4910) <= not a or b;
    layer2_outputs(4911) <= 1'b0;
    layer2_outputs(4912) <= not a or b;
    layer2_outputs(4913) <= a and b;
    layer2_outputs(4914) <= 1'b0;
    layer2_outputs(4915) <= 1'b1;
    layer2_outputs(4916) <= not a or b;
    layer2_outputs(4917) <= a;
    layer2_outputs(4918) <= 1'b1;
    layer2_outputs(4919) <= a or b;
    layer2_outputs(4920) <= not (a or b);
    layer2_outputs(4921) <= a and not b;
    layer2_outputs(4922) <= a xor b;
    layer2_outputs(4923) <= a;
    layer2_outputs(4924) <= not a or b;
    layer2_outputs(4925) <= not b;
    layer2_outputs(4926) <= not a;
    layer2_outputs(4927) <= a and not b;
    layer2_outputs(4928) <= a and b;
    layer2_outputs(4929) <= a and not b;
    layer2_outputs(4930) <= not a or b;
    layer2_outputs(4931) <= 1'b1;
    layer2_outputs(4932) <= b;
    layer2_outputs(4933) <= not a or b;
    layer2_outputs(4934) <= b;
    layer2_outputs(4935) <= not a or b;
    layer2_outputs(4936) <= a and not b;
    layer2_outputs(4937) <= not a or b;
    layer2_outputs(4938) <= not a;
    layer2_outputs(4939) <= b;
    layer2_outputs(4940) <= not (a or b);
    layer2_outputs(4941) <= not (a and b);
    layer2_outputs(4942) <= not b;
    layer2_outputs(4943) <= not b or a;
    layer2_outputs(4944) <= not (a and b);
    layer2_outputs(4945) <= b;
    layer2_outputs(4946) <= b and not a;
    layer2_outputs(4947) <= not b or a;
    layer2_outputs(4948) <= not a or b;
    layer2_outputs(4949) <= not (a or b);
    layer2_outputs(4950) <= not a;
    layer2_outputs(4951) <= not b or a;
    layer2_outputs(4952) <= not b or a;
    layer2_outputs(4953) <= not b or a;
    layer2_outputs(4954) <= not a;
    layer2_outputs(4955) <= 1'b0;
    layer2_outputs(4956) <= 1'b0;
    layer2_outputs(4957) <= not (a xor b);
    layer2_outputs(4958) <= a and b;
    layer2_outputs(4959) <= b;
    layer2_outputs(4960) <= 1'b0;
    layer2_outputs(4961) <= not a or b;
    layer2_outputs(4962) <= not b or a;
    layer2_outputs(4963) <= 1'b0;
    layer2_outputs(4964) <= a xor b;
    layer2_outputs(4965) <= 1'b0;
    layer2_outputs(4966) <= b and not a;
    layer2_outputs(4967) <= not a;
    layer2_outputs(4968) <= b;
    layer2_outputs(4969) <= 1'b1;
    layer2_outputs(4970) <= not a;
    layer2_outputs(4971) <= 1'b0;
    layer2_outputs(4972) <= not a;
    layer2_outputs(4973) <= b and not a;
    layer2_outputs(4974) <= not (a or b);
    layer2_outputs(4975) <= not b;
    layer2_outputs(4976) <= 1'b0;
    layer2_outputs(4977) <= a;
    layer2_outputs(4978) <= not (a or b);
    layer2_outputs(4979) <= b and not a;
    layer2_outputs(4980) <= a;
    layer2_outputs(4981) <= not a;
    layer2_outputs(4982) <= a and b;
    layer2_outputs(4983) <= a and not b;
    layer2_outputs(4984) <= a or b;
    layer2_outputs(4985) <= 1'b0;
    layer2_outputs(4986) <= b and not a;
    layer2_outputs(4987) <= 1'b0;
    layer2_outputs(4988) <= a and not b;
    layer2_outputs(4989) <= not (a and b);
    layer2_outputs(4990) <= a and not b;
    layer2_outputs(4991) <= not b or a;
    layer2_outputs(4992) <= not a or b;
    layer2_outputs(4993) <= not (a or b);
    layer2_outputs(4994) <= b and not a;
    layer2_outputs(4995) <= not a or b;
    layer2_outputs(4996) <= a;
    layer2_outputs(4997) <= b;
    layer2_outputs(4998) <= 1'b1;
    layer2_outputs(4999) <= not (a and b);
    layer2_outputs(5000) <= 1'b1;
    layer2_outputs(5001) <= a or b;
    layer2_outputs(5002) <= b and not a;
    layer2_outputs(5003) <= b and not a;
    layer2_outputs(5004) <= b and not a;
    layer2_outputs(5005) <= 1'b1;
    layer2_outputs(5006) <= a xor b;
    layer2_outputs(5007) <= b and not a;
    layer2_outputs(5008) <= a or b;
    layer2_outputs(5009) <= a;
    layer2_outputs(5010) <= not a;
    layer2_outputs(5011) <= not a or b;
    layer2_outputs(5012) <= 1'b0;
    layer2_outputs(5013) <= not b or a;
    layer2_outputs(5014) <= not b or a;
    layer2_outputs(5015) <= a;
    layer2_outputs(5016) <= a and b;
    layer2_outputs(5017) <= not b or a;
    layer2_outputs(5018) <= not b or a;
    layer2_outputs(5019) <= 1'b1;
    layer2_outputs(5020) <= 1'b0;
    layer2_outputs(5021) <= b;
    layer2_outputs(5022) <= a and b;
    layer2_outputs(5023) <= not a;
    layer2_outputs(5024) <= 1'b1;
    layer2_outputs(5025) <= a and b;
    layer2_outputs(5026) <= a and not b;
    layer2_outputs(5027) <= not (a and b);
    layer2_outputs(5028) <= not b or a;
    layer2_outputs(5029) <= b;
    layer2_outputs(5030) <= 1'b0;
    layer2_outputs(5031) <= not a;
    layer2_outputs(5032) <= not a;
    layer2_outputs(5033) <= 1'b0;
    layer2_outputs(5034) <= a and b;
    layer2_outputs(5035) <= not a or b;
    layer2_outputs(5036) <= b and not a;
    layer2_outputs(5037) <= not a;
    layer2_outputs(5038) <= a;
    layer2_outputs(5039) <= not b or a;
    layer2_outputs(5040) <= a and b;
    layer2_outputs(5041) <= not (a or b);
    layer2_outputs(5042) <= 1'b0;
    layer2_outputs(5043) <= not (a and b);
    layer2_outputs(5044) <= 1'b0;
    layer2_outputs(5045) <= not (a or b);
    layer2_outputs(5046) <= not (a or b);
    layer2_outputs(5047) <= not b or a;
    layer2_outputs(5048) <= not (a or b);
    layer2_outputs(5049) <= not a or b;
    layer2_outputs(5050) <= a and not b;
    layer2_outputs(5051) <= not (a or b);
    layer2_outputs(5052) <= a or b;
    layer2_outputs(5053) <= a;
    layer2_outputs(5054) <= not (a or b);
    layer2_outputs(5055) <= a xor b;
    layer2_outputs(5056) <= a and not b;
    layer2_outputs(5057) <= a and b;
    layer2_outputs(5058) <= b;
    layer2_outputs(5059) <= not b or a;
    layer2_outputs(5060) <= b and not a;
    layer2_outputs(5061) <= b;
    layer2_outputs(5062) <= not a;
    layer2_outputs(5063) <= b;
    layer2_outputs(5064) <= not a;
    layer2_outputs(5065) <= not (a or b);
    layer2_outputs(5066) <= 1'b0;
    layer2_outputs(5067) <= b;
    layer2_outputs(5068) <= a or b;
    layer2_outputs(5069) <= not b;
    layer2_outputs(5070) <= not (a or b);
    layer2_outputs(5071) <= a and not b;
    layer2_outputs(5072) <= not (a or b);
    layer2_outputs(5073) <= 1'b1;
    layer2_outputs(5074) <= not a;
    layer2_outputs(5075) <= b and not a;
    layer2_outputs(5076) <= not (a and b);
    layer2_outputs(5077) <= 1'b0;
    layer2_outputs(5078) <= a xor b;
    layer2_outputs(5079) <= not b;
    layer2_outputs(5080) <= 1'b0;
    layer2_outputs(5081) <= a xor b;
    layer2_outputs(5082) <= not b;
    layer2_outputs(5083) <= a xor b;
    layer2_outputs(5084) <= not a or b;
    layer2_outputs(5085) <= a and not b;
    layer2_outputs(5086) <= a and b;
    layer2_outputs(5087) <= a and not b;
    layer2_outputs(5088) <= 1'b0;
    layer2_outputs(5089) <= not a;
    layer2_outputs(5090) <= b;
    layer2_outputs(5091) <= 1'b0;
    layer2_outputs(5092) <= not (a or b);
    layer2_outputs(5093) <= a and not b;
    layer2_outputs(5094) <= not (a xor b);
    layer2_outputs(5095) <= a and not b;
    layer2_outputs(5096) <= b and not a;
    layer2_outputs(5097) <= not b;
    layer2_outputs(5098) <= not a or b;
    layer2_outputs(5099) <= a and b;
    layer2_outputs(5100) <= not a or b;
    layer2_outputs(5101) <= a or b;
    layer2_outputs(5102) <= 1'b0;
    layer2_outputs(5103) <= not (a xor b);
    layer2_outputs(5104) <= b;
    layer2_outputs(5105) <= not (a and b);
    layer2_outputs(5106) <= not (a and b);
    layer2_outputs(5107) <= a or b;
    layer2_outputs(5108) <= a or b;
    layer2_outputs(5109) <= not b;
    layer2_outputs(5110) <= not (a and b);
    layer2_outputs(5111) <= not (a or b);
    layer2_outputs(5112) <= not a;
    layer2_outputs(5113) <= not b;
    layer2_outputs(5114) <= not b;
    layer2_outputs(5115) <= a and not b;
    layer2_outputs(5116) <= a or b;
    layer2_outputs(5117) <= not (a or b);
    layer2_outputs(5118) <= not a or b;
    layer2_outputs(5119) <= not (a or b);
    layer2_outputs(5120) <= a and not b;
    layer2_outputs(5121) <= not (a and b);
    layer2_outputs(5122) <= not b;
    layer2_outputs(5123) <= not (a or b);
    layer2_outputs(5124) <= not b or a;
    layer2_outputs(5125) <= a or b;
    layer2_outputs(5126) <= not b;
    layer2_outputs(5127) <= a;
    layer2_outputs(5128) <= not (a xor b);
    layer2_outputs(5129) <= a and b;
    layer2_outputs(5130) <= 1'b1;
    layer2_outputs(5131) <= a and b;
    layer2_outputs(5132) <= b;
    layer2_outputs(5133) <= 1'b1;
    layer2_outputs(5134) <= a and b;
    layer2_outputs(5135) <= a and not b;
    layer2_outputs(5136) <= not a or b;
    layer2_outputs(5137) <= 1'b0;
    layer2_outputs(5138) <= a and b;
    layer2_outputs(5139) <= a xor b;
    layer2_outputs(5140) <= not a or b;
    layer2_outputs(5141) <= 1'b0;
    layer2_outputs(5142) <= b and not a;
    layer2_outputs(5143) <= a and b;
    layer2_outputs(5144) <= not a;
    layer2_outputs(5145) <= a and b;
    layer2_outputs(5146) <= not a or b;
    layer2_outputs(5147) <= not b;
    layer2_outputs(5148) <= b;
    layer2_outputs(5149) <= a and b;
    layer2_outputs(5150) <= a and not b;
    layer2_outputs(5151) <= a and b;
    layer2_outputs(5152) <= not b or a;
    layer2_outputs(5153) <= not (a and b);
    layer2_outputs(5154) <= not (a and b);
    layer2_outputs(5155) <= a and b;
    layer2_outputs(5156) <= 1'b0;
    layer2_outputs(5157) <= 1'b1;
    layer2_outputs(5158) <= b and not a;
    layer2_outputs(5159) <= a xor b;
    layer2_outputs(5160) <= not b or a;
    layer2_outputs(5161) <= b;
    layer2_outputs(5162) <= 1'b1;
    layer2_outputs(5163) <= 1'b0;
    layer2_outputs(5164) <= 1'b1;
    layer2_outputs(5165) <= 1'b0;
    layer2_outputs(5166) <= 1'b1;
    layer2_outputs(5167) <= not b;
    layer2_outputs(5168) <= not b;
    layer2_outputs(5169) <= 1'b1;
    layer2_outputs(5170) <= 1'b1;
    layer2_outputs(5171) <= b and not a;
    layer2_outputs(5172) <= not (a xor b);
    layer2_outputs(5173) <= 1'b0;
    layer2_outputs(5174) <= 1'b0;
    layer2_outputs(5175) <= not a;
    layer2_outputs(5176) <= not b or a;
    layer2_outputs(5177) <= a;
    layer2_outputs(5178) <= 1'b0;
    layer2_outputs(5179) <= not b or a;
    layer2_outputs(5180) <= not b;
    layer2_outputs(5181) <= not b;
    layer2_outputs(5182) <= a and not b;
    layer2_outputs(5183) <= not a;
    layer2_outputs(5184) <= 1'b0;
    layer2_outputs(5185) <= 1'b1;
    layer2_outputs(5186) <= not a;
    layer2_outputs(5187) <= a or b;
    layer2_outputs(5188) <= 1'b0;
    layer2_outputs(5189) <= a and not b;
    layer2_outputs(5190) <= not b;
    layer2_outputs(5191) <= 1'b1;
    layer2_outputs(5192) <= 1'b0;
    layer2_outputs(5193) <= 1'b1;
    layer2_outputs(5194) <= a or b;
    layer2_outputs(5195) <= not a;
    layer2_outputs(5196) <= 1'b1;
    layer2_outputs(5197) <= a and not b;
    layer2_outputs(5198) <= a or b;
    layer2_outputs(5199) <= 1'b1;
    layer2_outputs(5200) <= a and not b;
    layer2_outputs(5201) <= not a;
    layer2_outputs(5202) <= not b;
    layer2_outputs(5203) <= b and not a;
    layer2_outputs(5204) <= a and not b;
    layer2_outputs(5205) <= 1'b0;
    layer2_outputs(5206) <= 1'b0;
    layer2_outputs(5207) <= not a;
    layer2_outputs(5208) <= b and not a;
    layer2_outputs(5209) <= b;
    layer2_outputs(5210) <= a xor b;
    layer2_outputs(5211) <= 1'b0;
    layer2_outputs(5212) <= a and b;
    layer2_outputs(5213) <= a and not b;
    layer2_outputs(5214) <= a and not b;
    layer2_outputs(5215) <= b and not a;
    layer2_outputs(5216) <= 1'b1;
    layer2_outputs(5217) <= not (a and b);
    layer2_outputs(5218) <= b;
    layer2_outputs(5219) <= a and b;
    layer2_outputs(5220) <= b and not a;
    layer2_outputs(5221) <= b;
    layer2_outputs(5222) <= not b;
    layer2_outputs(5223) <= not a;
    layer2_outputs(5224) <= b and not a;
    layer2_outputs(5225) <= not a or b;
    layer2_outputs(5226) <= a and b;
    layer2_outputs(5227) <= not b or a;
    layer2_outputs(5228) <= b and not a;
    layer2_outputs(5229) <= a and not b;
    layer2_outputs(5230) <= a;
    layer2_outputs(5231) <= a;
    layer2_outputs(5232) <= not (a and b);
    layer2_outputs(5233) <= 1'b0;
    layer2_outputs(5234) <= a and b;
    layer2_outputs(5235) <= 1'b0;
    layer2_outputs(5236) <= not (a or b);
    layer2_outputs(5237) <= not (a or b);
    layer2_outputs(5238) <= not a or b;
    layer2_outputs(5239) <= not b;
    layer2_outputs(5240) <= 1'b1;
    layer2_outputs(5241) <= b and not a;
    layer2_outputs(5242) <= 1'b0;
    layer2_outputs(5243) <= 1'b0;
    layer2_outputs(5244) <= a;
    layer2_outputs(5245) <= a;
    layer2_outputs(5246) <= not a or b;
    layer2_outputs(5247) <= 1'b0;
    layer2_outputs(5248) <= b;
    layer2_outputs(5249) <= 1'b1;
    layer2_outputs(5250) <= b and not a;
    layer2_outputs(5251) <= a and b;
    layer2_outputs(5252) <= a and b;
    layer2_outputs(5253) <= b;
    layer2_outputs(5254) <= a xor b;
    layer2_outputs(5255) <= a and b;
    layer2_outputs(5256) <= a or b;
    layer2_outputs(5257) <= b and not a;
    layer2_outputs(5258) <= a;
    layer2_outputs(5259) <= a or b;
    layer2_outputs(5260) <= 1'b0;
    layer2_outputs(5261) <= not a;
    layer2_outputs(5262) <= not a;
    layer2_outputs(5263) <= b;
    layer2_outputs(5264) <= a;
    layer2_outputs(5265) <= b and not a;
    layer2_outputs(5266) <= 1'b1;
    layer2_outputs(5267) <= b and not a;
    layer2_outputs(5268) <= not b or a;
    layer2_outputs(5269) <= not a or b;
    layer2_outputs(5270) <= a and b;
    layer2_outputs(5271) <= not b or a;
    layer2_outputs(5272) <= not (a or b);
    layer2_outputs(5273) <= not b or a;
    layer2_outputs(5274) <= a or b;
    layer2_outputs(5275) <= not b;
    layer2_outputs(5276) <= 1'b0;
    layer2_outputs(5277) <= 1'b1;
    layer2_outputs(5278) <= not b or a;
    layer2_outputs(5279) <= not (a or b);
    layer2_outputs(5280) <= 1'b1;
    layer2_outputs(5281) <= not a or b;
    layer2_outputs(5282) <= not a;
    layer2_outputs(5283) <= not (a xor b);
    layer2_outputs(5284) <= b;
    layer2_outputs(5285) <= 1'b0;
    layer2_outputs(5286) <= not b or a;
    layer2_outputs(5287) <= a and b;
    layer2_outputs(5288) <= 1'b1;
    layer2_outputs(5289) <= not (a xor b);
    layer2_outputs(5290) <= 1'b0;
    layer2_outputs(5291) <= 1'b1;
    layer2_outputs(5292) <= 1'b1;
    layer2_outputs(5293) <= not a;
    layer2_outputs(5294) <= a;
    layer2_outputs(5295) <= not a;
    layer2_outputs(5296) <= not b or a;
    layer2_outputs(5297) <= b;
    layer2_outputs(5298) <= a;
    layer2_outputs(5299) <= a;
    layer2_outputs(5300) <= not b or a;
    layer2_outputs(5301) <= not a;
    layer2_outputs(5302) <= a and not b;
    layer2_outputs(5303) <= a and b;
    layer2_outputs(5304) <= not a;
    layer2_outputs(5305) <= not a;
    layer2_outputs(5306) <= 1'b1;
    layer2_outputs(5307) <= a and not b;
    layer2_outputs(5308) <= a and not b;
    layer2_outputs(5309) <= not (a or b);
    layer2_outputs(5310) <= a;
    layer2_outputs(5311) <= 1'b0;
    layer2_outputs(5312) <= not (a xor b);
    layer2_outputs(5313) <= b and not a;
    layer2_outputs(5314) <= 1'b1;
    layer2_outputs(5315) <= a xor b;
    layer2_outputs(5316) <= a and b;
    layer2_outputs(5317) <= not (a xor b);
    layer2_outputs(5318) <= a and not b;
    layer2_outputs(5319) <= not a;
    layer2_outputs(5320) <= a;
    layer2_outputs(5321) <= not b;
    layer2_outputs(5322) <= not (a and b);
    layer2_outputs(5323) <= b;
    layer2_outputs(5324) <= a and not b;
    layer2_outputs(5325) <= a;
    layer2_outputs(5326) <= a and not b;
    layer2_outputs(5327) <= a and b;
    layer2_outputs(5328) <= not b or a;
    layer2_outputs(5329) <= not (a and b);
    layer2_outputs(5330) <= not b or a;
    layer2_outputs(5331) <= a and b;
    layer2_outputs(5332) <= not (a and b);
    layer2_outputs(5333) <= not (a and b);
    layer2_outputs(5334) <= not (a and b);
    layer2_outputs(5335) <= not a;
    layer2_outputs(5336) <= not b;
    layer2_outputs(5337) <= 1'b0;
    layer2_outputs(5338) <= 1'b1;
    layer2_outputs(5339) <= not (a and b);
    layer2_outputs(5340) <= a;
    layer2_outputs(5341) <= not (a xor b);
    layer2_outputs(5342) <= 1'b1;
    layer2_outputs(5343) <= not b or a;
    layer2_outputs(5344) <= a or b;
    layer2_outputs(5345) <= 1'b0;
    layer2_outputs(5346) <= b and not a;
    layer2_outputs(5347) <= a and b;
    layer2_outputs(5348) <= not (a xor b);
    layer2_outputs(5349) <= b and not a;
    layer2_outputs(5350) <= not b or a;
    layer2_outputs(5351) <= not b or a;
    layer2_outputs(5352) <= a and not b;
    layer2_outputs(5353) <= not a;
    layer2_outputs(5354) <= not (a xor b);
    layer2_outputs(5355) <= 1'b0;
    layer2_outputs(5356) <= a and not b;
    layer2_outputs(5357) <= a and b;
    layer2_outputs(5358) <= a or b;
    layer2_outputs(5359) <= b and not a;
    layer2_outputs(5360) <= a;
    layer2_outputs(5361) <= 1'b0;
    layer2_outputs(5362) <= 1'b0;
    layer2_outputs(5363) <= not (a or b);
    layer2_outputs(5364) <= 1'b1;
    layer2_outputs(5365) <= not b;
    layer2_outputs(5366) <= 1'b1;
    layer2_outputs(5367) <= 1'b1;
    layer2_outputs(5368) <= a and b;
    layer2_outputs(5369) <= b;
    layer2_outputs(5370) <= 1'b0;
    layer2_outputs(5371) <= not a;
    layer2_outputs(5372) <= b and not a;
    layer2_outputs(5373) <= not (a or b);
    layer2_outputs(5374) <= a or b;
    layer2_outputs(5375) <= b;
    layer2_outputs(5376) <= a and b;
    layer2_outputs(5377) <= not b;
    layer2_outputs(5378) <= not b or a;
    layer2_outputs(5379) <= not b;
    layer2_outputs(5380) <= a;
    layer2_outputs(5381) <= b and not a;
    layer2_outputs(5382) <= b;
    layer2_outputs(5383) <= b and not a;
    layer2_outputs(5384) <= a and b;
    layer2_outputs(5385) <= b;
    layer2_outputs(5386) <= not (a or b);
    layer2_outputs(5387) <= not b or a;
    layer2_outputs(5388) <= not b or a;
    layer2_outputs(5389) <= not a or b;
    layer2_outputs(5390) <= not a or b;
    layer2_outputs(5391) <= a and not b;
    layer2_outputs(5392) <= not (a or b);
    layer2_outputs(5393) <= 1'b0;
    layer2_outputs(5394) <= not b or a;
    layer2_outputs(5395) <= a;
    layer2_outputs(5396) <= b;
    layer2_outputs(5397) <= not a;
    layer2_outputs(5398) <= a and b;
    layer2_outputs(5399) <= not a or b;
    layer2_outputs(5400) <= b;
    layer2_outputs(5401) <= a or b;
    layer2_outputs(5402) <= a and not b;
    layer2_outputs(5403) <= a and b;
    layer2_outputs(5404) <= 1'b1;
    layer2_outputs(5405) <= a;
    layer2_outputs(5406) <= a;
    layer2_outputs(5407) <= not a;
    layer2_outputs(5408) <= not (a or b);
    layer2_outputs(5409) <= a and not b;
    layer2_outputs(5410) <= a and not b;
    layer2_outputs(5411) <= a and b;
    layer2_outputs(5412) <= 1'b0;
    layer2_outputs(5413) <= not (a or b);
    layer2_outputs(5414) <= b;
    layer2_outputs(5415) <= not a;
    layer2_outputs(5416) <= a and b;
    layer2_outputs(5417) <= b and not a;
    layer2_outputs(5418) <= 1'b0;
    layer2_outputs(5419) <= 1'b1;
    layer2_outputs(5420) <= not b or a;
    layer2_outputs(5421) <= b;
    layer2_outputs(5422) <= a and b;
    layer2_outputs(5423) <= not (a or b);
    layer2_outputs(5424) <= a and not b;
    layer2_outputs(5425) <= a or b;
    layer2_outputs(5426) <= b and not a;
    layer2_outputs(5427) <= not a or b;
    layer2_outputs(5428) <= b and not a;
    layer2_outputs(5429) <= b and not a;
    layer2_outputs(5430) <= not (a and b);
    layer2_outputs(5431) <= not (a xor b);
    layer2_outputs(5432) <= not b;
    layer2_outputs(5433) <= a and not b;
    layer2_outputs(5434) <= not (a and b);
    layer2_outputs(5435) <= not a;
    layer2_outputs(5436) <= 1'b1;
    layer2_outputs(5437) <= 1'b1;
    layer2_outputs(5438) <= 1'b1;
    layer2_outputs(5439) <= a xor b;
    layer2_outputs(5440) <= 1'b1;
    layer2_outputs(5441) <= b and not a;
    layer2_outputs(5442) <= a or b;
    layer2_outputs(5443) <= not (a or b);
    layer2_outputs(5444) <= a and b;
    layer2_outputs(5445) <= a xor b;
    layer2_outputs(5446) <= not (a or b);
    layer2_outputs(5447) <= a and b;
    layer2_outputs(5448) <= a and not b;
    layer2_outputs(5449) <= a or b;
    layer2_outputs(5450) <= not (a and b);
    layer2_outputs(5451) <= a and b;
    layer2_outputs(5452) <= not a or b;
    layer2_outputs(5453) <= a and not b;
    layer2_outputs(5454) <= 1'b1;
    layer2_outputs(5455) <= 1'b1;
    layer2_outputs(5456) <= b and not a;
    layer2_outputs(5457) <= not (a xor b);
    layer2_outputs(5458) <= a;
    layer2_outputs(5459) <= a;
    layer2_outputs(5460) <= a;
    layer2_outputs(5461) <= a and not b;
    layer2_outputs(5462) <= not b or a;
    layer2_outputs(5463) <= 1'b1;
    layer2_outputs(5464) <= not a or b;
    layer2_outputs(5465) <= b;
    layer2_outputs(5466) <= a and b;
    layer2_outputs(5467) <= a and not b;
    layer2_outputs(5468) <= not a or b;
    layer2_outputs(5469) <= a and b;
    layer2_outputs(5470) <= not b;
    layer2_outputs(5471) <= not (a or b);
    layer2_outputs(5472) <= not b or a;
    layer2_outputs(5473) <= 1'b1;
    layer2_outputs(5474) <= a and b;
    layer2_outputs(5475) <= 1'b0;
    layer2_outputs(5476) <= a and b;
    layer2_outputs(5477) <= not (a and b);
    layer2_outputs(5478) <= not (a or b);
    layer2_outputs(5479) <= not a or b;
    layer2_outputs(5480) <= a and not b;
    layer2_outputs(5481) <= a and b;
    layer2_outputs(5482) <= not (a or b);
    layer2_outputs(5483) <= not (a and b);
    layer2_outputs(5484) <= a and not b;
    layer2_outputs(5485) <= 1'b1;
    layer2_outputs(5486) <= a and b;
    layer2_outputs(5487) <= not b or a;
    layer2_outputs(5488) <= not a;
    layer2_outputs(5489) <= not b or a;
    layer2_outputs(5490) <= 1'b0;
    layer2_outputs(5491) <= not b or a;
    layer2_outputs(5492) <= a and not b;
    layer2_outputs(5493) <= 1'b1;
    layer2_outputs(5494) <= not (a and b);
    layer2_outputs(5495) <= b and not a;
    layer2_outputs(5496) <= not b or a;
    layer2_outputs(5497) <= a and not b;
    layer2_outputs(5498) <= 1'b1;
    layer2_outputs(5499) <= a or b;
    layer2_outputs(5500) <= not (a and b);
    layer2_outputs(5501) <= a and b;
    layer2_outputs(5502) <= not b or a;
    layer2_outputs(5503) <= not a or b;
    layer2_outputs(5504) <= not (a or b);
    layer2_outputs(5505) <= a and b;
    layer2_outputs(5506) <= 1'b1;
    layer2_outputs(5507) <= not (a and b);
    layer2_outputs(5508) <= a and not b;
    layer2_outputs(5509) <= a or b;
    layer2_outputs(5510) <= b;
    layer2_outputs(5511) <= not (a and b);
    layer2_outputs(5512) <= not (a and b);
    layer2_outputs(5513) <= not (a and b);
    layer2_outputs(5514) <= 1'b0;
    layer2_outputs(5515) <= a and not b;
    layer2_outputs(5516) <= a or b;
    layer2_outputs(5517) <= b;
    layer2_outputs(5518) <= not b;
    layer2_outputs(5519) <= 1'b0;
    layer2_outputs(5520) <= not a or b;
    layer2_outputs(5521) <= 1'b0;
    layer2_outputs(5522) <= b and not a;
    layer2_outputs(5523) <= a and b;
    layer2_outputs(5524) <= not a;
    layer2_outputs(5525) <= a;
    layer2_outputs(5526) <= a or b;
    layer2_outputs(5527) <= a or b;
    layer2_outputs(5528) <= not a;
    layer2_outputs(5529) <= a and not b;
    layer2_outputs(5530) <= b and not a;
    layer2_outputs(5531) <= 1'b1;
    layer2_outputs(5532) <= a or b;
    layer2_outputs(5533) <= not (a or b);
    layer2_outputs(5534) <= not b;
    layer2_outputs(5535) <= not a or b;
    layer2_outputs(5536) <= b and not a;
    layer2_outputs(5537) <= not b;
    layer2_outputs(5538) <= not b;
    layer2_outputs(5539) <= b;
    layer2_outputs(5540) <= 1'b1;
    layer2_outputs(5541) <= not (a and b);
    layer2_outputs(5542) <= a and b;
    layer2_outputs(5543) <= not a or b;
    layer2_outputs(5544) <= not a;
    layer2_outputs(5545) <= not (a or b);
    layer2_outputs(5546) <= a and not b;
    layer2_outputs(5547) <= not a;
    layer2_outputs(5548) <= not b;
    layer2_outputs(5549) <= not (a and b);
    layer2_outputs(5550) <= not a or b;
    layer2_outputs(5551) <= a and b;
    layer2_outputs(5552) <= not (a and b);
    layer2_outputs(5553) <= not a;
    layer2_outputs(5554) <= 1'b0;
    layer2_outputs(5555) <= a and not b;
    layer2_outputs(5556) <= not a or b;
    layer2_outputs(5557) <= b and not a;
    layer2_outputs(5558) <= not (a and b);
    layer2_outputs(5559) <= 1'b1;
    layer2_outputs(5560) <= a and not b;
    layer2_outputs(5561) <= not a or b;
    layer2_outputs(5562) <= a and b;
    layer2_outputs(5563) <= 1'b0;
    layer2_outputs(5564) <= b and not a;
    layer2_outputs(5565) <= not (a and b);
    layer2_outputs(5566) <= not (a or b);
    layer2_outputs(5567) <= not (a or b);
    layer2_outputs(5568) <= 1'b1;
    layer2_outputs(5569) <= 1'b1;
    layer2_outputs(5570) <= 1'b1;
    layer2_outputs(5571) <= not a;
    layer2_outputs(5572) <= b;
    layer2_outputs(5573) <= a and not b;
    layer2_outputs(5574) <= not a or b;
    layer2_outputs(5575) <= not a;
    layer2_outputs(5576) <= b;
    layer2_outputs(5577) <= a or b;
    layer2_outputs(5578) <= not b or a;
    layer2_outputs(5579) <= a and not b;
    layer2_outputs(5580) <= not (a or b);
    layer2_outputs(5581) <= b;
    layer2_outputs(5582) <= not a;
    layer2_outputs(5583) <= not a;
    layer2_outputs(5584) <= not (a and b);
    layer2_outputs(5585) <= not a or b;
    layer2_outputs(5586) <= a;
    layer2_outputs(5587) <= a or b;
    layer2_outputs(5588) <= a and b;
    layer2_outputs(5589) <= not b or a;
    layer2_outputs(5590) <= not a;
    layer2_outputs(5591) <= not (a or b);
    layer2_outputs(5592) <= b;
    layer2_outputs(5593) <= not (a or b);
    layer2_outputs(5594) <= b and not a;
    layer2_outputs(5595) <= not a or b;
    layer2_outputs(5596) <= b;
    layer2_outputs(5597) <= not b or a;
    layer2_outputs(5598) <= 1'b0;
    layer2_outputs(5599) <= a or b;
    layer2_outputs(5600) <= a and b;
    layer2_outputs(5601) <= not (a or b);
    layer2_outputs(5602) <= not b or a;
    layer2_outputs(5603) <= not b;
    layer2_outputs(5604) <= not a or b;
    layer2_outputs(5605) <= b and not a;
    layer2_outputs(5606) <= 1'b1;
    layer2_outputs(5607) <= b and not a;
    layer2_outputs(5608) <= b;
    layer2_outputs(5609) <= a xor b;
    layer2_outputs(5610) <= 1'b0;
    layer2_outputs(5611) <= a;
    layer2_outputs(5612) <= a;
    layer2_outputs(5613) <= not a or b;
    layer2_outputs(5614) <= not (a and b);
    layer2_outputs(5615) <= b;
    layer2_outputs(5616) <= 1'b0;
    layer2_outputs(5617) <= not b;
    layer2_outputs(5618) <= 1'b0;
    layer2_outputs(5619) <= 1'b1;
    layer2_outputs(5620) <= 1'b1;
    layer2_outputs(5621) <= not (a or b);
    layer2_outputs(5622) <= 1'b0;
    layer2_outputs(5623) <= not (a xor b);
    layer2_outputs(5624) <= a and b;
    layer2_outputs(5625) <= a;
    layer2_outputs(5626) <= b;
    layer2_outputs(5627) <= 1'b0;
    layer2_outputs(5628) <= not (a and b);
    layer2_outputs(5629) <= not (a and b);
    layer2_outputs(5630) <= b and not a;
    layer2_outputs(5631) <= 1'b1;
    layer2_outputs(5632) <= not b;
    layer2_outputs(5633) <= not b;
    layer2_outputs(5634) <= b;
    layer2_outputs(5635) <= a and not b;
    layer2_outputs(5636) <= not b;
    layer2_outputs(5637) <= b and not a;
    layer2_outputs(5638) <= not (a or b);
    layer2_outputs(5639) <= 1'b0;
    layer2_outputs(5640) <= b;
    layer2_outputs(5641) <= not b or a;
    layer2_outputs(5642) <= a;
    layer2_outputs(5643) <= not b or a;
    layer2_outputs(5644) <= not (a and b);
    layer2_outputs(5645) <= a;
    layer2_outputs(5646) <= not b or a;
    layer2_outputs(5647) <= a and b;
    layer2_outputs(5648) <= a or b;
    layer2_outputs(5649) <= 1'b1;
    layer2_outputs(5650) <= 1'b0;
    layer2_outputs(5651) <= not b or a;
    layer2_outputs(5652) <= a or b;
    layer2_outputs(5653) <= a and not b;
    layer2_outputs(5654) <= not a or b;
    layer2_outputs(5655) <= 1'b1;
    layer2_outputs(5656) <= a;
    layer2_outputs(5657) <= not b or a;
    layer2_outputs(5658) <= not (a xor b);
    layer2_outputs(5659) <= 1'b0;
    layer2_outputs(5660) <= not b;
    layer2_outputs(5661) <= 1'b0;
    layer2_outputs(5662) <= not a or b;
    layer2_outputs(5663) <= not (a and b);
    layer2_outputs(5664) <= a;
    layer2_outputs(5665) <= a and b;
    layer2_outputs(5666) <= a and not b;
    layer2_outputs(5667) <= 1'b1;
    layer2_outputs(5668) <= a;
    layer2_outputs(5669) <= a and b;
    layer2_outputs(5670) <= a or b;
    layer2_outputs(5671) <= b and not a;
    layer2_outputs(5672) <= a and b;
    layer2_outputs(5673) <= b and not a;
    layer2_outputs(5674) <= a and b;
    layer2_outputs(5675) <= a or b;
    layer2_outputs(5676) <= 1'b0;
    layer2_outputs(5677) <= a xor b;
    layer2_outputs(5678) <= not a;
    layer2_outputs(5679) <= 1'b1;
    layer2_outputs(5680) <= 1'b1;
    layer2_outputs(5681) <= not b;
    layer2_outputs(5682) <= not a or b;
    layer2_outputs(5683) <= not b;
    layer2_outputs(5684) <= a and not b;
    layer2_outputs(5685) <= a and b;
    layer2_outputs(5686) <= b and not a;
    layer2_outputs(5687) <= not b or a;
    layer2_outputs(5688) <= a and b;
    layer2_outputs(5689) <= a;
    layer2_outputs(5690) <= b and not a;
    layer2_outputs(5691) <= not (a or b);
    layer2_outputs(5692) <= a and not b;
    layer2_outputs(5693) <= not (a and b);
    layer2_outputs(5694) <= not b or a;
    layer2_outputs(5695) <= a and b;
    layer2_outputs(5696) <= 1'b0;
    layer2_outputs(5697) <= a;
    layer2_outputs(5698) <= not a;
    layer2_outputs(5699) <= a and b;
    layer2_outputs(5700) <= 1'b1;
    layer2_outputs(5701) <= a and b;
    layer2_outputs(5702) <= 1'b0;
    layer2_outputs(5703) <= not a or b;
    layer2_outputs(5704) <= not b;
    layer2_outputs(5705) <= not a;
    layer2_outputs(5706) <= 1'b0;
    layer2_outputs(5707) <= 1'b1;
    layer2_outputs(5708) <= not a or b;
    layer2_outputs(5709) <= a and b;
    layer2_outputs(5710) <= not b or a;
    layer2_outputs(5711) <= not (a and b);
    layer2_outputs(5712) <= not a or b;
    layer2_outputs(5713) <= b and not a;
    layer2_outputs(5714) <= a or b;
    layer2_outputs(5715) <= a xor b;
    layer2_outputs(5716) <= not a;
    layer2_outputs(5717) <= not a or b;
    layer2_outputs(5718) <= not b or a;
    layer2_outputs(5719) <= 1'b1;
    layer2_outputs(5720) <= 1'b1;
    layer2_outputs(5721) <= not a or b;
    layer2_outputs(5722) <= not a or b;
    layer2_outputs(5723) <= a or b;
    layer2_outputs(5724) <= a and b;
    layer2_outputs(5725) <= not a;
    layer2_outputs(5726) <= a and not b;
    layer2_outputs(5727) <= 1'b1;
    layer2_outputs(5728) <= not a or b;
    layer2_outputs(5729) <= 1'b0;
    layer2_outputs(5730) <= 1'b1;
    layer2_outputs(5731) <= not (a and b);
    layer2_outputs(5732) <= b and not a;
    layer2_outputs(5733) <= a or b;
    layer2_outputs(5734) <= a and b;
    layer2_outputs(5735) <= a or b;
    layer2_outputs(5736) <= not b;
    layer2_outputs(5737) <= b;
    layer2_outputs(5738) <= not (a and b);
    layer2_outputs(5739) <= b;
    layer2_outputs(5740) <= a xor b;
    layer2_outputs(5741) <= not a or b;
    layer2_outputs(5742) <= a;
    layer2_outputs(5743) <= a and b;
    layer2_outputs(5744) <= not a;
    layer2_outputs(5745) <= a;
    layer2_outputs(5746) <= b and not a;
    layer2_outputs(5747) <= a xor b;
    layer2_outputs(5748) <= b;
    layer2_outputs(5749) <= not a or b;
    layer2_outputs(5750) <= not (a and b);
    layer2_outputs(5751) <= 1'b1;
    layer2_outputs(5752) <= a and not b;
    layer2_outputs(5753) <= a and b;
    layer2_outputs(5754) <= a xor b;
    layer2_outputs(5755) <= not (a or b);
    layer2_outputs(5756) <= a and not b;
    layer2_outputs(5757) <= not a;
    layer2_outputs(5758) <= not b or a;
    layer2_outputs(5759) <= 1'b0;
    layer2_outputs(5760) <= a and b;
    layer2_outputs(5761) <= a xor b;
    layer2_outputs(5762) <= 1'b1;
    layer2_outputs(5763) <= a and not b;
    layer2_outputs(5764) <= not (a and b);
    layer2_outputs(5765) <= 1'b1;
    layer2_outputs(5766) <= not a;
    layer2_outputs(5767) <= not b or a;
    layer2_outputs(5768) <= a;
    layer2_outputs(5769) <= a;
    layer2_outputs(5770) <= not a;
    layer2_outputs(5771) <= not b or a;
    layer2_outputs(5772) <= 1'b0;
    layer2_outputs(5773) <= b;
    layer2_outputs(5774) <= 1'b1;
    layer2_outputs(5775) <= not b or a;
    layer2_outputs(5776) <= not a;
    layer2_outputs(5777) <= 1'b1;
    layer2_outputs(5778) <= b;
    layer2_outputs(5779) <= not b;
    layer2_outputs(5780) <= not a or b;
    layer2_outputs(5781) <= not b;
    layer2_outputs(5782) <= a and not b;
    layer2_outputs(5783) <= a and not b;
    layer2_outputs(5784) <= a or b;
    layer2_outputs(5785) <= not b or a;
    layer2_outputs(5786) <= 1'b1;
    layer2_outputs(5787) <= not (a xor b);
    layer2_outputs(5788) <= not (a and b);
    layer2_outputs(5789) <= a and b;
    layer2_outputs(5790) <= 1'b0;
    layer2_outputs(5791) <= not (a xor b);
    layer2_outputs(5792) <= not b or a;
    layer2_outputs(5793) <= 1'b0;
    layer2_outputs(5794) <= a and not b;
    layer2_outputs(5795) <= not b or a;
    layer2_outputs(5796) <= b and not a;
    layer2_outputs(5797) <= not b or a;
    layer2_outputs(5798) <= not (a xor b);
    layer2_outputs(5799) <= not a;
    layer2_outputs(5800) <= a xor b;
    layer2_outputs(5801) <= a;
    layer2_outputs(5802) <= a;
    layer2_outputs(5803) <= not a or b;
    layer2_outputs(5804) <= a and b;
    layer2_outputs(5805) <= a and b;
    layer2_outputs(5806) <= not b or a;
    layer2_outputs(5807) <= not b or a;
    layer2_outputs(5808) <= not b;
    layer2_outputs(5809) <= b and not a;
    layer2_outputs(5810) <= not b;
    layer2_outputs(5811) <= a and not b;
    layer2_outputs(5812) <= not a or b;
    layer2_outputs(5813) <= a and not b;
    layer2_outputs(5814) <= b and not a;
    layer2_outputs(5815) <= not (a xor b);
    layer2_outputs(5816) <= not b or a;
    layer2_outputs(5817) <= b;
    layer2_outputs(5818) <= a and not b;
    layer2_outputs(5819) <= a and not b;
    layer2_outputs(5820) <= not b;
    layer2_outputs(5821) <= not (a xor b);
    layer2_outputs(5822) <= 1'b0;
    layer2_outputs(5823) <= 1'b0;
    layer2_outputs(5824) <= a;
    layer2_outputs(5825) <= b;
    layer2_outputs(5826) <= not b;
    layer2_outputs(5827) <= not b or a;
    layer2_outputs(5828) <= a and not b;
    layer2_outputs(5829) <= a or b;
    layer2_outputs(5830) <= not b;
    layer2_outputs(5831) <= b and not a;
    layer2_outputs(5832) <= a or b;
    layer2_outputs(5833) <= a and b;
    layer2_outputs(5834) <= b and not a;
    layer2_outputs(5835) <= not b;
    layer2_outputs(5836) <= b;
    layer2_outputs(5837) <= not b or a;
    layer2_outputs(5838) <= not a;
    layer2_outputs(5839) <= a and b;
    layer2_outputs(5840) <= 1'b0;
    layer2_outputs(5841) <= not (a or b);
    layer2_outputs(5842) <= a and not b;
    layer2_outputs(5843) <= not b or a;
    layer2_outputs(5844) <= b;
    layer2_outputs(5845) <= not a or b;
    layer2_outputs(5846) <= not b or a;
    layer2_outputs(5847) <= not b;
    layer2_outputs(5848) <= 1'b0;
    layer2_outputs(5849) <= a or b;
    layer2_outputs(5850) <= b;
    layer2_outputs(5851) <= not (a and b);
    layer2_outputs(5852) <= 1'b1;
    layer2_outputs(5853) <= 1'b0;
    layer2_outputs(5854) <= a or b;
    layer2_outputs(5855) <= b;
    layer2_outputs(5856) <= not (a and b);
    layer2_outputs(5857) <= a and not b;
    layer2_outputs(5858) <= not (a or b);
    layer2_outputs(5859) <= not (a and b);
    layer2_outputs(5860) <= b and not a;
    layer2_outputs(5861) <= a;
    layer2_outputs(5862) <= a and not b;
    layer2_outputs(5863) <= not b;
    layer2_outputs(5864) <= not (a or b);
    layer2_outputs(5865) <= not a;
    layer2_outputs(5866) <= a or b;
    layer2_outputs(5867) <= b;
    layer2_outputs(5868) <= not b;
    layer2_outputs(5869) <= a xor b;
    layer2_outputs(5870) <= not b;
    layer2_outputs(5871) <= not a or b;
    layer2_outputs(5872) <= a or b;
    layer2_outputs(5873) <= not (a and b);
    layer2_outputs(5874) <= not a or b;
    layer2_outputs(5875) <= a;
    layer2_outputs(5876) <= a and not b;
    layer2_outputs(5877) <= a and not b;
    layer2_outputs(5878) <= a and not b;
    layer2_outputs(5879) <= 1'b0;
    layer2_outputs(5880) <= not (a or b);
    layer2_outputs(5881) <= not (a xor b);
    layer2_outputs(5882) <= a and not b;
    layer2_outputs(5883) <= not (a xor b);
    layer2_outputs(5884) <= a or b;
    layer2_outputs(5885) <= a xor b;
    layer2_outputs(5886) <= b and not a;
    layer2_outputs(5887) <= b and not a;
    layer2_outputs(5888) <= not (a and b);
    layer2_outputs(5889) <= a or b;
    layer2_outputs(5890) <= not a;
    layer2_outputs(5891) <= a and b;
    layer2_outputs(5892) <= not a or b;
    layer2_outputs(5893) <= not (a xor b);
    layer2_outputs(5894) <= 1'b0;
    layer2_outputs(5895) <= not b;
    layer2_outputs(5896) <= not b or a;
    layer2_outputs(5897) <= a or b;
    layer2_outputs(5898) <= 1'b1;
    layer2_outputs(5899) <= b and not a;
    layer2_outputs(5900) <= a and not b;
    layer2_outputs(5901) <= a and not b;
    layer2_outputs(5902) <= not (a and b);
    layer2_outputs(5903) <= not a;
    layer2_outputs(5904) <= 1'b0;
    layer2_outputs(5905) <= a xor b;
    layer2_outputs(5906) <= not a;
    layer2_outputs(5907) <= a and b;
    layer2_outputs(5908) <= b;
    layer2_outputs(5909) <= a;
    layer2_outputs(5910) <= 1'b1;
    layer2_outputs(5911) <= not (a or b);
    layer2_outputs(5912) <= not (a and b);
    layer2_outputs(5913) <= 1'b1;
    layer2_outputs(5914) <= a xor b;
    layer2_outputs(5915) <= a;
    layer2_outputs(5916) <= not a or b;
    layer2_outputs(5917) <= a;
    layer2_outputs(5918) <= not b;
    layer2_outputs(5919) <= not b;
    layer2_outputs(5920) <= b;
    layer2_outputs(5921) <= not a;
    layer2_outputs(5922) <= 1'b1;
    layer2_outputs(5923) <= not (a or b);
    layer2_outputs(5924) <= a xor b;
    layer2_outputs(5925) <= not b or a;
    layer2_outputs(5926) <= a and b;
    layer2_outputs(5927) <= b and not a;
    layer2_outputs(5928) <= b and not a;
    layer2_outputs(5929) <= a and b;
    layer2_outputs(5930) <= not (a or b);
    layer2_outputs(5931) <= 1'b0;
    layer2_outputs(5932) <= a and not b;
    layer2_outputs(5933) <= not a;
    layer2_outputs(5934) <= b;
    layer2_outputs(5935) <= not a;
    layer2_outputs(5936) <= b;
    layer2_outputs(5937) <= not a;
    layer2_outputs(5938) <= b;
    layer2_outputs(5939) <= not b or a;
    layer2_outputs(5940) <= 1'b1;
    layer2_outputs(5941) <= not (a or b);
    layer2_outputs(5942) <= b and not a;
    layer2_outputs(5943) <= not (a or b);
    layer2_outputs(5944) <= b;
    layer2_outputs(5945) <= not (a and b);
    layer2_outputs(5946) <= not b or a;
    layer2_outputs(5947) <= 1'b0;
    layer2_outputs(5948) <= not (a or b);
    layer2_outputs(5949) <= not b or a;
    layer2_outputs(5950) <= a or b;
    layer2_outputs(5951) <= not a;
    layer2_outputs(5952) <= a and b;
    layer2_outputs(5953) <= a;
    layer2_outputs(5954) <= 1'b0;
    layer2_outputs(5955) <= b;
    layer2_outputs(5956) <= 1'b0;
    layer2_outputs(5957) <= not (a and b);
    layer2_outputs(5958) <= a or b;
    layer2_outputs(5959) <= a or b;
    layer2_outputs(5960) <= 1'b1;
    layer2_outputs(5961) <= not a or b;
    layer2_outputs(5962) <= not (a xor b);
    layer2_outputs(5963) <= 1'b1;
    layer2_outputs(5964) <= not (a and b);
    layer2_outputs(5965) <= not b;
    layer2_outputs(5966) <= not (a and b);
    layer2_outputs(5967) <= b and not a;
    layer2_outputs(5968) <= not (a and b);
    layer2_outputs(5969) <= not (a and b);
    layer2_outputs(5970) <= b and not a;
    layer2_outputs(5971) <= b and not a;
    layer2_outputs(5972) <= a or b;
    layer2_outputs(5973) <= 1'b0;
    layer2_outputs(5974) <= 1'b1;
    layer2_outputs(5975) <= b;
    layer2_outputs(5976) <= a xor b;
    layer2_outputs(5977) <= not b or a;
    layer2_outputs(5978) <= not (a and b);
    layer2_outputs(5979) <= a;
    layer2_outputs(5980) <= a or b;
    layer2_outputs(5981) <= a;
    layer2_outputs(5982) <= b and not a;
    layer2_outputs(5983) <= not b or a;
    layer2_outputs(5984) <= not (a xor b);
    layer2_outputs(5985) <= not (a or b);
    layer2_outputs(5986) <= not (a or b);
    layer2_outputs(5987) <= not a or b;
    layer2_outputs(5988) <= not b or a;
    layer2_outputs(5989) <= not a or b;
    layer2_outputs(5990) <= a and b;
    layer2_outputs(5991) <= not (a and b);
    layer2_outputs(5992) <= a and not b;
    layer2_outputs(5993) <= not b or a;
    layer2_outputs(5994) <= not b;
    layer2_outputs(5995) <= b and not a;
    layer2_outputs(5996) <= not a or b;
    layer2_outputs(5997) <= not a or b;
    layer2_outputs(5998) <= not (a and b);
    layer2_outputs(5999) <= not (a or b);
    layer2_outputs(6000) <= not b;
    layer2_outputs(6001) <= 1'b0;
    layer2_outputs(6002) <= not b;
    layer2_outputs(6003) <= not a or b;
    layer2_outputs(6004) <= not b;
    layer2_outputs(6005) <= not (a xor b);
    layer2_outputs(6006) <= a;
    layer2_outputs(6007) <= not (a and b);
    layer2_outputs(6008) <= a;
    layer2_outputs(6009) <= a or b;
    layer2_outputs(6010) <= a and not b;
    layer2_outputs(6011) <= b and not a;
    layer2_outputs(6012) <= a;
    layer2_outputs(6013) <= a and not b;
    layer2_outputs(6014) <= not a or b;
    layer2_outputs(6015) <= a;
    layer2_outputs(6016) <= b;
    layer2_outputs(6017) <= not a or b;
    layer2_outputs(6018) <= not b;
    layer2_outputs(6019) <= b and not a;
    layer2_outputs(6020) <= not a;
    layer2_outputs(6021) <= 1'b0;
    layer2_outputs(6022) <= 1'b0;
    layer2_outputs(6023) <= a or b;
    layer2_outputs(6024) <= not (a or b);
    layer2_outputs(6025) <= not (a or b);
    layer2_outputs(6026) <= not (a and b);
    layer2_outputs(6027) <= not b or a;
    layer2_outputs(6028) <= b and not a;
    layer2_outputs(6029) <= not (a or b);
    layer2_outputs(6030) <= b;
    layer2_outputs(6031) <= a and b;
    layer2_outputs(6032) <= a;
    layer2_outputs(6033) <= not (a or b);
    layer2_outputs(6034) <= not b or a;
    layer2_outputs(6035) <= 1'b1;
    layer2_outputs(6036) <= 1'b0;
    layer2_outputs(6037) <= not (a and b);
    layer2_outputs(6038) <= 1'b0;
    layer2_outputs(6039) <= a or b;
    layer2_outputs(6040) <= a xor b;
    layer2_outputs(6041) <= not b or a;
    layer2_outputs(6042) <= not b or a;
    layer2_outputs(6043) <= not (a or b);
    layer2_outputs(6044) <= not (a xor b);
    layer2_outputs(6045) <= 1'b1;
    layer2_outputs(6046) <= a and not b;
    layer2_outputs(6047) <= not a or b;
    layer2_outputs(6048) <= not a;
    layer2_outputs(6049) <= not a;
    layer2_outputs(6050) <= not (a or b);
    layer2_outputs(6051) <= b and not a;
    layer2_outputs(6052) <= b;
    layer2_outputs(6053) <= 1'b1;
    layer2_outputs(6054) <= not (a or b);
    layer2_outputs(6055) <= b;
    layer2_outputs(6056) <= 1'b0;
    layer2_outputs(6057) <= a or b;
    layer2_outputs(6058) <= 1'b0;
    layer2_outputs(6059) <= not b or a;
    layer2_outputs(6060) <= not a;
    layer2_outputs(6061) <= 1'b1;
    layer2_outputs(6062) <= a and not b;
    layer2_outputs(6063) <= not (a or b);
    layer2_outputs(6064) <= a;
    layer2_outputs(6065) <= a;
    layer2_outputs(6066) <= a or b;
    layer2_outputs(6067) <= not a or b;
    layer2_outputs(6068) <= not a;
    layer2_outputs(6069) <= not b or a;
    layer2_outputs(6070) <= b;
    layer2_outputs(6071) <= 1'b0;
    layer2_outputs(6072) <= a and b;
    layer2_outputs(6073) <= 1'b1;
    layer2_outputs(6074) <= not (a xor b);
    layer2_outputs(6075) <= a or b;
    layer2_outputs(6076) <= 1'b1;
    layer2_outputs(6077) <= not (a and b);
    layer2_outputs(6078) <= 1'b0;
    layer2_outputs(6079) <= not b or a;
    layer2_outputs(6080) <= not b or a;
    layer2_outputs(6081) <= not (a and b);
    layer2_outputs(6082) <= b;
    layer2_outputs(6083) <= not b;
    layer2_outputs(6084) <= not b or a;
    layer2_outputs(6085) <= not b;
    layer2_outputs(6086) <= a and not b;
    layer2_outputs(6087) <= a or b;
    layer2_outputs(6088) <= not b;
    layer2_outputs(6089) <= a and not b;
    layer2_outputs(6090) <= not (a xor b);
    layer2_outputs(6091) <= a and not b;
    layer2_outputs(6092) <= a;
    layer2_outputs(6093) <= not (a and b);
    layer2_outputs(6094) <= not (a or b);
    layer2_outputs(6095) <= not a or b;
    layer2_outputs(6096) <= a or b;
    layer2_outputs(6097) <= a;
    layer2_outputs(6098) <= a and not b;
    layer2_outputs(6099) <= a and b;
    layer2_outputs(6100) <= 1'b0;
    layer2_outputs(6101) <= not (a or b);
    layer2_outputs(6102) <= a and not b;
    layer2_outputs(6103) <= not a;
    layer2_outputs(6104) <= a;
    layer2_outputs(6105) <= 1'b0;
    layer2_outputs(6106) <= not (a or b);
    layer2_outputs(6107) <= b;
    layer2_outputs(6108) <= not b or a;
    layer2_outputs(6109) <= 1'b0;
    layer2_outputs(6110) <= 1'b0;
    layer2_outputs(6111) <= 1'b1;
    layer2_outputs(6112) <= not a or b;
    layer2_outputs(6113) <= a or b;
    layer2_outputs(6114) <= 1'b1;
    layer2_outputs(6115) <= not b;
    layer2_outputs(6116) <= a or b;
    layer2_outputs(6117) <= not (a or b);
    layer2_outputs(6118) <= b;
    layer2_outputs(6119) <= not b or a;
    layer2_outputs(6120) <= not a;
    layer2_outputs(6121) <= b;
    layer2_outputs(6122) <= a and b;
    layer2_outputs(6123) <= a and b;
    layer2_outputs(6124) <= a;
    layer2_outputs(6125) <= not (a or b);
    layer2_outputs(6126) <= 1'b1;
    layer2_outputs(6127) <= not (a and b);
    layer2_outputs(6128) <= b;
    layer2_outputs(6129) <= a;
    layer2_outputs(6130) <= a or b;
    layer2_outputs(6131) <= not (a and b);
    layer2_outputs(6132) <= not b or a;
    layer2_outputs(6133) <= not (a or b);
    layer2_outputs(6134) <= 1'b0;
    layer2_outputs(6135) <= not b;
    layer2_outputs(6136) <= not b or a;
    layer2_outputs(6137) <= not (a or b);
    layer2_outputs(6138) <= 1'b1;
    layer2_outputs(6139) <= 1'b1;
    layer2_outputs(6140) <= not b;
    layer2_outputs(6141) <= not a;
    layer2_outputs(6142) <= not a;
    layer2_outputs(6143) <= not b;
    layer2_outputs(6144) <= a and b;
    layer2_outputs(6145) <= a;
    layer2_outputs(6146) <= 1'b0;
    layer2_outputs(6147) <= not b or a;
    layer2_outputs(6148) <= not b;
    layer2_outputs(6149) <= not (a and b);
    layer2_outputs(6150) <= a and not b;
    layer2_outputs(6151) <= a or b;
    layer2_outputs(6152) <= 1'b0;
    layer2_outputs(6153) <= not b;
    layer2_outputs(6154) <= a or b;
    layer2_outputs(6155) <= a and not b;
    layer2_outputs(6156) <= not b or a;
    layer2_outputs(6157) <= b and not a;
    layer2_outputs(6158) <= 1'b0;
    layer2_outputs(6159) <= not (a xor b);
    layer2_outputs(6160) <= 1'b0;
    layer2_outputs(6161) <= not b;
    layer2_outputs(6162) <= not b;
    layer2_outputs(6163) <= a and b;
    layer2_outputs(6164) <= a or b;
    layer2_outputs(6165) <= not a or b;
    layer2_outputs(6166) <= a;
    layer2_outputs(6167) <= not a;
    layer2_outputs(6168) <= not (a or b);
    layer2_outputs(6169) <= a and b;
    layer2_outputs(6170) <= a;
    layer2_outputs(6171) <= a;
    layer2_outputs(6172) <= not (a and b);
    layer2_outputs(6173) <= not a;
    layer2_outputs(6174) <= a xor b;
    layer2_outputs(6175) <= a and not b;
    layer2_outputs(6176) <= not (a and b);
    layer2_outputs(6177) <= a;
    layer2_outputs(6178) <= 1'b1;
    layer2_outputs(6179) <= a or b;
    layer2_outputs(6180) <= not (a and b);
    layer2_outputs(6181) <= not a or b;
    layer2_outputs(6182) <= a and b;
    layer2_outputs(6183) <= 1'b0;
    layer2_outputs(6184) <= b and not a;
    layer2_outputs(6185) <= 1'b0;
    layer2_outputs(6186) <= a;
    layer2_outputs(6187) <= 1'b1;
    layer2_outputs(6188) <= a xor b;
    layer2_outputs(6189) <= a xor b;
    layer2_outputs(6190) <= b;
    layer2_outputs(6191) <= a;
    layer2_outputs(6192) <= b;
    layer2_outputs(6193) <= not (a or b);
    layer2_outputs(6194) <= not b;
    layer2_outputs(6195) <= a;
    layer2_outputs(6196) <= b and not a;
    layer2_outputs(6197) <= not a;
    layer2_outputs(6198) <= a and b;
    layer2_outputs(6199) <= not b or a;
    layer2_outputs(6200) <= not b;
    layer2_outputs(6201) <= a and b;
    layer2_outputs(6202) <= not b or a;
    layer2_outputs(6203) <= a and not b;
    layer2_outputs(6204) <= 1'b1;
    layer2_outputs(6205) <= not a;
    layer2_outputs(6206) <= a;
    layer2_outputs(6207) <= b and not a;
    layer2_outputs(6208) <= not b;
    layer2_outputs(6209) <= 1'b0;
    layer2_outputs(6210) <= b;
    layer2_outputs(6211) <= not b or a;
    layer2_outputs(6212) <= not b or a;
    layer2_outputs(6213) <= a;
    layer2_outputs(6214) <= not b;
    layer2_outputs(6215) <= not b;
    layer2_outputs(6216) <= a and b;
    layer2_outputs(6217) <= not (a and b);
    layer2_outputs(6218) <= not a or b;
    layer2_outputs(6219) <= not (a and b);
    layer2_outputs(6220) <= b and not a;
    layer2_outputs(6221) <= not a;
    layer2_outputs(6222) <= 1'b1;
    layer2_outputs(6223) <= b and not a;
    layer2_outputs(6224) <= not (a and b);
    layer2_outputs(6225) <= 1'b0;
    layer2_outputs(6226) <= a and b;
    layer2_outputs(6227) <= not a or b;
    layer2_outputs(6228) <= b;
    layer2_outputs(6229) <= 1'b1;
    layer2_outputs(6230) <= b;
    layer2_outputs(6231) <= not (a or b);
    layer2_outputs(6232) <= 1'b0;
    layer2_outputs(6233) <= not b or a;
    layer2_outputs(6234) <= not (a or b);
    layer2_outputs(6235) <= a xor b;
    layer2_outputs(6236) <= not b;
    layer2_outputs(6237) <= b and not a;
    layer2_outputs(6238) <= a or b;
    layer2_outputs(6239) <= not (a and b);
    layer2_outputs(6240) <= not a;
    layer2_outputs(6241) <= b and not a;
    layer2_outputs(6242) <= a and b;
    layer2_outputs(6243) <= not (a and b);
    layer2_outputs(6244) <= 1'b1;
    layer2_outputs(6245) <= a;
    layer2_outputs(6246) <= b;
    layer2_outputs(6247) <= not b or a;
    layer2_outputs(6248) <= a;
    layer2_outputs(6249) <= b;
    layer2_outputs(6250) <= a or b;
    layer2_outputs(6251) <= a and b;
    layer2_outputs(6252) <= not (a or b);
    layer2_outputs(6253) <= b;
    layer2_outputs(6254) <= not b;
    layer2_outputs(6255) <= 1'b0;
    layer2_outputs(6256) <= not (a or b);
    layer2_outputs(6257) <= 1'b1;
    layer2_outputs(6258) <= not (a or b);
    layer2_outputs(6259) <= not a;
    layer2_outputs(6260) <= 1'b0;
    layer2_outputs(6261) <= not a or b;
    layer2_outputs(6262) <= a;
    layer2_outputs(6263) <= 1'b1;
    layer2_outputs(6264) <= 1'b0;
    layer2_outputs(6265) <= b;
    layer2_outputs(6266) <= a;
    layer2_outputs(6267) <= b;
    layer2_outputs(6268) <= not (a or b);
    layer2_outputs(6269) <= b and not a;
    layer2_outputs(6270) <= a or b;
    layer2_outputs(6271) <= b and not a;
    layer2_outputs(6272) <= b;
    layer2_outputs(6273) <= a;
    layer2_outputs(6274) <= not a;
    layer2_outputs(6275) <= a and b;
    layer2_outputs(6276) <= 1'b0;
    layer2_outputs(6277) <= a and b;
    layer2_outputs(6278) <= not (a and b);
    layer2_outputs(6279) <= a or b;
    layer2_outputs(6280) <= a and b;
    layer2_outputs(6281) <= not b or a;
    layer2_outputs(6282) <= a xor b;
    layer2_outputs(6283) <= not a;
    layer2_outputs(6284) <= b and not a;
    layer2_outputs(6285) <= not (a and b);
    layer2_outputs(6286) <= a and not b;
    layer2_outputs(6287) <= not b;
    layer2_outputs(6288) <= a or b;
    layer2_outputs(6289) <= not a or b;
    layer2_outputs(6290) <= 1'b1;
    layer2_outputs(6291) <= not b or a;
    layer2_outputs(6292) <= b;
    layer2_outputs(6293) <= not b;
    layer2_outputs(6294) <= 1'b0;
    layer2_outputs(6295) <= a;
    layer2_outputs(6296) <= b;
    layer2_outputs(6297) <= a or b;
    layer2_outputs(6298) <= not (a or b);
    layer2_outputs(6299) <= not a or b;
    layer2_outputs(6300) <= not (a xor b);
    layer2_outputs(6301) <= a;
    layer2_outputs(6302) <= 1'b0;
    layer2_outputs(6303) <= 1'b0;
    layer2_outputs(6304) <= not (a or b);
    layer2_outputs(6305) <= a and b;
    layer2_outputs(6306) <= 1'b1;
    layer2_outputs(6307) <= not (a or b);
    layer2_outputs(6308) <= b;
    layer2_outputs(6309) <= not a;
    layer2_outputs(6310) <= a and not b;
    layer2_outputs(6311) <= not a;
    layer2_outputs(6312) <= 1'b0;
    layer2_outputs(6313) <= 1'b1;
    layer2_outputs(6314) <= not (a and b);
    layer2_outputs(6315) <= a and b;
    layer2_outputs(6316) <= not a or b;
    layer2_outputs(6317) <= 1'b0;
    layer2_outputs(6318) <= not (a or b);
    layer2_outputs(6319) <= not (a and b);
    layer2_outputs(6320) <= a and b;
    layer2_outputs(6321) <= a and b;
    layer2_outputs(6322) <= not (a or b);
    layer2_outputs(6323) <= a and not b;
    layer2_outputs(6324) <= not a;
    layer2_outputs(6325) <= not b or a;
    layer2_outputs(6326) <= not (a xor b);
    layer2_outputs(6327) <= 1'b0;
    layer2_outputs(6328) <= 1'b1;
    layer2_outputs(6329) <= a and b;
    layer2_outputs(6330) <= 1'b1;
    layer2_outputs(6331) <= a;
    layer2_outputs(6332) <= not b;
    layer2_outputs(6333) <= not (a xor b);
    layer2_outputs(6334) <= b;
    layer2_outputs(6335) <= a;
    layer2_outputs(6336) <= b and not a;
    layer2_outputs(6337) <= a and b;
    layer2_outputs(6338) <= a;
    layer2_outputs(6339) <= a or b;
    layer2_outputs(6340) <= a or b;
    layer2_outputs(6341) <= not (a and b);
    layer2_outputs(6342) <= a and b;
    layer2_outputs(6343) <= a and not b;
    layer2_outputs(6344) <= b;
    layer2_outputs(6345) <= not a or b;
    layer2_outputs(6346) <= not (a and b);
    layer2_outputs(6347) <= not (a or b);
    layer2_outputs(6348) <= 1'b0;
    layer2_outputs(6349) <= a and b;
    layer2_outputs(6350) <= not b or a;
    layer2_outputs(6351) <= a or b;
    layer2_outputs(6352) <= a;
    layer2_outputs(6353) <= not a;
    layer2_outputs(6354) <= not a;
    layer2_outputs(6355) <= a;
    layer2_outputs(6356) <= not b or a;
    layer2_outputs(6357) <= a;
    layer2_outputs(6358) <= b;
    layer2_outputs(6359) <= b and not a;
    layer2_outputs(6360) <= 1'b1;
    layer2_outputs(6361) <= not b or a;
    layer2_outputs(6362) <= 1'b1;
    layer2_outputs(6363) <= not (a and b);
    layer2_outputs(6364) <= 1'b1;
    layer2_outputs(6365) <= a and b;
    layer2_outputs(6366) <= 1'b0;
    layer2_outputs(6367) <= a and b;
    layer2_outputs(6368) <= a and b;
    layer2_outputs(6369) <= not b or a;
    layer2_outputs(6370) <= not (a and b);
    layer2_outputs(6371) <= not (a or b);
    layer2_outputs(6372) <= not b or a;
    layer2_outputs(6373) <= not b or a;
    layer2_outputs(6374) <= a and b;
    layer2_outputs(6375) <= b and not a;
    layer2_outputs(6376) <= not b;
    layer2_outputs(6377) <= a and not b;
    layer2_outputs(6378) <= b and not a;
    layer2_outputs(6379) <= not (a or b);
    layer2_outputs(6380) <= a and not b;
    layer2_outputs(6381) <= 1'b1;
    layer2_outputs(6382) <= not (a and b);
    layer2_outputs(6383) <= not a or b;
    layer2_outputs(6384) <= not (a and b);
    layer2_outputs(6385) <= a and not b;
    layer2_outputs(6386) <= a and b;
    layer2_outputs(6387) <= a or b;
    layer2_outputs(6388) <= 1'b1;
    layer2_outputs(6389) <= b and not a;
    layer2_outputs(6390) <= a xor b;
    layer2_outputs(6391) <= not (a or b);
    layer2_outputs(6392) <= not (a and b);
    layer2_outputs(6393) <= 1'b1;
    layer2_outputs(6394) <= a and not b;
    layer2_outputs(6395) <= 1'b1;
    layer2_outputs(6396) <= not (a or b);
    layer2_outputs(6397) <= not (a or b);
    layer2_outputs(6398) <= b and not a;
    layer2_outputs(6399) <= a;
    layer2_outputs(6400) <= 1'b0;
    layer2_outputs(6401) <= not (a and b);
    layer2_outputs(6402) <= not a or b;
    layer2_outputs(6403) <= not b or a;
    layer2_outputs(6404) <= 1'b1;
    layer2_outputs(6405) <= not a;
    layer2_outputs(6406) <= not a or b;
    layer2_outputs(6407) <= not a;
    layer2_outputs(6408) <= a and b;
    layer2_outputs(6409) <= a or b;
    layer2_outputs(6410) <= b;
    layer2_outputs(6411) <= not b or a;
    layer2_outputs(6412) <= 1'b0;
    layer2_outputs(6413) <= 1'b1;
    layer2_outputs(6414) <= a;
    layer2_outputs(6415) <= not (a or b);
    layer2_outputs(6416) <= a or b;
    layer2_outputs(6417) <= not (a xor b);
    layer2_outputs(6418) <= a;
    layer2_outputs(6419) <= not (a and b);
    layer2_outputs(6420) <= a or b;
    layer2_outputs(6421) <= not b;
    layer2_outputs(6422) <= b;
    layer2_outputs(6423) <= b and not a;
    layer2_outputs(6424) <= a and not b;
    layer2_outputs(6425) <= a or b;
    layer2_outputs(6426) <= a or b;
    layer2_outputs(6427) <= not b;
    layer2_outputs(6428) <= not b or a;
    layer2_outputs(6429) <= 1'b1;
    layer2_outputs(6430) <= 1'b0;
    layer2_outputs(6431) <= not a;
    layer2_outputs(6432) <= 1'b0;
    layer2_outputs(6433) <= not (a and b);
    layer2_outputs(6434) <= b;
    layer2_outputs(6435) <= not b or a;
    layer2_outputs(6436) <= 1'b0;
    layer2_outputs(6437) <= not a or b;
    layer2_outputs(6438) <= b and not a;
    layer2_outputs(6439) <= not (a or b);
    layer2_outputs(6440) <= not (a and b);
    layer2_outputs(6441) <= a and b;
    layer2_outputs(6442) <= a and not b;
    layer2_outputs(6443) <= not (a and b);
    layer2_outputs(6444) <= not a;
    layer2_outputs(6445) <= not (a and b);
    layer2_outputs(6446) <= not a or b;
    layer2_outputs(6447) <= 1'b1;
    layer2_outputs(6448) <= a and not b;
    layer2_outputs(6449) <= not (a and b);
    layer2_outputs(6450) <= b;
    layer2_outputs(6451) <= a or b;
    layer2_outputs(6452) <= a xor b;
    layer2_outputs(6453) <= b and not a;
    layer2_outputs(6454) <= not b;
    layer2_outputs(6455) <= a xor b;
    layer2_outputs(6456) <= 1'b1;
    layer2_outputs(6457) <= a and b;
    layer2_outputs(6458) <= not a or b;
    layer2_outputs(6459) <= b and not a;
    layer2_outputs(6460) <= b and not a;
    layer2_outputs(6461) <= a;
    layer2_outputs(6462) <= not b;
    layer2_outputs(6463) <= a and not b;
    layer2_outputs(6464) <= 1'b1;
    layer2_outputs(6465) <= not (a and b);
    layer2_outputs(6466) <= not (a and b);
    layer2_outputs(6467) <= a and b;
    layer2_outputs(6468) <= a and b;
    layer2_outputs(6469) <= not (a and b);
    layer2_outputs(6470) <= a and b;
    layer2_outputs(6471) <= 1'b1;
    layer2_outputs(6472) <= a or b;
    layer2_outputs(6473) <= not a or b;
    layer2_outputs(6474) <= not (a or b);
    layer2_outputs(6475) <= 1'b0;
    layer2_outputs(6476) <= not (a and b);
    layer2_outputs(6477) <= not (a and b);
    layer2_outputs(6478) <= b;
    layer2_outputs(6479) <= a;
    layer2_outputs(6480) <= 1'b0;
    layer2_outputs(6481) <= not a;
    layer2_outputs(6482) <= a or b;
    layer2_outputs(6483) <= a and b;
    layer2_outputs(6484) <= a;
    layer2_outputs(6485) <= not (a and b);
    layer2_outputs(6486) <= 1'b1;
    layer2_outputs(6487) <= not b or a;
    layer2_outputs(6488) <= not a or b;
    layer2_outputs(6489) <= a or b;
    layer2_outputs(6490) <= b and not a;
    layer2_outputs(6491) <= 1'b1;
    layer2_outputs(6492) <= not a or b;
    layer2_outputs(6493) <= not a;
    layer2_outputs(6494) <= 1'b1;
    layer2_outputs(6495) <= not (a xor b);
    layer2_outputs(6496) <= b and not a;
    layer2_outputs(6497) <= not b;
    layer2_outputs(6498) <= a or b;
    layer2_outputs(6499) <= 1'b1;
    layer2_outputs(6500) <= not a;
    layer2_outputs(6501) <= b and not a;
    layer2_outputs(6502) <= not (a xor b);
    layer2_outputs(6503) <= 1'b1;
    layer2_outputs(6504) <= b and not a;
    layer2_outputs(6505) <= not (a or b);
    layer2_outputs(6506) <= not (a xor b);
    layer2_outputs(6507) <= 1'b1;
    layer2_outputs(6508) <= not a or b;
    layer2_outputs(6509) <= 1'b0;
    layer2_outputs(6510) <= not b or a;
    layer2_outputs(6511) <= a and not b;
    layer2_outputs(6512) <= not b or a;
    layer2_outputs(6513) <= a;
    layer2_outputs(6514) <= b and not a;
    layer2_outputs(6515) <= not a;
    layer2_outputs(6516) <= b;
    layer2_outputs(6517) <= not a;
    layer2_outputs(6518) <= 1'b1;
    layer2_outputs(6519) <= not (a and b);
    layer2_outputs(6520) <= a and b;
    layer2_outputs(6521) <= b;
    layer2_outputs(6522) <= not a;
    layer2_outputs(6523) <= not (a or b);
    layer2_outputs(6524) <= not (a and b);
    layer2_outputs(6525) <= a and not b;
    layer2_outputs(6526) <= not (a xor b);
    layer2_outputs(6527) <= 1'b0;
    layer2_outputs(6528) <= not b or a;
    layer2_outputs(6529) <= 1'b1;
    layer2_outputs(6530) <= not (a xor b);
    layer2_outputs(6531) <= a;
    layer2_outputs(6532) <= b and not a;
    layer2_outputs(6533) <= a and not b;
    layer2_outputs(6534) <= not a;
    layer2_outputs(6535) <= a;
    layer2_outputs(6536) <= b;
    layer2_outputs(6537) <= b;
    layer2_outputs(6538) <= not (a and b);
    layer2_outputs(6539) <= a and b;
    layer2_outputs(6540) <= a and b;
    layer2_outputs(6541) <= not (a and b);
    layer2_outputs(6542) <= not (a or b);
    layer2_outputs(6543) <= b;
    layer2_outputs(6544) <= b and not a;
    layer2_outputs(6545) <= a and b;
    layer2_outputs(6546) <= not a;
    layer2_outputs(6547) <= not a;
    layer2_outputs(6548) <= b;
    layer2_outputs(6549) <= a or b;
    layer2_outputs(6550) <= 1'b0;
    layer2_outputs(6551) <= a and not b;
    layer2_outputs(6552) <= b and not a;
    layer2_outputs(6553) <= a;
    layer2_outputs(6554) <= 1'b0;
    layer2_outputs(6555) <= not b or a;
    layer2_outputs(6556) <= a and not b;
    layer2_outputs(6557) <= not a;
    layer2_outputs(6558) <= 1'b0;
    layer2_outputs(6559) <= not a or b;
    layer2_outputs(6560) <= a and not b;
    layer2_outputs(6561) <= not b or a;
    layer2_outputs(6562) <= a or b;
    layer2_outputs(6563) <= a or b;
    layer2_outputs(6564) <= not a;
    layer2_outputs(6565) <= a;
    layer2_outputs(6566) <= a;
    layer2_outputs(6567) <= b and not a;
    layer2_outputs(6568) <= b and not a;
    layer2_outputs(6569) <= b and not a;
    layer2_outputs(6570) <= b and not a;
    layer2_outputs(6571) <= not (a or b);
    layer2_outputs(6572) <= a;
    layer2_outputs(6573) <= 1'b0;
    layer2_outputs(6574) <= not a or b;
    layer2_outputs(6575) <= not a or b;
    layer2_outputs(6576) <= b;
    layer2_outputs(6577) <= a and not b;
    layer2_outputs(6578) <= a or b;
    layer2_outputs(6579) <= 1'b0;
    layer2_outputs(6580) <= not a or b;
    layer2_outputs(6581) <= a or b;
    layer2_outputs(6582) <= 1'b1;
    layer2_outputs(6583) <= a and not b;
    layer2_outputs(6584) <= not (a and b);
    layer2_outputs(6585) <= not (a or b);
    layer2_outputs(6586) <= a or b;
    layer2_outputs(6587) <= 1'b1;
    layer2_outputs(6588) <= not b or a;
    layer2_outputs(6589) <= not (a or b);
    layer2_outputs(6590) <= a and b;
    layer2_outputs(6591) <= not (a and b);
    layer2_outputs(6592) <= 1'b1;
    layer2_outputs(6593) <= b;
    layer2_outputs(6594) <= a;
    layer2_outputs(6595) <= 1'b1;
    layer2_outputs(6596) <= not a or b;
    layer2_outputs(6597) <= 1'b0;
    layer2_outputs(6598) <= 1'b1;
    layer2_outputs(6599) <= not a;
    layer2_outputs(6600) <= not b;
    layer2_outputs(6601) <= not (a and b);
    layer2_outputs(6602) <= not (a and b);
    layer2_outputs(6603) <= b and not a;
    layer2_outputs(6604) <= not (a xor b);
    layer2_outputs(6605) <= not b;
    layer2_outputs(6606) <= 1'b0;
    layer2_outputs(6607) <= 1'b1;
    layer2_outputs(6608) <= a and not b;
    layer2_outputs(6609) <= not b or a;
    layer2_outputs(6610) <= not b;
    layer2_outputs(6611) <= 1'b0;
    layer2_outputs(6612) <= a or b;
    layer2_outputs(6613) <= a and not b;
    layer2_outputs(6614) <= not a;
    layer2_outputs(6615) <= not (a or b);
    layer2_outputs(6616) <= not (a and b);
    layer2_outputs(6617) <= a and b;
    layer2_outputs(6618) <= not a;
    layer2_outputs(6619) <= a and b;
    layer2_outputs(6620) <= 1'b1;
    layer2_outputs(6621) <= b and not a;
    layer2_outputs(6622) <= a or b;
    layer2_outputs(6623) <= not (a xor b);
    layer2_outputs(6624) <= b;
    layer2_outputs(6625) <= not (a and b);
    layer2_outputs(6626) <= a or b;
    layer2_outputs(6627) <= a and b;
    layer2_outputs(6628) <= a and not b;
    layer2_outputs(6629) <= 1'b0;
    layer2_outputs(6630) <= a or b;
    layer2_outputs(6631) <= a;
    layer2_outputs(6632) <= 1'b0;
    layer2_outputs(6633) <= a and b;
    layer2_outputs(6634) <= 1'b1;
    layer2_outputs(6635) <= not a;
    layer2_outputs(6636) <= not b;
    layer2_outputs(6637) <= not b or a;
    layer2_outputs(6638) <= b and not a;
    layer2_outputs(6639) <= a and b;
    layer2_outputs(6640) <= 1'b0;
    layer2_outputs(6641) <= a and b;
    layer2_outputs(6642) <= b and not a;
    layer2_outputs(6643) <= a;
    layer2_outputs(6644) <= a and b;
    layer2_outputs(6645) <= not (a or b);
    layer2_outputs(6646) <= 1'b1;
    layer2_outputs(6647) <= not (a and b);
    layer2_outputs(6648) <= not (a or b);
    layer2_outputs(6649) <= 1'b1;
    layer2_outputs(6650) <= not (a and b);
    layer2_outputs(6651) <= a and not b;
    layer2_outputs(6652) <= a or b;
    layer2_outputs(6653) <= b and not a;
    layer2_outputs(6654) <= a;
    layer2_outputs(6655) <= not a;
    layer2_outputs(6656) <= a or b;
    layer2_outputs(6657) <= a;
    layer2_outputs(6658) <= b and not a;
    layer2_outputs(6659) <= not b;
    layer2_outputs(6660) <= not b;
    layer2_outputs(6661) <= 1'b0;
    layer2_outputs(6662) <= not b or a;
    layer2_outputs(6663) <= not b or a;
    layer2_outputs(6664) <= not b;
    layer2_outputs(6665) <= not a;
    layer2_outputs(6666) <= not b or a;
    layer2_outputs(6667) <= not b;
    layer2_outputs(6668) <= a and b;
    layer2_outputs(6669) <= a and b;
    layer2_outputs(6670) <= a and not b;
    layer2_outputs(6671) <= 1'b0;
    layer2_outputs(6672) <= b and not a;
    layer2_outputs(6673) <= not a or b;
    layer2_outputs(6674) <= 1'b0;
    layer2_outputs(6675) <= 1'b0;
    layer2_outputs(6676) <= 1'b1;
    layer2_outputs(6677) <= 1'b1;
    layer2_outputs(6678) <= a;
    layer2_outputs(6679) <= 1'b0;
    layer2_outputs(6680) <= 1'b1;
    layer2_outputs(6681) <= not a or b;
    layer2_outputs(6682) <= not a or b;
    layer2_outputs(6683) <= a;
    layer2_outputs(6684) <= a and not b;
    layer2_outputs(6685) <= a or b;
    layer2_outputs(6686) <= not b or a;
    layer2_outputs(6687) <= 1'b1;
    layer2_outputs(6688) <= a and b;
    layer2_outputs(6689) <= 1'b0;
    layer2_outputs(6690) <= not b;
    layer2_outputs(6691) <= b and not a;
    layer2_outputs(6692) <= a and b;
    layer2_outputs(6693) <= not (a and b);
    layer2_outputs(6694) <= b;
    layer2_outputs(6695) <= b and not a;
    layer2_outputs(6696) <= b and not a;
    layer2_outputs(6697) <= not a or b;
    layer2_outputs(6698) <= a and not b;
    layer2_outputs(6699) <= a and not b;
    layer2_outputs(6700) <= not a or b;
    layer2_outputs(6701) <= 1'b1;
    layer2_outputs(6702) <= not (a and b);
    layer2_outputs(6703) <= b and not a;
    layer2_outputs(6704) <= b;
    layer2_outputs(6705) <= b and not a;
    layer2_outputs(6706) <= b and not a;
    layer2_outputs(6707) <= 1'b0;
    layer2_outputs(6708) <= 1'b0;
    layer2_outputs(6709) <= not b;
    layer2_outputs(6710) <= 1'b0;
    layer2_outputs(6711) <= not (a or b);
    layer2_outputs(6712) <= not b;
    layer2_outputs(6713) <= a and b;
    layer2_outputs(6714) <= not a;
    layer2_outputs(6715) <= not b or a;
    layer2_outputs(6716) <= 1'b1;
    layer2_outputs(6717) <= 1'b1;
    layer2_outputs(6718) <= 1'b0;
    layer2_outputs(6719) <= a and not b;
    layer2_outputs(6720) <= not a;
    layer2_outputs(6721) <= not a or b;
    layer2_outputs(6722) <= 1'b0;
    layer2_outputs(6723) <= not a;
    layer2_outputs(6724) <= not (a or b);
    layer2_outputs(6725) <= 1'b0;
    layer2_outputs(6726) <= not b;
    layer2_outputs(6727) <= b and not a;
    layer2_outputs(6728) <= not a or b;
    layer2_outputs(6729) <= not b or a;
    layer2_outputs(6730) <= a;
    layer2_outputs(6731) <= b and not a;
    layer2_outputs(6732) <= 1'b0;
    layer2_outputs(6733) <= a or b;
    layer2_outputs(6734) <= not a or b;
    layer2_outputs(6735) <= b;
    layer2_outputs(6736) <= a and b;
    layer2_outputs(6737) <= not a;
    layer2_outputs(6738) <= not b;
    layer2_outputs(6739) <= not b or a;
    layer2_outputs(6740) <= a or b;
    layer2_outputs(6741) <= not (a or b);
    layer2_outputs(6742) <= not (a and b);
    layer2_outputs(6743) <= a;
    layer2_outputs(6744) <= a or b;
    layer2_outputs(6745) <= a and b;
    layer2_outputs(6746) <= 1'b1;
    layer2_outputs(6747) <= a or b;
    layer2_outputs(6748) <= not b or a;
    layer2_outputs(6749) <= not a or b;
    layer2_outputs(6750) <= not (a or b);
    layer2_outputs(6751) <= a or b;
    layer2_outputs(6752) <= not a or b;
    layer2_outputs(6753) <= 1'b1;
    layer2_outputs(6754) <= not b or a;
    layer2_outputs(6755) <= not b or a;
    layer2_outputs(6756) <= a xor b;
    layer2_outputs(6757) <= not b;
    layer2_outputs(6758) <= not (a xor b);
    layer2_outputs(6759) <= a and not b;
    layer2_outputs(6760) <= not a or b;
    layer2_outputs(6761) <= 1'b1;
    layer2_outputs(6762) <= a;
    layer2_outputs(6763) <= a and not b;
    layer2_outputs(6764) <= 1'b1;
    layer2_outputs(6765) <= 1'b1;
    layer2_outputs(6766) <= a or b;
    layer2_outputs(6767) <= 1'b0;
    layer2_outputs(6768) <= not (a and b);
    layer2_outputs(6769) <= 1'b1;
    layer2_outputs(6770) <= a and b;
    layer2_outputs(6771) <= a or b;
    layer2_outputs(6772) <= a;
    layer2_outputs(6773) <= not (a or b);
    layer2_outputs(6774) <= a or b;
    layer2_outputs(6775) <= not b or a;
    layer2_outputs(6776) <= not (a and b);
    layer2_outputs(6777) <= 1'b0;
    layer2_outputs(6778) <= not a;
    layer2_outputs(6779) <= 1'b1;
    layer2_outputs(6780) <= not (a and b);
    layer2_outputs(6781) <= b and not a;
    layer2_outputs(6782) <= b and not a;
    layer2_outputs(6783) <= not b or a;
    layer2_outputs(6784) <= not b or a;
    layer2_outputs(6785) <= a xor b;
    layer2_outputs(6786) <= not a or b;
    layer2_outputs(6787) <= not b or a;
    layer2_outputs(6788) <= not (a and b);
    layer2_outputs(6789) <= not a;
    layer2_outputs(6790) <= a or b;
    layer2_outputs(6791) <= a and b;
    layer2_outputs(6792) <= a or b;
    layer2_outputs(6793) <= not a;
    layer2_outputs(6794) <= 1'b0;
    layer2_outputs(6795) <= not (a and b);
    layer2_outputs(6796) <= 1'b1;
    layer2_outputs(6797) <= a and b;
    layer2_outputs(6798) <= 1'b0;
    layer2_outputs(6799) <= 1'b1;
    layer2_outputs(6800) <= 1'b1;
    layer2_outputs(6801) <= a and not b;
    layer2_outputs(6802) <= a or b;
    layer2_outputs(6803) <= a and b;
    layer2_outputs(6804) <= not b;
    layer2_outputs(6805) <= b and not a;
    layer2_outputs(6806) <= b;
    layer2_outputs(6807) <= not (a xor b);
    layer2_outputs(6808) <= not (a or b);
    layer2_outputs(6809) <= not (a xor b);
    layer2_outputs(6810) <= 1'b0;
    layer2_outputs(6811) <= not (a and b);
    layer2_outputs(6812) <= a and b;
    layer2_outputs(6813) <= 1'b1;
    layer2_outputs(6814) <= 1'b1;
    layer2_outputs(6815) <= a and b;
    layer2_outputs(6816) <= not b;
    layer2_outputs(6817) <= a;
    layer2_outputs(6818) <= 1'b0;
    layer2_outputs(6819) <= not a;
    layer2_outputs(6820) <= not b or a;
    layer2_outputs(6821) <= 1'b1;
    layer2_outputs(6822) <= not b;
    layer2_outputs(6823) <= not (a and b);
    layer2_outputs(6824) <= 1'b0;
    layer2_outputs(6825) <= b;
    layer2_outputs(6826) <= not b or a;
    layer2_outputs(6827) <= not b;
    layer2_outputs(6828) <= not (a and b);
    layer2_outputs(6829) <= not a;
    layer2_outputs(6830) <= not (a and b);
    layer2_outputs(6831) <= a and b;
    layer2_outputs(6832) <= 1'b1;
    layer2_outputs(6833) <= a and not b;
    layer2_outputs(6834) <= a and not b;
    layer2_outputs(6835) <= 1'b1;
    layer2_outputs(6836) <= 1'b1;
    layer2_outputs(6837) <= b and not a;
    layer2_outputs(6838) <= not (a xor b);
    layer2_outputs(6839) <= a;
    layer2_outputs(6840) <= not a;
    layer2_outputs(6841) <= not (a and b);
    layer2_outputs(6842) <= not (a xor b);
    layer2_outputs(6843) <= a and b;
    layer2_outputs(6844) <= not (a and b);
    layer2_outputs(6845) <= b and not a;
    layer2_outputs(6846) <= b;
    layer2_outputs(6847) <= not (a and b);
    layer2_outputs(6848) <= not a or b;
    layer2_outputs(6849) <= 1'b0;
    layer2_outputs(6850) <= a and not b;
    layer2_outputs(6851) <= b and not a;
    layer2_outputs(6852) <= b and not a;
    layer2_outputs(6853) <= a and b;
    layer2_outputs(6854) <= b;
    layer2_outputs(6855) <= 1'b1;
    layer2_outputs(6856) <= not a or b;
    layer2_outputs(6857) <= a;
    layer2_outputs(6858) <= a or b;
    layer2_outputs(6859) <= a and not b;
    layer2_outputs(6860) <= not b;
    layer2_outputs(6861) <= a and b;
    layer2_outputs(6862) <= not a;
    layer2_outputs(6863) <= not a or b;
    layer2_outputs(6864) <= not b;
    layer2_outputs(6865) <= 1'b0;
    layer2_outputs(6866) <= not b;
    layer2_outputs(6867) <= not b;
    layer2_outputs(6868) <= a and b;
    layer2_outputs(6869) <= not a or b;
    layer2_outputs(6870) <= not b or a;
    layer2_outputs(6871) <= not (a or b);
    layer2_outputs(6872) <= b and not a;
    layer2_outputs(6873) <= not b;
    layer2_outputs(6874) <= not a or b;
    layer2_outputs(6875) <= b;
    layer2_outputs(6876) <= a and not b;
    layer2_outputs(6877) <= not (a xor b);
    layer2_outputs(6878) <= not a;
    layer2_outputs(6879) <= not a or b;
    layer2_outputs(6880) <= a and b;
    layer2_outputs(6881) <= not (a or b);
    layer2_outputs(6882) <= not a;
    layer2_outputs(6883) <= not a or b;
    layer2_outputs(6884) <= not (a and b);
    layer2_outputs(6885) <= b and not a;
    layer2_outputs(6886) <= not b;
    layer2_outputs(6887) <= a and b;
    layer2_outputs(6888) <= not b or a;
    layer2_outputs(6889) <= not b or a;
    layer2_outputs(6890) <= not b;
    layer2_outputs(6891) <= not (a or b);
    layer2_outputs(6892) <= a;
    layer2_outputs(6893) <= not (a and b);
    layer2_outputs(6894) <= not (a and b);
    layer2_outputs(6895) <= 1'b1;
    layer2_outputs(6896) <= a and not b;
    layer2_outputs(6897) <= 1'b1;
    layer2_outputs(6898) <= a and not b;
    layer2_outputs(6899) <= a and not b;
    layer2_outputs(6900) <= b and not a;
    layer2_outputs(6901) <= a and b;
    layer2_outputs(6902) <= b and not a;
    layer2_outputs(6903) <= not a or b;
    layer2_outputs(6904) <= 1'b0;
    layer2_outputs(6905) <= 1'b0;
    layer2_outputs(6906) <= a or b;
    layer2_outputs(6907) <= 1'b1;
    layer2_outputs(6908) <= a or b;
    layer2_outputs(6909) <= not b or a;
    layer2_outputs(6910) <= not a;
    layer2_outputs(6911) <= not (a xor b);
    layer2_outputs(6912) <= 1'b1;
    layer2_outputs(6913) <= not a or b;
    layer2_outputs(6914) <= a and not b;
    layer2_outputs(6915) <= not (a and b);
    layer2_outputs(6916) <= a and b;
    layer2_outputs(6917) <= a or b;
    layer2_outputs(6918) <= 1'b1;
    layer2_outputs(6919) <= 1'b0;
    layer2_outputs(6920) <= a and not b;
    layer2_outputs(6921) <= 1'b0;
    layer2_outputs(6922) <= a;
    layer2_outputs(6923) <= 1'b0;
    layer2_outputs(6924) <= not b or a;
    layer2_outputs(6925) <= a;
    layer2_outputs(6926) <= not a or b;
    layer2_outputs(6927) <= a and not b;
    layer2_outputs(6928) <= 1'b0;
    layer2_outputs(6929) <= not b or a;
    layer2_outputs(6930) <= b and not a;
    layer2_outputs(6931) <= not a or b;
    layer2_outputs(6932) <= 1'b1;
    layer2_outputs(6933) <= a and not b;
    layer2_outputs(6934) <= a or b;
    layer2_outputs(6935) <= a and b;
    layer2_outputs(6936) <= not (a and b);
    layer2_outputs(6937) <= b and not a;
    layer2_outputs(6938) <= 1'b0;
    layer2_outputs(6939) <= not b or a;
    layer2_outputs(6940) <= not (a or b);
    layer2_outputs(6941) <= not b or a;
    layer2_outputs(6942) <= a and not b;
    layer2_outputs(6943) <= not (a and b);
    layer2_outputs(6944) <= not a;
    layer2_outputs(6945) <= not a or b;
    layer2_outputs(6946) <= not b;
    layer2_outputs(6947) <= a and b;
    layer2_outputs(6948) <= a xor b;
    layer2_outputs(6949) <= a and not b;
    layer2_outputs(6950) <= a and b;
    layer2_outputs(6951) <= 1'b1;
    layer2_outputs(6952) <= not (a and b);
    layer2_outputs(6953) <= not b or a;
    layer2_outputs(6954) <= not b or a;
    layer2_outputs(6955) <= a and not b;
    layer2_outputs(6956) <= 1'b1;
    layer2_outputs(6957) <= not (a and b);
    layer2_outputs(6958) <= not (a or b);
    layer2_outputs(6959) <= not a or b;
    layer2_outputs(6960) <= 1'b1;
    layer2_outputs(6961) <= 1'b1;
    layer2_outputs(6962) <= a;
    layer2_outputs(6963) <= not (a or b);
    layer2_outputs(6964) <= a and b;
    layer2_outputs(6965) <= not (a xor b);
    layer2_outputs(6966) <= a and b;
    layer2_outputs(6967) <= a and not b;
    layer2_outputs(6968) <= a;
    layer2_outputs(6969) <= not (a or b);
    layer2_outputs(6970) <= not a or b;
    layer2_outputs(6971) <= not a;
    layer2_outputs(6972) <= b and not a;
    layer2_outputs(6973) <= not b or a;
    layer2_outputs(6974) <= not b;
    layer2_outputs(6975) <= b;
    layer2_outputs(6976) <= not a;
    layer2_outputs(6977) <= a or b;
    layer2_outputs(6978) <= 1'b0;
    layer2_outputs(6979) <= b;
    layer2_outputs(6980) <= 1'b1;
    layer2_outputs(6981) <= 1'b0;
    layer2_outputs(6982) <= not b or a;
    layer2_outputs(6983) <= not (a or b);
    layer2_outputs(6984) <= a and b;
    layer2_outputs(6985) <= not a;
    layer2_outputs(6986) <= b;
    layer2_outputs(6987) <= not a or b;
    layer2_outputs(6988) <= not b or a;
    layer2_outputs(6989) <= not (a and b);
    layer2_outputs(6990) <= 1'b0;
    layer2_outputs(6991) <= a and b;
    layer2_outputs(6992) <= not a;
    layer2_outputs(6993) <= not b or a;
    layer2_outputs(6994) <= not (a and b);
    layer2_outputs(6995) <= b and not a;
    layer2_outputs(6996) <= not (a xor b);
    layer2_outputs(6997) <= 1'b0;
    layer2_outputs(6998) <= not (a and b);
    layer2_outputs(6999) <= a and not b;
    layer2_outputs(7000) <= a and b;
    layer2_outputs(7001) <= not (a xor b);
    layer2_outputs(7002) <= not (a or b);
    layer2_outputs(7003) <= 1'b0;
    layer2_outputs(7004) <= not (a or b);
    layer2_outputs(7005) <= a;
    layer2_outputs(7006) <= b and not a;
    layer2_outputs(7007) <= b and not a;
    layer2_outputs(7008) <= a and b;
    layer2_outputs(7009) <= not (a or b);
    layer2_outputs(7010) <= 1'b1;
    layer2_outputs(7011) <= a and not b;
    layer2_outputs(7012) <= not a;
    layer2_outputs(7013) <= a or b;
    layer2_outputs(7014) <= not a or b;
    layer2_outputs(7015) <= a and not b;
    layer2_outputs(7016) <= 1'b0;
    layer2_outputs(7017) <= a or b;
    layer2_outputs(7018) <= 1'b1;
    layer2_outputs(7019) <= not a;
    layer2_outputs(7020) <= 1'b0;
    layer2_outputs(7021) <= a or b;
    layer2_outputs(7022) <= not b or a;
    layer2_outputs(7023) <= b;
    layer2_outputs(7024) <= not (a or b);
    layer2_outputs(7025) <= not (a and b);
    layer2_outputs(7026) <= not (a or b);
    layer2_outputs(7027) <= not a or b;
    layer2_outputs(7028) <= a and not b;
    layer2_outputs(7029) <= 1'b1;
    layer2_outputs(7030) <= not b or a;
    layer2_outputs(7031) <= not (a and b);
    layer2_outputs(7032) <= not a or b;
    layer2_outputs(7033) <= a and b;
    layer2_outputs(7034) <= not a or b;
    layer2_outputs(7035) <= 1'b0;
    layer2_outputs(7036) <= a or b;
    layer2_outputs(7037) <= not a or b;
    layer2_outputs(7038) <= 1'b1;
    layer2_outputs(7039) <= not b or a;
    layer2_outputs(7040) <= not b;
    layer2_outputs(7041) <= 1'b0;
    layer2_outputs(7042) <= 1'b1;
    layer2_outputs(7043) <= not (a or b);
    layer2_outputs(7044) <= 1'b1;
    layer2_outputs(7045) <= a;
    layer2_outputs(7046) <= a and not b;
    layer2_outputs(7047) <= not a;
    layer2_outputs(7048) <= not a;
    layer2_outputs(7049) <= not a or b;
    layer2_outputs(7050) <= not a;
    layer2_outputs(7051) <= not b or a;
    layer2_outputs(7052) <= a or b;
    layer2_outputs(7053) <= 1'b1;
    layer2_outputs(7054) <= not (a xor b);
    layer2_outputs(7055) <= not b;
    layer2_outputs(7056) <= not b or a;
    layer2_outputs(7057) <= b and not a;
    layer2_outputs(7058) <= not a;
    layer2_outputs(7059) <= not (a or b);
    layer2_outputs(7060) <= not b or a;
    layer2_outputs(7061) <= a and not b;
    layer2_outputs(7062) <= a and not b;
    layer2_outputs(7063) <= a;
    layer2_outputs(7064) <= a;
    layer2_outputs(7065) <= 1'b0;
    layer2_outputs(7066) <= not a or b;
    layer2_outputs(7067) <= a and b;
    layer2_outputs(7068) <= 1'b1;
    layer2_outputs(7069) <= not a;
    layer2_outputs(7070) <= 1'b0;
    layer2_outputs(7071) <= a or b;
    layer2_outputs(7072) <= a or b;
    layer2_outputs(7073) <= b and not a;
    layer2_outputs(7074) <= b;
    layer2_outputs(7075) <= not b;
    layer2_outputs(7076) <= not (a or b);
    layer2_outputs(7077) <= 1'b0;
    layer2_outputs(7078) <= a and b;
    layer2_outputs(7079) <= not b or a;
    layer2_outputs(7080) <= a;
    layer2_outputs(7081) <= a and b;
    layer2_outputs(7082) <= a and b;
    layer2_outputs(7083) <= b and not a;
    layer2_outputs(7084) <= b and not a;
    layer2_outputs(7085) <= a and b;
    layer2_outputs(7086) <= not b;
    layer2_outputs(7087) <= not (a or b);
    layer2_outputs(7088) <= not b or a;
    layer2_outputs(7089) <= a and not b;
    layer2_outputs(7090) <= b and not a;
    layer2_outputs(7091) <= not (a and b);
    layer2_outputs(7092) <= not b or a;
    layer2_outputs(7093) <= a and b;
    layer2_outputs(7094) <= a or b;
    layer2_outputs(7095) <= 1'b0;
    layer2_outputs(7096) <= not (a or b);
    layer2_outputs(7097) <= b;
    layer2_outputs(7098) <= a or b;
    layer2_outputs(7099) <= not b or a;
    layer2_outputs(7100) <= not (a and b);
    layer2_outputs(7101) <= not b or a;
    layer2_outputs(7102) <= 1'b0;
    layer2_outputs(7103) <= a and b;
    layer2_outputs(7104) <= a or b;
    layer2_outputs(7105) <= not a or b;
    layer2_outputs(7106) <= b;
    layer2_outputs(7107) <= not a;
    layer2_outputs(7108) <= b;
    layer2_outputs(7109) <= not a;
    layer2_outputs(7110) <= b;
    layer2_outputs(7111) <= 1'b1;
    layer2_outputs(7112) <= not b or a;
    layer2_outputs(7113) <= a and not b;
    layer2_outputs(7114) <= not a or b;
    layer2_outputs(7115) <= not (a and b);
    layer2_outputs(7116) <= not a or b;
    layer2_outputs(7117) <= not a or b;
    layer2_outputs(7118) <= a xor b;
    layer2_outputs(7119) <= a xor b;
    layer2_outputs(7120) <= 1'b1;
    layer2_outputs(7121) <= b and not a;
    layer2_outputs(7122) <= a;
    layer2_outputs(7123) <= not a or b;
    layer2_outputs(7124) <= b;
    layer2_outputs(7125) <= b;
    layer2_outputs(7126) <= a;
    layer2_outputs(7127) <= not b or a;
    layer2_outputs(7128) <= not (a and b);
    layer2_outputs(7129) <= a and not b;
    layer2_outputs(7130) <= a and not b;
    layer2_outputs(7131) <= 1'b0;
    layer2_outputs(7132) <= a;
    layer2_outputs(7133) <= b and not a;
    layer2_outputs(7134) <= 1'b1;
    layer2_outputs(7135) <= 1'b1;
    layer2_outputs(7136) <= a and not b;
    layer2_outputs(7137) <= not b;
    layer2_outputs(7138) <= b;
    layer2_outputs(7139) <= not a or b;
    layer2_outputs(7140) <= not b;
    layer2_outputs(7141) <= a and not b;
    layer2_outputs(7142) <= b and not a;
    layer2_outputs(7143) <= not a;
    layer2_outputs(7144) <= not b or a;
    layer2_outputs(7145) <= b and not a;
    layer2_outputs(7146) <= not a or b;
    layer2_outputs(7147) <= not a or b;
    layer2_outputs(7148) <= a and not b;
    layer2_outputs(7149) <= not b;
    layer2_outputs(7150) <= not b;
    layer2_outputs(7151) <= not a;
    layer2_outputs(7152) <= 1'b1;
    layer2_outputs(7153) <= not a;
    layer2_outputs(7154) <= b and not a;
    layer2_outputs(7155) <= not b or a;
    layer2_outputs(7156) <= 1'b1;
    layer2_outputs(7157) <= not (a or b);
    layer2_outputs(7158) <= not a;
    layer2_outputs(7159) <= 1'b0;
    layer2_outputs(7160) <= 1'b0;
    layer2_outputs(7161) <= not b or a;
    layer2_outputs(7162) <= b and not a;
    layer2_outputs(7163) <= not a;
    layer2_outputs(7164) <= not a;
    layer2_outputs(7165) <= a;
    layer2_outputs(7166) <= 1'b1;
    layer2_outputs(7167) <= b and not a;
    layer2_outputs(7168) <= not (a or b);
    layer2_outputs(7169) <= a or b;
    layer2_outputs(7170) <= a and not b;
    layer2_outputs(7171) <= a or b;
    layer2_outputs(7172) <= 1'b1;
    layer2_outputs(7173) <= not a;
    layer2_outputs(7174) <= not a or b;
    layer2_outputs(7175) <= not (a and b);
    layer2_outputs(7176) <= a and not b;
    layer2_outputs(7177) <= not b or a;
    layer2_outputs(7178) <= a and not b;
    layer2_outputs(7179) <= not a;
    layer2_outputs(7180) <= not a or b;
    layer2_outputs(7181) <= not (a and b);
    layer2_outputs(7182) <= not (a xor b);
    layer2_outputs(7183) <= not a or b;
    layer2_outputs(7184) <= 1'b0;
    layer2_outputs(7185) <= not a;
    layer2_outputs(7186) <= not a or b;
    layer2_outputs(7187) <= 1'b0;
    layer2_outputs(7188) <= not (a and b);
    layer2_outputs(7189) <= a and b;
    layer2_outputs(7190) <= a and b;
    layer2_outputs(7191) <= not (a or b);
    layer2_outputs(7192) <= not (a or b);
    layer2_outputs(7193) <= not a or b;
    layer2_outputs(7194) <= not b;
    layer2_outputs(7195) <= a or b;
    layer2_outputs(7196) <= 1'b0;
    layer2_outputs(7197) <= not b;
    layer2_outputs(7198) <= a or b;
    layer2_outputs(7199) <= a and b;
    layer2_outputs(7200) <= not a or b;
    layer2_outputs(7201) <= not (a or b);
    layer2_outputs(7202) <= 1'b1;
    layer2_outputs(7203) <= not (a and b);
    layer2_outputs(7204) <= 1'b1;
    layer2_outputs(7205) <= not (a or b);
    layer2_outputs(7206) <= 1'b0;
    layer2_outputs(7207) <= b;
    layer2_outputs(7208) <= 1'b0;
    layer2_outputs(7209) <= 1'b0;
    layer2_outputs(7210) <= not a;
    layer2_outputs(7211) <= 1'b0;
    layer2_outputs(7212) <= a or b;
    layer2_outputs(7213) <= not (a or b);
    layer2_outputs(7214) <= not (a and b);
    layer2_outputs(7215) <= not (a xor b);
    layer2_outputs(7216) <= 1'b1;
    layer2_outputs(7217) <= not b;
    layer2_outputs(7218) <= b and not a;
    layer2_outputs(7219) <= a and not b;
    layer2_outputs(7220) <= b and not a;
    layer2_outputs(7221) <= a and not b;
    layer2_outputs(7222) <= not (a or b);
    layer2_outputs(7223) <= not (a or b);
    layer2_outputs(7224) <= a and b;
    layer2_outputs(7225) <= not b or a;
    layer2_outputs(7226) <= a;
    layer2_outputs(7227) <= a;
    layer2_outputs(7228) <= 1'b1;
    layer2_outputs(7229) <= 1'b0;
    layer2_outputs(7230) <= a and b;
    layer2_outputs(7231) <= a;
    layer2_outputs(7232) <= a and not b;
    layer2_outputs(7233) <= not (a or b);
    layer2_outputs(7234) <= 1'b1;
    layer2_outputs(7235) <= a xor b;
    layer2_outputs(7236) <= not (a and b);
    layer2_outputs(7237) <= not b;
    layer2_outputs(7238) <= a or b;
    layer2_outputs(7239) <= b;
    layer2_outputs(7240) <= not b;
    layer2_outputs(7241) <= not a or b;
    layer2_outputs(7242) <= 1'b1;
    layer2_outputs(7243) <= a;
    layer2_outputs(7244) <= not b or a;
    layer2_outputs(7245) <= not (a or b);
    layer2_outputs(7246) <= a and not b;
    layer2_outputs(7247) <= not a;
    layer2_outputs(7248) <= not a or b;
    layer2_outputs(7249) <= not a or b;
    layer2_outputs(7250) <= a xor b;
    layer2_outputs(7251) <= b and not a;
    layer2_outputs(7252) <= 1'b0;
    layer2_outputs(7253) <= not (a and b);
    layer2_outputs(7254) <= not a;
    layer2_outputs(7255) <= not b or a;
    layer2_outputs(7256) <= 1'b0;
    layer2_outputs(7257) <= not a;
    layer2_outputs(7258) <= 1'b1;
    layer2_outputs(7259) <= 1'b1;
    layer2_outputs(7260) <= a;
    layer2_outputs(7261) <= a or b;
    layer2_outputs(7262) <= not b or a;
    layer2_outputs(7263) <= not a or b;
    layer2_outputs(7264) <= not (a or b);
    layer2_outputs(7265) <= 1'b0;
    layer2_outputs(7266) <= not (a and b);
    layer2_outputs(7267) <= not a;
    layer2_outputs(7268) <= not a or b;
    layer2_outputs(7269) <= not a;
    layer2_outputs(7270) <= b;
    layer2_outputs(7271) <= not (a or b);
    layer2_outputs(7272) <= b and not a;
    layer2_outputs(7273) <= a xor b;
    layer2_outputs(7274) <= a xor b;
    layer2_outputs(7275) <= 1'b0;
    layer2_outputs(7276) <= b and not a;
    layer2_outputs(7277) <= not (a or b);
    layer2_outputs(7278) <= not (a or b);
    layer2_outputs(7279) <= b;
    layer2_outputs(7280) <= not (a and b);
    layer2_outputs(7281) <= 1'b1;
    layer2_outputs(7282) <= not (a or b);
    layer2_outputs(7283) <= a and b;
    layer2_outputs(7284) <= a and not b;
    layer2_outputs(7285) <= a and not b;
    layer2_outputs(7286) <= not a or b;
    layer2_outputs(7287) <= not a or b;
    layer2_outputs(7288) <= not (a or b);
    layer2_outputs(7289) <= b and not a;
    layer2_outputs(7290) <= not (a or b);
    layer2_outputs(7291) <= a and not b;
    layer2_outputs(7292) <= a xor b;
    layer2_outputs(7293) <= b;
    layer2_outputs(7294) <= not b;
    layer2_outputs(7295) <= not a or b;
    layer2_outputs(7296) <= a and b;
    layer2_outputs(7297) <= not (a and b);
    layer2_outputs(7298) <= a or b;
    layer2_outputs(7299) <= not (a and b);
    layer2_outputs(7300) <= a;
    layer2_outputs(7301) <= not a or b;
    layer2_outputs(7302) <= 1'b1;
    layer2_outputs(7303) <= b;
    layer2_outputs(7304) <= a and b;
    layer2_outputs(7305) <= 1'b1;
    layer2_outputs(7306) <= a and b;
    layer2_outputs(7307) <= 1'b0;
    layer2_outputs(7308) <= b;
    layer2_outputs(7309) <= a or b;
    layer2_outputs(7310) <= not a or b;
    layer2_outputs(7311) <= a or b;
    layer2_outputs(7312) <= not (a and b);
    layer2_outputs(7313) <= not (a and b);
    layer2_outputs(7314) <= 1'b0;
    layer2_outputs(7315) <= b and not a;
    layer2_outputs(7316) <= 1'b1;
    layer2_outputs(7317) <= a and not b;
    layer2_outputs(7318) <= 1'b1;
    layer2_outputs(7319) <= not b;
    layer2_outputs(7320) <= a;
    layer2_outputs(7321) <= 1'b1;
    layer2_outputs(7322) <= not b;
    layer2_outputs(7323) <= not b;
    layer2_outputs(7324) <= not b or a;
    layer2_outputs(7325) <= 1'b1;
    layer2_outputs(7326) <= not (a or b);
    layer2_outputs(7327) <= not b or a;
    layer2_outputs(7328) <= a;
    layer2_outputs(7329) <= not (a or b);
    layer2_outputs(7330) <= b and not a;
    layer2_outputs(7331) <= a and not b;
    layer2_outputs(7332) <= not a;
    layer2_outputs(7333) <= a and b;
    layer2_outputs(7334) <= 1'b0;
    layer2_outputs(7335) <= a xor b;
    layer2_outputs(7336) <= not (a xor b);
    layer2_outputs(7337) <= 1'b1;
    layer2_outputs(7338) <= 1'b0;
    layer2_outputs(7339) <= not a;
    layer2_outputs(7340) <= not (a or b);
    layer2_outputs(7341) <= not a;
    layer2_outputs(7342) <= 1'b0;
    layer2_outputs(7343) <= 1'b0;
    layer2_outputs(7344) <= a or b;
    layer2_outputs(7345) <= not b;
    layer2_outputs(7346) <= a;
    layer2_outputs(7347) <= b and not a;
    layer2_outputs(7348) <= not (a xor b);
    layer2_outputs(7349) <= 1'b1;
    layer2_outputs(7350) <= b;
    layer2_outputs(7351) <= not b;
    layer2_outputs(7352) <= b;
    layer2_outputs(7353) <= not b;
    layer2_outputs(7354) <= not a;
    layer2_outputs(7355) <= not b;
    layer2_outputs(7356) <= 1'b1;
    layer2_outputs(7357) <= 1'b0;
    layer2_outputs(7358) <= not a or b;
    layer2_outputs(7359) <= a and b;
    layer2_outputs(7360) <= b and not a;
    layer2_outputs(7361) <= not a;
    layer2_outputs(7362) <= not b or a;
    layer2_outputs(7363) <= not b or a;
    layer2_outputs(7364) <= b and not a;
    layer2_outputs(7365) <= b and not a;
    layer2_outputs(7366) <= 1'b0;
    layer2_outputs(7367) <= a;
    layer2_outputs(7368) <= not (a and b);
    layer2_outputs(7369) <= b;
    layer2_outputs(7370) <= b;
    layer2_outputs(7371) <= not (a and b);
    layer2_outputs(7372) <= not (a and b);
    layer2_outputs(7373) <= a or b;
    layer2_outputs(7374) <= a;
    layer2_outputs(7375) <= 1'b1;
    layer2_outputs(7376) <= not b;
    layer2_outputs(7377) <= a or b;
    layer2_outputs(7378) <= 1'b0;
    layer2_outputs(7379) <= a;
    layer2_outputs(7380) <= 1'b0;
    layer2_outputs(7381) <= 1'b1;
    layer2_outputs(7382) <= a or b;
    layer2_outputs(7383) <= a or b;
    layer2_outputs(7384) <= not b or a;
    layer2_outputs(7385) <= 1'b1;
    layer2_outputs(7386) <= not (a or b);
    layer2_outputs(7387) <= a and b;
    layer2_outputs(7388) <= 1'b0;
    layer2_outputs(7389) <= b;
    layer2_outputs(7390) <= 1'b1;
    layer2_outputs(7391) <= not a;
    layer2_outputs(7392) <= 1'b1;
    layer2_outputs(7393) <= b;
    layer2_outputs(7394) <= not (a and b);
    layer2_outputs(7395) <= not (a or b);
    layer2_outputs(7396) <= a;
    layer2_outputs(7397) <= a;
    layer2_outputs(7398) <= not b or a;
    layer2_outputs(7399) <= a;
    layer2_outputs(7400) <= a;
    layer2_outputs(7401) <= a and b;
    layer2_outputs(7402) <= a;
    layer2_outputs(7403) <= not a;
    layer2_outputs(7404) <= not b or a;
    layer2_outputs(7405) <= not a or b;
    layer2_outputs(7406) <= 1'b0;
    layer2_outputs(7407) <= b and not a;
    layer2_outputs(7408) <= not (a or b);
    layer2_outputs(7409) <= 1'b0;
    layer2_outputs(7410) <= a and not b;
    layer2_outputs(7411) <= not b;
    layer2_outputs(7412) <= not a;
    layer2_outputs(7413) <= a xor b;
    layer2_outputs(7414) <= b;
    layer2_outputs(7415) <= 1'b0;
    layer2_outputs(7416) <= not (a or b);
    layer2_outputs(7417) <= not b or a;
    layer2_outputs(7418) <= 1'b1;
    layer2_outputs(7419) <= 1'b0;
    layer2_outputs(7420) <= 1'b0;
    layer2_outputs(7421) <= a and not b;
    layer2_outputs(7422) <= a or b;
    layer2_outputs(7423) <= not a or b;
    layer2_outputs(7424) <= not a or b;
    layer2_outputs(7425) <= b and not a;
    layer2_outputs(7426) <= not a or b;
    layer2_outputs(7427) <= a xor b;
    layer2_outputs(7428) <= 1'b0;
    layer2_outputs(7429) <= b;
    layer2_outputs(7430) <= not b;
    layer2_outputs(7431) <= a;
    layer2_outputs(7432) <= a and b;
    layer2_outputs(7433) <= not a or b;
    layer2_outputs(7434) <= a and not b;
    layer2_outputs(7435) <= not a;
    layer2_outputs(7436) <= 1'b1;
    layer2_outputs(7437) <= 1'b0;
    layer2_outputs(7438) <= 1'b0;
    layer2_outputs(7439) <= 1'b1;
    layer2_outputs(7440) <= a and b;
    layer2_outputs(7441) <= not a;
    layer2_outputs(7442) <= 1'b1;
    layer2_outputs(7443) <= not a;
    layer2_outputs(7444) <= b;
    layer2_outputs(7445) <= not b or a;
    layer2_outputs(7446) <= 1'b1;
    layer2_outputs(7447) <= a and b;
    layer2_outputs(7448) <= a and b;
    layer2_outputs(7449) <= a and not b;
    layer2_outputs(7450) <= not (a xor b);
    layer2_outputs(7451) <= a or b;
    layer2_outputs(7452) <= not (a or b);
    layer2_outputs(7453) <= a;
    layer2_outputs(7454) <= not (a and b);
    layer2_outputs(7455) <= not a or b;
    layer2_outputs(7456) <= not b or a;
    layer2_outputs(7457) <= 1'b1;
    layer2_outputs(7458) <= b;
    layer2_outputs(7459) <= a;
    layer2_outputs(7460) <= 1'b1;
    layer2_outputs(7461) <= not a;
    layer2_outputs(7462) <= b;
    layer2_outputs(7463) <= b;
    layer2_outputs(7464) <= b and not a;
    layer2_outputs(7465) <= a and b;
    layer2_outputs(7466) <= a or b;
    layer2_outputs(7467) <= not a or b;
    layer2_outputs(7468) <= not b or a;
    layer2_outputs(7469) <= 1'b1;
    layer2_outputs(7470) <= a and not b;
    layer2_outputs(7471) <= not (a and b);
    layer2_outputs(7472) <= b;
    layer2_outputs(7473) <= not b or a;
    layer2_outputs(7474) <= not b or a;
    layer2_outputs(7475) <= not b or a;
    layer2_outputs(7476) <= a or b;
    layer2_outputs(7477) <= a or b;
    layer2_outputs(7478) <= not (a and b);
    layer2_outputs(7479) <= not b or a;
    layer2_outputs(7480) <= a or b;
    layer2_outputs(7481) <= not (a and b);
    layer2_outputs(7482) <= a and b;
    layer2_outputs(7483) <= not (a or b);
    layer2_outputs(7484) <= not a or b;
    layer2_outputs(7485) <= 1'b1;
    layer2_outputs(7486) <= not (a or b);
    layer2_outputs(7487) <= not (a xor b);
    layer2_outputs(7488) <= not a or b;
    layer2_outputs(7489) <= not (a or b);
    layer2_outputs(7490) <= not b or a;
    layer2_outputs(7491) <= not b;
    layer2_outputs(7492) <= not a;
    layer2_outputs(7493) <= 1'b1;
    layer2_outputs(7494) <= a and b;
    layer2_outputs(7495) <= 1'b0;
    layer2_outputs(7496) <= not b or a;
    layer2_outputs(7497) <= not a or b;
    layer2_outputs(7498) <= 1'b1;
    layer2_outputs(7499) <= not b or a;
    layer2_outputs(7500) <= 1'b1;
    layer2_outputs(7501) <= b and not a;
    layer2_outputs(7502) <= a and not b;
    layer2_outputs(7503) <= 1'b0;
    layer2_outputs(7504) <= 1'b1;
    layer2_outputs(7505) <= not (a or b);
    layer2_outputs(7506) <= a or b;
    layer2_outputs(7507) <= a and b;
    layer2_outputs(7508) <= not (a and b);
    layer2_outputs(7509) <= not b or a;
    layer2_outputs(7510) <= not (a and b);
    layer2_outputs(7511) <= b and not a;
    layer2_outputs(7512) <= not b;
    layer2_outputs(7513) <= 1'b1;
    layer2_outputs(7514) <= a or b;
    layer2_outputs(7515) <= b and not a;
    layer2_outputs(7516) <= a;
    layer2_outputs(7517) <= a and b;
    layer2_outputs(7518) <= not b or a;
    layer2_outputs(7519) <= a or b;
    layer2_outputs(7520) <= not (a and b);
    layer2_outputs(7521) <= a and not b;
    layer2_outputs(7522) <= 1'b1;
    layer2_outputs(7523) <= a;
    layer2_outputs(7524) <= 1'b1;
    layer2_outputs(7525) <= not b;
    layer2_outputs(7526) <= a;
    layer2_outputs(7527) <= a;
    layer2_outputs(7528) <= not b or a;
    layer2_outputs(7529) <= 1'b1;
    layer2_outputs(7530) <= not b;
    layer2_outputs(7531) <= not a or b;
    layer2_outputs(7532) <= a;
    layer2_outputs(7533) <= not (a xor b);
    layer2_outputs(7534) <= 1'b1;
    layer2_outputs(7535) <= 1'b0;
    layer2_outputs(7536) <= not b or a;
    layer2_outputs(7537) <= not a;
    layer2_outputs(7538) <= b and not a;
    layer2_outputs(7539) <= not (a xor b);
    layer2_outputs(7540) <= 1'b0;
    layer2_outputs(7541) <= not (a or b);
    layer2_outputs(7542) <= not (a and b);
    layer2_outputs(7543) <= not a or b;
    layer2_outputs(7544) <= a xor b;
    layer2_outputs(7545) <= b;
    layer2_outputs(7546) <= 1'b0;
    layer2_outputs(7547) <= 1'b0;
    layer2_outputs(7548) <= not b or a;
    layer2_outputs(7549) <= b;
    layer2_outputs(7550) <= not b or a;
    layer2_outputs(7551) <= b;
    layer2_outputs(7552) <= not (a and b);
    layer2_outputs(7553) <= not a or b;
    layer2_outputs(7554) <= 1'b1;
    layer2_outputs(7555) <= b and not a;
    layer2_outputs(7556) <= not b;
    layer2_outputs(7557) <= a and not b;
    layer2_outputs(7558) <= a;
    layer2_outputs(7559) <= not (a or b);
    layer2_outputs(7560) <= b;
    layer2_outputs(7561) <= b and not a;
    layer2_outputs(7562) <= a xor b;
    layer2_outputs(7563) <= not b;
    layer2_outputs(7564) <= not a or b;
    layer2_outputs(7565) <= 1'b1;
    layer2_outputs(7566) <= not (a and b);
    layer2_outputs(7567) <= not a;
    layer2_outputs(7568) <= 1'b0;
    layer2_outputs(7569) <= not (a or b);
    layer2_outputs(7570) <= b and not a;
    layer2_outputs(7571) <= 1'b1;
    layer2_outputs(7572) <= not b or a;
    layer2_outputs(7573) <= b and not a;
    layer2_outputs(7574) <= a xor b;
    layer2_outputs(7575) <= a or b;
    layer2_outputs(7576) <= b;
    layer2_outputs(7577) <= a and not b;
    layer2_outputs(7578) <= b and not a;
    layer2_outputs(7579) <= not b;
    layer2_outputs(7580) <= not (a or b);
    layer2_outputs(7581) <= a and not b;
    layer2_outputs(7582) <= not a;
    layer2_outputs(7583) <= not (a and b);
    layer2_outputs(7584) <= 1'b0;
    layer2_outputs(7585) <= not (a and b);
    layer2_outputs(7586) <= b and not a;
    layer2_outputs(7587) <= not b;
    layer2_outputs(7588) <= b and not a;
    layer2_outputs(7589) <= not b or a;
    layer2_outputs(7590) <= a or b;
    layer2_outputs(7591) <= a and b;
    layer2_outputs(7592) <= not (a or b);
    layer2_outputs(7593) <= not (a and b);
    layer2_outputs(7594) <= not a or b;
    layer2_outputs(7595) <= not a;
    layer2_outputs(7596) <= 1'b1;
    layer2_outputs(7597) <= a xor b;
    layer2_outputs(7598) <= a and not b;
    layer2_outputs(7599) <= a and b;
    layer2_outputs(7600) <= a;
    layer2_outputs(7601) <= b;
    layer2_outputs(7602) <= 1'b0;
    layer2_outputs(7603) <= not a;
    layer2_outputs(7604) <= b and not a;
    layer2_outputs(7605) <= 1'b1;
    layer2_outputs(7606) <= 1'b0;
    layer2_outputs(7607) <= not (a or b);
    layer2_outputs(7608) <= not a;
    layer2_outputs(7609) <= not b;
    layer2_outputs(7610) <= a;
    layer2_outputs(7611) <= a or b;
    layer2_outputs(7612) <= not b;
    layer2_outputs(7613) <= b;
    layer2_outputs(7614) <= a or b;
    layer2_outputs(7615) <= 1'b1;
    layer2_outputs(7616) <= not (a and b);
    layer2_outputs(7617) <= not (a and b);
    layer2_outputs(7618) <= a and not b;
    layer2_outputs(7619) <= a and b;
    layer2_outputs(7620) <= 1'b0;
    layer2_outputs(7621) <= not (a or b);
    layer2_outputs(7622) <= not (a or b);
    layer2_outputs(7623) <= b;
    layer2_outputs(7624) <= not (a and b);
    layer2_outputs(7625) <= not a;
    layer2_outputs(7626) <= not b;
    layer2_outputs(7627) <= not (a and b);
    layer2_outputs(7628) <= not a or b;
    layer2_outputs(7629) <= not (a and b);
    layer2_outputs(7630) <= not b or a;
    layer2_outputs(7631) <= 1'b0;
    layer2_outputs(7632) <= b;
    layer2_outputs(7633) <= 1'b1;
    layer2_outputs(7634) <= a or b;
    layer2_outputs(7635) <= 1'b0;
    layer2_outputs(7636) <= a or b;
    layer2_outputs(7637) <= not a or b;
    layer2_outputs(7638) <= not a or b;
    layer2_outputs(7639) <= 1'b1;
    layer2_outputs(7640) <= a or b;
    layer2_outputs(7641) <= not a or b;
    layer2_outputs(7642) <= a xor b;
    layer2_outputs(7643) <= not (a xor b);
    layer2_outputs(7644) <= not a or b;
    layer2_outputs(7645) <= not (a and b);
    layer2_outputs(7646) <= 1'b1;
    layer2_outputs(7647) <= not (a and b);
    layer2_outputs(7648) <= not (a and b);
    layer2_outputs(7649) <= a and not b;
    layer2_outputs(7650) <= not (a or b);
    layer2_outputs(7651) <= not b;
    layer2_outputs(7652) <= not (a xor b);
    layer2_outputs(7653) <= not b or a;
    layer2_outputs(7654) <= not a;
    layer2_outputs(7655) <= 1'b1;
    layer2_outputs(7656) <= b and not a;
    layer2_outputs(7657) <= a xor b;
    layer2_outputs(7658) <= not (a or b);
    layer2_outputs(7659) <= b and not a;
    layer2_outputs(7660) <= b;
    layer2_outputs(7661) <= not b;
    layer2_outputs(7662) <= not a;
    layer2_outputs(7663) <= a or b;
    layer2_outputs(7664) <= not b or a;
    layer2_outputs(7665) <= a;
    layer2_outputs(7666) <= 1'b0;
    layer2_outputs(7667) <= a and not b;
    layer2_outputs(7668) <= 1'b1;
    layer2_outputs(7669) <= not a or b;
    layer2_outputs(7670) <= not (a and b);
    layer2_outputs(7671) <= not b;
    layer2_outputs(7672) <= a and not b;
    layer2_outputs(7673) <= not b or a;
    layer2_outputs(7674) <= not (a or b);
    layer2_outputs(7675) <= not (a and b);
    layer2_outputs(7676) <= not (a or b);
    layer2_outputs(7677) <= not a or b;
    layer2_outputs(7678) <= a;
    layer2_outputs(7679) <= a and b;
    layer2_outputs(7680) <= 1'b1;
    layer2_outputs(7681) <= not a;
    layer2_outputs(7682) <= not b or a;
    layer2_outputs(7683) <= a and b;
    layer2_outputs(7684) <= not (a or b);
    layer2_outputs(7685) <= a;
    layer2_outputs(7686) <= not a or b;
    layer2_outputs(7687) <= not (a or b);
    layer2_outputs(7688) <= not (a or b);
    layer2_outputs(7689) <= 1'b1;
    layer2_outputs(7690) <= not (a or b);
    layer2_outputs(7691) <= b;
    layer2_outputs(7692) <= not a or b;
    layer2_outputs(7693) <= not (a and b);
    layer2_outputs(7694) <= not b or a;
    layer2_outputs(7695) <= not a;
    layer2_outputs(7696) <= a or b;
    layer2_outputs(7697) <= a;
    layer2_outputs(7698) <= a and b;
    layer2_outputs(7699) <= a and b;
    layer2_outputs(7700) <= a and not b;
    layer2_outputs(7701) <= b;
    layer2_outputs(7702) <= not a;
    layer2_outputs(7703) <= a;
    layer2_outputs(7704) <= 1'b1;
    layer2_outputs(7705) <= not (a or b);
    layer2_outputs(7706) <= a or b;
    layer2_outputs(7707) <= b and not a;
    layer2_outputs(7708) <= b;
    layer2_outputs(7709) <= 1'b0;
    layer2_outputs(7710) <= not a or b;
    layer2_outputs(7711) <= 1'b0;
    layer2_outputs(7712) <= 1'b1;
    layer2_outputs(7713) <= a and b;
    layer2_outputs(7714) <= not b;
    layer2_outputs(7715) <= b and not a;
    layer2_outputs(7716) <= a;
    layer2_outputs(7717) <= not b;
    layer2_outputs(7718) <= a or b;
    layer2_outputs(7719) <= not b;
    layer2_outputs(7720) <= not b;
    layer2_outputs(7721) <= not b or a;
    layer2_outputs(7722) <= not (a or b);
    layer2_outputs(7723) <= a or b;
    layer2_outputs(7724) <= a and b;
    layer2_outputs(7725) <= 1'b0;
    layer2_outputs(7726) <= not (a or b);
    layer2_outputs(7727) <= not a;
    layer2_outputs(7728) <= a;
    layer2_outputs(7729) <= not b;
    layer2_outputs(7730) <= a and b;
    layer2_outputs(7731) <= not a or b;
    layer2_outputs(7732) <= not b or a;
    layer2_outputs(7733) <= not (a and b);
    layer2_outputs(7734) <= a or b;
    layer2_outputs(7735) <= not a;
    layer2_outputs(7736) <= a;
    layer2_outputs(7737) <= not a;
    layer2_outputs(7738) <= not (a xor b);
    layer2_outputs(7739) <= a and b;
    layer2_outputs(7740) <= not b or a;
    layer2_outputs(7741) <= not (a and b);
    layer2_outputs(7742) <= not (a and b);
    layer2_outputs(7743) <= not a;
    layer2_outputs(7744) <= not b or a;
    layer2_outputs(7745) <= a and b;
    layer2_outputs(7746) <= not a;
    layer2_outputs(7747) <= b;
    layer2_outputs(7748) <= a or b;
    layer2_outputs(7749) <= not a or b;
    layer2_outputs(7750) <= b and not a;
    layer2_outputs(7751) <= not a;
    layer2_outputs(7752) <= b;
    layer2_outputs(7753) <= a or b;
    layer2_outputs(7754) <= a and b;
    layer2_outputs(7755) <= not a or b;
    layer2_outputs(7756) <= 1'b0;
    layer2_outputs(7757) <= b and not a;
    layer2_outputs(7758) <= a;
    layer2_outputs(7759) <= a and b;
    layer2_outputs(7760) <= not a or b;
    layer2_outputs(7761) <= a or b;
    layer2_outputs(7762) <= not (a and b);
    layer2_outputs(7763) <= not (a or b);
    layer2_outputs(7764) <= a and b;
    layer2_outputs(7765) <= not b;
    layer2_outputs(7766) <= b;
    layer2_outputs(7767) <= 1'b0;
    layer2_outputs(7768) <= b and not a;
    layer2_outputs(7769) <= 1'b1;
    layer2_outputs(7770) <= b and not a;
    layer2_outputs(7771) <= not (a and b);
    layer2_outputs(7772) <= a;
    layer2_outputs(7773) <= a and not b;
    layer2_outputs(7774) <= b and not a;
    layer2_outputs(7775) <= a and not b;
    layer2_outputs(7776) <= a xor b;
    layer2_outputs(7777) <= b and not a;
    layer2_outputs(7778) <= a and b;
    layer2_outputs(7779) <= not b or a;
    layer2_outputs(7780) <= b;
    layer2_outputs(7781) <= not b;
    layer2_outputs(7782) <= 1'b1;
    layer2_outputs(7783) <= a and not b;
    layer2_outputs(7784) <= not b or a;
    layer2_outputs(7785) <= 1'b0;
    layer2_outputs(7786) <= not (a or b);
    layer2_outputs(7787) <= b and not a;
    layer2_outputs(7788) <= a and not b;
    layer2_outputs(7789) <= not b;
    layer2_outputs(7790) <= a;
    layer2_outputs(7791) <= not (a and b);
    layer2_outputs(7792) <= 1'b1;
    layer2_outputs(7793) <= not (a and b);
    layer2_outputs(7794) <= a or b;
    layer2_outputs(7795) <= b and not a;
    layer2_outputs(7796) <= not b;
    layer2_outputs(7797) <= not a;
    layer2_outputs(7798) <= b and not a;
    layer2_outputs(7799) <= not (a xor b);
    layer2_outputs(7800) <= a and not b;
    layer2_outputs(7801) <= not a or b;
    layer2_outputs(7802) <= a and not b;
    layer2_outputs(7803) <= a and b;
    layer2_outputs(7804) <= a or b;
    layer2_outputs(7805) <= 1'b0;
    layer2_outputs(7806) <= not (a or b);
    layer2_outputs(7807) <= not (a xor b);
    layer2_outputs(7808) <= a and not b;
    layer2_outputs(7809) <= 1'b0;
    layer2_outputs(7810) <= a or b;
    layer2_outputs(7811) <= a and not b;
    layer2_outputs(7812) <= 1'b1;
    layer2_outputs(7813) <= not b;
    layer2_outputs(7814) <= not (a xor b);
    layer2_outputs(7815) <= b;
    layer2_outputs(7816) <= b;
    layer2_outputs(7817) <= a;
    layer2_outputs(7818) <= a or b;
    layer2_outputs(7819) <= a and not b;
    layer2_outputs(7820) <= a or b;
    layer2_outputs(7821) <= a and not b;
    layer2_outputs(7822) <= b;
    layer2_outputs(7823) <= a and not b;
    layer2_outputs(7824) <= not a or b;
    layer2_outputs(7825) <= a and b;
    layer2_outputs(7826) <= not a or b;
    layer2_outputs(7827) <= not (a or b);
    layer2_outputs(7828) <= a and not b;
    layer2_outputs(7829) <= 1'b1;
    layer2_outputs(7830) <= a and b;
    layer2_outputs(7831) <= b;
    layer2_outputs(7832) <= not (a or b);
    layer2_outputs(7833) <= 1'b0;
    layer2_outputs(7834) <= not (a and b);
    layer2_outputs(7835) <= b and not a;
    layer2_outputs(7836) <= not a;
    layer2_outputs(7837) <= not (a or b);
    layer2_outputs(7838) <= b and not a;
    layer2_outputs(7839) <= b and not a;
    layer2_outputs(7840) <= not a;
    layer2_outputs(7841) <= b and not a;
    layer2_outputs(7842) <= not a;
    layer2_outputs(7843) <= not a or b;
    layer2_outputs(7844) <= not (a or b);
    layer2_outputs(7845) <= not (a or b);
    layer2_outputs(7846) <= b and not a;
    layer2_outputs(7847) <= 1'b1;
    layer2_outputs(7848) <= not b;
    layer2_outputs(7849) <= 1'b1;
    layer2_outputs(7850) <= a and b;
    layer2_outputs(7851) <= b;
    layer2_outputs(7852) <= not (a or b);
    layer2_outputs(7853) <= not (a and b);
    layer2_outputs(7854) <= 1'b0;
    layer2_outputs(7855) <= a and b;
    layer2_outputs(7856) <= b and not a;
    layer2_outputs(7857) <= not a;
    layer2_outputs(7858) <= a or b;
    layer2_outputs(7859) <= not (a and b);
    layer2_outputs(7860) <= not b or a;
    layer2_outputs(7861) <= not (a or b);
    layer2_outputs(7862) <= not a or b;
    layer2_outputs(7863) <= not (a or b);
    layer2_outputs(7864) <= not b or a;
    layer2_outputs(7865) <= a or b;
    layer2_outputs(7866) <= not b;
    layer2_outputs(7867) <= not a;
    layer2_outputs(7868) <= a and not b;
    layer2_outputs(7869) <= not a;
    layer2_outputs(7870) <= 1'b0;
    layer2_outputs(7871) <= not (a and b);
    layer2_outputs(7872) <= not a or b;
    layer2_outputs(7873) <= not (a and b);
    layer2_outputs(7874) <= 1'b1;
    layer2_outputs(7875) <= not (a or b);
    layer2_outputs(7876) <= a;
    layer2_outputs(7877) <= a;
    layer2_outputs(7878) <= not (a or b);
    layer2_outputs(7879) <= a;
    layer2_outputs(7880) <= a xor b;
    layer2_outputs(7881) <= not (a and b);
    layer2_outputs(7882) <= not b or a;
    layer2_outputs(7883) <= a and b;
    layer2_outputs(7884) <= not b;
    layer2_outputs(7885) <= not a or b;
    layer2_outputs(7886) <= a and b;
    layer2_outputs(7887) <= not (a and b);
    layer2_outputs(7888) <= b;
    layer2_outputs(7889) <= not b or a;
    layer2_outputs(7890) <= a and b;
    layer2_outputs(7891) <= not (a and b);
    layer2_outputs(7892) <= not (a or b);
    layer2_outputs(7893) <= a and b;
    layer2_outputs(7894) <= not (a or b);
    layer2_outputs(7895) <= not (a and b);
    layer2_outputs(7896) <= not b or a;
    layer2_outputs(7897) <= a and b;
    layer2_outputs(7898) <= not b;
    layer2_outputs(7899) <= a and not b;
    layer2_outputs(7900) <= not (a xor b);
    layer2_outputs(7901) <= a;
    layer2_outputs(7902) <= not a or b;
    layer2_outputs(7903) <= a;
    layer2_outputs(7904) <= a xor b;
    layer2_outputs(7905) <= not b or a;
    layer2_outputs(7906) <= a and b;
    layer2_outputs(7907) <= not (a or b);
    layer2_outputs(7908) <= not b or a;
    layer2_outputs(7909) <= b;
    layer2_outputs(7910) <= b and not a;
    layer2_outputs(7911) <= a;
    layer2_outputs(7912) <= not (a and b);
    layer2_outputs(7913) <= b and not a;
    layer2_outputs(7914) <= b and not a;
    layer2_outputs(7915) <= not (a or b);
    layer2_outputs(7916) <= a and b;
    layer2_outputs(7917) <= 1'b1;
    layer2_outputs(7918) <= 1'b0;
    layer2_outputs(7919) <= not (a and b);
    layer2_outputs(7920) <= 1'b0;
    layer2_outputs(7921) <= not (a and b);
    layer2_outputs(7922) <= a and b;
    layer2_outputs(7923) <= a;
    layer2_outputs(7924) <= a and not b;
    layer2_outputs(7925) <= not (a and b);
    layer2_outputs(7926) <= a xor b;
    layer2_outputs(7927) <= not a or b;
    layer2_outputs(7928) <= not a;
    layer2_outputs(7929) <= not (a or b);
    layer2_outputs(7930) <= 1'b1;
    layer2_outputs(7931) <= b and not a;
    layer2_outputs(7932) <= b;
    layer2_outputs(7933) <= not (a xor b);
    layer2_outputs(7934) <= a and b;
    layer2_outputs(7935) <= 1'b0;
    layer2_outputs(7936) <= a or b;
    layer2_outputs(7937) <= 1'b1;
    layer2_outputs(7938) <= 1'b1;
    layer2_outputs(7939) <= a or b;
    layer2_outputs(7940) <= 1'b0;
    layer2_outputs(7941) <= not b or a;
    layer2_outputs(7942) <= not b or a;
    layer2_outputs(7943) <= b;
    layer2_outputs(7944) <= not (a and b);
    layer2_outputs(7945) <= a xor b;
    layer2_outputs(7946) <= 1'b1;
    layer2_outputs(7947) <= not a or b;
    layer2_outputs(7948) <= 1'b0;
    layer2_outputs(7949) <= 1'b0;
    layer2_outputs(7950) <= 1'b1;
    layer2_outputs(7951) <= a and not b;
    layer2_outputs(7952) <= a and b;
    layer2_outputs(7953) <= not b or a;
    layer2_outputs(7954) <= 1'b1;
    layer2_outputs(7955) <= not a or b;
    layer2_outputs(7956) <= a and not b;
    layer2_outputs(7957) <= b;
    layer2_outputs(7958) <= not b;
    layer2_outputs(7959) <= not b or a;
    layer2_outputs(7960) <= not (a and b);
    layer2_outputs(7961) <= not (a and b);
    layer2_outputs(7962) <= not (a or b);
    layer2_outputs(7963) <= a;
    layer2_outputs(7964) <= 1'b0;
    layer2_outputs(7965) <= not b;
    layer2_outputs(7966) <= b and not a;
    layer2_outputs(7967) <= 1'b0;
    layer2_outputs(7968) <= not (a or b);
    layer2_outputs(7969) <= a and b;
    layer2_outputs(7970) <= b and not a;
    layer2_outputs(7971) <= not (a and b);
    layer2_outputs(7972) <= not (a xor b);
    layer2_outputs(7973) <= 1'b0;
    layer2_outputs(7974) <= not (a and b);
    layer2_outputs(7975) <= not b or a;
    layer2_outputs(7976) <= 1'b1;
    layer2_outputs(7977) <= b and not a;
    layer2_outputs(7978) <= not b;
    layer2_outputs(7979) <= a;
    layer2_outputs(7980) <= not a;
    layer2_outputs(7981) <= not b;
    layer2_outputs(7982) <= a xor b;
    layer2_outputs(7983) <= not (a or b);
    layer2_outputs(7984) <= not b or a;
    layer2_outputs(7985) <= 1'b1;
    layer2_outputs(7986) <= not (a or b);
    layer2_outputs(7987) <= a and not b;
    layer2_outputs(7988) <= not (a and b);
    layer2_outputs(7989) <= not (a or b);
    layer2_outputs(7990) <= 1'b0;
    layer2_outputs(7991) <= a or b;
    layer2_outputs(7992) <= a or b;
    layer2_outputs(7993) <= not a;
    layer2_outputs(7994) <= a or b;
    layer2_outputs(7995) <= 1'b1;
    layer2_outputs(7996) <= a and b;
    layer2_outputs(7997) <= a;
    layer2_outputs(7998) <= b and not a;
    layer2_outputs(7999) <= a;
    layer2_outputs(8000) <= not a;
    layer2_outputs(8001) <= not b or a;
    layer2_outputs(8002) <= 1'b1;
    layer2_outputs(8003) <= b;
    layer2_outputs(8004) <= b;
    layer2_outputs(8005) <= not a or b;
    layer2_outputs(8006) <= not (a xor b);
    layer2_outputs(8007) <= a;
    layer2_outputs(8008) <= b;
    layer2_outputs(8009) <= not (a or b);
    layer2_outputs(8010) <= a and b;
    layer2_outputs(8011) <= not (a and b);
    layer2_outputs(8012) <= a and b;
    layer2_outputs(8013) <= b and not a;
    layer2_outputs(8014) <= not b or a;
    layer2_outputs(8015) <= 1'b0;
    layer2_outputs(8016) <= b;
    layer2_outputs(8017) <= 1'b1;
    layer2_outputs(8018) <= not b or a;
    layer2_outputs(8019) <= a;
    layer2_outputs(8020) <= not a or b;
    layer2_outputs(8021) <= 1'b0;
    layer2_outputs(8022) <= not b;
    layer2_outputs(8023) <= a or b;
    layer2_outputs(8024) <= not (a or b);
    layer2_outputs(8025) <= a and not b;
    layer2_outputs(8026) <= 1'b0;
    layer2_outputs(8027) <= 1'b1;
    layer2_outputs(8028) <= not (a or b);
    layer2_outputs(8029) <= a and b;
    layer2_outputs(8030) <= not b;
    layer2_outputs(8031) <= b and not a;
    layer2_outputs(8032) <= b and not a;
    layer2_outputs(8033) <= a or b;
    layer2_outputs(8034) <= b;
    layer2_outputs(8035) <= b and not a;
    layer2_outputs(8036) <= not a or b;
    layer2_outputs(8037) <= b and not a;
    layer2_outputs(8038) <= not b;
    layer2_outputs(8039) <= not (a or b);
    layer2_outputs(8040) <= not (a or b);
    layer2_outputs(8041) <= a and b;
    layer2_outputs(8042) <= 1'b0;
    layer2_outputs(8043) <= b and not a;
    layer2_outputs(8044) <= a and b;
    layer2_outputs(8045) <= 1'b0;
    layer2_outputs(8046) <= not (a or b);
    layer2_outputs(8047) <= not a or b;
    layer2_outputs(8048) <= 1'b1;
    layer2_outputs(8049) <= b;
    layer2_outputs(8050) <= a;
    layer2_outputs(8051) <= a and not b;
    layer2_outputs(8052) <= b and not a;
    layer2_outputs(8053) <= not (a or b);
    layer2_outputs(8054) <= a or b;
    layer2_outputs(8055) <= not (a and b);
    layer2_outputs(8056) <= not b;
    layer2_outputs(8057) <= a or b;
    layer2_outputs(8058) <= a or b;
    layer2_outputs(8059) <= not b;
    layer2_outputs(8060) <= 1'b1;
    layer2_outputs(8061) <= not a or b;
    layer2_outputs(8062) <= not b or a;
    layer2_outputs(8063) <= 1'b1;
    layer2_outputs(8064) <= a and not b;
    layer2_outputs(8065) <= b and not a;
    layer2_outputs(8066) <= 1'b0;
    layer2_outputs(8067) <= a or b;
    layer2_outputs(8068) <= 1'b0;
    layer2_outputs(8069) <= b;
    layer2_outputs(8070) <= not b;
    layer2_outputs(8071) <= a or b;
    layer2_outputs(8072) <= not (a and b);
    layer2_outputs(8073) <= a xor b;
    layer2_outputs(8074) <= a and b;
    layer2_outputs(8075) <= b and not a;
    layer2_outputs(8076) <= 1'b0;
    layer2_outputs(8077) <= b;
    layer2_outputs(8078) <= not b or a;
    layer2_outputs(8079) <= a;
    layer2_outputs(8080) <= not b;
    layer2_outputs(8081) <= not (a and b);
    layer2_outputs(8082) <= a and b;
    layer2_outputs(8083) <= b and not a;
    layer2_outputs(8084) <= b and not a;
    layer2_outputs(8085) <= a or b;
    layer2_outputs(8086) <= 1'b0;
    layer2_outputs(8087) <= not (a or b);
    layer2_outputs(8088) <= not b;
    layer2_outputs(8089) <= a or b;
    layer2_outputs(8090) <= not b;
    layer2_outputs(8091) <= not b;
    layer2_outputs(8092) <= not a or b;
    layer2_outputs(8093) <= a;
    layer2_outputs(8094) <= not a;
    layer2_outputs(8095) <= a;
    layer2_outputs(8096) <= a and b;
    layer2_outputs(8097) <= a and b;
    layer2_outputs(8098) <= not a;
    layer2_outputs(8099) <= a and b;
    layer2_outputs(8100) <= a and b;
    layer2_outputs(8101) <= not (a and b);
    layer2_outputs(8102) <= b and not a;
    layer2_outputs(8103) <= a;
    layer2_outputs(8104) <= not (a and b);
    layer2_outputs(8105) <= b and not a;
    layer2_outputs(8106) <= a and b;
    layer2_outputs(8107) <= 1'b1;
    layer2_outputs(8108) <= a and not b;
    layer2_outputs(8109) <= a and not b;
    layer2_outputs(8110) <= 1'b1;
    layer2_outputs(8111) <= b and not a;
    layer2_outputs(8112) <= 1'b1;
    layer2_outputs(8113) <= not b;
    layer2_outputs(8114) <= not (a and b);
    layer2_outputs(8115) <= b;
    layer2_outputs(8116) <= b;
    layer2_outputs(8117) <= a or b;
    layer2_outputs(8118) <= 1'b1;
    layer2_outputs(8119) <= not b or a;
    layer2_outputs(8120) <= a and b;
    layer2_outputs(8121) <= not (a and b);
    layer2_outputs(8122) <= not b;
    layer2_outputs(8123) <= b and not a;
    layer2_outputs(8124) <= 1'b1;
    layer2_outputs(8125) <= not b;
    layer2_outputs(8126) <= not (a or b);
    layer2_outputs(8127) <= a and not b;
    layer2_outputs(8128) <= a;
    layer2_outputs(8129) <= a xor b;
    layer2_outputs(8130) <= not (a or b);
    layer2_outputs(8131) <= a and b;
    layer2_outputs(8132) <= not (a and b);
    layer2_outputs(8133) <= a;
    layer2_outputs(8134) <= not (a and b);
    layer2_outputs(8135) <= not (a xor b);
    layer2_outputs(8136) <= a;
    layer2_outputs(8137) <= a and b;
    layer2_outputs(8138) <= 1'b1;
    layer2_outputs(8139) <= a;
    layer2_outputs(8140) <= not a or b;
    layer2_outputs(8141) <= not b;
    layer2_outputs(8142) <= 1'b1;
    layer2_outputs(8143) <= b;
    layer2_outputs(8144) <= not (a or b);
    layer2_outputs(8145) <= not a;
    layer2_outputs(8146) <= not a or b;
    layer2_outputs(8147) <= 1'b1;
    layer2_outputs(8148) <= not (a and b);
    layer2_outputs(8149) <= b;
    layer2_outputs(8150) <= a;
    layer2_outputs(8151) <= not (a or b);
    layer2_outputs(8152) <= not (a and b);
    layer2_outputs(8153) <= b and not a;
    layer2_outputs(8154) <= a and not b;
    layer2_outputs(8155) <= 1'b1;
    layer2_outputs(8156) <= not b or a;
    layer2_outputs(8157) <= b and not a;
    layer2_outputs(8158) <= not b;
    layer2_outputs(8159) <= a and not b;
    layer2_outputs(8160) <= b and not a;
    layer2_outputs(8161) <= 1'b1;
    layer2_outputs(8162) <= not (a or b);
    layer2_outputs(8163) <= a or b;
    layer2_outputs(8164) <= not b;
    layer2_outputs(8165) <= 1'b0;
    layer2_outputs(8166) <= a and not b;
    layer2_outputs(8167) <= not (a and b);
    layer2_outputs(8168) <= not b;
    layer2_outputs(8169) <= not b;
    layer2_outputs(8170) <= a xor b;
    layer2_outputs(8171) <= a or b;
    layer2_outputs(8172) <= a and not b;
    layer2_outputs(8173) <= b;
    layer2_outputs(8174) <= a or b;
    layer2_outputs(8175) <= a and b;
    layer2_outputs(8176) <= 1'b1;
    layer2_outputs(8177) <= not a or b;
    layer2_outputs(8178) <= not a;
    layer2_outputs(8179) <= 1'b0;
    layer2_outputs(8180) <= not b;
    layer2_outputs(8181) <= a and not b;
    layer2_outputs(8182) <= not a or b;
    layer2_outputs(8183) <= not b;
    layer2_outputs(8184) <= a or b;
    layer2_outputs(8185) <= 1'b0;
    layer2_outputs(8186) <= not b or a;
    layer2_outputs(8187) <= 1'b0;
    layer2_outputs(8188) <= not (a or b);
    layer2_outputs(8189) <= not (a xor b);
    layer2_outputs(8190) <= a and b;
    layer2_outputs(8191) <= a or b;
    layer2_outputs(8192) <= not a or b;
    layer2_outputs(8193) <= a and b;
    layer2_outputs(8194) <= not a or b;
    layer2_outputs(8195) <= not a or b;
    layer2_outputs(8196) <= b;
    layer2_outputs(8197) <= a and not b;
    layer2_outputs(8198) <= not b or a;
    layer2_outputs(8199) <= not (a xor b);
    layer2_outputs(8200) <= not a or b;
    layer2_outputs(8201) <= a and b;
    layer2_outputs(8202) <= b;
    layer2_outputs(8203) <= not b;
    layer2_outputs(8204) <= not a or b;
    layer2_outputs(8205) <= b;
    layer2_outputs(8206) <= b and not a;
    layer2_outputs(8207) <= a and b;
    layer2_outputs(8208) <= 1'b0;
    layer2_outputs(8209) <= not b;
    layer2_outputs(8210) <= a and b;
    layer2_outputs(8211) <= not (a and b);
    layer2_outputs(8212) <= not (a xor b);
    layer2_outputs(8213) <= 1'b0;
    layer2_outputs(8214) <= not (a or b);
    layer2_outputs(8215) <= a and b;
    layer2_outputs(8216) <= 1'b1;
    layer2_outputs(8217) <= 1'b1;
    layer2_outputs(8218) <= a and b;
    layer2_outputs(8219) <= b and not a;
    layer2_outputs(8220) <= not a or b;
    layer2_outputs(8221) <= 1'b0;
    layer2_outputs(8222) <= a and b;
    layer2_outputs(8223) <= 1'b1;
    layer2_outputs(8224) <= a or b;
    layer2_outputs(8225) <= not (a xor b);
    layer2_outputs(8226) <= a and b;
    layer2_outputs(8227) <= not b;
    layer2_outputs(8228) <= b;
    layer2_outputs(8229) <= b and not a;
    layer2_outputs(8230) <= a;
    layer2_outputs(8231) <= 1'b1;
    layer2_outputs(8232) <= not a or b;
    layer2_outputs(8233) <= 1'b0;
    layer2_outputs(8234) <= not (a and b);
    layer2_outputs(8235) <= not a;
    layer2_outputs(8236) <= b;
    layer2_outputs(8237) <= not b;
    layer2_outputs(8238) <= not a or b;
    layer2_outputs(8239) <= b;
    layer2_outputs(8240) <= 1'b0;
    layer2_outputs(8241) <= a;
    layer2_outputs(8242) <= not b or a;
    layer2_outputs(8243) <= a and not b;
    layer2_outputs(8244) <= 1'b1;
    layer2_outputs(8245) <= not b or a;
    layer2_outputs(8246) <= a and not b;
    layer2_outputs(8247) <= not b or a;
    layer2_outputs(8248) <= b and not a;
    layer2_outputs(8249) <= a and b;
    layer2_outputs(8250) <= not (a xor b);
    layer2_outputs(8251) <= a and not b;
    layer2_outputs(8252) <= not (a or b);
    layer2_outputs(8253) <= not (a and b);
    layer2_outputs(8254) <= 1'b1;
    layer2_outputs(8255) <= 1'b0;
    layer2_outputs(8256) <= 1'b0;
    layer2_outputs(8257) <= not b;
    layer2_outputs(8258) <= a or b;
    layer2_outputs(8259) <= not a or b;
    layer2_outputs(8260) <= not b;
    layer2_outputs(8261) <= not b;
    layer2_outputs(8262) <= not a or b;
    layer2_outputs(8263) <= not (a xor b);
    layer2_outputs(8264) <= not a or b;
    layer2_outputs(8265) <= b;
    layer2_outputs(8266) <= 1'b0;
    layer2_outputs(8267) <= b;
    layer2_outputs(8268) <= not b;
    layer2_outputs(8269) <= not b or a;
    layer2_outputs(8270) <= a and b;
    layer2_outputs(8271) <= 1'b1;
    layer2_outputs(8272) <= a and b;
    layer2_outputs(8273) <= not b;
    layer2_outputs(8274) <= a and not b;
    layer2_outputs(8275) <= a or b;
    layer2_outputs(8276) <= not (a or b);
    layer2_outputs(8277) <= not b;
    layer2_outputs(8278) <= a or b;
    layer2_outputs(8279) <= a and not b;
    layer2_outputs(8280) <= b and not a;
    layer2_outputs(8281) <= not a;
    layer2_outputs(8282) <= not (a or b);
    layer2_outputs(8283) <= not b;
    layer2_outputs(8284) <= not (a xor b);
    layer2_outputs(8285) <= not (a xor b);
    layer2_outputs(8286) <= not (a or b);
    layer2_outputs(8287) <= 1'b0;
    layer2_outputs(8288) <= 1'b0;
    layer2_outputs(8289) <= not a;
    layer2_outputs(8290) <= not a or b;
    layer2_outputs(8291) <= a or b;
    layer2_outputs(8292) <= not b;
    layer2_outputs(8293) <= not (a xor b);
    layer2_outputs(8294) <= 1'b0;
    layer2_outputs(8295) <= not (a and b);
    layer2_outputs(8296) <= not (a and b);
    layer2_outputs(8297) <= a and b;
    layer2_outputs(8298) <= b and not a;
    layer2_outputs(8299) <= 1'b0;
    layer2_outputs(8300) <= 1'b0;
    layer2_outputs(8301) <= b;
    layer2_outputs(8302) <= a or b;
    layer2_outputs(8303) <= 1'b1;
    layer2_outputs(8304) <= not a or b;
    layer2_outputs(8305) <= 1'b1;
    layer2_outputs(8306) <= b;
    layer2_outputs(8307) <= b and not a;
    layer2_outputs(8308) <= a and b;
    layer2_outputs(8309) <= 1'b1;
    layer2_outputs(8310) <= 1'b1;
    layer2_outputs(8311) <= b;
    layer2_outputs(8312) <= not b or a;
    layer2_outputs(8313) <= a or b;
    layer2_outputs(8314) <= not a;
    layer2_outputs(8315) <= b and not a;
    layer2_outputs(8316) <= not a or b;
    layer2_outputs(8317) <= b and not a;
    layer2_outputs(8318) <= a and b;
    layer2_outputs(8319) <= a or b;
    layer2_outputs(8320) <= not a;
    layer2_outputs(8321) <= 1'b0;
    layer2_outputs(8322) <= b and not a;
    layer2_outputs(8323) <= a and b;
    layer2_outputs(8324) <= a;
    layer2_outputs(8325) <= 1'b1;
    layer2_outputs(8326) <= a or b;
    layer2_outputs(8327) <= not (a or b);
    layer2_outputs(8328) <= 1'b1;
    layer2_outputs(8329) <= 1'b1;
    layer2_outputs(8330) <= a or b;
    layer2_outputs(8331) <= not b;
    layer2_outputs(8332) <= a xor b;
    layer2_outputs(8333) <= 1'b1;
    layer2_outputs(8334) <= a;
    layer2_outputs(8335) <= 1'b1;
    layer2_outputs(8336) <= 1'b0;
    layer2_outputs(8337) <= a xor b;
    layer2_outputs(8338) <= not a or b;
    layer2_outputs(8339) <= a and b;
    layer2_outputs(8340) <= not a or b;
    layer2_outputs(8341) <= not b or a;
    layer2_outputs(8342) <= not b;
    layer2_outputs(8343) <= 1'b1;
    layer2_outputs(8344) <= a;
    layer2_outputs(8345) <= b;
    layer2_outputs(8346) <= b and not a;
    layer2_outputs(8347) <= not a;
    layer2_outputs(8348) <= 1'b1;
    layer2_outputs(8349) <= not (a or b);
    layer2_outputs(8350) <= 1'b0;
    layer2_outputs(8351) <= 1'b1;
    layer2_outputs(8352) <= not b or a;
    layer2_outputs(8353) <= b and not a;
    layer2_outputs(8354) <= b;
    layer2_outputs(8355) <= a and not b;
    layer2_outputs(8356) <= 1'b1;
    layer2_outputs(8357) <= a;
    layer2_outputs(8358) <= not (a and b);
    layer2_outputs(8359) <= 1'b1;
    layer2_outputs(8360) <= not (a xor b);
    layer2_outputs(8361) <= not b;
    layer2_outputs(8362) <= not b;
    layer2_outputs(8363) <= 1'b1;
    layer2_outputs(8364) <= b;
    layer2_outputs(8365) <= not b;
    layer2_outputs(8366) <= a;
    layer2_outputs(8367) <= 1'b0;
    layer2_outputs(8368) <= not a or b;
    layer2_outputs(8369) <= not (a or b);
    layer2_outputs(8370) <= not a or b;
    layer2_outputs(8371) <= a and not b;
    layer2_outputs(8372) <= 1'b0;
    layer2_outputs(8373) <= not a or b;
    layer2_outputs(8374) <= not a or b;
    layer2_outputs(8375) <= 1'b1;
    layer2_outputs(8376) <= not a;
    layer2_outputs(8377) <= 1'b1;
    layer2_outputs(8378) <= not (a xor b);
    layer2_outputs(8379) <= a and b;
    layer2_outputs(8380) <= a and not b;
    layer2_outputs(8381) <= not (a or b);
    layer2_outputs(8382) <= not (a and b);
    layer2_outputs(8383) <= not b;
    layer2_outputs(8384) <= a and b;
    layer2_outputs(8385) <= a and not b;
    layer2_outputs(8386) <= not b;
    layer2_outputs(8387) <= b and not a;
    layer2_outputs(8388) <= a and not b;
    layer2_outputs(8389) <= a or b;
    layer2_outputs(8390) <= a and b;
    layer2_outputs(8391) <= a;
    layer2_outputs(8392) <= not a or b;
    layer2_outputs(8393) <= a;
    layer2_outputs(8394) <= not b or a;
    layer2_outputs(8395) <= b and not a;
    layer2_outputs(8396) <= not b;
    layer2_outputs(8397) <= not b;
    layer2_outputs(8398) <= not (a and b);
    layer2_outputs(8399) <= not (a or b);
    layer2_outputs(8400) <= not (a or b);
    layer2_outputs(8401) <= b and not a;
    layer2_outputs(8402) <= 1'b1;
    layer2_outputs(8403) <= a and not b;
    layer2_outputs(8404) <= not b or a;
    layer2_outputs(8405) <= a or b;
    layer2_outputs(8406) <= not (a or b);
    layer2_outputs(8407) <= not b;
    layer2_outputs(8408) <= not b or a;
    layer2_outputs(8409) <= not b;
    layer2_outputs(8410) <= not b or a;
    layer2_outputs(8411) <= a and not b;
    layer2_outputs(8412) <= not b or a;
    layer2_outputs(8413) <= a and b;
    layer2_outputs(8414) <= b and not a;
    layer2_outputs(8415) <= not b or a;
    layer2_outputs(8416) <= not b or a;
    layer2_outputs(8417) <= not a or b;
    layer2_outputs(8418) <= not a;
    layer2_outputs(8419) <= a or b;
    layer2_outputs(8420) <= not (a or b);
    layer2_outputs(8421) <= b and not a;
    layer2_outputs(8422) <= b;
    layer2_outputs(8423) <= not b or a;
    layer2_outputs(8424) <= not (a or b);
    layer2_outputs(8425) <= 1'b1;
    layer2_outputs(8426) <= 1'b1;
    layer2_outputs(8427) <= a or b;
    layer2_outputs(8428) <= a and not b;
    layer2_outputs(8429) <= not b;
    layer2_outputs(8430) <= not a;
    layer2_outputs(8431) <= b and not a;
    layer2_outputs(8432) <= a and not b;
    layer2_outputs(8433) <= a or b;
    layer2_outputs(8434) <= not a or b;
    layer2_outputs(8435) <= a and not b;
    layer2_outputs(8436) <= b and not a;
    layer2_outputs(8437) <= not (a and b);
    layer2_outputs(8438) <= not a;
    layer2_outputs(8439) <= a and b;
    layer2_outputs(8440) <= not (a and b);
    layer2_outputs(8441) <= not a;
    layer2_outputs(8442) <= b and not a;
    layer2_outputs(8443) <= a and b;
    layer2_outputs(8444) <= not (a and b);
    layer2_outputs(8445) <= a or b;
    layer2_outputs(8446) <= a and b;
    layer2_outputs(8447) <= a or b;
    layer2_outputs(8448) <= a;
    layer2_outputs(8449) <= not (a and b);
    layer2_outputs(8450) <= not b;
    layer2_outputs(8451) <= 1'b0;
    layer2_outputs(8452) <= a xor b;
    layer2_outputs(8453) <= not a;
    layer2_outputs(8454) <= 1'b1;
    layer2_outputs(8455) <= 1'b1;
    layer2_outputs(8456) <= a and b;
    layer2_outputs(8457) <= not (a and b);
    layer2_outputs(8458) <= not (a or b);
    layer2_outputs(8459) <= b and not a;
    layer2_outputs(8460) <= not (a or b);
    layer2_outputs(8461) <= not b or a;
    layer2_outputs(8462) <= b;
    layer2_outputs(8463) <= not b;
    layer2_outputs(8464) <= 1'b0;
    layer2_outputs(8465) <= 1'b1;
    layer2_outputs(8466) <= 1'b1;
    layer2_outputs(8467) <= b and not a;
    layer2_outputs(8468) <= 1'b1;
    layer2_outputs(8469) <= a and b;
    layer2_outputs(8470) <= not b or a;
    layer2_outputs(8471) <= a or b;
    layer2_outputs(8472) <= not b;
    layer2_outputs(8473) <= not (a and b);
    layer2_outputs(8474) <= 1'b1;
    layer2_outputs(8475) <= a and not b;
    layer2_outputs(8476) <= not b or a;
    layer2_outputs(8477) <= not a;
    layer2_outputs(8478) <= 1'b1;
    layer2_outputs(8479) <= a;
    layer2_outputs(8480) <= not b or a;
    layer2_outputs(8481) <= a;
    layer2_outputs(8482) <= a and b;
    layer2_outputs(8483) <= 1'b0;
    layer2_outputs(8484) <= a;
    layer2_outputs(8485) <= 1'b0;
    layer2_outputs(8486) <= 1'b1;
    layer2_outputs(8487) <= b;
    layer2_outputs(8488) <= a;
    layer2_outputs(8489) <= a and b;
    layer2_outputs(8490) <= not a;
    layer2_outputs(8491) <= b;
    layer2_outputs(8492) <= not b;
    layer2_outputs(8493) <= a and not b;
    layer2_outputs(8494) <= b and not a;
    layer2_outputs(8495) <= not b;
    layer2_outputs(8496) <= not a;
    layer2_outputs(8497) <= not b;
    layer2_outputs(8498) <= 1'b0;
    layer2_outputs(8499) <= a and b;
    layer2_outputs(8500) <= not (a xor b);
    layer2_outputs(8501) <= a and not b;
    layer2_outputs(8502) <= 1'b0;
    layer2_outputs(8503) <= not b or a;
    layer2_outputs(8504) <= not a or b;
    layer2_outputs(8505) <= 1'b0;
    layer2_outputs(8506) <= a;
    layer2_outputs(8507) <= not (a or b);
    layer2_outputs(8508) <= not (a or b);
    layer2_outputs(8509) <= not (a and b);
    layer2_outputs(8510) <= not (a and b);
    layer2_outputs(8511) <= not (a xor b);
    layer2_outputs(8512) <= a and b;
    layer2_outputs(8513) <= not b;
    layer2_outputs(8514) <= not b;
    layer2_outputs(8515) <= not b or a;
    layer2_outputs(8516) <= not a;
    layer2_outputs(8517) <= a or b;
    layer2_outputs(8518) <= a or b;
    layer2_outputs(8519) <= b;
    layer2_outputs(8520) <= not (a and b);
    layer2_outputs(8521) <= not b or a;
    layer2_outputs(8522) <= not b;
    layer2_outputs(8523) <= b;
    layer2_outputs(8524) <= not (a or b);
    layer2_outputs(8525) <= b and not a;
    layer2_outputs(8526) <= a and b;
    layer2_outputs(8527) <= not a;
    layer2_outputs(8528) <= not a or b;
    layer2_outputs(8529) <= not a;
    layer2_outputs(8530) <= a or b;
    layer2_outputs(8531) <= a or b;
    layer2_outputs(8532) <= a and not b;
    layer2_outputs(8533) <= a or b;
    layer2_outputs(8534) <= not (a or b);
    layer2_outputs(8535) <= a and b;
    layer2_outputs(8536) <= a;
    layer2_outputs(8537) <= a;
    layer2_outputs(8538) <= a and not b;
    layer2_outputs(8539) <= b and not a;
    layer2_outputs(8540) <= not b or a;
    layer2_outputs(8541) <= not (a or b);
    layer2_outputs(8542) <= a xor b;
    layer2_outputs(8543) <= a and not b;
    layer2_outputs(8544) <= 1'b0;
    layer2_outputs(8545) <= 1'b1;
    layer2_outputs(8546) <= b;
    layer2_outputs(8547) <= a xor b;
    layer2_outputs(8548) <= a;
    layer2_outputs(8549) <= not b or a;
    layer2_outputs(8550) <= not a or b;
    layer2_outputs(8551) <= not b or a;
    layer2_outputs(8552) <= a or b;
    layer2_outputs(8553) <= not a;
    layer2_outputs(8554) <= not (a and b);
    layer2_outputs(8555) <= not a or b;
    layer2_outputs(8556) <= b;
    layer2_outputs(8557) <= 1'b0;
    layer2_outputs(8558) <= a xor b;
    layer2_outputs(8559) <= not (a or b);
    layer2_outputs(8560) <= 1'b1;
    layer2_outputs(8561) <= a and b;
    layer2_outputs(8562) <= not (a and b);
    layer2_outputs(8563) <= a and b;
    layer2_outputs(8564) <= b and not a;
    layer2_outputs(8565) <= a;
    layer2_outputs(8566) <= not (a xor b);
    layer2_outputs(8567) <= not (a and b);
    layer2_outputs(8568) <= a or b;
    layer2_outputs(8569) <= not a or b;
    layer2_outputs(8570) <= a and b;
    layer2_outputs(8571) <= a and b;
    layer2_outputs(8572) <= 1'b0;
    layer2_outputs(8573) <= not (a and b);
    layer2_outputs(8574) <= 1'b1;
    layer2_outputs(8575) <= 1'b0;
    layer2_outputs(8576) <= not a;
    layer2_outputs(8577) <= not (a and b);
    layer2_outputs(8578) <= a and b;
    layer2_outputs(8579) <= not b or a;
    layer2_outputs(8580) <= a and b;
    layer2_outputs(8581) <= 1'b0;
    layer2_outputs(8582) <= a and b;
    layer2_outputs(8583) <= a xor b;
    layer2_outputs(8584) <= not (a and b);
    layer2_outputs(8585) <= not b or a;
    layer2_outputs(8586) <= not a;
    layer2_outputs(8587) <= 1'b0;
    layer2_outputs(8588) <= 1'b1;
    layer2_outputs(8589) <= not (a or b);
    layer2_outputs(8590) <= a and not b;
    layer2_outputs(8591) <= a and not b;
    layer2_outputs(8592) <= not (a or b);
    layer2_outputs(8593) <= 1'b0;
    layer2_outputs(8594) <= not a;
    layer2_outputs(8595) <= a or b;
    layer2_outputs(8596) <= a and not b;
    layer2_outputs(8597) <= b and not a;
    layer2_outputs(8598) <= not a or b;
    layer2_outputs(8599) <= not b or a;
    layer2_outputs(8600) <= not (a and b);
    layer2_outputs(8601) <= a and b;
    layer2_outputs(8602) <= b and not a;
    layer2_outputs(8603) <= a and not b;
    layer2_outputs(8604) <= a or b;
    layer2_outputs(8605) <= not b;
    layer2_outputs(8606) <= not (a and b);
    layer2_outputs(8607) <= 1'b0;
    layer2_outputs(8608) <= not b or a;
    layer2_outputs(8609) <= a and b;
    layer2_outputs(8610) <= b;
    layer2_outputs(8611) <= not b;
    layer2_outputs(8612) <= b and not a;
    layer2_outputs(8613) <= a or b;
    layer2_outputs(8614) <= a or b;
    layer2_outputs(8615) <= 1'b1;
    layer2_outputs(8616) <= not (a or b);
    layer2_outputs(8617) <= b;
    layer2_outputs(8618) <= 1'b0;
    layer2_outputs(8619) <= 1'b0;
    layer2_outputs(8620) <= a;
    layer2_outputs(8621) <= not (a or b);
    layer2_outputs(8622) <= not (a or b);
    layer2_outputs(8623) <= b and not a;
    layer2_outputs(8624) <= a xor b;
    layer2_outputs(8625) <= b and not a;
    layer2_outputs(8626) <= a and b;
    layer2_outputs(8627) <= not a or b;
    layer2_outputs(8628) <= not (a and b);
    layer2_outputs(8629) <= b and not a;
    layer2_outputs(8630) <= not b or a;
    layer2_outputs(8631) <= b and not a;
    layer2_outputs(8632) <= not a;
    layer2_outputs(8633) <= a and b;
    layer2_outputs(8634) <= 1'b0;
    layer2_outputs(8635) <= a and not b;
    layer2_outputs(8636) <= not (a or b);
    layer2_outputs(8637) <= a;
    layer2_outputs(8638) <= not b or a;
    layer2_outputs(8639) <= 1'b1;
    layer2_outputs(8640) <= 1'b1;
    layer2_outputs(8641) <= not (a xor b);
    layer2_outputs(8642) <= a and not b;
    layer2_outputs(8643) <= not a or b;
    layer2_outputs(8644) <= 1'b0;
    layer2_outputs(8645) <= not (a and b);
    layer2_outputs(8646) <= a;
    layer2_outputs(8647) <= a;
    layer2_outputs(8648) <= a;
    layer2_outputs(8649) <= not b;
    layer2_outputs(8650) <= not b or a;
    layer2_outputs(8651) <= b and not a;
    layer2_outputs(8652) <= not a or b;
    layer2_outputs(8653) <= not (a and b);
    layer2_outputs(8654) <= not (a and b);
    layer2_outputs(8655) <= not (a xor b);
    layer2_outputs(8656) <= a and b;
    layer2_outputs(8657) <= not (a and b);
    layer2_outputs(8658) <= not a;
    layer2_outputs(8659) <= b and not a;
    layer2_outputs(8660) <= a or b;
    layer2_outputs(8661) <= not (a xor b);
    layer2_outputs(8662) <= 1'b0;
    layer2_outputs(8663) <= not b or a;
    layer2_outputs(8664) <= a xor b;
    layer2_outputs(8665) <= not b or a;
    layer2_outputs(8666) <= 1'b1;
    layer2_outputs(8667) <= 1'b1;
    layer2_outputs(8668) <= not (a xor b);
    layer2_outputs(8669) <= 1'b1;
    layer2_outputs(8670) <= 1'b0;
    layer2_outputs(8671) <= a;
    layer2_outputs(8672) <= a;
    layer2_outputs(8673) <= not (a or b);
    layer2_outputs(8674) <= b and not a;
    layer2_outputs(8675) <= 1'b1;
    layer2_outputs(8676) <= a and not b;
    layer2_outputs(8677) <= not a or b;
    layer2_outputs(8678) <= 1'b1;
    layer2_outputs(8679) <= not (a and b);
    layer2_outputs(8680) <= not (a or b);
    layer2_outputs(8681) <= a and not b;
    layer2_outputs(8682) <= a and b;
    layer2_outputs(8683) <= 1'b0;
    layer2_outputs(8684) <= not (a xor b);
    layer2_outputs(8685) <= b;
    layer2_outputs(8686) <= not (a and b);
    layer2_outputs(8687) <= not b or a;
    layer2_outputs(8688) <= not (a and b);
    layer2_outputs(8689) <= b;
    layer2_outputs(8690) <= not b;
    layer2_outputs(8691) <= not b;
    layer2_outputs(8692) <= 1'b1;
    layer2_outputs(8693) <= a or b;
    layer2_outputs(8694) <= not a;
    layer2_outputs(8695) <= not a;
    layer2_outputs(8696) <= b and not a;
    layer2_outputs(8697) <= 1'b1;
    layer2_outputs(8698) <= a;
    layer2_outputs(8699) <= not (a or b);
    layer2_outputs(8700) <= b;
    layer2_outputs(8701) <= not b or a;
    layer2_outputs(8702) <= not b;
    layer2_outputs(8703) <= a and not b;
    layer2_outputs(8704) <= 1'b0;
    layer2_outputs(8705) <= b and not a;
    layer2_outputs(8706) <= not b or a;
    layer2_outputs(8707) <= 1'b1;
    layer2_outputs(8708) <= 1'b0;
    layer2_outputs(8709) <= not b;
    layer2_outputs(8710) <= a or b;
    layer2_outputs(8711) <= not (a and b);
    layer2_outputs(8712) <= not a or b;
    layer2_outputs(8713) <= not b or a;
    layer2_outputs(8714) <= not b;
    layer2_outputs(8715) <= a and not b;
    layer2_outputs(8716) <= 1'b0;
    layer2_outputs(8717) <= a and b;
    layer2_outputs(8718) <= not a;
    layer2_outputs(8719) <= b and not a;
    layer2_outputs(8720) <= 1'b0;
    layer2_outputs(8721) <= not b;
    layer2_outputs(8722) <= 1'b0;
    layer2_outputs(8723) <= b;
    layer2_outputs(8724) <= a and not b;
    layer2_outputs(8725) <= not (a and b);
    layer2_outputs(8726) <= a and b;
    layer2_outputs(8727) <= 1'b1;
    layer2_outputs(8728) <= not a or b;
    layer2_outputs(8729) <= 1'b1;
    layer2_outputs(8730) <= a or b;
    layer2_outputs(8731) <= a and not b;
    layer2_outputs(8732) <= not (a or b);
    layer2_outputs(8733) <= b and not a;
    layer2_outputs(8734) <= not b or a;
    layer2_outputs(8735) <= not (a or b);
    layer2_outputs(8736) <= not a;
    layer2_outputs(8737) <= a;
    layer2_outputs(8738) <= not (a or b);
    layer2_outputs(8739) <= not (a and b);
    layer2_outputs(8740) <= b and not a;
    layer2_outputs(8741) <= a;
    layer2_outputs(8742) <= a;
    layer2_outputs(8743) <= not (a and b);
    layer2_outputs(8744) <= a;
    layer2_outputs(8745) <= b;
    layer2_outputs(8746) <= 1'b0;
    layer2_outputs(8747) <= not a or b;
    layer2_outputs(8748) <= not b;
    layer2_outputs(8749) <= a or b;
    layer2_outputs(8750) <= b;
    layer2_outputs(8751) <= b and not a;
    layer2_outputs(8752) <= a;
    layer2_outputs(8753) <= 1'b0;
    layer2_outputs(8754) <= b and not a;
    layer2_outputs(8755) <= not (a xor b);
    layer2_outputs(8756) <= b;
    layer2_outputs(8757) <= not b or a;
    layer2_outputs(8758) <= a and not b;
    layer2_outputs(8759) <= not (a or b);
    layer2_outputs(8760) <= a and not b;
    layer2_outputs(8761) <= not b or a;
    layer2_outputs(8762) <= not a;
    layer2_outputs(8763) <= not a;
    layer2_outputs(8764) <= b;
    layer2_outputs(8765) <= not a or b;
    layer2_outputs(8766) <= a and b;
    layer2_outputs(8767) <= not b;
    layer2_outputs(8768) <= b and not a;
    layer2_outputs(8769) <= not a;
    layer2_outputs(8770) <= not a;
    layer2_outputs(8771) <= 1'b1;
    layer2_outputs(8772) <= a;
    layer2_outputs(8773) <= not a or b;
    layer2_outputs(8774) <= not a;
    layer2_outputs(8775) <= 1'b1;
    layer2_outputs(8776) <= not (a xor b);
    layer2_outputs(8777) <= 1'b1;
    layer2_outputs(8778) <= b;
    layer2_outputs(8779) <= not a;
    layer2_outputs(8780) <= 1'b0;
    layer2_outputs(8781) <= 1'b1;
    layer2_outputs(8782) <= a and not b;
    layer2_outputs(8783) <= 1'b0;
    layer2_outputs(8784) <= a;
    layer2_outputs(8785) <= 1'b0;
    layer2_outputs(8786) <= b;
    layer2_outputs(8787) <= not b;
    layer2_outputs(8788) <= b and not a;
    layer2_outputs(8789) <= not a or b;
    layer2_outputs(8790) <= not b or a;
    layer2_outputs(8791) <= b and not a;
    layer2_outputs(8792) <= b and not a;
    layer2_outputs(8793) <= 1'b1;
    layer2_outputs(8794) <= b and not a;
    layer2_outputs(8795) <= a and not b;
    layer2_outputs(8796) <= a;
    layer2_outputs(8797) <= not (a xor b);
    layer2_outputs(8798) <= a;
    layer2_outputs(8799) <= not b;
    layer2_outputs(8800) <= b and not a;
    layer2_outputs(8801) <= b and not a;
    layer2_outputs(8802) <= not (a and b);
    layer2_outputs(8803) <= not a;
    layer2_outputs(8804) <= a or b;
    layer2_outputs(8805) <= not b;
    layer2_outputs(8806) <= 1'b1;
    layer2_outputs(8807) <= not (a or b);
    layer2_outputs(8808) <= b and not a;
    layer2_outputs(8809) <= a and not b;
    layer2_outputs(8810) <= 1'b0;
    layer2_outputs(8811) <= not a or b;
    layer2_outputs(8812) <= b;
    layer2_outputs(8813) <= 1'b0;
    layer2_outputs(8814) <= a;
    layer2_outputs(8815) <= a and not b;
    layer2_outputs(8816) <= not b;
    layer2_outputs(8817) <= a or b;
    layer2_outputs(8818) <= not (a and b);
    layer2_outputs(8819) <= not b;
    layer2_outputs(8820) <= a and b;
    layer2_outputs(8821) <= not (a or b);
    layer2_outputs(8822) <= a or b;
    layer2_outputs(8823) <= a;
    layer2_outputs(8824) <= not (a and b);
    layer2_outputs(8825) <= 1'b0;
    layer2_outputs(8826) <= 1'b1;
    layer2_outputs(8827) <= a and not b;
    layer2_outputs(8828) <= not a;
    layer2_outputs(8829) <= not a;
    layer2_outputs(8830) <= a;
    layer2_outputs(8831) <= not b;
    layer2_outputs(8832) <= not b or a;
    layer2_outputs(8833) <= a;
    layer2_outputs(8834) <= not b or a;
    layer2_outputs(8835) <= 1'b0;
    layer2_outputs(8836) <= a or b;
    layer2_outputs(8837) <= not a or b;
    layer2_outputs(8838) <= a and b;
    layer2_outputs(8839) <= a and b;
    layer2_outputs(8840) <= not a or b;
    layer2_outputs(8841) <= not b;
    layer2_outputs(8842) <= a or b;
    layer2_outputs(8843) <= a or b;
    layer2_outputs(8844) <= a or b;
    layer2_outputs(8845) <= a and b;
    layer2_outputs(8846) <= b;
    layer2_outputs(8847) <= 1'b0;
    layer2_outputs(8848) <= b;
    layer2_outputs(8849) <= a and b;
    layer2_outputs(8850) <= 1'b1;
    layer2_outputs(8851) <= not (a and b);
    layer2_outputs(8852) <= not a;
    layer2_outputs(8853) <= a and b;
    layer2_outputs(8854) <= b and not a;
    layer2_outputs(8855) <= not (a or b);
    layer2_outputs(8856) <= not (a and b);
    layer2_outputs(8857) <= not (a xor b);
    layer2_outputs(8858) <= b and not a;
    layer2_outputs(8859) <= not b or a;
    layer2_outputs(8860) <= 1'b1;
    layer2_outputs(8861) <= a and b;
    layer2_outputs(8862) <= a;
    layer2_outputs(8863) <= not b or a;
    layer2_outputs(8864) <= not (a or b);
    layer2_outputs(8865) <= a or b;
    layer2_outputs(8866) <= not b or a;
    layer2_outputs(8867) <= b;
    layer2_outputs(8868) <= b;
    layer2_outputs(8869) <= a and b;
    layer2_outputs(8870) <= not (a and b);
    layer2_outputs(8871) <= not a or b;
    layer2_outputs(8872) <= 1'b1;
    layer2_outputs(8873) <= b;
    layer2_outputs(8874) <= not (a and b);
    layer2_outputs(8875) <= not b;
    layer2_outputs(8876) <= 1'b0;
    layer2_outputs(8877) <= a or b;
    layer2_outputs(8878) <= b and not a;
    layer2_outputs(8879) <= not b;
    layer2_outputs(8880) <= a and b;
    layer2_outputs(8881) <= a and not b;
    layer2_outputs(8882) <= a and not b;
    layer2_outputs(8883) <= not a or b;
    layer2_outputs(8884) <= a;
    layer2_outputs(8885) <= a and not b;
    layer2_outputs(8886) <= a;
    layer2_outputs(8887) <= not a;
    layer2_outputs(8888) <= not (a and b);
    layer2_outputs(8889) <= not b or a;
    layer2_outputs(8890) <= not b or a;
    layer2_outputs(8891) <= not a or b;
    layer2_outputs(8892) <= b and not a;
    layer2_outputs(8893) <= not (a xor b);
    layer2_outputs(8894) <= not b;
    layer2_outputs(8895) <= not (a and b);
    layer2_outputs(8896) <= b and not a;
    layer2_outputs(8897) <= a;
    layer2_outputs(8898) <= b;
    layer2_outputs(8899) <= b and not a;
    layer2_outputs(8900) <= 1'b1;
    layer2_outputs(8901) <= a and not b;
    layer2_outputs(8902) <= not b or a;
    layer2_outputs(8903) <= not a or b;
    layer2_outputs(8904) <= 1'b0;
    layer2_outputs(8905) <= a and not b;
    layer2_outputs(8906) <= not (a or b);
    layer2_outputs(8907) <= a and not b;
    layer2_outputs(8908) <= a and b;
    layer2_outputs(8909) <= not a or b;
    layer2_outputs(8910) <= not (a or b);
    layer2_outputs(8911) <= not b or a;
    layer2_outputs(8912) <= a or b;
    layer2_outputs(8913) <= not b or a;
    layer2_outputs(8914) <= a;
    layer2_outputs(8915) <= not (a or b);
    layer2_outputs(8916) <= 1'b1;
    layer2_outputs(8917) <= not a;
    layer2_outputs(8918) <= a or b;
    layer2_outputs(8919) <= 1'b1;
    layer2_outputs(8920) <= not a;
    layer2_outputs(8921) <= 1'b1;
    layer2_outputs(8922) <= a or b;
    layer2_outputs(8923) <= not a or b;
    layer2_outputs(8924) <= not (a and b);
    layer2_outputs(8925) <= not b or a;
    layer2_outputs(8926) <= a;
    layer2_outputs(8927) <= not b;
    layer2_outputs(8928) <= not (a and b);
    layer2_outputs(8929) <= b;
    layer2_outputs(8930) <= 1'b1;
    layer2_outputs(8931) <= b;
    layer2_outputs(8932) <= a xor b;
    layer2_outputs(8933) <= not (a or b);
    layer2_outputs(8934) <= b;
    layer2_outputs(8935) <= a;
    layer2_outputs(8936) <= not (a and b);
    layer2_outputs(8937) <= not b or a;
    layer2_outputs(8938) <= 1'b0;
    layer2_outputs(8939) <= not (a and b);
    layer2_outputs(8940) <= b;
    layer2_outputs(8941) <= 1'b0;
    layer2_outputs(8942) <= a and not b;
    layer2_outputs(8943) <= b;
    layer2_outputs(8944) <= not (a and b);
    layer2_outputs(8945) <= not a or b;
    layer2_outputs(8946) <= a xor b;
    layer2_outputs(8947) <= 1'b1;
    layer2_outputs(8948) <= not b;
    layer2_outputs(8949) <= a and b;
    layer2_outputs(8950) <= b and not a;
    layer2_outputs(8951) <= not a or b;
    layer2_outputs(8952) <= not a;
    layer2_outputs(8953) <= not b;
    layer2_outputs(8954) <= 1'b1;
    layer2_outputs(8955) <= a or b;
    layer2_outputs(8956) <= 1'b0;
    layer2_outputs(8957) <= b and not a;
    layer2_outputs(8958) <= a and not b;
    layer2_outputs(8959) <= 1'b0;
    layer2_outputs(8960) <= 1'b1;
    layer2_outputs(8961) <= not a or b;
    layer2_outputs(8962) <= 1'b1;
    layer2_outputs(8963) <= not (a or b);
    layer2_outputs(8964) <= a;
    layer2_outputs(8965) <= not a;
    layer2_outputs(8966) <= not b or a;
    layer2_outputs(8967) <= 1'b0;
    layer2_outputs(8968) <= b and not a;
    layer2_outputs(8969) <= not b;
    layer2_outputs(8970) <= not a;
    layer2_outputs(8971) <= a xor b;
    layer2_outputs(8972) <= a and b;
    layer2_outputs(8973) <= a and b;
    layer2_outputs(8974) <= not (a and b);
    layer2_outputs(8975) <= not (a and b);
    layer2_outputs(8976) <= a and not b;
    layer2_outputs(8977) <= not (a and b);
    layer2_outputs(8978) <= a and not b;
    layer2_outputs(8979) <= 1'b1;
    layer2_outputs(8980) <= a;
    layer2_outputs(8981) <= not (a and b);
    layer2_outputs(8982) <= a;
    layer2_outputs(8983) <= not a or b;
    layer2_outputs(8984) <= b;
    layer2_outputs(8985) <= not (a xor b);
    layer2_outputs(8986) <= 1'b1;
    layer2_outputs(8987) <= not (a and b);
    layer2_outputs(8988) <= not b;
    layer2_outputs(8989) <= not (a and b);
    layer2_outputs(8990) <= a xor b;
    layer2_outputs(8991) <= a xor b;
    layer2_outputs(8992) <= not a;
    layer2_outputs(8993) <= a and b;
    layer2_outputs(8994) <= 1'b0;
    layer2_outputs(8995) <= not (a or b);
    layer2_outputs(8996) <= a or b;
    layer2_outputs(8997) <= a and not b;
    layer2_outputs(8998) <= b and not a;
    layer2_outputs(8999) <= b;
    layer2_outputs(9000) <= b;
    layer2_outputs(9001) <= not (a and b);
    layer2_outputs(9002) <= not (a and b);
    layer2_outputs(9003) <= a and not b;
    layer2_outputs(9004) <= not b or a;
    layer2_outputs(9005) <= a and b;
    layer2_outputs(9006) <= 1'b1;
    layer2_outputs(9007) <= a or b;
    layer2_outputs(9008) <= not b;
    layer2_outputs(9009) <= a or b;
    layer2_outputs(9010) <= not b or a;
    layer2_outputs(9011) <= not a or b;
    layer2_outputs(9012) <= a and b;
    layer2_outputs(9013) <= 1'b1;
    layer2_outputs(9014) <= not (a and b);
    layer2_outputs(9015) <= a;
    layer2_outputs(9016) <= not b;
    layer2_outputs(9017) <= 1'b1;
    layer2_outputs(9018) <= a and not b;
    layer2_outputs(9019) <= a and not b;
    layer2_outputs(9020) <= b and not a;
    layer2_outputs(9021) <= b;
    layer2_outputs(9022) <= 1'b0;
    layer2_outputs(9023) <= not b;
    layer2_outputs(9024) <= a and b;
    layer2_outputs(9025) <= not b;
    layer2_outputs(9026) <= a xor b;
    layer2_outputs(9027) <= not b or a;
    layer2_outputs(9028) <= a and not b;
    layer2_outputs(9029) <= b and not a;
    layer2_outputs(9030) <= 1'b0;
    layer2_outputs(9031) <= a and not b;
    layer2_outputs(9032) <= a or b;
    layer2_outputs(9033) <= not a;
    layer2_outputs(9034) <= a or b;
    layer2_outputs(9035) <= 1'b0;
    layer2_outputs(9036) <= not (a and b);
    layer2_outputs(9037) <= a or b;
    layer2_outputs(9038) <= not (a or b);
    layer2_outputs(9039) <= not b;
    layer2_outputs(9040) <= 1'b0;
    layer2_outputs(9041) <= not (a or b);
    layer2_outputs(9042) <= a xor b;
    layer2_outputs(9043) <= a and b;
    layer2_outputs(9044) <= 1'b0;
    layer2_outputs(9045) <= not (a and b);
    layer2_outputs(9046) <= 1'b1;
    layer2_outputs(9047) <= a xor b;
    layer2_outputs(9048) <= not (a and b);
    layer2_outputs(9049) <= b;
    layer2_outputs(9050) <= not a;
    layer2_outputs(9051) <= not (a or b);
    layer2_outputs(9052) <= b and not a;
    layer2_outputs(9053) <= b;
    layer2_outputs(9054) <= 1'b1;
    layer2_outputs(9055) <= a and not b;
    layer2_outputs(9056) <= not (a xor b);
    layer2_outputs(9057) <= a or b;
    layer2_outputs(9058) <= not (a or b);
    layer2_outputs(9059) <= a xor b;
    layer2_outputs(9060) <= not b;
    layer2_outputs(9061) <= a or b;
    layer2_outputs(9062) <= not (a or b);
    layer2_outputs(9063) <= not b or a;
    layer2_outputs(9064) <= a and b;
    layer2_outputs(9065) <= a and b;
    layer2_outputs(9066) <= not (a or b);
    layer2_outputs(9067) <= not (a and b);
    layer2_outputs(9068) <= not b;
    layer2_outputs(9069) <= a and not b;
    layer2_outputs(9070) <= a xor b;
    layer2_outputs(9071) <= not a;
    layer2_outputs(9072) <= b and not a;
    layer2_outputs(9073) <= not (a xor b);
    layer2_outputs(9074) <= not a or b;
    layer2_outputs(9075) <= a;
    layer2_outputs(9076) <= a and not b;
    layer2_outputs(9077) <= not (a and b);
    layer2_outputs(9078) <= not b or a;
    layer2_outputs(9079) <= 1'b0;
    layer2_outputs(9080) <= a and not b;
    layer2_outputs(9081) <= a and not b;
    layer2_outputs(9082) <= a and b;
    layer2_outputs(9083) <= a and not b;
    layer2_outputs(9084) <= b and not a;
    layer2_outputs(9085) <= a or b;
    layer2_outputs(9086) <= a and not b;
    layer2_outputs(9087) <= a;
    layer2_outputs(9088) <= not b;
    layer2_outputs(9089) <= not b or a;
    layer2_outputs(9090) <= not (a and b);
    layer2_outputs(9091) <= not (a and b);
    layer2_outputs(9092) <= 1'b1;
    layer2_outputs(9093) <= a or b;
    layer2_outputs(9094) <= b;
    layer2_outputs(9095) <= not a;
    layer2_outputs(9096) <= b and not a;
    layer2_outputs(9097) <= a;
    layer2_outputs(9098) <= 1'b1;
    layer2_outputs(9099) <= 1'b1;
    layer2_outputs(9100) <= 1'b1;
    layer2_outputs(9101) <= a or b;
    layer2_outputs(9102) <= a xor b;
    layer2_outputs(9103) <= not b;
    layer2_outputs(9104) <= 1'b1;
    layer2_outputs(9105) <= a and b;
    layer2_outputs(9106) <= b;
    layer2_outputs(9107) <= a or b;
    layer2_outputs(9108) <= a or b;
    layer2_outputs(9109) <= not b;
    layer2_outputs(9110) <= 1'b0;
    layer2_outputs(9111) <= not (a or b);
    layer2_outputs(9112) <= a and b;
    layer2_outputs(9113) <= 1'b1;
    layer2_outputs(9114) <= not b or a;
    layer2_outputs(9115) <= not a;
    layer2_outputs(9116) <= a and b;
    layer2_outputs(9117) <= not a;
    layer2_outputs(9118) <= a;
    layer2_outputs(9119) <= a and not b;
    layer2_outputs(9120) <= b and not a;
    layer2_outputs(9121) <= a xor b;
    layer2_outputs(9122) <= not (a or b);
    layer2_outputs(9123) <= a and b;
    layer2_outputs(9124) <= not (a and b);
    layer2_outputs(9125) <= not (a or b);
    layer2_outputs(9126) <= 1'b1;
    layer2_outputs(9127) <= 1'b1;
    layer2_outputs(9128) <= not (a and b);
    layer2_outputs(9129) <= b and not a;
    layer2_outputs(9130) <= 1'b1;
    layer2_outputs(9131) <= a and not b;
    layer2_outputs(9132) <= not a;
    layer2_outputs(9133) <= a and not b;
    layer2_outputs(9134) <= not b or a;
    layer2_outputs(9135) <= a or b;
    layer2_outputs(9136) <= 1'b0;
    layer2_outputs(9137) <= b and not a;
    layer2_outputs(9138) <= a or b;
    layer2_outputs(9139) <= not b or a;
    layer2_outputs(9140) <= 1'b0;
    layer2_outputs(9141) <= 1'b0;
    layer2_outputs(9142) <= not a;
    layer2_outputs(9143) <= a and b;
    layer2_outputs(9144) <= not (a or b);
    layer2_outputs(9145) <= a;
    layer2_outputs(9146) <= not b;
    layer2_outputs(9147) <= 1'b0;
    layer2_outputs(9148) <= 1'b1;
    layer2_outputs(9149) <= not (a and b);
    layer2_outputs(9150) <= a and b;
    layer2_outputs(9151) <= b and not a;
    layer2_outputs(9152) <= not a or b;
    layer2_outputs(9153) <= not a;
    layer2_outputs(9154) <= 1'b1;
    layer2_outputs(9155) <= not (a xor b);
    layer2_outputs(9156) <= b and not a;
    layer2_outputs(9157) <= 1'b1;
    layer2_outputs(9158) <= not a or b;
    layer2_outputs(9159) <= not a or b;
    layer2_outputs(9160) <= a or b;
    layer2_outputs(9161) <= a or b;
    layer2_outputs(9162) <= not (a xor b);
    layer2_outputs(9163) <= not (a or b);
    layer2_outputs(9164) <= not b or a;
    layer2_outputs(9165) <= not b;
    layer2_outputs(9166) <= b;
    layer2_outputs(9167) <= not (a or b);
    layer2_outputs(9168) <= a or b;
    layer2_outputs(9169) <= 1'b0;
    layer2_outputs(9170) <= b and not a;
    layer2_outputs(9171) <= not b or a;
    layer2_outputs(9172) <= a or b;
    layer2_outputs(9173) <= b;
    layer2_outputs(9174) <= a and b;
    layer2_outputs(9175) <= not a or b;
    layer2_outputs(9176) <= not a or b;
    layer2_outputs(9177) <= 1'b0;
    layer2_outputs(9178) <= 1'b1;
    layer2_outputs(9179) <= a and b;
    layer2_outputs(9180) <= b and not a;
    layer2_outputs(9181) <= not a or b;
    layer2_outputs(9182) <= not a;
    layer2_outputs(9183) <= a and b;
    layer2_outputs(9184) <= not (a and b);
    layer2_outputs(9185) <= a or b;
    layer2_outputs(9186) <= not (a and b);
    layer2_outputs(9187) <= a and not b;
    layer2_outputs(9188) <= a or b;
    layer2_outputs(9189) <= b;
    layer2_outputs(9190) <= 1'b1;
    layer2_outputs(9191) <= b;
    layer2_outputs(9192) <= not (a xor b);
    layer2_outputs(9193) <= not b or a;
    layer2_outputs(9194) <= not a or b;
    layer2_outputs(9195) <= not (a or b);
    layer2_outputs(9196) <= not b;
    layer2_outputs(9197) <= not b;
    layer2_outputs(9198) <= not a or b;
    layer2_outputs(9199) <= b and not a;
    layer2_outputs(9200) <= b;
    layer2_outputs(9201) <= a or b;
    layer2_outputs(9202) <= not a or b;
    layer2_outputs(9203) <= not a;
    layer2_outputs(9204) <= b and not a;
    layer2_outputs(9205) <= a;
    layer2_outputs(9206) <= 1'b0;
    layer2_outputs(9207) <= a;
    layer2_outputs(9208) <= a;
    layer2_outputs(9209) <= b;
    layer2_outputs(9210) <= not b or a;
    layer2_outputs(9211) <= a and not b;
    layer2_outputs(9212) <= not b;
    layer2_outputs(9213) <= not a;
    layer2_outputs(9214) <= a or b;
    layer2_outputs(9215) <= not a or b;
    layer2_outputs(9216) <= not (a and b);
    layer2_outputs(9217) <= 1'b1;
    layer2_outputs(9218) <= b;
    layer2_outputs(9219) <= not (a and b);
    layer2_outputs(9220) <= 1'b0;
    layer2_outputs(9221) <= a;
    layer2_outputs(9222) <= 1'b0;
    layer2_outputs(9223) <= a and not b;
    layer2_outputs(9224) <= a and b;
    layer2_outputs(9225) <= 1'b0;
    layer2_outputs(9226) <= 1'b1;
    layer2_outputs(9227) <= not a;
    layer2_outputs(9228) <= 1'b1;
    layer2_outputs(9229) <= a and not b;
    layer2_outputs(9230) <= not a or b;
    layer2_outputs(9231) <= a;
    layer2_outputs(9232) <= not a or b;
    layer2_outputs(9233) <= 1'b0;
    layer2_outputs(9234) <= 1'b1;
    layer2_outputs(9235) <= b;
    layer2_outputs(9236) <= b and not a;
    layer2_outputs(9237) <= b;
    layer2_outputs(9238) <= not b or a;
    layer2_outputs(9239) <= b;
    layer2_outputs(9240) <= a and not b;
    layer2_outputs(9241) <= 1'b1;
    layer2_outputs(9242) <= not a;
    layer2_outputs(9243) <= not a;
    layer2_outputs(9244) <= a;
    layer2_outputs(9245) <= 1'b0;
    layer2_outputs(9246) <= not a or b;
    layer2_outputs(9247) <= a and b;
    layer2_outputs(9248) <= not (a xor b);
    layer2_outputs(9249) <= a or b;
    layer2_outputs(9250) <= a and b;
    layer2_outputs(9251) <= b;
    layer2_outputs(9252) <= not (a and b);
    layer2_outputs(9253) <= not (a and b);
    layer2_outputs(9254) <= a and not b;
    layer2_outputs(9255) <= a and not b;
    layer2_outputs(9256) <= not (a and b);
    layer2_outputs(9257) <= not (a and b);
    layer2_outputs(9258) <= 1'b1;
    layer2_outputs(9259) <= not a;
    layer2_outputs(9260) <= not b or a;
    layer2_outputs(9261) <= a or b;
    layer2_outputs(9262) <= a;
    layer2_outputs(9263) <= not (a and b);
    layer2_outputs(9264) <= not a or b;
    layer2_outputs(9265) <= b and not a;
    layer2_outputs(9266) <= not b;
    layer2_outputs(9267) <= 1'b0;
    layer2_outputs(9268) <= not a;
    layer2_outputs(9269) <= a and not b;
    layer2_outputs(9270) <= b;
    layer2_outputs(9271) <= not (a xor b);
    layer2_outputs(9272) <= a and b;
    layer2_outputs(9273) <= not (a and b);
    layer2_outputs(9274) <= not b;
    layer2_outputs(9275) <= not b;
    layer2_outputs(9276) <= a and not b;
    layer2_outputs(9277) <= not b or a;
    layer2_outputs(9278) <= 1'b0;
    layer2_outputs(9279) <= not b;
    layer2_outputs(9280) <= not a or b;
    layer2_outputs(9281) <= a and b;
    layer2_outputs(9282) <= 1'b1;
    layer2_outputs(9283) <= not (a or b);
    layer2_outputs(9284) <= not b;
    layer2_outputs(9285) <= not b or a;
    layer2_outputs(9286) <= b;
    layer2_outputs(9287) <= 1'b0;
    layer2_outputs(9288) <= b and not a;
    layer2_outputs(9289) <= a or b;
    layer2_outputs(9290) <= not (a and b);
    layer2_outputs(9291) <= not a;
    layer2_outputs(9292) <= b;
    layer2_outputs(9293) <= a and not b;
    layer2_outputs(9294) <= a or b;
    layer2_outputs(9295) <= not (a and b);
    layer2_outputs(9296) <= a;
    layer2_outputs(9297) <= 1'b1;
    layer2_outputs(9298) <= not a or b;
    layer2_outputs(9299) <= not (a or b);
    layer2_outputs(9300) <= not b or a;
    layer2_outputs(9301) <= 1'b0;
    layer2_outputs(9302) <= not (a or b);
    layer2_outputs(9303) <= b and not a;
    layer2_outputs(9304) <= not a or b;
    layer2_outputs(9305) <= b;
    layer2_outputs(9306) <= a and not b;
    layer2_outputs(9307) <= not (a or b);
    layer2_outputs(9308) <= 1'b1;
    layer2_outputs(9309) <= 1'b0;
    layer2_outputs(9310) <= b and not a;
    layer2_outputs(9311) <= not (a or b);
    layer2_outputs(9312) <= not a;
    layer2_outputs(9313) <= a and not b;
    layer2_outputs(9314) <= not b;
    layer2_outputs(9315) <= 1'b1;
    layer2_outputs(9316) <= b and not a;
    layer2_outputs(9317) <= not a;
    layer2_outputs(9318) <= 1'b1;
    layer2_outputs(9319) <= a and b;
    layer2_outputs(9320) <= 1'b1;
    layer2_outputs(9321) <= not a;
    layer2_outputs(9322) <= not a or b;
    layer2_outputs(9323) <= b and not a;
    layer2_outputs(9324) <= a or b;
    layer2_outputs(9325) <= not (a xor b);
    layer2_outputs(9326) <= a or b;
    layer2_outputs(9327) <= a or b;
    layer2_outputs(9328) <= not a or b;
    layer2_outputs(9329) <= 1'b0;
    layer2_outputs(9330) <= not (a or b);
    layer2_outputs(9331) <= not a or b;
    layer2_outputs(9332) <= b and not a;
    layer2_outputs(9333) <= a xor b;
    layer2_outputs(9334) <= a and not b;
    layer2_outputs(9335) <= not b or a;
    layer2_outputs(9336) <= not b;
    layer2_outputs(9337) <= b and not a;
    layer2_outputs(9338) <= a and not b;
    layer2_outputs(9339) <= a;
    layer2_outputs(9340) <= not a or b;
    layer2_outputs(9341) <= not b;
    layer2_outputs(9342) <= a and not b;
    layer2_outputs(9343) <= not (a or b);
    layer2_outputs(9344) <= a and b;
    layer2_outputs(9345) <= not b;
    layer2_outputs(9346) <= not (a and b);
    layer2_outputs(9347) <= a or b;
    layer2_outputs(9348) <= not b;
    layer2_outputs(9349) <= not a;
    layer2_outputs(9350) <= b;
    layer2_outputs(9351) <= not (a xor b);
    layer2_outputs(9352) <= not b or a;
    layer2_outputs(9353) <= b and not a;
    layer2_outputs(9354) <= a and b;
    layer2_outputs(9355) <= 1'b1;
    layer2_outputs(9356) <= not (a xor b);
    layer2_outputs(9357) <= b;
    layer2_outputs(9358) <= a or b;
    layer2_outputs(9359) <= not a;
    layer2_outputs(9360) <= not a or b;
    layer2_outputs(9361) <= not (a and b);
    layer2_outputs(9362) <= 1'b0;
    layer2_outputs(9363) <= a xor b;
    layer2_outputs(9364) <= not a or b;
    layer2_outputs(9365) <= a;
    layer2_outputs(9366) <= a;
    layer2_outputs(9367) <= not a;
    layer2_outputs(9368) <= b and not a;
    layer2_outputs(9369) <= not b;
    layer2_outputs(9370) <= 1'b0;
    layer2_outputs(9371) <= 1'b0;
    layer2_outputs(9372) <= not (a or b);
    layer2_outputs(9373) <= b;
    layer2_outputs(9374) <= not a;
    layer2_outputs(9375) <= not (a or b);
    layer2_outputs(9376) <= not (a or b);
    layer2_outputs(9377) <= a or b;
    layer2_outputs(9378) <= a and not b;
    layer2_outputs(9379) <= a and b;
    layer2_outputs(9380) <= 1'b0;
    layer2_outputs(9381) <= not (a xor b);
    layer2_outputs(9382) <= 1'b1;
    layer2_outputs(9383) <= not a;
    layer2_outputs(9384) <= not (a or b);
    layer2_outputs(9385) <= not (a xor b);
    layer2_outputs(9386) <= 1'b0;
    layer2_outputs(9387) <= not a or b;
    layer2_outputs(9388) <= not (a and b);
    layer2_outputs(9389) <= not (a and b);
    layer2_outputs(9390) <= 1'b0;
    layer2_outputs(9391) <= a or b;
    layer2_outputs(9392) <= not b;
    layer2_outputs(9393) <= 1'b1;
    layer2_outputs(9394) <= not a;
    layer2_outputs(9395) <= not (a or b);
    layer2_outputs(9396) <= a and b;
    layer2_outputs(9397) <= 1'b0;
    layer2_outputs(9398) <= a or b;
    layer2_outputs(9399) <= b;
    layer2_outputs(9400) <= b and not a;
    layer2_outputs(9401) <= not a;
    layer2_outputs(9402) <= not (a or b);
    layer2_outputs(9403) <= 1'b0;
    layer2_outputs(9404) <= not (a or b);
    layer2_outputs(9405) <= 1'b0;
    layer2_outputs(9406) <= 1'b1;
    layer2_outputs(9407) <= b and not a;
    layer2_outputs(9408) <= 1'b1;
    layer2_outputs(9409) <= not a or b;
    layer2_outputs(9410) <= a or b;
    layer2_outputs(9411) <= a and not b;
    layer2_outputs(9412) <= a and not b;
    layer2_outputs(9413) <= not b;
    layer2_outputs(9414) <= 1'b1;
    layer2_outputs(9415) <= not b or a;
    layer2_outputs(9416) <= not (a and b);
    layer2_outputs(9417) <= b;
    layer2_outputs(9418) <= not b;
    layer2_outputs(9419) <= not a or b;
    layer2_outputs(9420) <= not a;
    layer2_outputs(9421) <= a xor b;
    layer2_outputs(9422) <= not a or b;
    layer2_outputs(9423) <= b;
    layer2_outputs(9424) <= b;
    layer2_outputs(9425) <= not a or b;
    layer2_outputs(9426) <= not b;
    layer2_outputs(9427) <= not b or a;
    layer2_outputs(9428) <= 1'b0;
    layer2_outputs(9429) <= a and not b;
    layer2_outputs(9430) <= b and not a;
    layer2_outputs(9431) <= 1'b0;
    layer2_outputs(9432) <= not b or a;
    layer2_outputs(9433) <= not a or b;
    layer2_outputs(9434) <= a and not b;
    layer2_outputs(9435) <= not b or a;
    layer2_outputs(9436) <= not (a or b);
    layer2_outputs(9437) <= not (a and b);
    layer2_outputs(9438) <= not (a or b);
    layer2_outputs(9439) <= 1'b0;
    layer2_outputs(9440) <= a or b;
    layer2_outputs(9441) <= a and b;
    layer2_outputs(9442) <= not b;
    layer2_outputs(9443) <= not a or b;
    layer2_outputs(9444) <= not b or a;
    layer2_outputs(9445) <= not a;
    layer2_outputs(9446) <= a and not b;
    layer2_outputs(9447) <= a or b;
    layer2_outputs(9448) <= not b;
    layer2_outputs(9449) <= not (a or b);
    layer2_outputs(9450) <= not b or a;
    layer2_outputs(9451) <= 1'b1;
    layer2_outputs(9452) <= b and not a;
    layer2_outputs(9453) <= 1'b1;
    layer2_outputs(9454) <= a and b;
    layer2_outputs(9455) <= 1'b0;
    layer2_outputs(9456) <= not a or b;
    layer2_outputs(9457) <= a and not b;
    layer2_outputs(9458) <= not b or a;
    layer2_outputs(9459) <= a and b;
    layer2_outputs(9460) <= not b or a;
    layer2_outputs(9461) <= not (a or b);
    layer2_outputs(9462) <= 1'b0;
    layer2_outputs(9463) <= 1'b0;
    layer2_outputs(9464) <= not a;
    layer2_outputs(9465) <= 1'b0;
    layer2_outputs(9466) <= b and not a;
    layer2_outputs(9467) <= 1'b1;
    layer2_outputs(9468) <= 1'b0;
    layer2_outputs(9469) <= b and not a;
    layer2_outputs(9470) <= 1'b0;
    layer2_outputs(9471) <= not b;
    layer2_outputs(9472) <= not a;
    layer2_outputs(9473) <= a;
    layer2_outputs(9474) <= not b or a;
    layer2_outputs(9475) <= not (a or b);
    layer2_outputs(9476) <= 1'b1;
    layer2_outputs(9477) <= not (a and b);
    layer2_outputs(9478) <= 1'b1;
    layer2_outputs(9479) <= not (a and b);
    layer2_outputs(9480) <= b;
    layer2_outputs(9481) <= 1'b1;
    layer2_outputs(9482) <= not a;
    layer2_outputs(9483) <= 1'b1;
    layer2_outputs(9484) <= a;
    layer2_outputs(9485) <= a or b;
    layer2_outputs(9486) <= a and b;
    layer2_outputs(9487) <= a or b;
    layer2_outputs(9488) <= 1'b0;
    layer2_outputs(9489) <= not b;
    layer2_outputs(9490) <= not b or a;
    layer2_outputs(9491) <= not a;
    layer2_outputs(9492) <= not a;
    layer2_outputs(9493) <= a and not b;
    layer2_outputs(9494) <= b;
    layer2_outputs(9495) <= a and b;
    layer2_outputs(9496) <= not (a or b);
    layer2_outputs(9497) <= a;
    layer2_outputs(9498) <= b;
    layer2_outputs(9499) <= not (a xor b);
    layer2_outputs(9500) <= b and not a;
    layer2_outputs(9501) <= b and not a;
    layer2_outputs(9502) <= b and not a;
    layer2_outputs(9503) <= not a;
    layer2_outputs(9504) <= a and not b;
    layer2_outputs(9505) <= not a or b;
    layer2_outputs(9506) <= 1'b1;
    layer2_outputs(9507) <= not a;
    layer2_outputs(9508) <= b;
    layer2_outputs(9509) <= b and not a;
    layer2_outputs(9510) <= a and not b;
    layer2_outputs(9511) <= not b;
    layer2_outputs(9512) <= a;
    layer2_outputs(9513) <= not a;
    layer2_outputs(9514) <= b and not a;
    layer2_outputs(9515) <= a and b;
    layer2_outputs(9516) <= not b or a;
    layer2_outputs(9517) <= a and b;
    layer2_outputs(9518) <= not a or b;
    layer2_outputs(9519) <= 1'b1;
    layer2_outputs(9520) <= a and b;
    layer2_outputs(9521) <= a or b;
    layer2_outputs(9522) <= not (a and b);
    layer2_outputs(9523) <= a and b;
    layer2_outputs(9524) <= a or b;
    layer2_outputs(9525) <= not (a and b);
    layer2_outputs(9526) <= not b;
    layer2_outputs(9527) <= not (a and b);
    layer2_outputs(9528) <= 1'b0;
    layer2_outputs(9529) <= not (a and b);
    layer2_outputs(9530) <= not a;
    layer2_outputs(9531) <= b;
    layer2_outputs(9532) <= not a or b;
    layer2_outputs(9533) <= not b or a;
    layer2_outputs(9534) <= not a or b;
    layer2_outputs(9535) <= not a or b;
    layer2_outputs(9536) <= not (a and b);
    layer2_outputs(9537) <= not b;
    layer2_outputs(9538) <= a and b;
    layer2_outputs(9539) <= b and not a;
    layer2_outputs(9540) <= not a;
    layer2_outputs(9541) <= 1'b0;
    layer2_outputs(9542) <= b;
    layer2_outputs(9543) <= not (a or b);
    layer2_outputs(9544) <= a;
    layer2_outputs(9545) <= b;
    layer2_outputs(9546) <= a xor b;
    layer2_outputs(9547) <= not a;
    layer2_outputs(9548) <= not b;
    layer2_outputs(9549) <= a and b;
    layer2_outputs(9550) <= a or b;
    layer2_outputs(9551) <= b and not a;
    layer2_outputs(9552) <= not a;
    layer2_outputs(9553) <= not (a or b);
    layer2_outputs(9554) <= 1'b1;
    layer2_outputs(9555) <= not b or a;
    layer2_outputs(9556) <= not a;
    layer2_outputs(9557) <= a;
    layer2_outputs(9558) <= b and not a;
    layer2_outputs(9559) <= a;
    layer2_outputs(9560) <= a and b;
    layer2_outputs(9561) <= not a;
    layer2_outputs(9562) <= not (a and b);
    layer2_outputs(9563) <= 1'b1;
    layer2_outputs(9564) <= b and not a;
    layer2_outputs(9565) <= not (a and b);
    layer2_outputs(9566) <= 1'b0;
    layer2_outputs(9567) <= 1'b1;
    layer2_outputs(9568) <= a or b;
    layer2_outputs(9569) <= not (a or b);
    layer2_outputs(9570) <= not a;
    layer2_outputs(9571) <= not (a or b);
    layer2_outputs(9572) <= a and not b;
    layer2_outputs(9573) <= a;
    layer2_outputs(9574) <= 1'b1;
    layer2_outputs(9575) <= a xor b;
    layer2_outputs(9576) <= b;
    layer2_outputs(9577) <= not (a or b);
    layer2_outputs(9578) <= a and not b;
    layer2_outputs(9579) <= not (a and b);
    layer2_outputs(9580) <= not a or b;
    layer2_outputs(9581) <= not b;
    layer2_outputs(9582) <= not (a xor b);
    layer2_outputs(9583) <= not (a and b);
    layer2_outputs(9584) <= 1'b0;
    layer2_outputs(9585) <= b and not a;
    layer2_outputs(9586) <= not (a or b);
    layer2_outputs(9587) <= b and not a;
    layer2_outputs(9588) <= a and not b;
    layer2_outputs(9589) <= a or b;
    layer2_outputs(9590) <= 1'b1;
    layer2_outputs(9591) <= 1'b1;
    layer2_outputs(9592) <= a or b;
    layer2_outputs(9593) <= not b or a;
    layer2_outputs(9594) <= 1'b1;
    layer2_outputs(9595) <= 1'b0;
    layer2_outputs(9596) <= a and b;
    layer2_outputs(9597) <= b;
    layer2_outputs(9598) <= b and not a;
    layer2_outputs(9599) <= a and not b;
    layer2_outputs(9600) <= a and b;
    layer2_outputs(9601) <= a and b;
    layer2_outputs(9602) <= a and not b;
    layer2_outputs(9603) <= not (a and b);
    layer2_outputs(9604) <= not b or a;
    layer2_outputs(9605) <= a;
    layer2_outputs(9606) <= not (a or b);
    layer2_outputs(9607) <= not (a and b);
    layer2_outputs(9608) <= 1'b0;
    layer2_outputs(9609) <= a and b;
    layer2_outputs(9610) <= a xor b;
    layer2_outputs(9611) <= a and not b;
    layer2_outputs(9612) <= b and not a;
    layer2_outputs(9613) <= not (a or b);
    layer2_outputs(9614) <= b and not a;
    layer2_outputs(9615) <= not b or a;
    layer2_outputs(9616) <= not b;
    layer2_outputs(9617) <= not b or a;
    layer2_outputs(9618) <= 1'b0;
    layer2_outputs(9619) <= 1'b0;
    layer2_outputs(9620) <= a or b;
    layer2_outputs(9621) <= a or b;
    layer2_outputs(9622) <= not b or a;
    layer2_outputs(9623) <= 1'b0;
    layer2_outputs(9624) <= not (a xor b);
    layer2_outputs(9625) <= not a;
    layer2_outputs(9626) <= b;
    layer2_outputs(9627) <= a and b;
    layer2_outputs(9628) <= b and not a;
    layer2_outputs(9629) <= 1'b1;
    layer2_outputs(9630) <= 1'b0;
    layer2_outputs(9631) <= not b or a;
    layer2_outputs(9632) <= a xor b;
    layer2_outputs(9633) <= not a;
    layer2_outputs(9634) <= not a or b;
    layer2_outputs(9635) <= not b or a;
    layer2_outputs(9636) <= 1'b0;
    layer2_outputs(9637) <= 1'b0;
    layer2_outputs(9638) <= a and not b;
    layer2_outputs(9639) <= not (a or b);
    layer2_outputs(9640) <= 1'b0;
    layer2_outputs(9641) <= a or b;
    layer2_outputs(9642) <= not (a and b);
    layer2_outputs(9643) <= not (a or b);
    layer2_outputs(9644) <= b;
    layer2_outputs(9645) <= b and not a;
    layer2_outputs(9646) <= not (a xor b);
    layer2_outputs(9647) <= not (a or b);
    layer2_outputs(9648) <= 1'b1;
    layer2_outputs(9649) <= not a or b;
    layer2_outputs(9650) <= a or b;
    layer2_outputs(9651) <= not (a or b);
    layer2_outputs(9652) <= not (a or b);
    layer2_outputs(9653) <= 1'b1;
    layer2_outputs(9654) <= b;
    layer2_outputs(9655) <= 1'b1;
    layer2_outputs(9656) <= 1'b0;
    layer2_outputs(9657) <= a or b;
    layer2_outputs(9658) <= a and not b;
    layer2_outputs(9659) <= 1'b1;
    layer2_outputs(9660) <= a and not b;
    layer2_outputs(9661) <= a and not b;
    layer2_outputs(9662) <= 1'b0;
    layer2_outputs(9663) <= a and not b;
    layer2_outputs(9664) <= not (a or b);
    layer2_outputs(9665) <= 1'b0;
    layer2_outputs(9666) <= not b;
    layer2_outputs(9667) <= a and b;
    layer2_outputs(9668) <= not a or b;
    layer2_outputs(9669) <= 1'b1;
    layer2_outputs(9670) <= a or b;
    layer2_outputs(9671) <= a and not b;
    layer2_outputs(9672) <= not a or b;
    layer2_outputs(9673) <= not (a and b);
    layer2_outputs(9674) <= a or b;
    layer2_outputs(9675) <= 1'b1;
    layer2_outputs(9676) <= not (a or b);
    layer2_outputs(9677) <= a xor b;
    layer2_outputs(9678) <= a and b;
    layer2_outputs(9679) <= not b or a;
    layer2_outputs(9680) <= b and not a;
    layer2_outputs(9681) <= 1'b1;
    layer2_outputs(9682) <= not b or a;
    layer2_outputs(9683) <= b and not a;
    layer2_outputs(9684) <= a and not b;
    layer2_outputs(9685) <= not a or b;
    layer2_outputs(9686) <= a or b;
    layer2_outputs(9687) <= 1'b1;
    layer2_outputs(9688) <= not (a or b);
    layer2_outputs(9689) <= not a;
    layer2_outputs(9690) <= b;
    layer2_outputs(9691) <= not a or b;
    layer2_outputs(9692) <= not (a xor b);
    layer2_outputs(9693) <= 1'b0;
    layer2_outputs(9694) <= not b;
    layer2_outputs(9695) <= not b;
    layer2_outputs(9696) <= not a;
    layer2_outputs(9697) <= not b or a;
    layer2_outputs(9698) <= not (a and b);
    layer2_outputs(9699) <= not a;
    layer2_outputs(9700) <= a or b;
    layer2_outputs(9701) <= a and b;
    layer2_outputs(9702) <= not a;
    layer2_outputs(9703) <= 1'b0;
    layer2_outputs(9704) <= a and b;
    layer2_outputs(9705) <= a or b;
    layer2_outputs(9706) <= not b or a;
    layer2_outputs(9707) <= not b or a;
    layer2_outputs(9708) <= not (a and b);
    layer2_outputs(9709) <= a xor b;
    layer2_outputs(9710) <= a or b;
    layer2_outputs(9711) <= not (a xor b);
    layer2_outputs(9712) <= b;
    layer2_outputs(9713) <= 1'b0;
    layer2_outputs(9714) <= a;
    layer2_outputs(9715) <= a xor b;
    layer2_outputs(9716) <= b and not a;
    layer2_outputs(9717) <= a and not b;
    layer2_outputs(9718) <= not a or b;
    layer2_outputs(9719) <= a;
    layer2_outputs(9720) <= a and b;
    layer2_outputs(9721) <= a and not b;
    layer2_outputs(9722) <= a or b;
    layer2_outputs(9723) <= not (a or b);
    layer2_outputs(9724) <= not a;
    layer2_outputs(9725) <= not b or a;
    layer2_outputs(9726) <= a and b;
    layer2_outputs(9727) <= not (a or b);
    layer2_outputs(9728) <= 1'b1;
    layer2_outputs(9729) <= b and not a;
    layer2_outputs(9730) <= a xor b;
    layer2_outputs(9731) <= not a;
    layer2_outputs(9732) <= b;
    layer2_outputs(9733) <= b and not a;
    layer2_outputs(9734) <= a and b;
    layer2_outputs(9735) <= b and not a;
    layer2_outputs(9736) <= a or b;
    layer2_outputs(9737) <= not (a or b);
    layer2_outputs(9738) <= a and b;
    layer2_outputs(9739) <= not (a and b);
    layer2_outputs(9740) <= a and b;
    layer2_outputs(9741) <= not b;
    layer2_outputs(9742) <= not b;
    layer2_outputs(9743) <= not (a and b);
    layer2_outputs(9744) <= not a or b;
    layer2_outputs(9745) <= a and not b;
    layer2_outputs(9746) <= a;
    layer2_outputs(9747) <= not a;
    layer2_outputs(9748) <= not a;
    layer2_outputs(9749) <= a and not b;
    layer2_outputs(9750) <= not a;
    layer2_outputs(9751) <= not b;
    layer2_outputs(9752) <= not b or a;
    layer2_outputs(9753) <= a and b;
    layer2_outputs(9754) <= a or b;
    layer2_outputs(9755) <= not b;
    layer2_outputs(9756) <= a and b;
    layer2_outputs(9757) <= b;
    layer2_outputs(9758) <= not (a and b);
    layer2_outputs(9759) <= b;
    layer2_outputs(9760) <= 1'b1;
    layer2_outputs(9761) <= a and b;
    layer2_outputs(9762) <= not b or a;
    layer2_outputs(9763) <= not (a or b);
    layer2_outputs(9764) <= not (a and b);
    layer2_outputs(9765) <= a and b;
    layer2_outputs(9766) <= a and b;
    layer2_outputs(9767) <= 1'b0;
    layer2_outputs(9768) <= a;
    layer2_outputs(9769) <= not b;
    layer2_outputs(9770) <= not b;
    layer2_outputs(9771) <= 1'b0;
    layer2_outputs(9772) <= not b or a;
    layer2_outputs(9773) <= not (a and b);
    layer2_outputs(9774) <= not b;
    layer2_outputs(9775) <= not a or b;
    layer2_outputs(9776) <= a;
    layer2_outputs(9777) <= b;
    layer2_outputs(9778) <= a xor b;
    layer2_outputs(9779) <= a;
    layer2_outputs(9780) <= not a;
    layer2_outputs(9781) <= not b or a;
    layer2_outputs(9782) <= not (a xor b);
    layer2_outputs(9783) <= a and not b;
    layer2_outputs(9784) <= not (a and b);
    layer2_outputs(9785) <= 1'b0;
    layer2_outputs(9786) <= a or b;
    layer2_outputs(9787) <= 1'b0;
    layer2_outputs(9788) <= a and not b;
    layer2_outputs(9789) <= 1'b0;
    layer2_outputs(9790) <= a;
    layer2_outputs(9791) <= not b;
    layer2_outputs(9792) <= a and not b;
    layer2_outputs(9793) <= not b;
    layer2_outputs(9794) <= not a or b;
    layer2_outputs(9795) <= 1'b1;
    layer2_outputs(9796) <= not b;
    layer2_outputs(9797) <= 1'b1;
    layer2_outputs(9798) <= b;
    layer2_outputs(9799) <= 1'b0;
    layer2_outputs(9800) <= not b or a;
    layer2_outputs(9801) <= 1'b0;
    layer2_outputs(9802) <= 1'b0;
    layer2_outputs(9803) <= 1'b1;
    layer2_outputs(9804) <= not b or a;
    layer2_outputs(9805) <= not (a xor b);
    layer2_outputs(9806) <= not b;
    layer2_outputs(9807) <= a and b;
    layer2_outputs(9808) <= 1'b1;
    layer2_outputs(9809) <= a and b;
    layer2_outputs(9810) <= b and not a;
    layer2_outputs(9811) <= not a;
    layer2_outputs(9812) <= 1'b0;
    layer2_outputs(9813) <= 1'b0;
    layer2_outputs(9814) <= a and b;
    layer2_outputs(9815) <= 1'b1;
    layer2_outputs(9816) <= a or b;
    layer2_outputs(9817) <= not (a or b);
    layer2_outputs(9818) <= not (a and b);
    layer2_outputs(9819) <= a and not b;
    layer2_outputs(9820) <= not (a and b);
    layer2_outputs(9821) <= not b or a;
    layer2_outputs(9822) <= 1'b0;
    layer2_outputs(9823) <= not (a xor b);
    layer2_outputs(9824) <= not b or a;
    layer2_outputs(9825) <= a and not b;
    layer2_outputs(9826) <= a;
    layer2_outputs(9827) <= a or b;
    layer2_outputs(9828) <= not (a and b);
    layer2_outputs(9829) <= not b;
    layer2_outputs(9830) <= a and b;
    layer2_outputs(9831) <= not b;
    layer2_outputs(9832) <= a and b;
    layer2_outputs(9833) <= 1'b1;
    layer2_outputs(9834) <= not a;
    layer2_outputs(9835) <= a;
    layer2_outputs(9836) <= not b;
    layer2_outputs(9837) <= a or b;
    layer2_outputs(9838) <= not (a and b);
    layer2_outputs(9839) <= 1'b0;
    layer2_outputs(9840) <= 1'b0;
    layer2_outputs(9841) <= a xor b;
    layer2_outputs(9842) <= a and b;
    layer2_outputs(9843) <= a and b;
    layer2_outputs(9844) <= 1'b0;
    layer2_outputs(9845) <= 1'b1;
    layer2_outputs(9846) <= a and b;
    layer2_outputs(9847) <= a;
    layer2_outputs(9848) <= not (a or b);
    layer2_outputs(9849) <= a xor b;
    layer2_outputs(9850) <= not (a or b);
    layer2_outputs(9851) <= a or b;
    layer2_outputs(9852) <= b;
    layer2_outputs(9853) <= a and b;
    layer2_outputs(9854) <= a and not b;
    layer2_outputs(9855) <= a;
    layer2_outputs(9856) <= not (a xor b);
    layer2_outputs(9857) <= not (a and b);
    layer2_outputs(9858) <= not a or b;
    layer2_outputs(9859) <= a;
    layer2_outputs(9860) <= b;
    layer2_outputs(9861) <= b and not a;
    layer2_outputs(9862) <= a xor b;
    layer2_outputs(9863) <= a or b;
    layer2_outputs(9864) <= a or b;
    layer2_outputs(9865) <= 1'b1;
    layer2_outputs(9866) <= b;
    layer2_outputs(9867) <= not b or a;
    layer2_outputs(9868) <= 1'b0;
    layer2_outputs(9869) <= not b or a;
    layer2_outputs(9870) <= not (a xor b);
    layer2_outputs(9871) <= a;
    layer2_outputs(9872) <= not (a or b);
    layer2_outputs(9873) <= not (a and b);
    layer2_outputs(9874) <= 1'b1;
    layer2_outputs(9875) <= not a or b;
    layer2_outputs(9876) <= 1'b1;
    layer2_outputs(9877) <= b;
    layer2_outputs(9878) <= not b;
    layer2_outputs(9879) <= a and b;
    layer2_outputs(9880) <= 1'b0;
    layer2_outputs(9881) <= 1'b0;
    layer2_outputs(9882) <= 1'b1;
    layer2_outputs(9883) <= a;
    layer2_outputs(9884) <= b and not a;
    layer2_outputs(9885) <= not a;
    layer2_outputs(9886) <= a and b;
    layer2_outputs(9887) <= a;
    layer2_outputs(9888) <= not (a or b);
    layer2_outputs(9889) <= 1'b0;
    layer2_outputs(9890) <= not a;
    layer2_outputs(9891) <= not a;
    layer2_outputs(9892) <= 1'b1;
    layer2_outputs(9893) <= a and not b;
    layer2_outputs(9894) <= a and b;
    layer2_outputs(9895) <= not a;
    layer2_outputs(9896) <= a and b;
    layer2_outputs(9897) <= not b;
    layer2_outputs(9898) <= not (a and b);
    layer2_outputs(9899) <= not a or b;
    layer2_outputs(9900) <= not a or b;
    layer2_outputs(9901) <= a and b;
    layer2_outputs(9902) <= not a or b;
    layer2_outputs(9903) <= not b;
    layer2_outputs(9904) <= 1'b0;
    layer2_outputs(9905) <= a and not b;
    layer2_outputs(9906) <= not (a or b);
    layer2_outputs(9907) <= a xor b;
    layer2_outputs(9908) <= a;
    layer2_outputs(9909) <= 1'b1;
    layer2_outputs(9910) <= 1'b1;
    layer2_outputs(9911) <= a and not b;
    layer2_outputs(9912) <= a and b;
    layer2_outputs(9913) <= a and not b;
    layer2_outputs(9914) <= a and b;
    layer2_outputs(9915) <= not (a and b);
    layer2_outputs(9916) <= a;
    layer2_outputs(9917) <= not a or b;
    layer2_outputs(9918) <= not b or a;
    layer2_outputs(9919) <= not b or a;
    layer2_outputs(9920) <= a and not b;
    layer2_outputs(9921) <= a or b;
    layer2_outputs(9922) <= a and b;
    layer2_outputs(9923) <= not b;
    layer2_outputs(9924) <= not b or a;
    layer2_outputs(9925) <= b;
    layer2_outputs(9926) <= not (a and b);
    layer2_outputs(9927) <= a or b;
    layer2_outputs(9928) <= not a;
    layer2_outputs(9929) <= not (a and b);
    layer2_outputs(9930) <= not b or a;
    layer2_outputs(9931) <= 1'b1;
    layer2_outputs(9932) <= a;
    layer2_outputs(9933) <= not a or b;
    layer2_outputs(9934) <= a and b;
    layer2_outputs(9935) <= not a or b;
    layer2_outputs(9936) <= a and not b;
    layer2_outputs(9937) <= a and not b;
    layer2_outputs(9938) <= not a or b;
    layer2_outputs(9939) <= a or b;
    layer2_outputs(9940) <= 1'b1;
    layer2_outputs(9941) <= 1'b0;
    layer2_outputs(9942) <= a or b;
    layer2_outputs(9943) <= not a;
    layer2_outputs(9944) <= 1'b0;
    layer2_outputs(9945) <= a and b;
    layer2_outputs(9946) <= not b;
    layer2_outputs(9947) <= not a;
    layer2_outputs(9948) <= not b or a;
    layer2_outputs(9949) <= not a;
    layer2_outputs(9950) <= b;
    layer2_outputs(9951) <= a or b;
    layer2_outputs(9952) <= 1'b0;
    layer2_outputs(9953) <= b and not a;
    layer2_outputs(9954) <= a and not b;
    layer2_outputs(9955) <= not a;
    layer2_outputs(9956) <= a and b;
    layer2_outputs(9957) <= a;
    layer2_outputs(9958) <= not a or b;
    layer2_outputs(9959) <= a and b;
    layer2_outputs(9960) <= 1'b1;
    layer2_outputs(9961) <= not a or b;
    layer2_outputs(9962) <= a and not b;
    layer2_outputs(9963) <= a and not b;
    layer2_outputs(9964) <= b;
    layer2_outputs(9965) <= 1'b1;
    layer2_outputs(9966) <= not (a xor b);
    layer2_outputs(9967) <= not a or b;
    layer2_outputs(9968) <= b and not a;
    layer2_outputs(9969) <= not (a and b);
    layer2_outputs(9970) <= not b or a;
    layer2_outputs(9971) <= 1'b1;
    layer2_outputs(9972) <= not b or a;
    layer2_outputs(9973) <= b;
    layer2_outputs(9974) <= a;
    layer2_outputs(9975) <= not b or a;
    layer2_outputs(9976) <= not b;
    layer2_outputs(9977) <= not a or b;
    layer2_outputs(9978) <= a and b;
    layer2_outputs(9979) <= a or b;
    layer2_outputs(9980) <= 1'b0;
    layer2_outputs(9981) <= not b;
    layer2_outputs(9982) <= 1'b0;
    layer2_outputs(9983) <= a or b;
    layer2_outputs(9984) <= b and not a;
    layer2_outputs(9985) <= 1'b0;
    layer2_outputs(9986) <= a xor b;
    layer2_outputs(9987) <= not (a and b);
    layer2_outputs(9988) <= a and not b;
    layer2_outputs(9989) <= a and not b;
    layer2_outputs(9990) <= not b;
    layer2_outputs(9991) <= b;
    layer2_outputs(9992) <= b and not a;
    layer2_outputs(9993) <= not a or b;
    layer2_outputs(9994) <= a and not b;
    layer2_outputs(9995) <= b;
    layer2_outputs(9996) <= not (a or b);
    layer2_outputs(9997) <= a;
    layer2_outputs(9998) <= a;
    layer2_outputs(9999) <= not (a xor b);
    layer2_outputs(10000) <= not (a or b);
    layer2_outputs(10001) <= a and not b;
    layer2_outputs(10002) <= a and b;
    layer2_outputs(10003) <= not a or b;
    layer2_outputs(10004) <= not a or b;
    layer2_outputs(10005) <= not (a or b);
    layer2_outputs(10006) <= 1'b0;
    layer2_outputs(10007) <= 1'b1;
    layer2_outputs(10008) <= not b or a;
    layer2_outputs(10009) <= 1'b1;
    layer2_outputs(10010) <= 1'b1;
    layer2_outputs(10011) <= b;
    layer2_outputs(10012) <= b and not a;
    layer2_outputs(10013) <= 1'b0;
    layer2_outputs(10014) <= a;
    layer2_outputs(10015) <= b and not a;
    layer2_outputs(10016) <= not (a and b);
    layer2_outputs(10017) <= 1'b0;
    layer2_outputs(10018) <= not a or b;
    layer2_outputs(10019) <= 1'b0;
    layer2_outputs(10020) <= a and not b;
    layer2_outputs(10021) <= a;
    layer2_outputs(10022) <= a or b;
    layer2_outputs(10023) <= a and not b;
    layer2_outputs(10024) <= not a or b;
    layer2_outputs(10025) <= 1'b1;
    layer2_outputs(10026) <= a or b;
    layer2_outputs(10027) <= a or b;
    layer2_outputs(10028) <= not (a and b);
    layer2_outputs(10029) <= not (a xor b);
    layer2_outputs(10030) <= not (a and b);
    layer2_outputs(10031) <= not b;
    layer2_outputs(10032) <= 1'b1;
    layer2_outputs(10033) <= 1'b1;
    layer2_outputs(10034) <= not (a and b);
    layer2_outputs(10035) <= a xor b;
    layer2_outputs(10036) <= 1'b1;
    layer2_outputs(10037) <= not a or b;
    layer2_outputs(10038) <= a xor b;
    layer2_outputs(10039) <= not (a and b);
    layer2_outputs(10040) <= b;
    layer2_outputs(10041) <= a and b;
    layer2_outputs(10042) <= a;
    layer2_outputs(10043) <= a;
    layer2_outputs(10044) <= not a or b;
    layer2_outputs(10045) <= 1'b0;
    layer2_outputs(10046) <= not a;
    layer2_outputs(10047) <= not b or a;
    layer2_outputs(10048) <= a and not b;
    layer2_outputs(10049) <= not b;
    layer2_outputs(10050) <= a;
    layer2_outputs(10051) <= 1'b1;
    layer2_outputs(10052) <= not a or b;
    layer2_outputs(10053) <= a;
    layer2_outputs(10054) <= b;
    layer2_outputs(10055) <= a;
    layer2_outputs(10056) <= a and not b;
    layer2_outputs(10057) <= not (a xor b);
    layer2_outputs(10058) <= a and not b;
    layer2_outputs(10059) <= not a or b;
    layer2_outputs(10060) <= 1'b0;
    layer2_outputs(10061) <= not (a and b);
    layer2_outputs(10062) <= 1'b0;
    layer2_outputs(10063) <= not b or a;
    layer2_outputs(10064) <= not (a xor b);
    layer2_outputs(10065) <= not (a xor b);
    layer2_outputs(10066) <= not (a or b);
    layer2_outputs(10067) <= not a;
    layer2_outputs(10068) <= not b;
    layer2_outputs(10069) <= not a;
    layer2_outputs(10070) <= b;
    layer2_outputs(10071) <= a or b;
    layer2_outputs(10072) <= a or b;
    layer2_outputs(10073) <= not (a xor b);
    layer2_outputs(10074) <= 1'b1;
    layer2_outputs(10075) <= not b;
    layer2_outputs(10076) <= a;
    layer2_outputs(10077) <= a;
    layer2_outputs(10078) <= not b;
    layer2_outputs(10079) <= not a;
    layer2_outputs(10080) <= not a or b;
    layer2_outputs(10081) <= not a or b;
    layer2_outputs(10082) <= not b or a;
    layer2_outputs(10083) <= not b or a;
    layer2_outputs(10084) <= not (a xor b);
    layer2_outputs(10085) <= not b;
    layer2_outputs(10086) <= not (a and b);
    layer2_outputs(10087) <= a or b;
    layer2_outputs(10088) <= 1'b1;
    layer2_outputs(10089) <= a;
    layer2_outputs(10090) <= a and b;
    layer2_outputs(10091) <= a or b;
    layer2_outputs(10092) <= 1'b1;
    layer2_outputs(10093) <= a and b;
    layer2_outputs(10094) <= a;
    layer2_outputs(10095) <= 1'b1;
    layer2_outputs(10096) <= not b;
    layer2_outputs(10097) <= a;
    layer2_outputs(10098) <= not b;
    layer2_outputs(10099) <= not (a and b);
    layer2_outputs(10100) <= 1'b1;
    layer2_outputs(10101) <= not b;
    layer2_outputs(10102) <= a and not b;
    layer2_outputs(10103) <= not b or a;
    layer2_outputs(10104) <= a and b;
    layer2_outputs(10105) <= a or b;
    layer2_outputs(10106) <= 1'b0;
    layer2_outputs(10107) <= 1'b0;
    layer2_outputs(10108) <= 1'b0;
    layer2_outputs(10109) <= a;
    layer2_outputs(10110) <= not a;
    layer2_outputs(10111) <= not a or b;
    layer2_outputs(10112) <= not b or a;
    layer2_outputs(10113) <= 1'b0;
    layer2_outputs(10114) <= b;
    layer2_outputs(10115) <= b and not a;
    layer2_outputs(10116) <= a and b;
    layer2_outputs(10117) <= b;
    layer2_outputs(10118) <= not b or a;
    layer2_outputs(10119) <= a and not b;
    layer2_outputs(10120) <= b;
    layer2_outputs(10121) <= b and not a;
    layer2_outputs(10122) <= not b;
    layer2_outputs(10123) <= b and not a;
    layer2_outputs(10124) <= b;
    layer2_outputs(10125) <= b and not a;
    layer2_outputs(10126) <= 1'b0;
    layer2_outputs(10127) <= a;
    layer2_outputs(10128) <= not a or b;
    layer2_outputs(10129) <= a or b;
    layer2_outputs(10130) <= not a;
    layer2_outputs(10131) <= a and not b;
    layer2_outputs(10132) <= not b or a;
    layer2_outputs(10133) <= a or b;
    layer2_outputs(10134) <= 1'b1;
    layer2_outputs(10135) <= not b or a;
    layer2_outputs(10136) <= not b;
    layer2_outputs(10137) <= not a;
    layer2_outputs(10138) <= a and b;
    layer2_outputs(10139) <= a or b;
    layer2_outputs(10140) <= not b or a;
    layer2_outputs(10141) <= b and not a;
    layer2_outputs(10142) <= not a or b;
    layer2_outputs(10143) <= a or b;
    layer2_outputs(10144) <= not (a or b);
    layer2_outputs(10145) <= not a;
    layer2_outputs(10146) <= a;
    layer2_outputs(10147) <= a and not b;
    layer2_outputs(10148) <= not a or b;
    layer2_outputs(10149) <= a xor b;
    layer2_outputs(10150) <= b;
    layer2_outputs(10151) <= not b;
    layer2_outputs(10152) <= a and not b;
    layer2_outputs(10153) <= 1'b1;
    layer2_outputs(10154) <= not a or b;
    layer2_outputs(10155) <= not a or b;
    layer2_outputs(10156) <= b;
    layer2_outputs(10157) <= 1'b0;
    layer2_outputs(10158) <= 1'b0;
    layer2_outputs(10159) <= not a or b;
    layer2_outputs(10160) <= 1'b0;
    layer2_outputs(10161) <= not b;
    layer2_outputs(10162) <= a and b;
    layer2_outputs(10163) <= not b or a;
    layer2_outputs(10164) <= not (a and b);
    layer2_outputs(10165) <= b;
    layer2_outputs(10166) <= not b or a;
    layer2_outputs(10167) <= 1'b0;
    layer2_outputs(10168) <= 1'b1;
    layer2_outputs(10169) <= a or b;
    layer2_outputs(10170) <= 1'b0;
    layer2_outputs(10171) <= 1'b1;
    layer2_outputs(10172) <= not (a or b);
    layer2_outputs(10173) <= 1'b1;
    layer2_outputs(10174) <= not b;
    layer2_outputs(10175) <= a or b;
    layer2_outputs(10176) <= not b;
    layer2_outputs(10177) <= b;
    layer2_outputs(10178) <= b and not a;
    layer2_outputs(10179) <= not (a or b);
    layer2_outputs(10180) <= 1'b1;
    layer2_outputs(10181) <= a;
    layer2_outputs(10182) <= a xor b;
    layer2_outputs(10183) <= not b;
    layer2_outputs(10184) <= not a;
    layer2_outputs(10185) <= b and not a;
    layer2_outputs(10186) <= a or b;
    layer2_outputs(10187) <= not a;
    layer2_outputs(10188) <= 1'b0;
    layer2_outputs(10189) <= a and b;
    layer2_outputs(10190) <= b;
    layer2_outputs(10191) <= not b;
    layer2_outputs(10192) <= not b;
    layer2_outputs(10193) <= 1'b1;
    layer2_outputs(10194) <= not b;
    layer2_outputs(10195) <= a and b;
    layer2_outputs(10196) <= not (a or b);
    layer2_outputs(10197) <= not a or b;
    layer2_outputs(10198) <= a;
    layer2_outputs(10199) <= 1'b1;
    layer2_outputs(10200) <= a and b;
    layer2_outputs(10201) <= a and b;
    layer2_outputs(10202) <= a and not b;
    layer2_outputs(10203) <= a or b;
    layer2_outputs(10204) <= not b;
    layer2_outputs(10205) <= not (a or b);
    layer2_outputs(10206) <= b;
    layer2_outputs(10207) <= not (a and b);
    layer2_outputs(10208) <= a;
    layer2_outputs(10209) <= not b;
    layer2_outputs(10210) <= not b;
    layer2_outputs(10211) <= a and b;
    layer2_outputs(10212) <= a and b;
    layer2_outputs(10213) <= 1'b0;
    layer2_outputs(10214) <= 1'b0;
    layer2_outputs(10215) <= 1'b0;
    layer2_outputs(10216) <= not a;
    layer2_outputs(10217) <= not b;
    layer2_outputs(10218) <= b and not a;
    layer2_outputs(10219) <= a or b;
    layer2_outputs(10220) <= 1'b0;
    layer2_outputs(10221) <= not (a and b);
    layer2_outputs(10222) <= not a;
    layer2_outputs(10223) <= 1'b1;
    layer2_outputs(10224) <= not a;
    layer2_outputs(10225) <= not b;
    layer2_outputs(10226) <= not (a or b);
    layer2_outputs(10227) <= a and not b;
    layer2_outputs(10228) <= a or b;
    layer2_outputs(10229) <= not b or a;
    layer2_outputs(10230) <= a;
    layer2_outputs(10231) <= a;
    layer2_outputs(10232) <= a or b;
    layer2_outputs(10233) <= not b or a;
    layer2_outputs(10234) <= not a or b;
    layer2_outputs(10235) <= a or b;
    layer2_outputs(10236) <= 1'b1;
    layer2_outputs(10237) <= b and not a;
    layer2_outputs(10238) <= a or b;
    layer2_outputs(10239) <= b;
    layer3_outputs(0) <= not b or a;
    layer3_outputs(1) <= not (a and b);
    layer3_outputs(2) <= not a or b;
    layer3_outputs(3) <= not b or a;
    layer3_outputs(4) <= a and not b;
    layer3_outputs(5) <= 1'b1;
    layer3_outputs(6) <= not (a and b);
    layer3_outputs(7) <= b;
    layer3_outputs(8) <= a or b;
    layer3_outputs(9) <= not a;
    layer3_outputs(10) <= not b or a;
    layer3_outputs(11) <= not a or b;
    layer3_outputs(12) <= a and b;
    layer3_outputs(13) <= not a or b;
    layer3_outputs(14) <= not (a or b);
    layer3_outputs(15) <= a;
    layer3_outputs(16) <= a and not b;
    layer3_outputs(17) <= not a or b;
    layer3_outputs(18) <= a and b;
    layer3_outputs(19) <= 1'b1;
    layer3_outputs(20) <= a;
    layer3_outputs(21) <= a xor b;
    layer3_outputs(22) <= b and not a;
    layer3_outputs(23) <= a and b;
    layer3_outputs(24) <= not (a or b);
    layer3_outputs(25) <= a or b;
    layer3_outputs(26) <= a and not b;
    layer3_outputs(27) <= a and b;
    layer3_outputs(28) <= not b;
    layer3_outputs(29) <= not b;
    layer3_outputs(30) <= b and not a;
    layer3_outputs(31) <= a or b;
    layer3_outputs(32) <= 1'b1;
    layer3_outputs(33) <= not a or b;
    layer3_outputs(34) <= a;
    layer3_outputs(35) <= 1'b1;
    layer3_outputs(36) <= not b or a;
    layer3_outputs(37) <= not (a or b);
    layer3_outputs(38) <= b and not a;
    layer3_outputs(39) <= b and not a;
    layer3_outputs(40) <= not a;
    layer3_outputs(41) <= a;
    layer3_outputs(42) <= b;
    layer3_outputs(43) <= not (a or b);
    layer3_outputs(44) <= a and b;
    layer3_outputs(45) <= not a or b;
    layer3_outputs(46) <= not (a and b);
    layer3_outputs(47) <= a;
    layer3_outputs(48) <= b and not a;
    layer3_outputs(49) <= not (a xor b);
    layer3_outputs(50) <= 1'b0;
    layer3_outputs(51) <= 1'b0;
    layer3_outputs(52) <= a or b;
    layer3_outputs(53) <= b and not a;
    layer3_outputs(54) <= not b or a;
    layer3_outputs(55) <= b;
    layer3_outputs(56) <= b;
    layer3_outputs(57) <= not (a and b);
    layer3_outputs(58) <= not (a xor b);
    layer3_outputs(59) <= not a or b;
    layer3_outputs(60) <= a and b;
    layer3_outputs(61) <= a;
    layer3_outputs(62) <= b;
    layer3_outputs(63) <= b;
    layer3_outputs(64) <= not a or b;
    layer3_outputs(65) <= a and b;
    layer3_outputs(66) <= a;
    layer3_outputs(67) <= not a;
    layer3_outputs(68) <= not b;
    layer3_outputs(69) <= a or b;
    layer3_outputs(70) <= a and not b;
    layer3_outputs(71) <= 1'b1;
    layer3_outputs(72) <= a xor b;
    layer3_outputs(73) <= b;
    layer3_outputs(74) <= a or b;
    layer3_outputs(75) <= not a;
    layer3_outputs(76) <= not a;
    layer3_outputs(77) <= a or b;
    layer3_outputs(78) <= not b;
    layer3_outputs(79) <= b;
    layer3_outputs(80) <= 1'b1;
    layer3_outputs(81) <= b and not a;
    layer3_outputs(82) <= not a;
    layer3_outputs(83) <= not (a and b);
    layer3_outputs(84) <= not b or a;
    layer3_outputs(85) <= 1'b1;
    layer3_outputs(86) <= a and not b;
    layer3_outputs(87) <= not (a or b);
    layer3_outputs(88) <= b;
    layer3_outputs(89) <= not a;
    layer3_outputs(90) <= not a;
    layer3_outputs(91) <= a;
    layer3_outputs(92) <= not a or b;
    layer3_outputs(93) <= b and not a;
    layer3_outputs(94) <= a and not b;
    layer3_outputs(95) <= a and not b;
    layer3_outputs(96) <= b;
    layer3_outputs(97) <= b and not a;
    layer3_outputs(98) <= a xor b;
    layer3_outputs(99) <= not (a and b);
    layer3_outputs(100) <= a;
    layer3_outputs(101) <= b and not a;
    layer3_outputs(102) <= 1'b0;
    layer3_outputs(103) <= a or b;
    layer3_outputs(104) <= 1'b0;
    layer3_outputs(105) <= not b or a;
    layer3_outputs(106) <= not a;
    layer3_outputs(107) <= a or b;
    layer3_outputs(108) <= a and not b;
    layer3_outputs(109) <= not b;
    layer3_outputs(110) <= 1'b0;
    layer3_outputs(111) <= 1'b0;
    layer3_outputs(112) <= 1'b1;
    layer3_outputs(113) <= a xor b;
    layer3_outputs(114) <= a;
    layer3_outputs(115) <= not a or b;
    layer3_outputs(116) <= not b or a;
    layer3_outputs(117) <= not b;
    layer3_outputs(118) <= 1'b0;
    layer3_outputs(119) <= a or b;
    layer3_outputs(120) <= not (a or b);
    layer3_outputs(121) <= 1'b0;
    layer3_outputs(122) <= a xor b;
    layer3_outputs(123) <= not b;
    layer3_outputs(124) <= a and not b;
    layer3_outputs(125) <= b and not a;
    layer3_outputs(126) <= b and not a;
    layer3_outputs(127) <= a or b;
    layer3_outputs(128) <= not a or b;
    layer3_outputs(129) <= not b or a;
    layer3_outputs(130) <= a and not b;
    layer3_outputs(131) <= not b;
    layer3_outputs(132) <= a and b;
    layer3_outputs(133) <= not b;
    layer3_outputs(134) <= not a;
    layer3_outputs(135) <= b and not a;
    layer3_outputs(136) <= 1'b1;
    layer3_outputs(137) <= not (a and b);
    layer3_outputs(138) <= 1'b0;
    layer3_outputs(139) <= not b;
    layer3_outputs(140) <= a or b;
    layer3_outputs(141) <= b;
    layer3_outputs(142) <= not (a or b);
    layer3_outputs(143) <= a xor b;
    layer3_outputs(144) <= not b or a;
    layer3_outputs(145) <= not a or b;
    layer3_outputs(146) <= b and not a;
    layer3_outputs(147) <= not a;
    layer3_outputs(148) <= not b or a;
    layer3_outputs(149) <= a;
    layer3_outputs(150) <= not (a and b);
    layer3_outputs(151) <= 1'b0;
    layer3_outputs(152) <= a or b;
    layer3_outputs(153) <= not b;
    layer3_outputs(154) <= a and b;
    layer3_outputs(155) <= not (a xor b);
    layer3_outputs(156) <= a and not b;
    layer3_outputs(157) <= b and not a;
    layer3_outputs(158) <= not (a or b);
    layer3_outputs(159) <= a xor b;
    layer3_outputs(160) <= b and not a;
    layer3_outputs(161) <= b and not a;
    layer3_outputs(162) <= a;
    layer3_outputs(163) <= a and b;
    layer3_outputs(164) <= not (a or b);
    layer3_outputs(165) <= 1'b0;
    layer3_outputs(166) <= b and not a;
    layer3_outputs(167) <= 1'b0;
    layer3_outputs(168) <= not (a or b);
    layer3_outputs(169) <= b;
    layer3_outputs(170) <= 1'b1;
    layer3_outputs(171) <= not b or a;
    layer3_outputs(172) <= not a;
    layer3_outputs(173) <= not (a and b);
    layer3_outputs(174) <= a;
    layer3_outputs(175) <= not a or b;
    layer3_outputs(176) <= not (a and b);
    layer3_outputs(177) <= b and not a;
    layer3_outputs(178) <= 1'b1;
    layer3_outputs(179) <= not a or b;
    layer3_outputs(180) <= not (a or b);
    layer3_outputs(181) <= b and not a;
    layer3_outputs(182) <= not (a or b);
    layer3_outputs(183) <= a or b;
    layer3_outputs(184) <= 1'b0;
    layer3_outputs(185) <= a and not b;
    layer3_outputs(186) <= not a;
    layer3_outputs(187) <= a and b;
    layer3_outputs(188) <= a;
    layer3_outputs(189) <= 1'b0;
    layer3_outputs(190) <= a or b;
    layer3_outputs(191) <= not a;
    layer3_outputs(192) <= b;
    layer3_outputs(193) <= not (a and b);
    layer3_outputs(194) <= a xor b;
    layer3_outputs(195) <= b;
    layer3_outputs(196) <= not b or a;
    layer3_outputs(197) <= a and not b;
    layer3_outputs(198) <= not a or b;
    layer3_outputs(199) <= not a;
    layer3_outputs(200) <= a;
    layer3_outputs(201) <= b and not a;
    layer3_outputs(202) <= not b or a;
    layer3_outputs(203) <= not b;
    layer3_outputs(204) <= not (a or b);
    layer3_outputs(205) <= 1'b0;
    layer3_outputs(206) <= a and b;
    layer3_outputs(207) <= b;
    layer3_outputs(208) <= b;
    layer3_outputs(209) <= a and not b;
    layer3_outputs(210) <= not (a and b);
    layer3_outputs(211) <= b and not a;
    layer3_outputs(212) <= a and b;
    layer3_outputs(213) <= b;
    layer3_outputs(214) <= 1'b0;
    layer3_outputs(215) <= b;
    layer3_outputs(216) <= not a or b;
    layer3_outputs(217) <= 1'b0;
    layer3_outputs(218) <= not (a xor b);
    layer3_outputs(219) <= a;
    layer3_outputs(220) <= 1'b1;
    layer3_outputs(221) <= a and b;
    layer3_outputs(222) <= a and not b;
    layer3_outputs(223) <= not (a and b);
    layer3_outputs(224) <= b;
    layer3_outputs(225) <= 1'b0;
    layer3_outputs(226) <= b and not a;
    layer3_outputs(227) <= not b;
    layer3_outputs(228) <= b and not a;
    layer3_outputs(229) <= not a or b;
    layer3_outputs(230) <= b and not a;
    layer3_outputs(231) <= not a or b;
    layer3_outputs(232) <= b;
    layer3_outputs(233) <= a or b;
    layer3_outputs(234) <= a xor b;
    layer3_outputs(235) <= 1'b1;
    layer3_outputs(236) <= not b or a;
    layer3_outputs(237) <= not (a or b);
    layer3_outputs(238) <= not (a or b);
    layer3_outputs(239) <= not b or a;
    layer3_outputs(240) <= 1'b0;
    layer3_outputs(241) <= not b or a;
    layer3_outputs(242) <= not (a and b);
    layer3_outputs(243) <= b;
    layer3_outputs(244) <= not b;
    layer3_outputs(245) <= not b or a;
    layer3_outputs(246) <= 1'b1;
    layer3_outputs(247) <= 1'b1;
    layer3_outputs(248) <= 1'b1;
    layer3_outputs(249) <= not a;
    layer3_outputs(250) <= not (a xor b);
    layer3_outputs(251) <= not b or a;
    layer3_outputs(252) <= not (a and b);
    layer3_outputs(253) <= 1'b1;
    layer3_outputs(254) <= not (a and b);
    layer3_outputs(255) <= 1'b1;
    layer3_outputs(256) <= b and not a;
    layer3_outputs(257) <= b and not a;
    layer3_outputs(258) <= b;
    layer3_outputs(259) <= a or b;
    layer3_outputs(260) <= a and not b;
    layer3_outputs(261) <= a and not b;
    layer3_outputs(262) <= not b or a;
    layer3_outputs(263) <= b and not a;
    layer3_outputs(264) <= not (a and b);
    layer3_outputs(265) <= not a;
    layer3_outputs(266) <= 1'b0;
    layer3_outputs(267) <= not a;
    layer3_outputs(268) <= 1'b1;
    layer3_outputs(269) <= not b or a;
    layer3_outputs(270) <= not b or a;
    layer3_outputs(271) <= not (a or b);
    layer3_outputs(272) <= not a or b;
    layer3_outputs(273) <= not b;
    layer3_outputs(274) <= 1'b1;
    layer3_outputs(275) <= not a;
    layer3_outputs(276) <= 1'b1;
    layer3_outputs(277) <= a xor b;
    layer3_outputs(278) <= 1'b0;
    layer3_outputs(279) <= a and b;
    layer3_outputs(280) <= 1'b1;
    layer3_outputs(281) <= a;
    layer3_outputs(282) <= not (a xor b);
    layer3_outputs(283) <= not a;
    layer3_outputs(284) <= not a;
    layer3_outputs(285) <= not a or b;
    layer3_outputs(286) <= not (a or b);
    layer3_outputs(287) <= b and not a;
    layer3_outputs(288) <= a or b;
    layer3_outputs(289) <= b;
    layer3_outputs(290) <= a and b;
    layer3_outputs(291) <= a and not b;
    layer3_outputs(292) <= b and not a;
    layer3_outputs(293) <= b and not a;
    layer3_outputs(294) <= not a or b;
    layer3_outputs(295) <= 1'b0;
    layer3_outputs(296) <= 1'b1;
    layer3_outputs(297) <= not (a and b);
    layer3_outputs(298) <= not b or a;
    layer3_outputs(299) <= not a or b;
    layer3_outputs(300) <= not (a or b);
    layer3_outputs(301) <= b and not a;
    layer3_outputs(302) <= a and b;
    layer3_outputs(303) <= not (a or b);
    layer3_outputs(304) <= not (a and b);
    layer3_outputs(305) <= not (a and b);
    layer3_outputs(306) <= not (a and b);
    layer3_outputs(307) <= not a;
    layer3_outputs(308) <= not (a xor b);
    layer3_outputs(309) <= 1'b1;
    layer3_outputs(310) <= a;
    layer3_outputs(311) <= a;
    layer3_outputs(312) <= not b;
    layer3_outputs(313) <= a and b;
    layer3_outputs(314) <= not (a or b);
    layer3_outputs(315) <= a;
    layer3_outputs(316) <= 1'b0;
    layer3_outputs(317) <= a and b;
    layer3_outputs(318) <= b;
    layer3_outputs(319) <= not (a xor b);
    layer3_outputs(320) <= not (a and b);
    layer3_outputs(321) <= a and b;
    layer3_outputs(322) <= a xor b;
    layer3_outputs(323) <= a and b;
    layer3_outputs(324) <= 1'b1;
    layer3_outputs(325) <= 1'b0;
    layer3_outputs(326) <= not (a or b);
    layer3_outputs(327) <= not (a or b);
    layer3_outputs(328) <= not a or b;
    layer3_outputs(329) <= 1'b0;
    layer3_outputs(330) <= not a;
    layer3_outputs(331) <= b and not a;
    layer3_outputs(332) <= a;
    layer3_outputs(333) <= a or b;
    layer3_outputs(334) <= b;
    layer3_outputs(335) <= not a or b;
    layer3_outputs(336) <= not (a and b);
    layer3_outputs(337) <= a and b;
    layer3_outputs(338) <= 1'b0;
    layer3_outputs(339) <= not (a and b);
    layer3_outputs(340) <= a or b;
    layer3_outputs(341) <= b and not a;
    layer3_outputs(342) <= 1'b0;
    layer3_outputs(343) <= a or b;
    layer3_outputs(344) <= b and not a;
    layer3_outputs(345) <= b;
    layer3_outputs(346) <= not (a and b);
    layer3_outputs(347) <= not (a and b);
    layer3_outputs(348) <= a xor b;
    layer3_outputs(349) <= a;
    layer3_outputs(350) <= 1'b0;
    layer3_outputs(351) <= 1'b1;
    layer3_outputs(352) <= not (a or b);
    layer3_outputs(353) <= a or b;
    layer3_outputs(354) <= b and not a;
    layer3_outputs(355) <= b;
    layer3_outputs(356) <= a or b;
    layer3_outputs(357) <= b and not a;
    layer3_outputs(358) <= not b or a;
    layer3_outputs(359) <= b and not a;
    layer3_outputs(360) <= 1'b1;
    layer3_outputs(361) <= not (a and b);
    layer3_outputs(362) <= b and not a;
    layer3_outputs(363) <= a and b;
    layer3_outputs(364) <= b;
    layer3_outputs(365) <= a;
    layer3_outputs(366) <= b and not a;
    layer3_outputs(367) <= a and not b;
    layer3_outputs(368) <= b;
    layer3_outputs(369) <= not a;
    layer3_outputs(370) <= a;
    layer3_outputs(371) <= 1'b0;
    layer3_outputs(372) <= b and not a;
    layer3_outputs(373) <= 1'b1;
    layer3_outputs(374) <= b and not a;
    layer3_outputs(375) <= not (a and b);
    layer3_outputs(376) <= a and b;
    layer3_outputs(377) <= a and b;
    layer3_outputs(378) <= a xor b;
    layer3_outputs(379) <= a and b;
    layer3_outputs(380) <= 1'b0;
    layer3_outputs(381) <= not (a and b);
    layer3_outputs(382) <= b;
    layer3_outputs(383) <= not (a or b);
    layer3_outputs(384) <= a xor b;
    layer3_outputs(385) <= a;
    layer3_outputs(386) <= b and not a;
    layer3_outputs(387) <= b;
    layer3_outputs(388) <= not b or a;
    layer3_outputs(389) <= a;
    layer3_outputs(390) <= not b or a;
    layer3_outputs(391) <= a and b;
    layer3_outputs(392) <= b and not a;
    layer3_outputs(393) <= not a or b;
    layer3_outputs(394) <= not a or b;
    layer3_outputs(395) <= not b or a;
    layer3_outputs(396) <= 1'b1;
    layer3_outputs(397) <= not a;
    layer3_outputs(398) <= not a;
    layer3_outputs(399) <= b;
    layer3_outputs(400) <= a and b;
    layer3_outputs(401) <= b;
    layer3_outputs(402) <= a or b;
    layer3_outputs(403) <= 1'b0;
    layer3_outputs(404) <= not (a and b);
    layer3_outputs(405) <= not a or b;
    layer3_outputs(406) <= b and not a;
    layer3_outputs(407) <= not a;
    layer3_outputs(408) <= 1'b1;
    layer3_outputs(409) <= b;
    layer3_outputs(410) <= a or b;
    layer3_outputs(411) <= a;
    layer3_outputs(412) <= 1'b0;
    layer3_outputs(413) <= a or b;
    layer3_outputs(414) <= b;
    layer3_outputs(415) <= 1'b0;
    layer3_outputs(416) <= b;
    layer3_outputs(417) <= not b;
    layer3_outputs(418) <= 1'b1;
    layer3_outputs(419) <= a and b;
    layer3_outputs(420) <= b and not a;
    layer3_outputs(421) <= not b or a;
    layer3_outputs(422) <= not (a or b);
    layer3_outputs(423) <= not (a and b);
    layer3_outputs(424) <= a or b;
    layer3_outputs(425) <= b;
    layer3_outputs(426) <= a or b;
    layer3_outputs(427) <= 1'b1;
    layer3_outputs(428) <= not (a or b);
    layer3_outputs(429) <= b and not a;
    layer3_outputs(430) <= a and not b;
    layer3_outputs(431) <= not b or a;
    layer3_outputs(432) <= not a;
    layer3_outputs(433) <= not b or a;
    layer3_outputs(434) <= 1'b1;
    layer3_outputs(435) <= a or b;
    layer3_outputs(436) <= b and not a;
    layer3_outputs(437) <= a and not b;
    layer3_outputs(438) <= not a or b;
    layer3_outputs(439) <= 1'b0;
    layer3_outputs(440) <= not b or a;
    layer3_outputs(441) <= not (a and b);
    layer3_outputs(442) <= 1'b1;
    layer3_outputs(443) <= not a;
    layer3_outputs(444) <= not b or a;
    layer3_outputs(445) <= not b;
    layer3_outputs(446) <= 1'b0;
    layer3_outputs(447) <= not a;
    layer3_outputs(448) <= not (a or b);
    layer3_outputs(449) <= not b;
    layer3_outputs(450) <= 1'b1;
    layer3_outputs(451) <= a;
    layer3_outputs(452) <= 1'b0;
    layer3_outputs(453) <= not a;
    layer3_outputs(454) <= not a;
    layer3_outputs(455) <= b;
    layer3_outputs(456) <= not a or b;
    layer3_outputs(457) <= not b;
    layer3_outputs(458) <= b;
    layer3_outputs(459) <= 1'b1;
    layer3_outputs(460) <= 1'b0;
    layer3_outputs(461) <= not b;
    layer3_outputs(462) <= 1'b0;
    layer3_outputs(463) <= a xor b;
    layer3_outputs(464) <= a and not b;
    layer3_outputs(465) <= a and not b;
    layer3_outputs(466) <= not (a and b);
    layer3_outputs(467) <= not b or a;
    layer3_outputs(468) <= not (a and b);
    layer3_outputs(469) <= 1'b1;
    layer3_outputs(470) <= a or b;
    layer3_outputs(471) <= not a;
    layer3_outputs(472) <= b;
    layer3_outputs(473) <= not b or a;
    layer3_outputs(474) <= 1'b1;
    layer3_outputs(475) <= 1'b0;
    layer3_outputs(476) <= not b;
    layer3_outputs(477) <= b;
    layer3_outputs(478) <= b;
    layer3_outputs(479) <= not b or a;
    layer3_outputs(480) <= a and b;
    layer3_outputs(481) <= a;
    layer3_outputs(482) <= b and not a;
    layer3_outputs(483) <= a and not b;
    layer3_outputs(484) <= not a;
    layer3_outputs(485) <= not (a xor b);
    layer3_outputs(486) <= not b or a;
    layer3_outputs(487) <= not (a or b);
    layer3_outputs(488) <= not (a and b);
    layer3_outputs(489) <= a and b;
    layer3_outputs(490) <= not (a xor b);
    layer3_outputs(491) <= b and not a;
    layer3_outputs(492) <= b and not a;
    layer3_outputs(493) <= 1'b1;
    layer3_outputs(494) <= 1'b0;
    layer3_outputs(495) <= a or b;
    layer3_outputs(496) <= not (a or b);
    layer3_outputs(497) <= not (a and b);
    layer3_outputs(498) <= a or b;
    layer3_outputs(499) <= not (a and b);
    layer3_outputs(500) <= not (a or b);
    layer3_outputs(501) <= 1'b1;
    layer3_outputs(502) <= 1'b0;
    layer3_outputs(503) <= a;
    layer3_outputs(504) <= 1'b0;
    layer3_outputs(505) <= not (a xor b);
    layer3_outputs(506) <= not (a xor b);
    layer3_outputs(507) <= not b or a;
    layer3_outputs(508) <= not b or a;
    layer3_outputs(509) <= not (a xor b);
    layer3_outputs(510) <= 1'b1;
    layer3_outputs(511) <= not (a and b);
    layer3_outputs(512) <= not b;
    layer3_outputs(513) <= b;
    layer3_outputs(514) <= b and not a;
    layer3_outputs(515) <= not b;
    layer3_outputs(516) <= a;
    layer3_outputs(517) <= not (a and b);
    layer3_outputs(518) <= not a;
    layer3_outputs(519) <= not a or b;
    layer3_outputs(520) <= not b;
    layer3_outputs(521) <= 1'b1;
    layer3_outputs(522) <= 1'b0;
    layer3_outputs(523) <= b;
    layer3_outputs(524) <= not a or b;
    layer3_outputs(525) <= a and b;
    layer3_outputs(526) <= a xor b;
    layer3_outputs(527) <= not a;
    layer3_outputs(528) <= b;
    layer3_outputs(529) <= b and not a;
    layer3_outputs(530) <= not a or b;
    layer3_outputs(531) <= not a;
    layer3_outputs(532) <= a;
    layer3_outputs(533) <= not (a and b);
    layer3_outputs(534) <= b;
    layer3_outputs(535) <= not a;
    layer3_outputs(536) <= not a;
    layer3_outputs(537) <= not b;
    layer3_outputs(538) <= 1'b1;
    layer3_outputs(539) <= not b;
    layer3_outputs(540) <= a;
    layer3_outputs(541) <= a and b;
    layer3_outputs(542) <= not a or b;
    layer3_outputs(543) <= 1'b1;
    layer3_outputs(544) <= not (a and b);
    layer3_outputs(545) <= 1'b1;
    layer3_outputs(546) <= a xor b;
    layer3_outputs(547) <= not b or a;
    layer3_outputs(548) <= not (a xor b);
    layer3_outputs(549) <= 1'b0;
    layer3_outputs(550) <= a;
    layer3_outputs(551) <= not b or a;
    layer3_outputs(552) <= a or b;
    layer3_outputs(553) <= not a or b;
    layer3_outputs(554) <= a or b;
    layer3_outputs(555) <= b;
    layer3_outputs(556) <= a;
    layer3_outputs(557) <= a and not b;
    layer3_outputs(558) <= not (a or b);
    layer3_outputs(559) <= not b;
    layer3_outputs(560) <= not a;
    layer3_outputs(561) <= not (a and b);
    layer3_outputs(562) <= not a;
    layer3_outputs(563) <= b;
    layer3_outputs(564) <= not a;
    layer3_outputs(565) <= not b;
    layer3_outputs(566) <= a and b;
    layer3_outputs(567) <= not b or a;
    layer3_outputs(568) <= not (a xor b);
    layer3_outputs(569) <= not a;
    layer3_outputs(570) <= a;
    layer3_outputs(571) <= not b;
    layer3_outputs(572) <= 1'b1;
    layer3_outputs(573) <= not (a or b);
    layer3_outputs(574) <= a and b;
    layer3_outputs(575) <= a and not b;
    layer3_outputs(576) <= not a or b;
    layer3_outputs(577) <= a and not b;
    layer3_outputs(578) <= a and b;
    layer3_outputs(579) <= a and b;
    layer3_outputs(580) <= not a or b;
    layer3_outputs(581) <= not (a or b);
    layer3_outputs(582) <= not b;
    layer3_outputs(583) <= a or b;
    layer3_outputs(584) <= a xor b;
    layer3_outputs(585) <= b and not a;
    layer3_outputs(586) <= b;
    layer3_outputs(587) <= a;
    layer3_outputs(588) <= a and b;
    layer3_outputs(589) <= not a;
    layer3_outputs(590) <= not (a or b);
    layer3_outputs(591) <= not (a or b);
    layer3_outputs(592) <= b;
    layer3_outputs(593) <= not (a and b);
    layer3_outputs(594) <= not a;
    layer3_outputs(595) <= not (a or b);
    layer3_outputs(596) <= not (a and b);
    layer3_outputs(597) <= a and b;
    layer3_outputs(598) <= b;
    layer3_outputs(599) <= not (a and b);
    layer3_outputs(600) <= b and not a;
    layer3_outputs(601) <= not b;
    layer3_outputs(602) <= b;
    layer3_outputs(603) <= not (a or b);
    layer3_outputs(604) <= not b or a;
    layer3_outputs(605) <= 1'b0;
    layer3_outputs(606) <= a and b;
    layer3_outputs(607) <= b and not a;
    layer3_outputs(608) <= b;
    layer3_outputs(609) <= 1'b0;
    layer3_outputs(610) <= not (a xor b);
    layer3_outputs(611) <= not (a and b);
    layer3_outputs(612) <= not (a and b);
    layer3_outputs(613) <= not b;
    layer3_outputs(614) <= b;
    layer3_outputs(615) <= 1'b1;
    layer3_outputs(616) <= not (a or b);
    layer3_outputs(617) <= 1'b1;
    layer3_outputs(618) <= 1'b1;
    layer3_outputs(619) <= not b or a;
    layer3_outputs(620) <= not (a or b);
    layer3_outputs(621) <= not b or a;
    layer3_outputs(622) <= 1'b1;
    layer3_outputs(623) <= a and b;
    layer3_outputs(624) <= b;
    layer3_outputs(625) <= a;
    layer3_outputs(626) <= b and not a;
    layer3_outputs(627) <= b;
    layer3_outputs(628) <= not b or a;
    layer3_outputs(629) <= not (a and b);
    layer3_outputs(630) <= not b;
    layer3_outputs(631) <= a or b;
    layer3_outputs(632) <= not (a and b);
    layer3_outputs(633) <= not a;
    layer3_outputs(634) <= a and b;
    layer3_outputs(635) <= not (a or b);
    layer3_outputs(636) <= b;
    layer3_outputs(637) <= b and not a;
    layer3_outputs(638) <= b;
    layer3_outputs(639) <= a or b;
    layer3_outputs(640) <= a xor b;
    layer3_outputs(641) <= not b;
    layer3_outputs(642) <= a or b;
    layer3_outputs(643) <= 1'b0;
    layer3_outputs(644) <= not a;
    layer3_outputs(645) <= not b or a;
    layer3_outputs(646) <= not (a or b);
    layer3_outputs(647) <= not b or a;
    layer3_outputs(648) <= b;
    layer3_outputs(649) <= not a or b;
    layer3_outputs(650) <= b;
    layer3_outputs(651) <= b and not a;
    layer3_outputs(652) <= b;
    layer3_outputs(653) <= a;
    layer3_outputs(654) <= not a or b;
    layer3_outputs(655) <= not (a or b);
    layer3_outputs(656) <= a;
    layer3_outputs(657) <= 1'b1;
    layer3_outputs(658) <= not a;
    layer3_outputs(659) <= 1'b0;
    layer3_outputs(660) <= not (a xor b);
    layer3_outputs(661) <= 1'b0;
    layer3_outputs(662) <= b;
    layer3_outputs(663) <= a and b;
    layer3_outputs(664) <= 1'b1;
    layer3_outputs(665) <= not (a and b);
    layer3_outputs(666) <= a;
    layer3_outputs(667) <= not a or b;
    layer3_outputs(668) <= b;
    layer3_outputs(669) <= not b or a;
    layer3_outputs(670) <= not b or a;
    layer3_outputs(671) <= 1'b1;
    layer3_outputs(672) <= not a or b;
    layer3_outputs(673) <= a and not b;
    layer3_outputs(674) <= a;
    layer3_outputs(675) <= 1'b1;
    layer3_outputs(676) <= 1'b1;
    layer3_outputs(677) <= not (a xor b);
    layer3_outputs(678) <= a or b;
    layer3_outputs(679) <= not a or b;
    layer3_outputs(680) <= 1'b0;
    layer3_outputs(681) <= 1'b0;
    layer3_outputs(682) <= not a or b;
    layer3_outputs(683) <= a;
    layer3_outputs(684) <= b;
    layer3_outputs(685) <= a xor b;
    layer3_outputs(686) <= 1'b0;
    layer3_outputs(687) <= not (a or b);
    layer3_outputs(688) <= not (a and b);
    layer3_outputs(689) <= a;
    layer3_outputs(690) <= 1'b0;
    layer3_outputs(691) <= not a or b;
    layer3_outputs(692) <= b;
    layer3_outputs(693) <= a and b;
    layer3_outputs(694) <= not a or b;
    layer3_outputs(695) <= not (a or b);
    layer3_outputs(696) <= not b or a;
    layer3_outputs(697) <= not (a xor b);
    layer3_outputs(698) <= a xor b;
    layer3_outputs(699) <= 1'b0;
    layer3_outputs(700) <= a and not b;
    layer3_outputs(701) <= a and not b;
    layer3_outputs(702) <= a;
    layer3_outputs(703) <= a xor b;
    layer3_outputs(704) <= a and b;
    layer3_outputs(705) <= a and b;
    layer3_outputs(706) <= not b or a;
    layer3_outputs(707) <= b;
    layer3_outputs(708) <= 1'b0;
    layer3_outputs(709) <= a;
    layer3_outputs(710) <= a or b;
    layer3_outputs(711) <= not b or a;
    layer3_outputs(712) <= a or b;
    layer3_outputs(713) <= not (a xor b);
    layer3_outputs(714) <= a or b;
    layer3_outputs(715) <= not (a and b);
    layer3_outputs(716) <= a;
    layer3_outputs(717) <= 1'b0;
    layer3_outputs(718) <= a or b;
    layer3_outputs(719) <= a or b;
    layer3_outputs(720) <= not b;
    layer3_outputs(721) <= not a or b;
    layer3_outputs(722) <= not (a or b);
    layer3_outputs(723) <= not b or a;
    layer3_outputs(724) <= a and not b;
    layer3_outputs(725) <= a;
    layer3_outputs(726) <= a;
    layer3_outputs(727) <= a and b;
    layer3_outputs(728) <= a or b;
    layer3_outputs(729) <= a;
    layer3_outputs(730) <= not (a or b);
    layer3_outputs(731) <= a and not b;
    layer3_outputs(732) <= a and not b;
    layer3_outputs(733) <= 1'b1;
    layer3_outputs(734) <= not (a and b);
    layer3_outputs(735) <= a;
    layer3_outputs(736) <= b;
    layer3_outputs(737) <= not b;
    layer3_outputs(738) <= not a;
    layer3_outputs(739) <= b and not a;
    layer3_outputs(740) <= not b or a;
    layer3_outputs(741) <= not (a or b);
    layer3_outputs(742) <= a and b;
    layer3_outputs(743) <= a and not b;
    layer3_outputs(744) <= not b or a;
    layer3_outputs(745) <= not a or b;
    layer3_outputs(746) <= not (a and b);
    layer3_outputs(747) <= not b;
    layer3_outputs(748) <= a and b;
    layer3_outputs(749) <= not (a and b);
    layer3_outputs(750) <= a;
    layer3_outputs(751) <= a and not b;
    layer3_outputs(752) <= not a;
    layer3_outputs(753) <= not a;
    layer3_outputs(754) <= b;
    layer3_outputs(755) <= not a;
    layer3_outputs(756) <= not a;
    layer3_outputs(757) <= 1'b0;
    layer3_outputs(758) <= b;
    layer3_outputs(759) <= a or b;
    layer3_outputs(760) <= not b or a;
    layer3_outputs(761) <= a and not b;
    layer3_outputs(762) <= a;
    layer3_outputs(763) <= 1'b1;
    layer3_outputs(764) <= a or b;
    layer3_outputs(765) <= 1'b1;
    layer3_outputs(766) <= a;
    layer3_outputs(767) <= not b;
    layer3_outputs(768) <= 1'b0;
    layer3_outputs(769) <= not a or b;
    layer3_outputs(770) <= a or b;
    layer3_outputs(771) <= not a or b;
    layer3_outputs(772) <= a and b;
    layer3_outputs(773) <= not (a or b);
    layer3_outputs(774) <= a or b;
    layer3_outputs(775) <= not b;
    layer3_outputs(776) <= a and not b;
    layer3_outputs(777) <= not (a or b);
    layer3_outputs(778) <= not b;
    layer3_outputs(779) <= not a or b;
    layer3_outputs(780) <= not (a and b);
    layer3_outputs(781) <= not (a and b);
    layer3_outputs(782) <= 1'b1;
    layer3_outputs(783) <= a xor b;
    layer3_outputs(784) <= 1'b1;
    layer3_outputs(785) <= a and b;
    layer3_outputs(786) <= b and not a;
    layer3_outputs(787) <= not a or b;
    layer3_outputs(788) <= a and b;
    layer3_outputs(789) <= a and b;
    layer3_outputs(790) <= not (a and b);
    layer3_outputs(791) <= not (a xor b);
    layer3_outputs(792) <= 1'b0;
    layer3_outputs(793) <= not a or b;
    layer3_outputs(794) <= a and b;
    layer3_outputs(795) <= not b;
    layer3_outputs(796) <= a or b;
    layer3_outputs(797) <= not a;
    layer3_outputs(798) <= a and not b;
    layer3_outputs(799) <= not b;
    layer3_outputs(800) <= not (a xor b);
    layer3_outputs(801) <= 1'b0;
    layer3_outputs(802) <= a and b;
    layer3_outputs(803) <= not a;
    layer3_outputs(804) <= b and not a;
    layer3_outputs(805) <= 1'b1;
    layer3_outputs(806) <= not a;
    layer3_outputs(807) <= not (a or b);
    layer3_outputs(808) <= not b;
    layer3_outputs(809) <= a;
    layer3_outputs(810) <= not b;
    layer3_outputs(811) <= 1'b1;
    layer3_outputs(812) <= not (a or b);
    layer3_outputs(813) <= b;
    layer3_outputs(814) <= not b or a;
    layer3_outputs(815) <= a;
    layer3_outputs(816) <= b and not a;
    layer3_outputs(817) <= not (a and b);
    layer3_outputs(818) <= not b;
    layer3_outputs(819) <= not (a or b);
    layer3_outputs(820) <= not (a and b);
    layer3_outputs(821) <= b and not a;
    layer3_outputs(822) <= a and b;
    layer3_outputs(823) <= not b or a;
    layer3_outputs(824) <= 1'b0;
    layer3_outputs(825) <= a or b;
    layer3_outputs(826) <= 1'b1;
    layer3_outputs(827) <= a and not b;
    layer3_outputs(828) <= not b;
    layer3_outputs(829) <= 1'b0;
    layer3_outputs(830) <= 1'b1;
    layer3_outputs(831) <= 1'b0;
    layer3_outputs(832) <= b;
    layer3_outputs(833) <= a;
    layer3_outputs(834) <= not (a and b);
    layer3_outputs(835) <= 1'b0;
    layer3_outputs(836) <= 1'b0;
    layer3_outputs(837) <= not b;
    layer3_outputs(838) <= not (a and b);
    layer3_outputs(839) <= a and b;
    layer3_outputs(840) <= a or b;
    layer3_outputs(841) <= a;
    layer3_outputs(842) <= a;
    layer3_outputs(843) <= a or b;
    layer3_outputs(844) <= a xor b;
    layer3_outputs(845) <= b and not a;
    layer3_outputs(846) <= b and not a;
    layer3_outputs(847) <= not a or b;
    layer3_outputs(848) <= not b;
    layer3_outputs(849) <= a or b;
    layer3_outputs(850) <= b;
    layer3_outputs(851) <= not (a and b);
    layer3_outputs(852) <= b and not a;
    layer3_outputs(853) <= not a;
    layer3_outputs(854) <= not (a xor b);
    layer3_outputs(855) <= not b or a;
    layer3_outputs(856) <= not a or b;
    layer3_outputs(857) <= not a or b;
    layer3_outputs(858) <= b;
    layer3_outputs(859) <= a;
    layer3_outputs(860) <= a and b;
    layer3_outputs(861) <= not (a or b);
    layer3_outputs(862) <= not b or a;
    layer3_outputs(863) <= not (a or b);
    layer3_outputs(864) <= not a;
    layer3_outputs(865) <= not b;
    layer3_outputs(866) <= not a or b;
    layer3_outputs(867) <= a or b;
    layer3_outputs(868) <= a;
    layer3_outputs(869) <= a xor b;
    layer3_outputs(870) <= a;
    layer3_outputs(871) <= not a or b;
    layer3_outputs(872) <= not b;
    layer3_outputs(873) <= a;
    layer3_outputs(874) <= 1'b0;
    layer3_outputs(875) <= not a;
    layer3_outputs(876) <= not (a and b);
    layer3_outputs(877) <= a xor b;
    layer3_outputs(878) <= not (a and b);
    layer3_outputs(879) <= not b;
    layer3_outputs(880) <= not a;
    layer3_outputs(881) <= not a;
    layer3_outputs(882) <= not b;
    layer3_outputs(883) <= a;
    layer3_outputs(884) <= a;
    layer3_outputs(885) <= 1'b1;
    layer3_outputs(886) <= not a;
    layer3_outputs(887) <= not b or a;
    layer3_outputs(888) <= not a;
    layer3_outputs(889) <= b;
    layer3_outputs(890) <= not (a or b);
    layer3_outputs(891) <= a and not b;
    layer3_outputs(892) <= b and not a;
    layer3_outputs(893) <= not a or b;
    layer3_outputs(894) <= a and not b;
    layer3_outputs(895) <= a and not b;
    layer3_outputs(896) <= a;
    layer3_outputs(897) <= not (a or b);
    layer3_outputs(898) <= 1'b0;
    layer3_outputs(899) <= a;
    layer3_outputs(900) <= a;
    layer3_outputs(901) <= 1'b1;
    layer3_outputs(902) <= b;
    layer3_outputs(903) <= a;
    layer3_outputs(904) <= b;
    layer3_outputs(905) <= not (a and b);
    layer3_outputs(906) <= not a;
    layer3_outputs(907) <= a;
    layer3_outputs(908) <= not a or b;
    layer3_outputs(909) <= not b;
    layer3_outputs(910) <= a;
    layer3_outputs(911) <= a;
    layer3_outputs(912) <= not b or a;
    layer3_outputs(913) <= not a or b;
    layer3_outputs(914) <= not (a or b);
    layer3_outputs(915) <= a;
    layer3_outputs(916) <= a or b;
    layer3_outputs(917) <= a and not b;
    layer3_outputs(918) <= a and b;
    layer3_outputs(919) <= a or b;
    layer3_outputs(920) <= not (a or b);
    layer3_outputs(921) <= not b;
    layer3_outputs(922) <= not a;
    layer3_outputs(923) <= not (a and b);
    layer3_outputs(924) <= a or b;
    layer3_outputs(925) <= not a or b;
    layer3_outputs(926) <= a;
    layer3_outputs(927) <= not a or b;
    layer3_outputs(928) <= 1'b0;
    layer3_outputs(929) <= not b or a;
    layer3_outputs(930) <= a and not b;
    layer3_outputs(931) <= a and not b;
    layer3_outputs(932) <= b and not a;
    layer3_outputs(933) <= not (a or b);
    layer3_outputs(934) <= not b;
    layer3_outputs(935) <= 1'b0;
    layer3_outputs(936) <= not b or a;
    layer3_outputs(937) <= a and not b;
    layer3_outputs(938) <= a or b;
    layer3_outputs(939) <= not (a and b);
    layer3_outputs(940) <= not a or b;
    layer3_outputs(941) <= not (a and b);
    layer3_outputs(942) <= b;
    layer3_outputs(943) <= a;
    layer3_outputs(944) <= not b;
    layer3_outputs(945) <= not b or a;
    layer3_outputs(946) <= not (a and b);
    layer3_outputs(947) <= a;
    layer3_outputs(948) <= not (a or b);
    layer3_outputs(949) <= a and not b;
    layer3_outputs(950) <= b and not a;
    layer3_outputs(951) <= not (a xor b);
    layer3_outputs(952) <= a and not b;
    layer3_outputs(953) <= not a or b;
    layer3_outputs(954) <= 1'b1;
    layer3_outputs(955) <= not (a and b);
    layer3_outputs(956) <= b;
    layer3_outputs(957) <= a or b;
    layer3_outputs(958) <= not b or a;
    layer3_outputs(959) <= not a or b;
    layer3_outputs(960) <= a and b;
    layer3_outputs(961) <= not (a or b);
    layer3_outputs(962) <= not a or b;
    layer3_outputs(963) <= not a;
    layer3_outputs(964) <= b;
    layer3_outputs(965) <= a and not b;
    layer3_outputs(966) <= b;
    layer3_outputs(967) <= 1'b1;
    layer3_outputs(968) <= 1'b1;
    layer3_outputs(969) <= a and b;
    layer3_outputs(970) <= not (a or b);
    layer3_outputs(971) <= not a;
    layer3_outputs(972) <= not a or b;
    layer3_outputs(973) <= not (a xor b);
    layer3_outputs(974) <= a or b;
    layer3_outputs(975) <= not b or a;
    layer3_outputs(976) <= not a;
    layer3_outputs(977) <= 1'b0;
    layer3_outputs(978) <= a and not b;
    layer3_outputs(979) <= not a or b;
    layer3_outputs(980) <= not b;
    layer3_outputs(981) <= not b;
    layer3_outputs(982) <= a and not b;
    layer3_outputs(983) <= a and b;
    layer3_outputs(984) <= a;
    layer3_outputs(985) <= not a;
    layer3_outputs(986) <= not (a and b);
    layer3_outputs(987) <= not (a or b);
    layer3_outputs(988) <= not (a and b);
    layer3_outputs(989) <= not b or a;
    layer3_outputs(990) <= not (a and b);
    layer3_outputs(991) <= a;
    layer3_outputs(992) <= b and not a;
    layer3_outputs(993) <= a xor b;
    layer3_outputs(994) <= not a or b;
    layer3_outputs(995) <= not a;
    layer3_outputs(996) <= not (a and b);
    layer3_outputs(997) <= not (a and b);
    layer3_outputs(998) <= a and not b;
    layer3_outputs(999) <= not (a and b);
    layer3_outputs(1000) <= not (a xor b);
    layer3_outputs(1001) <= not b;
    layer3_outputs(1002) <= a;
    layer3_outputs(1003) <= not b;
    layer3_outputs(1004) <= not b or a;
    layer3_outputs(1005) <= not (a or b);
    layer3_outputs(1006) <= b;
    layer3_outputs(1007) <= not (a and b);
    layer3_outputs(1008) <= not (a and b);
    layer3_outputs(1009) <= 1'b0;
    layer3_outputs(1010) <= a xor b;
    layer3_outputs(1011) <= a and not b;
    layer3_outputs(1012) <= 1'b1;
    layer3_outputs(1013) <= 1'b0;
    layer3_outputs(1014) <= not (a and b);
    layer3_outputs(1015) <= not (a and b);
    layer3_outputs(1016) <= 1'b1;
    layer3_outputs(1017) <= a;
    layer3_outputs(1018) <= b;
    layer3_outputs(1019) <= not (a xor b);
    layer3_outputs(1020) <= b and not a;
    layer3_outputs(1021) <= not a;
    layer3_outputs(1022) <= b and not a;
    layer3_outputs(1023) <= not (a and b);
    layer3_outputs(1024) <= a and b;
    layer3_outputs(1025) <= not b;
    layer3_outputs(1026) <= b;
    layer3_outputs(1027) <= not a or b;
    layer3_outputs(1028) <= a and b;
    layer3_outputs(1029) <= a or b;
    layer3_outputs(1030) <= not b;
    layer3_outputs(1031) <= not b;
    layer3_outputs(1032) <= not (a or b);
    layer3_outputs(1033) <= a or b;
    layer3_outputs(1034) <= not b;
    layer3_outputs(1035) <= not (a and b);
    layer3_outputs(1036) <= a and b;
    layer3_outputs(1037) <= 1'b0;
    layer3_outputs(1038) <= a;
    layer3_outputs(1039) <= not a;
    layer3_outputs(1040) <= 1'b0;
    layer3_outputs(1041) <= a and not b;
    layer3_outputs(1042) <= a or b;
    layer3_outputs(1043) <= 1'b1;
    layer3_outputs(1044) <= b and not a;
    layer3_outputs(1045) <= not b;
    layer3_outputs(1046) <= b and not a;
    layer3_outputs(1047) <= not a;
    layer3_outputs(1048) <= not a or b;
    layer3_outputs(1049) <= a and b;
    layer3_outputs(1050) <= b and not a;
    layer3_outputs(1051) <= a;
    layer3_outputs(1052) <= not b;
    layer3_outputs(1053) <= a and not b;
    layer3_outputs(1054) <= a and not b;
    layer3_outputs(1055) <= not b or a;
    layer3_outputs(1056) <= a or b;
    layer3_outputs(1057) <= not b or a;
    layer3_outputs(1058) <= b and not a;
    layer3_outputs(1059) <= not (a and b);
    layer3_outputs(1060) <= a and not b;
    layer3_outputs(1061) <= a;
    layer3_outputs(1062) <= 1'b0;
    layer3_outputs(1063) <= b;
    layer3_outputs(1064) <= 1'b1;
    layer3_outputs(1065) <= not b or a;
    layer3_outputs(1066) <= 1'b0;
    layer3_outputs(1067) <= b and not a;
    layer3_outputs(1068) <= a or b;
    layer3_outputs(1069) <= not b;
    layer3_outputs(1070) <= b;
    layer3_outputs(1071) <= not a or b;
    layer3_outputs(1072) <= not a;
    layer3_outputs(1073) <= a and b;
    layer3_outputs(1074) <= a and b;
    layer3_outputs(1075) <= not (a and b);
    layer3_outputs(1076) <= not a;
    layer3_outputs(1077) <= a xor b;
    layer3_outputs(1078) <= a or b;
    layer3_outputs(1079) <= not a or b;
    layer3_outputs(1080) <= not b;
    layer3_outputs(1081) <= not (a and b);
    layer3_outputs(1082) <= b;
    layer3_outputs(1083) <= b;
    layer3_outputs(1084) <= 1'b1;
    layer3_outputs(1085) <= 1'b0;
    layer3_outputs(1086) <= a and not b;
    layer3_outputs(1087) <= b;
    layer3_outputs(1088) <= not (a and b);
    layer3_outputs(1089) <= a and b;
    layer3_outputs(1090) <= not a or b;
    layer3_outputs(1091) <= not a;
    layer3_outputs(1092) <= not a or b;
    layer3_outputs(1093) <= a and not b;
    layer3_outputs(1094) <= b;
    layer3_outputs(1095) <= 1'b0;
    layer3_outputs(1096) <= not (a and b);
    layer3_outputs(1097) <= 1'b0;
    layer3_outputs(1098) <= 1'b1;
    layer3_outputs(1099) <= 1'b1;
    layer3_outputs(1100) <= not a;
    layer3_outputs(1101) <= a or b;
    layer3_outputs(1102) <= a;
    layer3_outputs(1103) <= not b;
    layer3_outputs(1104) <= b;
    layer3_outputs(1105) <= not (a and b);
    layer3_outputs(1106) <= 1'b1;
    layer3_outputs(1107) <= not a;
    layer3_outputs(1108) <= 1'b1;
    layer3_outputs(1109) <= b;
    layer3_outputs(1110) <= a and not b;
    layer3_outputs(1111) <= not a;
    layer3_outputs(1112) <= not (a and b);
    layer3_outputs(1113) <= 1'b1;
    layer3_outputs(1114) <= a;
    layer3_outputs(1115) <= a or b;
    layer3_outputs(1116) <= a and b;
    layer3_outputs(1117) <= not a;
    layer3_outputs(1118) <= a and b;
    layer3_outputs(1119) <= 1'b1;
    layer3_outputs(1120) <= b and not a;
    layer3_outputs(1121) <= not a;
    layer3_outputs(1122) <= not (a or b);
    layer3_outputs(1123) <= a or b;
    layer3_outputs(1124) <= b;
    layer3_outputs(1125) <= a;
    layer3_outputs(1126) <= not a;
    layer3_outputs(1127) <= 1'b0;
    layer3_outputs(1128) <= 1'b0;
    layer3_outputs(1129) <= not b or a;
    layer3_outputs(1130) <= a;
    layer3_outputs(1131) <= not a or b;
    layer3_outputs(1132) <= not (a and b);
    layer3_outputs(1133) <= a;
    layer3_outputs(1134) <= a and not b;
    layer3_outputs(1135) <= not (a or b);
    layer3_outputs(1136) <= not b;
    layer3_outputs(1137) <= 1'b1;
    layer3_outputs(1138) <= 1'b1;
    layer3_outputs(1139) <= not (a and b);
    layer3_outputs(1140) <= not a or b;
    layer3_outputs(1141) <= not a;
    layer3_outputs(1142) <= a and not b;
    layer3_outputs(1143) <= not a;
    layer3_outputs(1144) <= 1'b0;
    layer3_outputs(1145) <= not b;
    layer3_outputs(1146) <= not (a and b);
    layer3_outputs(1147) <= a and not b;
    layer3_outputs(1148) <= 1'b0;
    layer3_outputs(1149) <= not a;
    layer3_outputs(1150) <= not (a or b);
    layer3_outputs(1151) <= not a;
    layer3_outputs(1152) <= a or b;
    layer3_outputs(1153) <= a and b;
    layer3_outputs(1154) <= not b;
    layer3_outputs(1155) <= a and not b;
    layer3_outputs(1156) <= a and b;
    layer3_outputs(1157) <= not (a or b);
    layer3_outputs(1158) <= 1'b1;
    layer3_outputs(1159) <= not b;
    layer3_outputs(1160) <= a and b;
    layer3_outputs(1161) <= a and not b;
    layer3_outputs(1162) <= not (a or b);
    layer3_outputs(1163) <= not a;
    layer3_outputs(1164) <= not (a xor b);
    layer3_outputs(1165) <= a and not b;
    layer3_outputs(1166) <= not a or b;
    layer3_outputs(1167) <= 1'b0;
    layer3_outputs(1168) <= a and b;
    layer3_outputs(1169) <= a and not b;
    layer3_outputs(1170) <= not (a or b);
    layer3_outputs(1171) <= a and b;
    layer3_outputs(1172) <= not (a or b);
    layer3_outputs(1173) <= 1'b0;
    layer3_outputs(1174) <= not a or b;
    layer3_outputs(1175) <= not a or b;
    layer3_outputs(1176) <= 1'b0;
    layer3_outputs(1177) <= 1'b1;
    layer3_outputs(1178) <= a;
    layer3_outputs(1179) <= 1'b1;
    layer3_outputs(1180) <= not (a and b);
    layer3_outputs(1181) <= not (a or b);
    layer3_outputs(1182) <= not b;
    layer3_outputs(1183) <= a or b;
    layer3_outputs(1184) <= not (a or b);
    layer3_outputs(1185) <= 1'b1;
    layer3_outputs(1186) <= not b;
    layer3_outputs(1187) <= b;
    layer3_outputs(1188) <= not a or b;
    layer3_outputs(1189) <= not b;
    layer3_outputs(1190) <= a and b;
    layer3_outputs(1191) <= a and not b;
    layer3_outputs(1192) <= a or b;
    layer3_outputs(1193) <= a and not b;
    layer3_outputs(1194) <= a;
    layer3_outputs(1195) <= a and not b;
    layer3_outputs(1196) <= not (a and b);
    layer3_outputs(1197) <= not a or b;
    layer3_outputs(1198) <= not a;
    layer3_outputs(1199) <= not a or b;
    layer3_outputs(1200) <= not b;
    layer3_outputs(1201) <= not a or b;
    layer3_outputs(1202) <= b;
    layer3_outputs(1203) <= not (a and b);
    layer3_outputs(1204) <= 1'b1;
    layer3_outputs(1205) <= not a or b;
    layer3_outputs(1206) <= a or b;
    layer3_outputs(1207) <= a and b;
    layer3_outputs(1208) <= 1'b1;
    layer3_outputs(1209) <= a xor b;
    layer3_outputs(1210) <= a and b;
    layer3_outputs(1211) <= 1'b1;
    layer3_outputs(1212) <= not (a or b);
    layer3_outputs(1213) <= not a;
    layer3_outputs(1214) <= b and not a;
    layer3_outputs(1215) <= a and not b;
    layer3_outputs(1216) <= 1'b1;
    layer3_outputs(1217) <= 1'b0;
    layer3_outputs(1218) <= not a;
    layer3_outputs(1219) <= 1'b0;
    layer3_outputs(1220) <= not (a or b);
    layer3_outputs(1221) <= not (a or b);
    layer3_outputs(1222) <= not b;
    layer3_outputs(1223) <= not b or a;
    layer3_outputs(1224) <= a or b;
    layer3_outputs(1225) <= not b or a;
    layer3_outputs(1226) <= not (a xor b);
    layer3_outputs(1227) <= 1'b1;
    layer3_outputs(1228) <= b;
    layer3_outputs(1229) <= 1'b1;
    layer3_outputs(1230) <= not b;
    layer3_outputs(1231) <= a and b;
    layer3_outputs(1232) <= 1'b1;
    layer3_outputs(1233) <= a and not b;
    layer3_outputs(1234) <= not a;
    layer3_outputs(1235) <= 1'b1;
    layer3_outputs(1236) <= not (a and b);
    layer3_outputs(1237) <= a or b;
    layer3_outputs(1238) <= 1'b0;
    layer3_outputs(1239) <= a;
    layer3_outputs(1240) <= a;
    layer3_outputs(1241) <= not a or b;
    layer3_outputs(1242) <= a or b;
    layer3_outputs(1243) <= b and not a;
    layer3_outputs(1244) <= a;
    layer3_outputs(1245) <= not (a and b);
    layer3_outputs(1246) <= a;
    layer3_outputs(1247) <= b and not a;
    layer3_outputs(1248) <= a and b;
    layer3_outputs(1249) <= b;
    layer3_outputs(1250) <= not (a or b);
    layer3_outputs(1251) <= a and b;
    layer3_outputs(1252) <= not a or b;
    layer3_outputs(1253) <= not (a and b);
    layer3_outputs(1254) <= 1'b1;
    layer3_outputs(1255) <= not b;
    layer3_outputs(1256) <= not a or b;
    layer3_outputs(1257) <= 1'b1;
    layer3_outputs(1258) <= not (a or b);
    layer3_outputs(1259) <= a or b;
    layer3_outputs(1260) <= a and b;
    layer3_outputs(1261) <= a and b;
    layer3_outputs(1262) <= 1'b0;
    layer3_outputs(1263) <= 1'b1;
    layer3_outputs(1264) <= not a;
    layer3_outputs(1265) <= not b or a;
    layer3_outputs(1266) <= 1'b1;
    layer3_outputs(1267) <= a;
    layer3_outputs(1268) <= not a;
    layer3_outputs(1269) <= not a or b;
    layer3_outputs(1270) <= a;
    layer3_outputs(1271) <= b;
    layer3_outputs(1272) <= a and not b;
    layer3_outputs(1273) <= a and b;
    layer3_outputs(1274) <= a and not b;
    layer3_outputs(1275) <= a and not b;
    layer3_outputs(1276) <= a;
    layer3_outputs(1277) <= a and b;
    layer3_outputs(1278) <= not (a or b);
    layer3_outputs(1279) <= 1'b1;
    layer3_outputs(1280) <= b;
    layer3_outputs(1281) <= 1'b1;
    layer3_outputs(1282) <= a and b;
    layer3_outputs(1283) <= 1'b1;
    layer3_outputs(1284) <= not b;
    layer3_outputs(1285) <= not a or b;
    layer3_outputs(1286) <= not a;
    layer3_outputs(1287) <= not (a or b);
    layer3_outputs(1288) <= not (a xor b);
    layer3_outputs(1289) <= a and not b;
    layer3_outputs(1290) <= b and not a;
    layer3_outputs(1291) <= a xor b;
    layer3_outputs(1292) <= 1'b1;
    layer3_outputs(1293) <= 1'b1;
    layer3_outputs(1294) <= a and b;
    layer3_outputs(1295) <= b and not a;
    layer3_outputs(1296) <= not b or a;
    layer3_outputs(1297) <= b and not a;
    layer3_outputs(1298) <= 1'b0;
    layer3_outputs(1299) <= a and not b;
    layer3_outputs(1300) <= not a;
    layer3_outputs(1301) <= a;
    layer3_outputs(1302) <= not b or a;
    layer3_outputs(1303) <= not (a or b);
    layer3_outputs(1304) <= not a or b;
    layer3_outputs(1305) <= not a or b;
    layer3_outputs(1306) <= not (a and b);
    layer3_outputs(1307) <= a or b;
    layer3_outputs(1308) <= a xor b;
    layer3_outputs(1309) <= not (a xor b);
    layer3_outputs(1310) <= 1'b0;
    layer3_outputs(1311) <= a;
    layer3_outputs(1312) <= not a;
    layer3_outputs(1313) <= b;
    layer3_outputs(1314) <= a or b;
    layer3_outputs(1315) <= 1'b0;
    layer3_outputs(1316) <= a or b;
    layer3_outputs(1317) <= not b or a;
    layer3_outputs(1318) <= a and not b;
    layer3_outputs(1319) <= 1'b1;
    layer3_outputs(1320) <= a and b;
    layer3_outputs(1321) <= not a or b;
    layer3_outputs(1322) <= 1'b0;
    layer3_outputs(1323) <= b and not a;
    layer3_outputs(1324) <= not (a xor b);
    layer3_outputs(1325) <= a and not b;
    layer3_outputs(1326) <= a;
    layer3_outputs(1327) <= a or b;
    layer3_outputs(1328) <= not a;
    layer3_outputs(1329) <= a;
    layer3_outputs(1330) <= not (a and b);
    layer3_outputs(1331) <= b;
    layer3_outputs(1332) <= a or b;
    layer3_outputs(1333) <= not b or a;
    layer3_outputs(1334) <= not (a or b);
    layer3_outputs(1335) <= not a or b;
    layer3_outputs(1336) <= 1'b0;
    layer3_outputs(1337) <= not (a xor b);
    layer3_outputs(1338) <= not b;
    layer3_outputs(1339) <= not b or a;
    layer3_outputs(1340) <= not a;
    layer3_outputs(1341) <= not (a xor b);
    layer3_outputs(1342) <= not (a and b);
    layer3_outputs(1343) <= a or b;
    layer3_outputs(1344) <= 1'b1;
    layer3_outputs(1345) <= a or b;
    layer3_outputs(1346) <= not (a or b);
    layer3_outputs(1347) <= 1'b0;
    layer3_outputs(1348) <= 1'b1;
    layer3_outputs(1349) <= not (a and b);
    layer3_outputs(1350) <= b and not a;
    layer3_outputs(1351) <= not b or a;
    layer3_outputs(1352) <= not a or b;
    layer3_outputs(1353) <= not b or a;
    layer3_outputs(1354) <= a and not b;
    layer3_outputs(1355) <= not (a or b);
    layer3_outputs(1356) <= not b;
    layer3_outputs(1357) <= not (a or b);
    layer3_outputs(1358) <= not (a or b);
    layer3_outputs(1359) <= a and b;
    layer3_outputs(1360) <= 1'b0;
    layer3_outputs(1361) <= not (a and b);
    layer3_outputs(1362) <= not (a and b);
    layer3_outputs(1363) <= a;
    layer3_outputs(1364) <= a;
    layer3_outputs(1365) <= a;
    layer3_outputs(1366) <= not (a or b);
    layer3_outputs(1367) <= not (a or b);
    layer3_outputs(1368) <= a and b;
    layer3_outputs(1369) <= b and not a;
    layer3_outputs(1370) <= a and not b;
    layer3_outputs(1371) <= not a or b;
    layer3_outputs(1372) <= 1'b1;
    layer3_outputs(1373) <= a or b;
    layer3_outputs(1374) <= not (a xor b);
    layer3_outputs(1375) <= not (a and b);
    layer3_outputs(1376) <= b;
    layer3_outputs(1377) <= not a;
    layer3_outputs(1378) <= not (a or b);
    layer3_outputs(1379) <= not a;
    layer3_outputs(1380) <= not (a xor b);
    layer3_outputs(1381) <= a;
    layer3_outputs(1382) <= not (a or b);
    layer3_outputs(1383) <= b and not a;
    layer3_outputs(1384) <= not b or a;
    layer3_outputs(1385) <= not b;
    layer3_outputs(1386) <= not (a and b);
    layer3_outputs(1387) <= a or b;
    layer3_outputs(1388) <= not a;
    layer3_outputs(1389) <= not b or a;
    layer3_outputs(1390) <= a;
    layer3_outputs(1391) <= not (a xor b);
    layer3_outputs(1392) <= not a or b;
    layer3_outputs(1393) <= not a;
    layer3_outputs(1394) <= b and not a;
    layer3_outputs(1395) <= b and not a;
    layer3_outputs(1396) <= b;
    layer3_outputs(1397) <= a;
    layer3_outputs(1398) <= not b or a;
    layer3_outputs(1399) <= not (a and b);
    layer3_outputs(1400) <= not a;
    layer3_outputs(1401) <= not (a and b);
    layer3_outputs(1402) <= not a or b;
    layer3_outputs(1403) <= b and not a;
    layer3_outputs(1404) <= not (a or b);
    layer3_outputs(1405) <= not a or b;
    layer3_outputs(1406) <= not a;
    layer3_outputs(1407) <= not b or a;
    layer3_outputs(1408) <= not b;
    layer3_outputs(1409) <= a and not b;
    layer3_outputs(1410) <= not b;
    layer3_outputs(1411) <= a or b;
    layer3_outputs(1412) <= not (a or b);
    layer3_outputs(1413) <= a or b;
    layer3_outputs(1414) <= not a;
    layer3_outputs(1415) <= b;
    layer3_outputs(1416) <= not b or a;
    layer3_outputs(1417) <= a;
    layer3_outputs(1418) <= a and not b;
    layer3_outputs(1419) <= a and b;
    layer3_outputs(1420) <= a and not b;
    layer3_outputs(1421) <= b and not a;
    layer3_outputs(1422) <= b;
    layer3_outputs(1423) <= a and b;
    layer3_outputs(1424) <= a and not b;
    layer3_outputs(1425) <= 1'b1;
    layer3_outputs(1426) <= 1'b1;
    layer3_outputs(1427) <= not (a or b);
    layer3_outputs(1428) <= a and not b;
    layer3_outputs(1429) <= not b;
    layer3_outputs(1430) <= b and not a;
    layer3_outputs(1431) <= not a or b;
    layer3_outputs(1432) <= b;
    layer3_outputs(1433) <= not b or a;
    layer3_outputs(1434) <= a and not b;
    layer3_outputs(1435) <= b and not a;
    layer3_outputs(1436) <= a;
    layer3_outputs(1437) <= not a or b;
    layer3_outputs(1438) <= not a or b;
    layer3_outputs(1439) <= not (a or b);
    layer3_outputs(1440) <= not b or a;
    layer3_outputs(1441) <= 1'b1;
    layer3_outputs(1442) <= 1'b1;
    layer3_outputs(1443) <= not a or b;
    layer3_outputs(1444) <= a and b;
    layer3_outputs(1445) <= b and not a;
    layer3_outputs(1446) <= not (a xor b);
    layer3_outputs(1447) <= a xor b;
    layer3_outputs(1448) <= a and b;
    layer3_outputs(1449) <= 1'b0;
    layer3_outputs(1450) <= not a or b;
    layer3_outputs(1451) <= a and b;
    layer3_outputs(1452) <= not (a and b);
    layer3_outputs(1453) <= a;
    layer3_outputs(1454) <= 1'b0;
    layer3_outputs(1455) <= not a;
    layer3_outputs(1456) <= not a;
    layer3_outputs(1457) <= a and b;
    layer3_outputs(1458) <= b;
    layer3_outputs(1459) <= a;
    layer3_outputs(1460) <= not b;
    layer3_outputs(1461) <= not a;
    layer3_outputs(1462) <= b;
    layer3_outputs(1463) <= b;
    layer3_outputs(1464) <= a;
    layer3_outputs(1465) <= b;
    layer3_outputs(1466) <= a or b;
    layer3_outputs(1467) <= not b or a;
    layer3_outputs(1468) <= 1'b1;
    layer3_outputs(1469) <= not a;
    layer3_outputs(1470) <= b and not a;
    layer3_outputs(1471) <= not a;
    layer3_outputs(1472) <= not (a and b);
    layer3_outputs(1473) <= not b or a;
    layer3_outputs(1474) <= a or b;
    layer3_outputs(1475) <= 1'b0;
    layer3_outputs(1476) <= not b;
    layer3_outputs(1477) <= not (a xor b);
    layer3_outputs(1478) <= b;
    layer3_outputs(1479) <= a;
    layer3_outputs(1480) <= b and not a;
    layer3_outputs(1481) <= 1'b1;
    layer3_outputs(1482) <= a and not b;
    layer3_outputs(1483) <= not b or a;
    layer3_outputs(1484) <= not b or a;
    layer3_outputs(1485) <= b;
    layer3_outputs(1486) <= not b or a;
    layer3_outputs(1487) <= not a;
    layer3_outputs(1488) <= not (a and b);
    layer3_outputs(1489) <= not (a or b);
    layer3_outputs(1490) <= not b;
    layer3_outputs(1491) <= a or b;
    layer3_outputs(1492) <= not (a or b);
    layer3_outputs(1493) <= 1'b1;
    layer3_outputs(1494) <= not b;
    layer3_outputs(1495) <= not (a or b);
    layer3_outputs(1496) <= not a;
    layer3_outputs(1497) <= a and b;
    layer3_outputs(1498) <= b and not a;
    layer3_outputs(1499) <= not a;
    layer3_outputs(1500) <= not (a and b);
    layer3_outputs(1501) <= not a;
    layer3_outputs(1502) <= not (a and b);
    layer3_outputs(1503) <= not a;
    layer3_outputs(1504) <= not (a and b);
    layer3_outputs(1505) <= not b or a;
    layer3_outputs(1506) <= not a;
    layer3_outputs(1507) <= a;
    layer3_outputs(1508) <= a;
    layer3_outputs(1509) <= a;
    layer3_outputs(1510) <= a and not b;
    layer3_outputs(1511) <= not a;
    layer3_outputs(1512) <= b and not a;
    layer3_outputs(1513) <= not a or b;
    layer3_outputs(1514) <= a or b;
    layer3_outputs(1515) <= not a;
    layer3_outputs(1516) <= b;
    layer3_outputs(1517) <= a and b;
    layer3_outputs(1518) <= not a or b;
    layer3_outputs(1519) <= not (a and b);
    layer3_outputs(1520) <= not b;
    layer3_outputs(1521) <= a and b;
    layer3_outputs(1522) <= not b;
    layer3_outputs(1523) <= a and not b;
    layer3_outputs(1524) <= 1'b0;
    layer3_outputs(1525) <= not (a xor b);
    layer3_outputs(1526) <= b;
    layer3_outputs(1527) <= not (a or b);
    layer3_outputs(1528) <= not (a and b);
    layer3_outputs(1529) <= not a;
    layer3_outputs(1530) <= not (a and b);
    layer3_outputs(1531) <= not b or a;
    layer3_outputs(1532) <= not a;
    layer3_outputs(1533) <= not a;
    layer3_outputs(1534) <= a and b;
    layer3_outputs(1535) <= not a or b;
    layer3_outputs(1536) <= not (a or b);
    layer3_outputs(1537) <= a;
    layer3_outputs(1538) <= not b or a;
    layer3_outputs(1539) <= 1'b0;
    layer3_outputs(1540) <= a and b;
    layer3_outputs(1541) <= a and b;
    layer3_outputs(1542) <= a or b;
    layer3_outputs(1543) <= a and not b;
    layer3_outputs(1544) <= b and not a;
    layer3_outputs(1545) <= 1'b1;
    layer3_outputs(1546) <= a or b;
    layer3_outputs(1547) <= 1'b0;
    layer3_outputs(1548) <= not (a or b);
    layer3_outputs(1549) <= b;
    layer3_outputs(1550) <= b;
    layer3_outputs(1551) <= a;
    layer3_outputs(1552) <= not b or a;
    layer3_outputs(1553) <= a and b;
    layer3_outputs(1554) <= not (a or b);
    layer3_outputs(1555) <= not b;
    layer3_outputs(1556) <= 1'b0;
    layer3_outputs(1557) <= b and not a;
    layer3_outputs(1558) <= not a;
    layer3_outputs(1559) <= not b;
    layer3_outputs(1560) <= 1'b0;
    layer3_outputs(1561) <= b;
    layer3_outputs(1562) <= 1'b1;
    layer3_outputs(1563) <= 1'b1;
    layer3_outputs(1564) <= b and not a;
    layer3_outputs(1565) <= not b;
    layer3_outputs(1566) <= not (a or b);
    layer3_outputs(1567) <= not b;
    layer3_outputs(1568) <= 1'b0;
    layer3_outputs(1569) <= not (a xor b);
    layer3_outputs(1570) <= b;
    layer3_outputs(1571) <= not b;
    layer3_outputs(1572) <= not a or b;
    layer3_outputs(1573) <= not a or b;
    layer3_outputs(1574) <= a or b;
    layer3_outputs(1575) <= not (a or b);
    layer3_outputs(1576) <= b and not a;
    layer3_outputs(1577) <= not (a and b);
    layer3_outputs(1578) <= 1'b1;
    layer3_outputs(1579) <= a or b;
    layer3_outputs(1580) <= not (a and b);
    layer3_outputs(1581) <= 1'b1;
    layer3_outputs(1582) <= a;
    layer3_outputs(1583) <= 1'b0;
    layer3_outputs(1584) <= a and not b;
    layer3_outputs(1585) <= 1'b1;
    layer3_outputs(1586) <= 1'b0;
    layer3_outputs(1587) <= a and not b;
    layer3_outputs(1588) <= a and b;
    layer3_outputs(1589) <= not a;
    layer3_outputs(1590) <= not a;
    layer3_outputs(1591) <= 1'b1;
    layer3_outputs(1592) <= not (a or b);
    layer3_outputs(1593) <= a and not b;
    layer3_outputs(1594) <= a and b;
    layer3_outputs(1595) <= 1'b0;
    layer3_outputs(1596) <= not (a or b);
    layer3_outputs(1597) <= not (a and b);
    layer3_outputs(1598) <= not (a or b);
    layer3_outputs(1599) <= b and not a;
    layer3_outputs(1600) <= not b or a;
    layer3_outputs(1601) <= a xor b;
    layer3_outputs(1602) <= a and b;
    layer3_outputs(1603) <= not (a and b);
    layer3_outputs(1604) <= a xor b;
    layer3_outputs(1605) <= 1'b1;
    layer3_outputs(1606) <= not (a or b);
    layer3_outputs(1607) <= 1'b0;
    layer3_outputs(1608) <= b and not a;
    layer3_outputs(1609) <= not (a and b);
    layer3_outputs(1610) <= not b;
    layer3_outputs(1611) <= a;
    layer3_outputs(1612) <= 1'b0;
    layer3_outputs(1613) <= not b;
    layer3_outputs(1614) <= not b or a;
    layer3_outputs(1615) <= a xor b;
    layer3_outputs(1616) <= not (a and b);
    layer3_outputs(1617) <= 1'b0;
    layer3_outputs(1618) <= 1'b1;
    layer3_outputs(1619) <= b and not a;
    layer3_outputs(1620) <= a;
    layer3_outputs(1621) <= not a or b;
    layer3_outputs(1622) <= not a;
    layer3_outputs(1623) <= b and not a;
    layer3_outputs(1624) <= not (a or b);
    layer3_outputs(1625) <= a and b;
    layer3_outputs(1626) <= not a;
    layer3_outputs(1627) <= not b;
    layer3_outputs(1628) <= a and b;
    layer3_outputs(1629) <= not a;
    layer3_outputs(1630) <= 1'b1;
    layer3_outputs(1631) <= a;
    layer3_outputs(1632) <= not (a xor b);
    layer3_outputs(1633) <= a and not b;
    layer3_outputs(1634) <= 1'b1;
    layer3_outputs(1635) <= b and not a;
    layer3_outputs(1636) <= a;
    layer3_outputs(1637) <= a and not b;
    layer3_outputs(1638) <= b;
    layer3_outputs(1639) <= not (a or b);
    layer3_outputs(1640) <= not (a or b);
    layer3_outputs(1641) <= not (a and b);
    layer3_outputs(1642) <= not a or b;
    layer3_outputs(1643) <= 1'b0;
    layer3_outputs(1644) <= a and not b;
    layer3_outputs(1645) <= not (a and b);
    layer3_outputs(1646) <= not (a and b);
    layer3_outputs(1647) <= a and not b;
    layer3_outputs(1648) <= 1'b0;
    layer3_outputs(1649) <= a and not b;
    layer3_outputs(1650) <= not a;
    layer3_outputs(1651) <= not (a or b);
    layer3_outputs(1652) <= 1'b0;
    layer3_outputs(1653) <= not (a or b);
    layer3_outputs(1654) <= a and b;
    layer3_outputs(1655) <= a;
    layer3_outputs(1656) <= not b or a;
    layer3_outputs(1657) <= not b or a;
    layer3_outputs(1658) <= 1'b1;
    layer3_outputs(1659) <= not (a or b);
    layer3_outputs(1660) <= a;
    layer3_outputs(1661) <= not a or b;
    layer3_outputs(1662) <= not b or a;
    layer3_outputs(1663) <= not b;
    layer3_outputs(1664) <= not (a and b);
    layer3_outputs(1665) <= b and not a;
    layer3_outputs(1666) <= not (a or b);
    layer3_outputs(1667) <= not b or a;
    layer3_outputs(1668) <= not a;
    layer3_outputs(1669) <= b and not a;
    layer3_outputs(1670) <= a or b;
    layer3_outputs(1671) <= not a;
    layer3_outputs(1672) <= a xor b;
    layer3_outputs(1673) <= 1'b1;
    layer3_outputs(1674) <= not b or a;
    layer3_outputs(1675) <= 1'b1;
    layer3_outputs(1676) <= not (a or b);
    layer3_outputs(1677) <= a and not b;
    layer3_outputs(1678) <= a and b;
    layer3_outputs(1679) <= b;
    layer3_outputs(1680) <= not b or a;
    layer3_outputs(1681) <= a;
    layer3_outputs(1682) <= b and not a;
    layer3_outputs(1683) <= not b;
    layer3_outputs(1684) <= 1'b1;
    layer3_outputs(1685) <= 1'b1;
    layer3_outputs(1686) <= not a;
    layer3_outputs(1687) <= a xor b;
    layer3_outputs(1688) <= b and not a;
    layer3_outputs(1689) <= a;
    layer3_outputs(1690) <= a and b;
    layer3_outputs(1691) <= not a;
    layer3_outputs(1692) <= a or b;
    layer3_outputs(1693) <= not (a xor b);
    layer3_outputs(1694) <= a;
    layer3_outputs(1695) <= not b or a;
    layer3_outputs(1696) <= a and b;
    layer3_outputs(1697) <= a xor b;
    layer3_outputs(1698) <= 1'b0;
    layer3_outputs(1699) <= 1'b1;
    layer3_outputs(1700) <= not a or b;
    layer3_outputs(1701) <= a;
    layer3_outputs(1702) <= not b;
    layer3_outputs(1703) <= not b;
    layer3_outputs(1704) <= a and b;
    layer3_outputs(1705) <= b;
    layer3_outputs(1706) <= not b;
    layer3_outputs(1707) <= not b or a;
    layer3_outputs(1708) <= not a;
    layer3_outputs(1709) <= not (a or b);
    layer3_outputs(1710) <= not (a or b);
    layer3_outputs(1711) <= not a or b;
    layer3_outputs(1712) <= 1'b1;
    layer3_outputs(1713) <= not (a or b);
    layer3_outputs(1714) <= not a or b;
    layer3_outputs(1715) <= b and not a;
    layer3_outputs(1716) <= b and not a;
    layer3_outputs(1717) <= a or b;
    layer3_outputs(1718) <= b and not a;
    layer3_outputs(1719) <= not (a or b);
    layer3_outputs(1720) <= a;
    layer3_outputs(1721) <= b;
    layer3_outputs(1722) <= 1'b1;
    layer3_outputs(1723) <= not b;
    layer3_outputs(1724) <= 1'b1;
    layer3_outputs(1725) <= not a;
    layer3_outputs(1726) <= a or b;
    layer3_outputs(1727) <= b;
    layer3_outputs(1728) <= not a;
    layer3_outputs(1729) <= not (a or b);
    layer3_outputs(1730) <= not (a and b);
    layer3_outputs(1731) <= 1'b1;
    layer3_outputs(1732) <= a;
    layer3_outputs(1733) <= not (a xor b);
    layer3_outputs(1734) <= not (a xor b);
    layer3_outputs(1735) <= not b;
    layer3_outputs(1736) <= not a;
    layer3_outputs(1737) <= not a;
    layer3_outputs(1738) <= a and b;
    layer3_outputs(1739) <= a xor b;
    layer3_outputs(1740) <= not b;
    layer3_outputs(1741) <= not a or b;
    layer3_outputs(1742) <= not b or a;
    layer3_outputs(1743) <= not a or b;
    layer3_outputs(1744) <= not (a and b);
    layer3_outputs(1745) <= not (a or b);
    layer3_outputs(1746) <= not b or a;
    layer3_outputs(1747) <= not a;
    layer3_outputs(1748) <= not b;
    layer3_outputs(1749) <= a and b;
    layer3_outputs(1750) <= a xor b;
    layer3_outputs(1751) <= not b or a;
    layer3_outputs(1752) <= not b;
    layer3_outputs(1753) <= a;
    layer3_outputs(1754) <= not (a xor b);
    layer3_outputs(1755) <= 1'b0;
    layer3_outputs(1756) <= not b or a;
    layer3_outputs(1757) <= b and not a;
    layer3_outputs(1758) <= not (a and b);
    layer3_outputs(1759) <= a and not b;
    layer3_outputs(1760) <= not (a and b);
    layer3_outputs(1761) <= b;
    layer3_outputs(1762) <= not b;
    layer3_outputs(1763) <= a or b;
    layer3_outputs(1764) <= b;
    layer3_outputs(1765) <= not a;
    layer3_outputs(1766) <= not b;
    layer3_outputs(1767) <= 1'b1;
    layer3_outputs(1768) <= a xor b;
    layer3_outputs(1769) <= a;
    layer3_outputs(1770) <= b and not a;
    layer3_outputs(1771) <= not (a and b);
    layer3_outputs(1772) <= b;
    layer3_outputs(1773) <= b;
    layer3_outputs(1774) <= not (a and b);
    layer3_outputs(1775) <= b;
    layer3_outputs(1776) <= not (a and b);
    layer3_outputs(1777) <= a or b;
    layer3_outputs(1778) <= not b or a;
    layer3_outputs(1779) <= not (a and b);
    layer3_outputs(1780) <= 1'b0;
    layer3_outputs(1781) <= a xor b;
    layer3_outputs(1782) <= a;
    layer3_outputs(1783) <= 1'b0;
    layer3_outputs(1784) <= not b or a;
    layer3_outputs(1785) <= not (a or b);
    layer3_outputs(1786) <= not b or a;
    layer3_outputs(1787) <= a and b;
    layer3_outputs(1788) <= a or b;
    layer3_outputs(1789) <= a;
    layer3_outputs(1790) <= a;
    layer3_outputs(1791) <= b;
    layer3_outputs(1792) <= a or b;
    layer3_outputs(1793) <= 1'b0;
    layer3_outputs(1794) <= a xor b;
    layer3_outputs(1795) <= a;
    layer3_outputs(1796) <= b;
    layer3_outputs(1797) <= 1'b1;
    layer3_outputs(1798) <= not a or b;
    layer3_outputs(1799) <= a;
    layer3_outputs(1800) <= not b;
    layer3_outputs(1801) <= not (a or b);
    layer3_outputs(1802) <= a xor b;
    layer3_outputs(1803) <= a and b;
    layer3_outputs(1804) <= b and not a;
    layer3_outputs(1805) <= not a or b;
    layer3_outputs(1806) <= b;
    layer3_outputs(1807) <= not b or a;
    layer3_outputs(1808) <= 1'b1;
    layer3_outputs(1809) <= b and not a;
    layer3_outputs(1810) <= not a or b;
    layer3_outputs(1811) <= b and not a;
    layer3_outputs(1812) <= 1'b0;
    layer3_outputs(1813) <= not (a xor b);
    layer3_outputs(1814) <= not (a and b);
    layer3_outputs(1815) <= a or b;
    layer3_outputs(1816) <= 1'b0;
    layer3_outputs(1817) <= 1'b0;
    layer3_outputs(1818) <= not b;
    layer3_outputs(1819) <= a and b;
    layer3_outputs(1820) <= b;
    layer3_outputs(1821) <= a;
    layer3_outputs(1822) <= a and not b;
    layer3_outputs(1823) <= a or b;
    layer3_outputs(1824) <= a and not b;
    layer3_outputs(1825) <= b and not a;
    layer3_outputs(1826) <= a and not b;
    layer3_outputs(1827) <= b;
    layer3_outputs(1828) <= a and not b;
    layer3_outputs(1829) <= not (a and b);
    layer3_outputs(1830) <= a or b;
    layer3_outputs(1831) <= a or b;
    layer3_outputs(1832) <= a and not b;
    layer3_outputs(1833) <= b;
    layer3_outputs(1834) <= a xor b;
    layer3_outputs(1835) <= a and b;
    layer3_outputs(1836) <= b;
    layer3_outputs(1837) <= a and b;
    layer3_outputs(1838) <= not a or b;
    layer3_outputs(1839) <= a;
    layer3_outputs(1840) <= a or b;
    layer3_outputs(1841) <= a;
    layer3_outputs(1842) <= a xor b;
    layer3_outputs(1843) <= b and not a;
    layer3_outputs(1844) <= b and not a;
    layer3_outputs(1845) <= b;
    layer3_outputs(1846) <= b;
    layer3_outputs(1847) <= not b;
    layer3_outputs(1848) <= 1'b1;
    layer3_outputs(1849) <= a;
    layer3_outputs(1850) <= not (a and b);
    layer3_outputs(1851) <= not a or b;
    layer3_outputs(1852) <= not (a or b);
    layer3_outputs(1853) <= b and not a;
    layer3_outputs(1854) <= not (a and b);
    layer3_outputs(1855) <= not (a and b);
    layer3_outputs(1856) <= 1'b1;
    layer3_outputs(1857) <= not (a and b);
    layer3_outputs(1858) <= not b or a;
    layer3_outputs(1859) <= not b;
    layer3_outputs(1860) <= a and not b;
    layer3_outputs(1861) <= not b;
    layer3_outputs(1862) <= 1'b0;
    layer3_outputs(1863) <= not (a and b);
    layer3_outputs(1864) <= not (a and b);
    layer3_outputs(1865) <= b;
    layer3_outputs(1866) <= not a;
    layer3_outputs(1867) <= not b or a;
    layer3_outputs(1868) <= not (a or b);
    layer3_outputs(1869) <= not (a or b);
    layer3_outputs(1870) <= not (a or b);
    layer3_outputs(1871) <= not a;
    layer3_outputs(1872) <= not b;
    layer3_outputs(1873) <= b and not a;
    layer3_outputs(1874) <= not b;
    layer3_outputs(1875) <= 1'b1;
    layer3_outputs(1876) <= not b;
    layer3_outputs(1877) <= not b or a;
    layer3_outputs(1878) <= not b or a;
    layer3_outputs(1879) <= not a;
    layer3_outputs(1880) <= not a or b;
    layer3_outputs(1881) <= not (a xor b);
    layer3_outputs(1882) <= not a;
    layer3_outputs(1883) <= a and b;
    layer3_outputs(1884) <= a and not b;
    layer3_outputs(1885) <= not b or a;
    layer3_outputs(1886) <= b and not a;
    layer3_outputs(1887) <= not (a and b);
    layer3_outputs(1888) <= not a or b;
    layer3_outputs(1889) <= not a;
    layer3_outputs(1890) <= a;
    layer3_outputs(1891) <= 1'b1;
    layer3_outputs(1892) <= a;
    layer3_outputs(1893) <= 1'b1;
    layer3_outputs(1894) <= 1'b0;
    layer3_outputs(1895) <= a or b;
    layer3_outputs(1896) <= not b;
    layer3_outputs(1897) <= not (a or b);
    layer3_outputs(1898) <= not b or a;
    layer3_outputs(1899) <= a and b;
    layer3_outputs(1900) <= 1'b1;
    layer3_outputs(1901) <= a and b;
    layer3_outputs(1902) <= b;
    layer3_outputs(1903) <= not a or b;
    layer3_outputs(1904) <= not a or b;
    layer3_outputs(1905) <= not b;
    layer3_outputs(1906) <= not a;
    layer3_outputs(1907) <= not a;
    layer3_outputs(1908) <= 1'b1;
    layer3_outputs(1909) <= not a;
    layer3_outputs(1910) <= 1'b1;
    layer3_outputs(1911) <= not a;
    layer3_outputs(1912) <= 1'b0;
    layer3_outputs(1913) <= not b;
    layer3_outputs(1914) <= a or b;
    layer3_outputs(1915) <= not a;
    layer3_outputs(1916) <= not a;
    layer3_outputs(1917) <= b and not a;
    layer3_outputs(1918) <= not (a and b);
    layer3_outputs(1919) <= b;
    layer3_outputs(1920) <= not b;
    layer3_outputs(1921) <= not (a or b);
    layer3_outputs(1922) <= 1'b0;
    layer3_outputs(1923) <= not a or b;
    layer3_outputs(1924) <= a or b;
    layer3_outputs(1925) <= a and not b;
    layer3_outputs(1926) <= not b or a;
    layer3_outputs(1927) <= not a;
    layer3_outputs(1928) <= b and not a;
    layer3_outputs(1929) <= 1'b0;
    layer3_outputs(1930) <= not b or a;
    layer3_outputs(1931) <= a and not b;
    layer3_outputs(1932) <= not a or b;
    layer3_outputs(1933) <= not b or a;
    layer3_outputs(1934) <= not (a xor b);
    layer3_outputs(1935) <= 1'b0;
    layer3_outputs(1936) <= 1'b0;
    layer3_outputs(1937) <= 1'b0;
    layer3_outputs(1938) <= not a;
    layer3_outputs(1939) <= b;
    layer3_outputs(1940) <= b and not a;
    layer3_outputs(1941) <= b and not a;
    layer3_outputs(1942) <= b;
    layer3_outputs(1943) <= b;
    layer3_outputs(1944) <= 1'b1;
    layer3_outputs(1945) <= 1'b0;
    layer3_outputs(1946) <= a and not b;
    layer3_outputs(1947) <= not b;
    layer3_outputs(1948) <= not a or b;
    layer3_outputs(1949) <= not b or a;
    layer3_outputs(1950) <= a and b;
    layer3_outputs(1951) <= 1'b1;
    layer3_outputs(1952) <= a;
    layer3_outputs(1953) <= a and not b;
    layer3_outputs(1954) <= not a or b;
    layer3_outputs(1955) <= b and not a;
    layer3_outputs(1956) <= not b or a;
    layer3_outputs(1957) <= a;
    layer3_outputs(1958) <= not (a or b);
    layer3_outputs(1959) <= not (a or b);
    layer3_outputs(1960) <= a;
    layer3_outputs(1961) <= not a or b;
    layer3_outputs(1962) <= 1'b1;
    layer3_outputs(1963) <= 1'b1;
    layer3_outputs(1964) <= 1'b1;
    layer3_outputs(1965) <= not a;
    layer3_outputs(1966) <= 1'b1;
    layer3_outputs(1967) <= not b or a;
    layer3_outputs(1968) <= a and not b;
    layer3_outputs(1969) <= a or b;
    layer3_outputs(1970) <= a xor b;
    layer3_outputs(1971) <= 1'b1;
    layer3_outputs(1972) <= not a;
    layer3_outputs(1973) <= b and not a;
    layer3_outputs(1974) <= a or b;
    layer3_outputs(1975) <= not b;
    layer3_outputs(1976) <= not (a xor b);
    layer3_outputs(1977) <= a and not b;
    layer3_outputs(1978) <= 1'b1;
    layer3_outputs(1979) <= a;
    layer3_outputs(1980) <= not (a and b);
    layer3_outputs(1981) <= a xor b;
    layer3_outputs(1982) <= a;
    layer3_outputs(1983) <= 1'b1;
    layer3_outputs(1984) <= a and not b;
    layer3_outputs(1985) <= a or b;
    layer3_outputs(1986) <= not (a or b);
    layer3_outputs(1987) <= a and not b;
    layer3_outputs(1988) <= a;
    layer3_outputs(1989) <= a;
    layer3_outputs(1990) <= a xor b;
    layer3_outputs(1991) <= not a or b;
    layer3_outputs(1992) <= not b or a;
    layer3_outputs(1993) <= not a or b;
    layer3_outputs(1994) <= 1'b1;
    layer3_outputs(1995) <= b and not a;
    layer3_outputs(1996) <= 1'b0;
    layer3_outputs(1997) <= not (a or b);
    layer3_outputs(1998) <= not a;
    layer3_outputs(1999) <= not a;
    layer3_outputs(2000) <= 1'b1;
    layer3_outputs(2001) <= 1'b1;
    layer3_outputs(2002) <= not (a xor b);
    layer3_outputs(2003) <= 1'b1;
    layer3_outputs(2004) <= not a;
    layer3_outputs(2005) <= a or b;
    layer3_outputs(2006) <= a and not b;
    layer3_outputs(2007) <= a and not b;
    layer3_outputs(2008) <= 1'b0;
    layer3_outputs(2009) <= 1'b1;
    layer3_outputs(2010) <= a and b;
    layer3_outputs(2011) <= not (a or b);
    layer3_outputs(2012) <= not a;
    layer3_outputs(2013) <= not a or b;
    layer3_outputs(2014) <= not a;
    layer3_outputs(2015) <= 1'b1;
    layer3_outputs(2016) <= not a;
    layer3_outputs(2017) <= not (a and b);
    layer3_outputs(2018) <= not (a xor b);
    layer3_outputs(2019) <= b;
    layer3_outputs(2020) <= 1'b1;
    layer3_outputs(2021) <= not (a and b);
    layer3_outputs(2022) <= not (a and b);
    layer3_outputs(2023) <= not b;
    layer3_outputs(2024) <= 1'b1;
    layer3_outputs(2025) <= a or b;
    layer3_outputs(2026) <= 1'b1;
    layer3_outputs(2027) <= not (a xor b);
    layer3_outputs(2028) <= not a;
    layer3_outputs(2029) <= b;
    layer3_outputs(2030) <= a and not b;
    layer3_outputs(2031) <= a or b;
    layer3_outputs(2032) <= a and b;
    layer3_outputs(2033) <= not b or a;
    layer3_outputs(2034) <= not a;
    layer3_outputs(2035) <= 1'b0;
    layer3_outputs(2036) <= 1'b0;
    layer3_outputs(2037) <= a;
    layer3_outputs(2038) <= a or b;
    layer3_outputs(2039) <= a or b;
    layer3_outputs(2040) <= b and not a;
    layer3_outputs(2041) <= a or b;
    layer3_outputs(2042) <= not b;
    layer3_outputs(2043) <= a and not b;
    layer3_outputs(2044) <= 1'b1;
    layer3_outputs(2045) <= b;
    layer3_outputs(2046) <= not (a and b);
    layer3_outputs(2047) <= a;
    layer3_outputs(2048) <= not b or a;
    layer3_outputs(2049) <= not a;
    layer3_outputs(2050) <= not a or b;
    layer3_outputs(2051) <= 1'b0;
    layer3_outputs(2052) <= not a;
    layer3_outputs(2053) <= not b;
    layer3_outputs(2054) <= a or b;
    layer3_outputs(2055) <= not b or a;
    layer3_outputs(2056) <= b and not a;
    layer3_outputs(2057) <= 1'b0;
    layer3_outputs(2058) <= not a;
    layer3_outputs(2059) <= not a;
    layer3_outputs(2060) <= a or b;
    layer3_outputs(2061) <= a and b;
    layer3_outputs(2062) <= b and not a;
    layer3_outputs(2063) <= b;
    layer3_outputs(2064) <= not a;
    layer3_outputs(2065) <= a;
    layer3_outputs(2066) <= not (a or b);
    layer3_outputs(2067) <= a and b;
    layer3_outputs(2068) <= 1'b1;
    layer3_outputs(2069) <= 1'b0;
    layer3_outputs(2070) <= not a or b;
    layer3_outputs(2071) <= not a or b;
    layer3_outputs(2072) <= not b;
    layer3_outputs(2073) <= a or b;
    layer3_outputs(2074) <= not a or b;
    layer3_outputs(2075) <= b and not a;
    layer3_outputs(2076) <= a and b;
    layer3_outputs(2077) <= a and not b;
    layer3_outputs(2078) <= b and not a;
    layer3_outputs(2079) <= a and b;
    layer3_outputs(2080) <= not b or a;
    layer3_outputs(2081) <= not b or a;
    layer3_outputs(2082) <= a;
    layer3_outputs(2083) <= a;
    layer3_outputs(2084) <= b and not a;
    layer3_outputs(2085) <= not b or a;
    layer3_outputs(2086) <= 1'b0;
    layer3_outputs(2087) <= a or b;
    layer3_outputs(2088) <= a;
    layer3_outputs(2089) <= not (a or b);
    layer3_outputs(2090) <= b;
    layer3_outputs(2091) <= not (a and b);
    layer3_outputs(2092) <= a and not b;
    layer3_outputs(2093) <= not a or b;
    layer3_outputs(2094) <= a or b;
    layer3_outputs(2095) <= not b;
    layer3_outputs(2096) <= a;
    layer3_outputs(2097) <= a and b;
    layer3_outputs(2098) <= 1'b1;
    layer3_outputs(2099) <= a and b;
    layer3_outputs(2100) <= b;
    layer3_outputs(2101) <= not (a and b);
    layer3_outputs(2102) <= not b or a;
    layer3_outputs(2103) <= not a or b;
    layer3_outputs(2104) <= a;
    layer3_outputs(2105) <= a;
    layer3_outputs(2106) <= not (a or b);
    layer3_outputs(2107) <= 1'b0;
    layer3_outputs(2108) <= not (a or b);
    layer3_outputs(2109) <= not b;
    layer3_outputs(2110) <= not (a or b);
    layer3_outputs(2111) <= a and not b;
    layer3_outputs(2112) <= 1'b1;
    layer3_outputs(2113) <= b and not a;
    layer3_outputs(2114) <= a and not b;
    layer3_outputs(2115) <= b and not a;
    layer3_outputs(2116) <= not a;
    layer3_outputs(2117) <= not a or b;
    layer3_outputs(2118) <= not (a and b);
    layer3_outputs(2119) <= not (a and b);
    layer3_outputs(2120) <= not a;
    layer3_outputs(2121) <= b and not a;
    layer3_outputs(2122) <= b and not a;
    layer3_outputs(2123) <= 1'b0;
    layer3_outputs(2124) <= a;
    layer3_outputs(2125) <= not b or a;
    layer3_outputs(2126) <= not a;
    layer3_outputs(2127) <= b;
    layer3_outputs(2128) <= not (a and b);
    layer3_outputs(2129) <= b and not a;
    layer3_outputs(2130) <= 1'b0;
    layer3_outputs(2131) <= not a or b;
    layer3_outputs(2132) <= b and not a;
    layer3_outputs(2133) <= a;
    layer3_outputs(2134) <= a or b;
    layer3_outputs(2135) <= a;
    layer3_outputs(2136) <= a;
    layer3_outputs(2137) <= not (a and b);
    layer3_outputs(2138) <= a and not b;
    layer3_outputs(2139) <= 1'b0;
    layer3_outputs(2140) <= 1'b1;
    layer3_outputs(2141) <= 1'b0;
    layer3_outputs(2142) <= not (a and b);
    layer3_outputs(2143) <= b;
    layer3_outputs(2144) <= not a or b;
    layer3_outputs(2145) <= a xor b;
    layer3_outputs(2146) <= b;
    layer3_outputs(2147) <= a and not b;
    layer3_outputs(2148) <= a;
    layer3_outputs(2149) <= a;
    layer3_outputs(2150) <= not a;
    layer3_outputs(2151) <= not (a and b);
    layer3_outputs(2152) <= not a or b;
    layer3_outputs(2153) <= a and not b;
    layer3_outputs(2154) <= not a;
    layer3_outputs(2155) <= not (a or b);
    layer3_outputs(2156) <= not b or a;
    layer3_outputs(2157) <= a and not b;
    layer3_outputs(2158) <= b;
    layer3_outputs(2159) <= 1'b0;
    layer3_outputs(2160) <= 1'b0;
    layer3_outputs(2161) <= not b or a;
    layer3_outputs(2162) <= not a;
    layer3_outputs(2163) <= not (a and b);
    layer3_outputs(2164) <= a or b;
    layer3_outputs(2165) <= not b or a;
    layer3_outputs(2166) <= a or b;
    layer3_outputs(2167) <= b and not a;
    layer3_outputs(2168) <= a;
    layer3_outputs(2169) <= a and b;
    layer3_outputs(2170) <= not (a or b);
    layer3_outputs(2171) <= b;
    layer3_outputs(2172) <= not a or b;
    layer3_outputs(2173) <= b and not a;
    layer3_outputs(2174) <= not (a xor b);
    layer3_outputs(2175) <= not b;
    layer3_outputs(2176) <= b;
    layer3_outputs(2177) <= a and not b;
    layer3_outputs(2178) <= a and b;
    layer3_outputs(2179) <= not b or a;
    layer3_outputs(2180) <= not a;
    layer3_outputs(2181) <= 1'b0;
    layer3_outputs(2182) <= a xor b;
    layer3_outputs(2183) <= 1'b1;
    layer3_outputs(2184) <= not a;
    layer3_outputs(2185) <= b and not a;
    layer3_outputs(2186) <= a or b;
    layer3_outputs(2187) <= not a;
    layer3_outputs(2188) <= a;
    layer3_outputs(2189) <= not b;
    layer3_outputs(2190) <= a and not b;
    layer3_outputs(2191) <= b and not a;
    layer3_outputs(2192) <= not (a and b);
    layer3_outputs(2193) <= a and b;
    layer3_outputs(2194) <= not (a xor b);
    layer3_outputs(2195) <= 1'b0;
    layer3_outputs(2196) <= 1'b1;
    layer3_outputs(2197) <= not a;
    layer3_outputs(2198) <= a and not b;
    layer3_outputs(2199) <= not (a and b);
    layer3_outputs(2200) <= 1'b0;
    layer3_outputs(2201) <= a;
    layer3_outputs(2202) <= a or b;
    layer3_outputs(2203) <= a;
    layer3_outputs(2204) <= not b;
    layer3_outputs(2205) <= not b or a;
    layer3_outputs(2206) <= not b or a;
    layer3_outputs(2207) <= not b;
    layer3_outputs(2208) <= not (a xor b);
    layer3_outputs(2209) <= not (a and b);
    layer3_outputs(2210) <= not a or b;
    layer3_outputs(2211) <= not b or a;
    layer3_outputs(2212) <= 1'b1;
    layer3_outputs(2213) <= not a or b;
    layer3_outputs(2214) <= a and not b;
    layer3_outputs(2215) <= a;
    layer3_outputs(2216) <= not (a xor b);
    layer3_outputs(2217) <= a;
    layer3_outputs(2218) <= not b;
    layer3_outputs(2219) <= not (a and b);
    layer3_outputs(2220) <= a and not b;
    layer3_outputs(2221) <= b;
    layer3_outputs(2222) <= a;
    layer3_outputs(2223) <= not a;
    layer3_outputs(2224) <= 1'b1;
    layer3_outputs(2225) <= not a or b;
    layer3_outputs(2226) <= a;
    layer3_outputs(2227) <= a or b;
    layer3_outputs(2228) <= 1'b0;
    layer3_outputs(2229) <= b and not a;
    layer3_outputs(2230) <= not a;
    layer3_outputs(2231) <= 1'b0;
    layer3_outputs(2232) <= not b;
    layer3_outputs(2233) <= not b or a;
    layer3_outputs(2234) <= a or b;
    layer3_outputs(2235) <= not a;
    layer3_outputs(2236) <= not (a or b);
    layer3_outputs(2237) <= not b or a;
    layer3_outputs(2238) <= 1'b1;
    layer3_outputs(2239) <= not (a or b);
    layer3_outputs(2240) <= b;
    layer3_outputs(2241) <= not b or a;
    layer3_outputs(2242) <= not (a and b);
    layer3_outputs(2243) <= not b or a;
    layer3_outputs(2244) <= not a;
    layer3_outputs(2245) <= not (a or b);
    layer3_outputs(2246) <= not b or a;
    layer3_outputs(2247) <= not a;
    layer3_outputs(2248) <= not b;
    layer3_outputs(2249) <= not a;
    layer3_outputs(2250) <= not b or a;
    layer3_outputs(2251) <= a or b;
    layer3_outputs(2252) <= 1'b1;
    layer3_outputs(2253) <= 1'b0;
    layer3_outputs(2254) <= 1'b0;
    layer3_outputs(2255) <= not b;
    layer3_outputs(2256) <= not b;
    layer3_outputs(2257) <= 1'b0;
    layer3_outputs(2258) <= b and not a;
    layer3_outputs(2259) <= not b;
    layer3_outputs(2260) <= a and not b;
    layer3_outputs(2261) <= not (a or b);
    layer3_outputs(2262) <= a and not b;
    layer3_outputs(2263) <= not b or a;
    layer3_outputs(2264) <= a and b;
    layer3_outputs(2265) <= not (a and b);
    layer3_outputs(2266) <= a and not b;
    layer3_outputs(2267) <= a and not b;
    layer3_outputs(2268) <= a or b;
    layer3_outputs(2269) <= 1'b0;
    layer3_outputs(2270) <= a or b;
    layer3_outputs(2271) <= not b;
    layer3_outputs(2272) <= b and not a;
    layer3_outputs(2273) <= not a or b;
    layer3_outputs(2274) <= a and b;
    layer3_outputs(2275) <= not (a xor b);
    layer3_outputs(2276) <= not (a and b);
    layer3_outputs(2277) <= 1'b0;
    layer3_outputs(2278) <= b and not a;
    layer3_outputs(2279) <= b and not a;
    layer3_outputs(2280) <= a or b;
    layer3_outputs(2281) <= b and not a;
    layer3_outputs(2282) <= a and not b;
    layer3_outputs(2283) <= not a;
    layer3_outputs(2284) <= b;
    layer3_outputs(2285) <= not (a xor b);
    layer3_outputs(2286) <= b;
    layer3_outputs(2287) <= b and not a;
    layer3_outputs(2288) <= not a or b;
    layer3_outputs(2289) <= 1'b0;
    layer3_outputs(2290) <= not (a or b);
    layer3_outputs(2291) <= 1'b1;
    layer3_outputs(2292) <= b;
    layer3_outputs(2293) <= not b or a;
    layer3_outputs(2294) <= a;
    layer3_outputs(2295) <= 1'b1;
    layer3_outputs(2296) <= a xor b;
    layer3_outputs(2297) <= not a or b;
    layer3_outputs(2298) <= a and b;
    layer3_outputs(2299) <= not b or a;
    layer3_outputs(2300) <= not a;
    layer3_outputs(2301) <= b and not a;
    layer3_outputs(2302) <= 1'b1;
    layer3_outputs(2303) <= not (a or b);
    layer3_outputs(2304) <= a and b;
    layer3_outputs(2305) <= not b or a;
    layer3_outputs(2306) <= 1'b1;
    layer3_outputs(2307) <= b and not a;
    layer3_outputs(2308) <= not b;
    layer3_outputs(2309) <= 1'b0;
    layer3_outputs(2310) <= b;
    layer3_outputs(2311) <= 1'b0;
    layer3_outputs(2312) <= a;
    layer3_outputs(2313) <= not a;
    layer3_outputs(2314) <= a xor b;
    layer3_outputs(2315) <= b and not a;
    layer3_outputs(2316) <= not a;
    layer3_outputs(2317) <= not (a and b);
    layer3_outputs(2318) <= a or b;
    layer3_outputs(2319) <= not b;
    layer3_outputs(2320) <= a and not b;
    layer3_outputs(2321) <= not (a or b);
    layer3_outputs(2322) <= not a;
    layer3_outputs(2323) <= b and not a;
    layer3_outputs(2324) <= b and not a;
    layer3_outputs(2325) <= 1'b0;
    layer3_outputs(2326) <= not a;
    layer3_outputs(2327) <= not b or a;
    layer3_outputs(2328) <= not (a xor b);
    layer3_outputs(2329) <= not a;
    layer3_outputs(2330) <= 1'b1;
    layer3_outputs(2331) <= 1'b0;
    layer3_outputs(2332) <= not (a and b);
    layer3_outputs(2333) <= not a or b;
    layer3_outputs(2334) <= not (a and b);
    layer3_outputs(2335) <= b;
    layer3_outputs(2336) <= a or b;
    layer3_outputs(2337) <= 1'b1;
    layer3_outputs(2338) <= 1'b0;
    layer3_outputs(2339) <= not b;
    layer3_outputs(2340) <= a;
    layer3_outputs(2341) <= not (a or b);
    layer3_outputs(2342) <= not (a or b);
    layer3_outputs(2343) <= a;
    layer3_outputs(2344) <= not b;
    layer3_outputs(2345) <= a or b;
    layer3_outputs(2346) <= a or b;
    layer3_outputs(2347) <= 1'b1;
    layer3_outputs(2348) <= a or b;
    layer3_outputs(2349) <= a;
    layer3_outputs(2350) <= not (a and b);
    layer3_outputs(2351) <= 1'b1;
    layer3_outputs(2352) <= 1'b0;
    layer3_outputs(2353) <= a xor b;
    layer3_outputs(2354) <= a and b;
    layer3_outputs(2355) <= not b;
    layer3_outputs(2356) <= b and not a;
    layer3_outputs(2357) <= 1'b0;
    layer3_outputs(2358) <= not a;
    layer3_outputs(2359) <= not a;
    layer3_outputs(2360) <= a;
    layer3_outputs(2361) <= not a;
    layer3_outputs(2362) <= not (a or b);
    layer3_outputs(2363) <= a;
    layer3_outputs(2364) <= 1'b0;
    layer3_outputs(2365) <= not b or a;
    layer3_outputs(2366) <= b and not a;
    layer3_outputs(2367) <= 1'b0;
    layer3_outputs(2368) <= not (a or b);
    layer3_outputs(2369) <= not b;
    layer3_outputs(2370) <= not a or b;
    layer3_outputs(2371) <= not a;
    layer3_outputs(2372) <= not a or b;
    layer3_outputs(2373) <= not a;
    layer3_outputs(2374) <= b and not a;
    layer3_outputs(2375) <= not b;
    layer3_outputs(2376) <= not a or b;
    layer3_outputs(2377) <= not b or a;
    layer3_outputs(2378) <= not a or b;
    layer3_outputs(2379) <= not (a and b);
    layer3_outputs(2380) <= a;
    layer3_outputs(2381) <= 1'b0;
    layer3_outputs(2382) <= not b or a;
    layer3_outputs(2383) <= not a;
    layer3_outputs(2384) <= not (a xor b);
    layer3_outputs(2385) <= b and not a;
    layer3_outputs(2386) <= not a or b;
    layer3_outputs(2387) <= not (a or b);
    layer3_outputs(2388) <= b and not a;
    layer3_outputs(2389) <= not b or a;
    layer3_outputs(2390) <= not b;
    layer3_outputs(2391) <= a and b;
    layer3_outputs(2392) <= a;
    layer3_outputs(2393) <= a xor b;
    layer3_outputs(2394) <= not (a or b);
    layer3_outputs(2395) <= a or b;
    layer3_outputs(2396) <= not a;
    layer3_outputs(2397) <= 1'b0;
    layer3_outputs(2398) <= not (a and b);
    layer3_outputs(2399) <= a and not b;
    layer3_outputs(2400) <= not (a and b);
    layer3_outputs(2401) <= not (a or b);
    layer3_outputs(2402) <= 1'b1;
    layer3_outputs(2403) <= not b;
    layer3_outputs(2404) <= not b or a;
    layer3_outputs(2405) <= not b;
    layer3_outputs(2406) <= a or b;
    layer3_outputs(2407) <= not (a and b);
    layer3_outputs(2408) <= not (a and b);
    layer3_outputs(2409) <= a;
    layer3_outputs(2410) <= a and b;
    layer3_outputs(2411) <= not a or b;
    layer3_outputs(2412) <= not (a or b);
    layer3_outputs(2413) <= not b;
    layer3_outputs(2414) <= not b or a;
    layer3_outputs(2415) <= a or b;
    layer3_outputs(2416) <= not b or a;
    layer3_outputs(2417) <= not (a xor b);
    layer3_outputs(2418) <= not a;
    layer3_outputs(2419) <= a and b;
    layer3_outputs(2420) <= a and not b;
    layer3_outputs(2421) <= not b or a;
    layer3_outputs(2422) <= a;
    layer3_outputs(2423) <= a and not b;
    layer3_outputs(2424) <= not (a and b);
    layer3_outputs(2425) <= not a;
    layer3_outputs(2426) <= a or b;
    layer3_outputs(2427) <= not (a and b);
    layer3_outputs(2428) <= a xor b;
    layer3_outputs(2429) <= not (a or b);
    layer3_outputs(2430) <= b;
    layer3_outputs(2431) <= not (a and b);
    layer3_outputs(2432) <= not b or a;
    layer3_outputs(2433) <= a and not b;
    layer3_outputs(2434) <= 1'b0;
    layer3_outputs(2435) <= not a or b;
    layer3_outputs(2436) <= a;
    layer3_outputs(2437) <= not (a or b);
    layer3_outputs(2438) <= not b;
    layer3_outputs(2439) <= not a;
    layer3_outputs(2440) <= a;
    layer3_outputs(2441) <= not a or b;
    layer3_outputs(2442) <= a and not b;
    layer3_outputs(2443) <= a and b;
    layer3_outputs(2444) <= not (a and b);
    layer3_outputs(2445) <= not a or b;
    layer3_outputs(2446) <= not b;
    layer3_outputs(2447) <= a and not b;
    layer3_outputs(2448) <= 1'b1;
    layer3_outputs(2449) <= a or b;
    layer3_outputs(2450) <= not b or a;
    layer3_outputs(2451) <= 1'b0;
    layer3_outputs(2452) <= not b;
    layer3_outputs(2453) <= not (a and b);
    layer3_outputs(2454) <= 1'b1;
    layer3_outputs(2455) <= b and not a;
    layer3_outputs(2456) <= b and not a;
    layer3_outputs(2457) <= b;
    layer3_outputs(2458) <= a and not b;
    layer3_outputs(2459) <= not (a or b);
    layer3_outputs(2460) <= not a;
    layer3_outputs(2461) <= b;
    layer3_outputs(2462) <= not b;
    layer3_outputs(2463) <= not (a or b);
    layer3_outputs(2464) <= not b;
    layer3_outputs(2465) <= not (a or b);
    layer3_outputs(2466) <= a or b;
    layer3_outputs(2467) <= not a or b;
    layer3_outputs(2468) <= not a;
    layer3_outputs(2469) <= not (a or b);
    layer3_outputs(2470) <= b and not a;
    layer3_outputs(2471) <= b;
    layer3_outputs(2472) <= b and not a;
    layer3_outputs(2473) <= a xor b;
    layer3_outputs(2474) <= b and not a;
    layer3_outputs(2475) <= 1'b1;
    layer3_outputs(2476) <= not a or b;
    layer3_outputs(2477) <= not b;
    layer3_outputs(2478) <= 1'b1;
    layer3_outputs(2479) <= not (a xor b);
    layer3_outputs(2480) <= not b or a;
    layer3_outputs(2481) <= a;
    layer3_outputs(2482) <= a;
    layer3_outputs(2483) <= not b;
    layer3_outputs(2484) <= b and not a;
    layer3_outputs(2485) <= not (a and b);
    layer3_outputs(2486) <= b;
    layer3_outputs(2487) <= not a or b;
    layer3_outputs(2488) <= b;
    layer3_outputs(2489) <= a and not b;
    layer3_outputs(2490) <= b;
    layer3_outputs(2491) <= not (a and b);
    layer3_outputs(2492) <= not a or b;
    layer3_outputs(2493) <= not (a or b);
    layer3_outputs(2494) <= not a;
    layer3_outputs(2495) <= b;
    layer3_outputs(2496) <= b and not a;
    layer3_outputs(2497) <= b;
    layer3_outputs(2498) <= a and not b;
    layer3_outputs(2499) <= a and not b;
    layer3_outputs(2500) <= not b or a;
    layer3_outputs(2501) <= not a or b;
    layer3_outputs(2502) <= not a;
    layer3_outputs(2503) <= b;
    layer3_outputs(2504) <= b;
    layer3_outputs(2505) <= a or b;
    layer3_outputs(2506) <= a;
    layer3_outputs(2507) <= not (a and b);
    layer3_outputs(2508) <= a and not b;
    layer3_outputs(2509) <= a and b;
    layer3_outputs(2510) <= 1'b0;
    layer3_outputs(2511) <= a and b;
    layer3_outputs(2512) <= not (a or b);
    layer3_outputs(2513) <= 1'b0;
    layer3_outputs(2514) <= b;
    layer3_outputs(2515) <= a and not b;
    layer3_outputs(2516) <= a or b;
    layer3_outputs(2517) <= a and not b;
    layer3_outputs(2518) <= a and not b;
    layer3_outputs(2519) <= b and not a;
    layer3_outputs(2520) <= b;
    layer3_outputs(2521) <= a and b;
    layer3_outputs(2522) <= not a;
    layer3_outputs(2523) <= not a or b;
    layer3_outputs(2524) <= not b;
    layer3_outputs(2525) <= b and not a;
    layer3_outputs(2526) <= a and not b;
    layer3_outputs(2527) <= not (a and b);
    layer3_outputs(2528) <= a or b;
    layer3_outputs(2529) <= a and not b;
    layer3_outputs(2530) <= not b;
    layer3_outputs(2531) <= b;
    layer3_outputs(2532) <= 1'b0;
    layer3_outputs(2533) <= a or b;
    layer3_outputs(2534) <= 1'b1;
    layer3_outputs(2535) <= not b;
    layer3_outputs(2536) <= 1'b1;
    layer3_outputs(2537) <= not a or b;
    layer3_outputs(2538) <= not (a or b);
    layer3_outputs(2539) <= not (a and b);
    layer3_outputs(2540) <= 1'b1;
    layer3_outputs(2541) <= not a or b;
    layer3_outputs(2542) <= not b;
    layer3_outputs(2543) <= a and b;
    layer3_outputs(2544) <= not b or a;
    layer3_outputs(2545) <= a or b;
    layer3_outputs(2546) <= a and b;
    layer3_outputs(2547) <= 1'b0;
    layer3_outputs(2548) <= 1'b0;
    layer3_outputs(2549) <= not (a and b);
    layer3_outputs(2550) <= 1'b1;
    layer3_outputs(2551) <= not (a and b);
    layer3_outputs(2552) <= a and not b;
    layer3_outputs(2553) <= 1'b0;
    layer3_outputs(2554) <= not (a and b);
    layer3_outputs(2555) <= b and not a;
    layer3_outputs(2556) <= b and not a;
    layer3_outputs(2557) <= not (a and b);
    layer3_outputs(2558) <= not b;
    layer3_outputs(2559) <= not a or b;
    layer3_outputs(2560) <= a;
    layer3_outputs(2561) <= not b or a;
    layer3_outputs(2562) <= b and not a;
    layer3_outputs(2563) <= b and not a;
    layer3_outputs(2564) <= 1'b0;
    layer3_outputs(2565) <= not b;
    layer3_outputs(2566) <= not a;
    layer3_outputs(2567) <= not b;
    layer3_outputs(2568) <= a;
    layer3_outputs(2569) <= not b;
    layer3_outputs(2570) <= 1'b1;
    layer3_outputs(2571) <= a and not b;
    layer3_outputs(2572) <= not (a or b);
    layer3_outputs(2573) <= not (a xor b);
    layer3_outputs(2574) <= b;
    layer3_outputs(2575) <= a xor b;
    layer3_outputs(2576) <= a;
    layer3_outputs(2577) <= not (a xor b);
    layer3_outputs(2578) <= not (a and b);
    layer3_outputs(2579) <= 1'b1;
    layer3_outputs(2580) <= b and not a;
    layer3_outputs(2581) <= not (a or b);
    layer3_outputs(2582) <= a and b;
    layer3_outputs(2583) <= not a;
    layer3_outputs(2584) <= a and not b;
    layer3_outputs(2585) <= b and not a;
    layer3_outputs(2586) <= a and b;
    layer3_outputs(2587) <= a and b;
    layer3_outputs(2588) <= not b or a;
    layer3_outputs(2589) <= 1'b1;
    layer3_outputs(2590) <= a;
    layer3_outputs(2591) <= not a or b;
    layer3_outputs(2592) <= 1'b1;
    layer3_outputs(2593) <= b;
    layer3_outputs(2594) <= not a;
    layer3_outputs(2595) <= not (a or b);
    layer3_outputs(2596) <= b;
    layer3_outputs(2597) <= not a;
    layer3_outputs(2598) <= not b;
    layer3_outputs(2599) <= not b;
    layer3_outputs(2600) <= not a;
    layer3_outputs(2601) <= 1'b0;
    layer3_outputs(2602) <= not a or b;
    layer3_outputs(2603) <= not b;
    layer3_outputs(2604) <= not (a and b);
    layer3_outputs(2605) <= b and not a;
    layer3_outputs(2606) <= not b;
    layer3_outputs(2607) <= not b;
    layer3_outputs(2608) <= a and not b;
    layer3_outputs(2609) <= 1'b0;
    layer3_outputs(2610) <= not (a or b);
    layer3_outputs(2611) <= b and not a;
    layer3_outputs(2612) <= a and not b;
    layer3_outputs(2613) <= b and not a;
    layer3_outputs(2614) <= not a;
    layer3_outputs(2615) <= a and not b;
    layer3_outputs(2616) <= b and not a;
    layer3_outputs(2617) <= 1'b1;
    layer3_outputs(2618) <= b;
    layer3_outputs(2619) <= a and not b;
    layer3_outputs(2620) <= a;
    layer3_outputs(2621) <= a and b;
    layer3_outputs(2622) <= b and not a;
    layer3_outputs(2623) <= 1'b1;
    layer3_outputs(2624) <= not (a xor b);
    layer3_outputs(2625) <= not b;
    layer3_outputs(2626) <= a and b;
    layer3_outputs(2627) <= b;
    layer3_outputs(2628) <= a and not b;
    layer3_outputs(2629) <= not a;
    layer3_outputs(2630) <= a or b;
    layer3_outputs(2631) <= 1'b1;
    layer3_outputs(2632) <= a;
    layer3_outputs(2633) <= b and not a;
    layer3_outputs(2634) <= a and not b;
    layer3_outputs(2635) <= a or b;
    layer3_outputs(2636) <= not (a or b);
    layer3_outputs(2637) <= not (a xor b);
    layer3_outputs(2638) <= not a or b;
    layer3_outputs(2639) <= a and b;
    layer3_outputs(2640) <= 1'b0;
    layer3_outputs(2641) <= not a or b;
    layer3_outputs(2642) <= a or b;
    layer3_outputs(2643) <= a and b;
    layer3_outputs(2644) <= b;
    layer3_outputs(2645) <= not a;
    layer3_outputs(2646) <= 1'b1;
    layer3_outputs(2647) <= 1'b0;
    layer3_outputs(2648) <= not b;
    layer3_outputs(2649) <= b;
    layer3_outputs(2650) <= not (a and b);
    layer3_outputs(2651) <= a and b;
    layer3_outputs(2652) <= a or b;
    layer3_outputs(2653) <= 1'b0;
    layer3_outputs(2654) <= a xor b;
    layer3_outputs(2655) <= not b;
    layer3_outputs(2656) <= a xor b;
    layer3_outputs(2657) <= b;
    layer3_outputs(2658) <= b;
    layer3_outputs(2659) <= 1'b1;
    layer3_outputs(2660) <= a and b;
    layer3_outputs(2661) <= a and b;
    layer3_outputs(2662) <= not a or b;
    layer3_outputs(2663) <= a and not b;
    layer3_outputs(2664) <= 1'b1;
    layer3_outputs(2665) <= a;
    layer3_outputs(2666) <= not b;
    layer3_outputs(2667) <= 1'b1;
    layer3_outputs(2668) <= a;
    layer3_outputs(2669) <= a and not b;
    layer3_outputs(2670) <= 1'b1;
    layer3_outputs(2671) <= not (a or b);
    layer3_outputs(2672) <= a or b;
    layer3_outputs(2673) <= not a;
    layer3_outputs(2674) <= a or b;
    layer3_outputs(2675) <= not a or b;
    layer3_outputs(2676) <= a or b;
    layer3_outputs(2677) <= a and b;
    layer3_outputs(2678) <= a and b;
    layer3_outputs(2679) <= b;
    layer3_outputs(2680) <= a and not b;
    layer3_outputs(2681) <= b and not a;
    layer3_outputs(2682) <= 1'b1;
    layer3_outputs(2683) <= b and not a;
    layer3_outputs(2684) <= not (a or b);
    layer3_outputs(2685) <= b and not a;
    layer3_outputs(2686) <= a or b;
    layer3_outputs(2687) <= not a or b;
    layer3_outputs(2688) <= not a or b;
    layer3_outputs(2689) <= not (a or b);
    layer3_outputs(2690) <= not a;
    layer3_outputs(2691) <= b and not a;
    layer3_outputs(2692) <= 1'b1;
    layer3_outputs(2693) <= not (a or b);
    layer3_outputs(2694) <= a and not b;
    layer3_outputs(2695) <= not a or b;
    layer3_outputs(2696) <= a xor b;
    layer3_outputs(2697) <= not b;
    layer3_outputs(2698) <= not (a and b);
    layer3_outputs(2699) <= a and not b;
    layer3_outputs(2700) <= 1'b0;
    layer3_outputs(2701) <= not b;
    layer3_outputs(2702) <= a;
    layer3_outputs(2703) <= 1'b1;
    layer3_outputs(2704) <= not (a or b);
    layer3_outputs(2705) <= not b or a;
    layer3_outputs(2706) <= a or b;
    layer3_outputs(2707) <= 1'b1;
    layer3_outputs(2708) <= a or b;
    layer3_outputs(2709) <= a or b;
    layer3_outputs(2710) <= not a or b;
    layer3_outputs(2711) <= not (a and b);
    layer3_outputs(2712) <= a;
    layer3_outputs(2713) <= a and not b;
    layer3_outputs(2714) <= b and not a;
    layer3_outputs(2715) <= a and not b;
    layer3_outputs(2716) <= b;
    layer3_outputs(2717) <= b;
    layer3_outputs(2718) <= not a or b;
    layer3_outputs(2719) <= not a;
    layer3_outputs(2720) <= b;
    layer3_outputs(2721) <= 1'b0;
    layer3_outputs(2722) <= a;
    layer3_outputs(2723) <= not b or a;
    layer3_outputs(2724) <= not (a xor b);
    layer3_outputs(2725) <= 1'b0;
    layer3_outputs(2726) <= b;
    layer3_outputs(2727) <= a and not b;
    layer3_outputs(2728) <= 1'b1;
    layer3_outputs(2729) <= not a or b;
    layer3_outputs(2730) <= a and b;
    layer3_outputs(2731) <= a and not b;
    layer3_outputs(2732) <= a and b;
    layer3_outputs(2733) <= not b;
    layer3_outputs(2734) <= a;
    layer3_outputs(2735) <= not (a xor b);
    layer3_outputs(2736) <= a or b;
    layer3_outputs(2737) <= a and b;
    layer3_outputs(2738) <= b and not a;
    layer3_outputs(2739) <= not (a or b);
    layer3_outputs(2740) <= not b;
    layer3_outputs(2741) <= a xor b;
    layer3_outputs(2742) <= b;
    layer3_outputs(2743) <= b and not a;
    layer3_outputs(2744) <= not (a and b);
    layer3_outputs(2745) <= a;
    layer3_outputs(2746) <= not (a and b);
    layer3_outputs(2747) <= not a;
    layer3_outputs(2748) <= a and b;
    layer3_outputs(2749) <= 1'b1;
    layer3_outputs(2750) <= b and not a;
    layer3_outputs(2751) <= a and not b;
    layer3_outputs(2752) <= b;
    layer3_outputs(2753) <= a and b;
    layer3_outputs(2754) <= b and not a;
    layer3_outputs(2755) <= b and not a;
    layer3_outputs(2756) <= a xor b;
    layer3_outputs(2757) <= b;
    layer3_outputs(2758) <= a and not b;
    layer3_outputs(2759) <= 1'b0;
    layer3_outputs(2760) <= 1'b1;
    layer3_outputs(2761) <= not b;
    layer3_outputs(2762) <= not (a or b);
    layer3_outputs(2763) <= b;
    layer3_outputs(2764) <= not a;
    layer3_outputs(2765) <= 1'b1;
    layer3_outputs(2766) <= a and not b;
    layer3_outputs(2767) <= b and not a;
    layer3_outputs(2768) <= not a or b;
    layer3_outputs(2769) <= not b or a;
    layer3_outputs(2770) <= not a or b;
    layer3_outputs(2771) <= not (a and b);
    layer3_outputs(2772) <= not b or a;
    layer3_outputs(2773) <= a;
    layer3_outputs(2774) <= a xor b;
    layer3_outputs(2775) <= not (a and b);
    layer3_outputs(2776) <= not a;
    layer3_outputs(2777) <= a and b;
    layer3_outputs(2778) <= not (a xor b);
    layer3_outputs(2779) <= not b;
    layer3_outputs(2780) <= a and b;
    layer3_outputs(2781) <= not b or a;
    layer3_outputs(2782) <= b;
    layer3_outputs(2783) <= a;
    layer3_outputs(2784) <= not (a or b);
    layer3_outputs(2785) <= not a;
    layer3_outputs(2786) <= not b;
    layer3_outputs(2787) <= not a;
    layer3_outputs(2788) <= not (a or b);
    layer3_outputs(2789) <= not (a or b);
    layer3_outputs(2790) <= b;
    layer3_outputs(2791) <= a and not b;
    layer3_outputs(2792) <= not b;
    layer3_outputs(2793) <= 1'b1;
    layer3_outputs(2794) <= not (a xor b);
    layer3_outputs(2795) <= not a;
    layer3_outputs(2796) <= not b;
    layer3_outputs(2797) <= not (a and b);
    layer3_outputs(2798) <= not a;
    layer3_outputs(2799) <= 1'b1;
    layer3_outputs(2800) <= 1'b0;
    layer3_outputs(2801) <= not a or b;
    layer3_outputs(2802) <= not (a and b);
    layer3_outputs(2803) <= b;
    layer3_outputs(2804) <= 1'b0;
    layer3_outputs(2805) <= a;
    layer3_outputs(2806) <= not b or a;
    layer3_outputs(2807) <= b;
    layer3_outputs(2808) <= not b or a;
    layer3_outputs(2809) <= not (a xor b);
    layer3_outputs(2810) <= not b or a;
    layer3_outputs(2811) <= a and not b;
    layer3_outputs(2812) <= a;
    layer3_outputs(2813) <= not b or a;
    layer3_outputs(2814) <= 1'b0;
    layer3_outputs(2815) <= not a;
    layer3_outputs(2816) <= a and not b;
    layer3_outputs(2817) <= b and not a;
    layer3_outputs(2818) <= a and b;
    layer3_outputs(2819) <= not b or a;
    layer3_outputs(2820) <= 1'b1;
    layer3_outputs(2821) <= not a or b;
    layer3_outputs(2822) <= not (a or b);
    layer3_outputs(2823) <= a xor b;
    layer3_outputs(2824) <= a or b;
    layer3_outputs(2825) <= not b or a;
    layer3_outputs(2826) <= not (a and b);
    layer3_outputs(2827) <= a and not b;
    layer3_outputs(2828) <= b;
    layer3_outputs(2829) <= a;
    layer3_outputs(2830) <= not b or a;
    layer3_outputs(2831) <= a or b;
    layer3_outputs(2832) <= not (a or b);
    layer3_outputs(2833) <= a and not b;
    layer3_outputs(2834) <= b;
    layer3_outputs(2835) <= not b;
    layer3_outputs(2836) <= not b;
    layer3_outputs(2837) <= a and b;
    layer3_outputs(2838) <= 1'b0;
    layer3_outputs(2839) <= a;
    layer3_outputs(2840) <= not (a and b);
    layer3_outputs(2841) <= 1'b0;
    layer3_outputs(2842) <= not a;
    layer3_outputs(2843) <= b and not a;
    layer3_outputs(2844) <= 1'b1;
    layer3_outputs(2845) <= b and not a;
    layer3_outputs(2846) <= a;
    layer3_outputs(2847) <= not (a and b);
    layer3_outputs(2848) <= not a or b;
    layer3_outputs(2849) <= 1'b0;
    layer3_outputs(2850) <= not a;
    layer3_outputs(2851) <= b;
    layer3_outputs(2852) <= not a;
    layer3_outputs(2853) <= not b;
    layer3_outputs(2854) <= not (a xor b);
    layer3_outputs(2855) <= b and not a;
    layer3_outputs(2856) <= not b or a;
    layer3_outputs(2857) <= 1'b0;
    layer3_outputs(2858) <= b and not a;
    layer3_outputs(2859) <= a;
    layer3_outputs(2860) <= a and not b;
    layer3_outputs(2861) <= not (a and b);
    layer3_outputs(2862) <= not (a and b);
    layer3_outputs(2863) <= a;
    layer3_outputs(2864) <= not (a or b);
    layer3_outputs(2865) <= not (a xor b);
    layer3_outputs(2866) <= not b or a;
    layer3_outputs(2867) <= not a;
    layer3_outputs(2868) <= 1'b1;
    layer3_outputs(2869) <= not b;
    layer3_outputs(2870) <= not a or b;
    layer3_outputs(2871) <= a or b;
    layer3_outputs(2872) <= a and not b;
    layer3_outputs(2873) <= not (a xor b);
    layer3_outputs(2874) <= not a;
    layer3_outputs(2875) <= not b;
    layer3_outputs(2876) <= b and not a;
    layer3_outputs(2877) <= a;
    layer3_outputs(2878) <= not (a and b);
    layer3_outputs(2879) <= not b;
    layer3_outputs(2880) <= b and not a;
    layer3_outputs(2881) <= a and b;
    layer3_outputs(2882) <= a or b;
    layer3_outputs(2883) <= not a;
    layer3_outputs(2884) <= a or b;
    layer3_outputs(2885) <= not (a and b);
    layer3_outputs(2886) <= 1'b0;
    layer3_outputs(2887) <= not b;
    layer3_outputs(2888) <= a;
    layer3_outputs(2889) <= 1'b0;
    layer3_outputs(2890) <= b and not a;
    layer3_outputs(2891) <= 1'b1;
    layer3_outputs(2892) <= a or b;
    layer3_outputs(2893) <= a and b;
    layer3_outputs(2894) <= b;
    layer3_outputs(2895) <= a;
    layer3_outputs(2896) <= not (a and b);
    layer3_outputs(2897) <= a;
    layer3_outputs(2898) <= 1'b1;
    layer3_outputs(2899) <= not a or b;
    layer3_outputs(2900) <= not a;
    layer3_outputs(2901) <= not b or a;
    layer3_outputs(2902) <= 1'b1;
    layer3_outputs(2903) <= not b;
    layer3_outputs(2904) <= not a or b;
    layer3_outputs(2905) <= not b or a;
    layer3_outputs(2906) <= b and not a;
    layer3_outputs(2907) <= not b or a;
    layer3_outputs(2908) <= 1'b1;
    layer3_outputs(2909) <= 1'b0;
    layer3_outputs(2910) <= not (a xor b);
    layer3_outputs(2911) <= not a or b;
    layer3_outputs(2912) <= a;
    layer3_outputs(2913) <= not (a or b);
    layer3_outputs(2914) <= a and not b;
    layer3_outputs(2915) <= a and b;
    layer3_outputs(2916) <= b;
    layer3_outputs(2917) <= a and not b;
    layer3_outputs(2918) <= a and b;
    layer3_outputs(2919) <= a and b;
    layer3_outputs(2920) <= not (a or b);
    layer3_outputs(2921) <= b;
    layer3_outputs(2922) <= not a or b;
    layer3_outputs(2923) <= a or b;
    layer3_outputs(2924) <= 1'b0;
    layer3_outputs(2925) <= b and not a;
    layer3_outputs(2926) <= b and not a;
    layer3_outputs(2927) <= 1'b1;
    layer3_outputs(2928) <= b and not a;
    layer3_outputs(2929) <= not (a or b);
    layer3_outputs(2930) <= not (a and b);
    layer3_outputs(2931) <= not a or b;
    layer3_outputs(2932) <= not b or a;
    layer3_outputs(2933) <= not (a or b);
    layer3_outputs(2934) <= not b;
    layer3_outputs(2935) <= 1'b0;
    layer3_outputs(2936) <= not b or a;
    layer3_outputs(2937) <= a or b;
    layer3_outputs(2938) <= 1'b1;
    layer3_outputs(2939) <= not a;
    layer3_outputs(2940) <= a and b;
    layer3_outputs(2941) <= not (a and b);
    layer3_outputs(2942) <= not b or a;
    layer3_outputs(2943) <= b and not a;
    layer3_outputs(2944) <= 1'b1;
    layer3_outputs(2945) <= a and not b;
    layer3_outputs(2946) <= not a;
    layer3_outputs(2947) <= 1'b0;
    layer3_outputs(2948) <= not (a or b);
    layer3_outputs(2949) <= not (a and b);
    layer3_outputs(2950) <= not (a or b);
    layer3_outputs(2951) <= 1'b1;
    layer3_outputs(2952) <= not a or b;
    layer3_outputs(2953) <= a or b;
    layer3_outputs(2954) <= not b or a;
    layer3_outputs(2955) <= a;
    layer3_outputs(2956) <= not (a and b);
    layer3_outputs(2957) <= not b;
    layer3_outputs(2958) <= a;
    layer3_outputs(2959) <= a or b;
    layer3_outputs(2960) <= not a or b;
    layer3_outputs(2961) <= 1'b0;
    layer3_outputs(2962) <= 1'b1;
    layer3_outputs(2963) <= not a or b;
    layer3_outputs(2964) <= b and not a;
    layer3_outputs(2965) <= 1'b1;
    layer3_outputs(2966) <= b;
    layer3_outputs(2967) <= not a;
    layer3_outputs(2968) <= not (a or b);
    layer3_outputs(2969) <= not (a or b);
    layer3_outputs(2970) <= not a or b;
    layer3_outputs(2971) <= 1'b0;
    layer3_outputs(2972) <= b and not a;
    layer3_outputs(2973) <= not (a and b);
    layer3_outputs(2974) <= not b;
    layer3_outputs(2975) <= a and b;
    layer3_outputs(2976) <= not (a or b);
    layer3_outputs(2977) <= a or b;
    layer3_outputs(2978) <= a and not b;
    layer3_outputs(2979) <= not a;
    layer3_outputs(2980) <= not b;
    layer3_outputs(2981) <= not (a or b);
    layer3_outputs(2982) <= b;
    layer3_outputs(2983) <= not b;
    layer3_outputs(2984) <= a and not b;
    layer3_outputs(2985) <= a and b;
    layer3_outputs(2986) <= not a;
    layer3_outputs(2987) <= not (a and b);
    layer3_outputs(2988) <= a;
    layer3_outputs(2989) <= not b or a;
    layer3_outputs(2990) <= not (a xor b);
    layer3_outputs(2991) <= 1'b0;
    layer3_outputs(2992) <= not (a and b);
    layer3_outputs(2993) <= b;
    layer3_outputs(2994) <= b;
    layer3_outputs(2995) <= a;
    layer3_outputs(2996) <= a;
    layer3_outputs(2997) <= not a;
    layer3_outputs(2998) <= b;
    layer3_outputs(2999) <= not a;
    layer3_outputs(3000) <= a and not b;
    layer3_outputs(3001) <= not (a xor b);
    layer3_outputs(3002) <= not (a and b);
    layer3_outputs(3003) <= a and b;
    layer3_outputs(3004) <= a and b;
    layer3_outputs(3005) <= a xor b;
    layer3_outputs(3006) <= a xor b;
    layer3_outputs(3007) <= a and not b;
    layer3_outputs(3008) <= not b;
    layer3_outputs(3009) <= b;
    layer3_outputs(3010) <= a and not b;
    layer3_outputs(3011) <= a and not b;
    layer3_outputs(3012) <= not a;
    layer3_outputs(3013) <= a or b;
    layer3_outputs(3014) <= not (a xor b);
    layer3_outputs(3015) <= a and b;
    layer3_outputs(3016) <= a or b;
    layer3_outputs(3017) <= not b;
    layer3_outputs(3018) <= a or b;
    layer3_outputs(3019) <= b and not a;
    layer3_outputs(3020) <= not b or a;
    layer3_outputs(3021) <= a or b;
    layer3_outputs(3022) <= a and b;
    layer3_outputs(3023) <= not (a and b);
    layer3_outputs(3024) <= a or b;
    layer3_outputs(3025) <= 1'b0;
    layer3_outputs(3026) <= not b;
    layer3_outputs(3027) <= a;
    layer3_outputs(3028) <= a;
    layer3_outputs(3029) <= not (a or b);
    layer3_outputs(3030) <= not (a or b);
    layer3_outputs(3031) <= not (a or b);
    layer3_outputs(3032) <= not a or b;
    layer3_outputs(3033) <= not a or b;
    layer3_outputs(3034) <= 1'b0;
    layer3_outputs(3035) <= not b or a;
    layer3_outputs(3036) <= not a or b;
    layer3_outputs(3037) <= not a or b;
    layer3_outputs(3038) <= not b or a;
    layer3_outputs(3039) <= not (a or b);
    layer3_outputs(3040) <= a and not b;
    layer3_outputs(3041) <= a and b;
    layer3_outputs(3042) <= a and b;
    layer3_outputs(3043) <= not b or a;
    layer3_outputs(3044) <= b and not a;
    layer3_outputs(3045) <= not (a or b);
    layer3_outputs(3046) <= b and not a;
    layer3_outputs(3047) <= not a;
    layer3_outputs(3048) <= a and not b;
    layer3_outputs(3049) <= 1'b0;
    layer3_outputs(3050) <= not a;
    layer3_outputs(3051) <= b;
    layer3_outputs(3052) <= not b or a;
    layer3_outputs(3053) <= a or b;
    layer3_outputs(3054) <= 1'b0;
    layer3_outputs(3055) <= a;
    layer3_outputs(3056) <= b and not a;
    layer3_outputs(3057) <= not a;
    layer3_outputs(3058) <= a;
    layer3_outputs(3059) <= a;
    layer3_outputs(3060) <= not a or b;
    layer3_outputs(3061) <= not (a and b);
    layer3_outputs(3062) <= a;
    layer3_outputs(3063) <= not (a or b);
    layer3_outputs(3064) <= not (a or b);
    layer3_outputs(3065) <= 1'b1;
    layer3_outputs(3066) <= b and not a;
    layer3_outputs(3067) <= b and not a;
    layer3_outputs(3068) <= 1'b1;
    layer3_outputs(3069) <= 1'b0;
    layer3_outputs(3070) <= not b or a;
    layer3_outputs(3071) <= not a or b;
    layer3_outputs(3072) <= not b;
    layer3_outputs(3073) <= a and b;
    layer3_outputs(3074) <= not (a xor b);
    layer3_outputs(3075) <= a or b;
    layer3_outputs(3076) <= a or b;
    layer3_outputs(3077) <= not a or b;
    layer3_outputs(3078) <= not a or b;
    layer3_outputs(3079) <= a;
    layer3_outputs(3080) <= b;
    layer3_outputs(3081) <= 1'b1;
    layer3_outputs(3082) <= 1'b0;
    layer3_outputs(3083) <= not a;
    layer3_outputs(3084) <= not a or b;
    layer3_outputs(3085) <= a or b;
    layer3_outputs(3086) <= b and not a;
    layer3_outputs(3087) <= a and not b;
    layer3_outputs(3088) <= not (a xor b);
    layer3_outputs(3089) <= a and b;
    layer3_outputs(3090) <= a and not b;
    layer3_outputs(3091) <= a xor b;
    layer3_outputs(3092) <= not a or b;
    layer3_outputs(3093) <= a and b;
    layer3_outputs(3094) <= b and not a;
    layer3_outputs(3095) <= not (a xor b);
    layer3_outputs(3096) <= a;
    layer3_outputs(3097) <= a or b;
    layer3_outputs(3098) <= not b or a;
    layer3_outputs(3099) <= not b;
    layer3_outputs(3100) <= 1'b1;
    layer3_outputs(3101) <= b and not a;
    layer3_outputs(3102) <= a;
    layer3_outputs(3103) <= not b;
    layer3_outputs(3104) <= a and b;
    layer3_outputs(3105) <= not a;
    layer3_outputs(3106) <= not a or b;
    layer3_outputs(3107) <= b;
    layer3_outputs(3108) <= not b;
    layer3_outputs(3109) <= a xor b;
    layer3_outputs(3110) <= 1'b0;
    layer3_outputs(3111) <= not (a xor b);
    layer3_outputs(3112) <= a and not b;
    layer3_outputs(3113) <= 1'b0;
    layer3_outputs(3114) <= a and b;
    layer3_outputs(3115) <= b and not a;
    layer3_outputs(3116) <= a and b;
    layer3_outputs(3117) <= a and not b;
    layer3_outputs(3118) <= a and b;
    layer3_outputs(3119) <= 1'b1;
    layer3_outputs(3120) <= b;
    layer3_outputs(3121) <= not b;
    layer3_outputs(3122) <= b and not a;
    layer3_outputs(3123) <= not (a and b);
    layer3_outputs(3124) <= a;
    layer3_outputs(3125) <= not (a and b);
    layer3_outputs(3126) <= not (a or b);
    layer3_outputs(3127) <= not a or b;
    layer3_outputs(3128) <= b and not a;
    layer3_outputs(3129) <= not a;
    layer3_outputs(3130) <= 1'b1;
    layer3_outputs(3131) <= b;
    layer3_outputs(3132) <= not a;
    layer3_outputs(3133) <= not b;
    layer3_outputs(3134) <= a;
    layer3_outputs(3135) <= b;
    layer3_outputs(3136) <= a and b;
    layer3_outputs(3137) <= 1'b0;
    layer3_outputs(3138) <= a and b;
    layer3_outputs(3139) <= a and not b;
    layer3_outputs(3140) <= not a;
    layer3_outputs(3141) <= a xor b;
    layer3_outputs(3142) <= a or b;
    layer3_outputs(3143) <= a and b;
    layer3_outputs(3144) <= 1'b1;
    layer3_outputs(3145) <= b;
    layer3_outputs(3146) <= not a;
    layer3_outputs(3147) <= not a or b;
    layer3_outputs(3148) <= 1'b0;
    layer3_outputs(3149) <= a or b;
    layer3_outputs(3150) <= not (a or b);
    layer3_outputs(3151) <= a and not b;
    layer3_outputs(3152) <= 1'b1;
    layer3_outputs(3153) <= not (a xor b);
    layer3_outputs(3154) <= not b or a;
    layer3_outputs(3155) <= not b or a;
    layer3_outputs(3156) <= 1'b1;
    layer3_outputs(3157) <= a xor b;
    layer3_outputs(3158) <= not b;
    layer3_outputs(3159) <= 1'b0;
    layer3_outputs(3160) <= a or b;
    layer3_outputs(3161) <= not (a and b);
    layer3_outputs(3162) <= a or b;
    layer3_outputs(3163) <= not (a xor b);
    layer3_outputs(3164) <= a and b;
    layer3_outputs(3165) <= b and not a;
    layer3_outputs(3166) <= 1'b1;
    layer3_outputs(3167) <= a or b;
    layer3_outputs(3168) <= 1'b1;
    layer3_outputs(3169) <= b;
    layer3_outputs(3170) <= not b or a;
    layer3_outputs(3171) <= a and not b;
    layer3_outputs(3172) <= a and not b;
    layer3_outputs(3173) <= 1'b0;
    layer3_outputs(3174) <= not a or b;
    layer3_outputs(3175) <= not (a or b);
    layer3_outputs(3176) <= a and b;
    layer3_outputs(3177) <= a and b;
    layer3_outputs(3178) <= 1'b1;
    layer3_outputs(3179) <= a and b;
    layer3_outputs(3180) <= 1'b0;
    layer3_outputs(3181) <= a;
    layer3_outputs(3182) <= a and b;
    layer3_outputs(3183) <= not (a xor b);
    layer3_outputs(3184) <= not b or a;
    layer3_outputs(3185) <= not a;
    layer3_outputs(3186) <= b and not a;
    layer3_outputs(3187) <= b;
    layer3_outputs(3188) <= b and not a;
    layer3_outputs(3189) <= not b;
    layer3_outputs(3190) <= not (a and b);
    layer3_outputs(3191) <= not (a or b);
    layer3_outputs(3192) <= a;
    layer3_outputs(3193) <= 1'b1;
    layer3_outputs(3194) <= 1'b0;
    layer3_outputs(3195) <= not a or b;
    layer3_outputs(3196) <= not a or b;
    layer3_outputs(3197) <= not a or b;
    layer3_outputs(3198) <= a;
    layer3_outputs(3199) <= a and b;
    layer3_outputs(3200) <= not (a and b);
    layer3_outputs(3201) <= not (a and b);
    layer3_outputs(3202) <= not (a or b);
    layer3_outputs(3203) <= b;
    layer3_outputs(3204) <= a xor b;
    layer3_outputs(3205) <= a and not b;
    layer3_outputs(3206) <= not (a or b);
    layer3_outputs(3207) <= not b;
    layer3_outputs(3208) <= a or b;
    layer3_outputs(3209) <= 1'b1;
    layer3_outputs(3210) <= not (a or b);
    layer3_outputs(3211) <= a and not b;
    layer3_outputs(3212) <= not a;
    layer3_outputs(3213) <= a;
    layer3_outputs(3214) <= not b or a;
    layer3_outputs(3215) <= not (a or b);
    layer3_outputs(3216) <= not (a or b);
    layer3_outputs(3217) <= 1'b0;
    layer3_outputs(3218) <= not b;
    layer3_outputs(3219) <= a and not b;
    layer3_outputs(3220) <= a;
    layer3_outputs(3221) <= not (a or b);
    layer3_outputs(3222) <= 1'b1;
    layer3_outputs(3223) <= b;
    layer3_outputs(3224) <= a and b;
    layer3_outputs(3225) <= not a;
    layer3_outputs(3226) <= b;
    layer3_outputs(3227) <= b and not a;
    layer3_outputs(3228) <= 1'b0;
    layer3_outputs(3229) <= not (a or b);
    layer3_outputs(3230) <= not a or b;
    layer3_outputs(3231) <= b;
    layer3_outputs(3232) <= 1'b0;
    layer3_outputs(3233) <= not (a or b);
    layer3_outputs(3234) <= not b;
    layer3_outputs(3235) <= a or b;
    layer3_outputs(3236) <= 1'b0;
    layer3_outputs(3237) <= 1'b1;
    layer3_outputs(3238) <= not b or a;
    layer3_outputs(3239) <= not a;
    layer3_outputs(3240) <= a or b;
    layer3_outputs(3241) <= 1'b1;
    layer3_outputs(3242) <= a;
    layer3_outputs(3243) <= not (a or b);
    layer3_outputs(3244) <= not a;
    layer3_outputs(3245) <= a;
    layer3_outputs(3246) <= 1'b1;
    layer3_outputs(3247) <= 1'b0;
    layer3_outputs(3248) <= a and b;
    layer3_outputs(3249) <= a or b;
    layer3_outputs(3250) <= b and not a;
    layer3_outputs(3251) <= a and b;
    layer3_outputs(3252) <= a and not b;
    layer3_outputs(3253) <= not b or a;
    layer3_outputs(3254) <= b and not a;
    layer3_outputs(3255) <= b;
    layer3_outputs(3256) <= 1'b1;
    layer3_outputs(3257) <= not b or a;
    layer3_outputs(3258) <= a and not b;
    layer3_outputs(3259) <= not (a and b);
    layer3_outputs(3260) <= not a or b;
    layer3_outputs(3261) <= not (a and b);
    layer3_outputs(3262) <= a and b;
    layer3_outputs(3263) <= 1'b1;
    layer3_outputs(3264) <= not a or b;
    layer3_outputs(3265) <= b;
    layer3_outputs(3266) <= 1'b1;
    layer3_outputs(3267) <= not b;
    layer3_outputs(3268) <= 1'b0;
    layer3_outputs(3269) <= a xor b;
    layer3_outputs(3270) <= 1'b1;
    layer3_outputs(3271) <= not (a or b);
    layer3_outputs(3272) <= not (a and b);
    layer3_outputs(3273) <= a or b;
    layer3_outputs(3274) <= b;
    layer3_outputs(3275) <= a or b;
    layer3_outputs(3276) <= not b;
    layer3_outputs(3277) <= b and not a;
    layer3_outputs(3278) <= not a or b;
    layer3_outputs(3279) <= a and b;
    layer3_outputs(3280) <= not b;
    layer3_outputs(3281) <= not b;
    layer3_outputs(3282) <= a or b;
    layer3_outputs(3283) <= b and not a;
    layer3_outputs(3284) <= 1'b1;
    layer3_outputs(3285) <= not a or b;
    layer3_outputs(3286) <= a;
    layer3_outputs(3287) <= not b;
    layer3_outputs(3288) <= not a or b;
    layer3_outputs(3289) <= a and b;
    layer3_outputs(3290) <= not b or a;
    layer3_outputs(3291) <= not a or b;
    layer3_outputs(3292) <= b and not a;
    layer3_outputs(3293) <= a and not b;
    layer3_outputs(3294) <= a or b;
    layer3_outputs(3295) <= a and not b;
    layer3_outputs(3296) <= not (a and b);
    layer3_outputs(3297) <= b;
    layer3_outputs(3298) <= a or b;
    layer3_outputs(3299) <= b;
    layer3_outputs(3300) <= not (a and b);
    layer3_outputs(3301) <= not (a and b);
    layer3_outputs(3302) <= not a;
    layer3_outputs(3303) <= not b or a;
    layer3_outputs(3304) <= b;
    layer3_outputs(3305) <= 1'b0;
    layer3_outputs(3306) <= not a;
    layer3_outputs(3307) <= not (a and b);
    layer3_outputs(3308) <= not (a xor b);
    layer3_outputs(3309) <= b and not a;
    layer3_outputs(3310) <= 1'b0;
    layer3_outputs(3311) <= 1'b0;
    layer3_outputs(3312) <= a and b;
    layer3_outputs(3313) <= a and not b;
    layer3_outputs(3314) <= not a or b;
    layer3_outputs(3315) <= b and not a;
    layer3_outputs(3316) <= a;
    layer3_outputs(3317) <= a and not b;
    layer3_outputs(3318) <= not (a and b);
    layer3_outputs(3319) <= 1'b1;
    layer3_outputs(3320) <= a or b;
    layer3_outputs(3321) <= b;
    layer3_outputs(3322) <= not (a or b);
    layer3_outputs(3323) <= 1'b1;
    layer3_outputs(3324) <= a;
    layer3_outputs(3325) <= not b or a;
    layer3_outputs(3326) <= not (a xor b);
    layer3_outputs(3327) <= not b;
    layer3_outputs(3328) <= 1'b1;
    layer3_outputs(3329) <= a or b;
    layer3_outputs(3330) <= b and not a;
    layer3_outputs(3331) <= a or b;
    layer3_outputs(3332) <= not a or b;
    layer3_outputs(3333) <= a and b;
    layer3_outputs(3334) <= not b;
    layer3_outputs(3335) <= a;
    layer3_outputs(3336) <= b;
    layer3_outputs(3337) <= 1'b0;
    layer3_outputs(3338) <= b and not a;
    layer3_outputs(3339) <= a xor b;
    layer3_outputs(3340) <= not (a and b);
    layer3_outputs(3341) <= a or b;
    layer3_outputs(3342) <= not (a and b);
    layer3_outputs(3343) <= not (a or b);
    layer3_outputs(3344) <= not a or b;
    layer3_outputs(3345) <= a xor b;
    layer3_outputs(3346) <= not a or b;
    layer3_outputs(3347) <= not a;
    layer3_outputs(3348) <= b;
    layer3_outputs(3349) <= a;
    layer3_outputs(3350) <= a;
    layer3_outputs(3351) <= not (a and b);
    layer3_outputs(3352) <= not b or a;
    layer3_outputs(3353) <= 1'b1;
    layer3_outputs(3354) <= a and not b;
    layer3_outputs(3355) <= not (a or b);
    layer3_outputs(3356) <= not b;
    layer3_outputs(3357) <= not (a or b);
    layer3_outputs(3358) <= 1'b0;
    layer3_outputs(3359) <= a and b;
    layer3_outputs(3360) <= a or b;
    layer3_outputs(3361) <= not a;
    layer3_outputs(3362) <= a;
    layer3_outputs(3363) <= 1'b0;
    layer3_outputs(3364) <= 1'b0;
    layer3_outputs(3365) <= not b or a;
    layer3_outputs(3366) <= 1'b1;
    layer3_outputs(3367) <= not a;
    layer3_outputs(3368) <= not (a and b);
    layer3_outputs(3369) <= a and b;
    layer3_outputs(3370) <= a and not b;
    layer3_outputs(3371) <= not b;
    layer3_outputs(3372) <= b and not a;
    layer3_outputs(3373) <= 1'b0;
    layer3_outputs(3374) <= 1'b0;
    layer3_outputs(3375) <= not (a or b);
    layer3_outputs(3376) <= b and not a;
    layer3_outputs(3377) <= 1'b0;
    layer3_outputs(3378) <= a and b;
    layer3_outputs(3379) <= b;
    layer3_outputs(3380) <= a or b;
    layer3_outputs(3381) <= a or b;
    layer3_outputs(3382) <= not a or b;
    layer3_outputs(3383) <= not (a and b);
    layer3_outputs(3384) <= not a;
    layer3_outputs(3385) <= a;
    layer3_outputs(3386) <= 1'b1;
    layer3_outputs(3387) <= not a or b;
    layer3_outputs(3388) <= not (a and b);
    layer3_outputs(3389) <= b and not a;
    layer3_outputs(3390) <= b and not a;
    layer3_outputs(3391) <= b;
    layer3_outputs(3392) <= a or b;
    layer3_outputs(3393) <= not b or a;
    layer3_outputs(3394) <= not a or b;
    layer3_outputs(3395) <= a and b;
    layer3_outputs(3396) <= 1'b1;
    layer3_outputs(3397) <= b;
    layer3_outputs(3398) <= not (a or b);
    layer3_outputs(3399) <= not b or a;
    layer3_outputs(3400) <= 1'b1;
    layer3_outputs(3401) <= 1'b1;
    layer3_outputs(3402) <= not a;
    layer3_outputs(3403) <= b;
    layer3_outputs(3404) <= not b or a;
    layer3_outputs(3405) <= a;
    layer3_outputs(3406) <= a and b;
    layer3_outputs(3407) <= a;
    layer3_outputs(3408) <= b and not a;
    layer3_outputs(3409) <= not b or a;
    layer3_outputs(3410) <= not b;
    layer3_outputs(3411) <= 1'b1;
    layer3_outputs(3412) <= not (a or b);
    layer3_outputs(3413) <= 1'b1;
    layer3_outputs(3414) <= not (a or b);
    layer3_outputs(3415) <= not (a and b);
    layer3_outputs(3416) <= a or b;
    layer3_outputs(3417) <= b;
    layer3_outputs(3418) <= b;
    layer3_outputs(3419) <= not b;
    layer3_outputs(3420) <= a and b;
    layer3_outputs(3421) <= not b or a;
    layer3_outputs(3422) <= a and not b;
    layer3_outputs(3423) <= not (a xor b);
    layer3_outputs(3424) <= not a or b;
    layer3_outputs(3425) <= a and not b;
    layer3_outputs(3426) <= not (a and b);
    layer3_outputs(3427) <= b and not a;
    layer3_outputs(3428) <= not (a or b);
    layer3_outputs(3429) <= a and not b;
    layer3_outputs(3430) <= 1'b1;
    layer3_outputs(3431) <= not (a and b);
    layer3_outputs(3432) <= 1'b1;
    layer3_outputs(3433) <= not b or a;
    layer3_outputs(3434) <= b and not a;
    layer3_outputs(3435) <= a and b;
    layer3_outputs(3436) <= not b;
    layer3_outputs(3437) <= a and not b;
    layer3_outputs(3438) <= 1'b0;
    layer3_outputs(3439) <= not a;
    layer3_outputs(3440) <= not (a and b);
    layer3_outputs(3441) <= 1'b1;
    layer3_outputs(3442) <= a;
    layer3_outputs(3443) <= not a;
    layer3_outputs(3444) <= b;
    layer3_outputs(3445) <= not a;
    layer3_outputs(3446) <= not a or b;
    layer3_outputs(3447) <= b and not a;
    layer3_outputs(3448) <= b;
    layer3_outputs(3449) <= b and not a;
    layer3_outputs(3450) <= a or b;
    layer3_outputs(3451) <= b;
    layer3_outputs(3452) <= a;
    layer3_outputs(3453) <= a and not b;
    layer3_outputs(3454) <= not a;
    layer3_outputs(3455) <= a and not b;
    layer3_outputs(3456) <= 1'b0;
    layer3_outputs(3457) <= a;
    layer3_outputs(3458) <= a and b;
    layer3_outputs(3459) <= a or b;
    layer3_outputs(3460) <= not a;
    layer3_outputs(3461) <= b;
    layer3_outputs(3462) <= a or b;
    layer3_outputs(3463) <= not a or b;
    layer3_outputs(3464) <= 1'b0;
    layer3_outputs(3465) <= not b or a;
    layer3_outputs(3466) <= not (a and b);
    layer3_outputs(3467) <= b and not a;
    layer3_outputs(3468) <= not b or a;
    layer3_outputs(3469) <= 1'b1;
    layer3_outputs(3470) <= b;
    layer3_outputs(3471) <= a;
    layer3_outputs(3472) <= not (a and b);
    layer3_outputs(3473) <= not a;
    layer3_outputs(3474) <= not (a xor b);
    layer3_outputs(3475) <= 1'b1;
    layer3_outputs(3476) <= a and not b;
    layer3_outputs(3477) <= a or b;
    layer3_outputs(3478) <= not (a xor b);
    layer3_outputs(3479) <= b and not a;
    layer3_outputs(3480) <= b and not a;
    layer3_outputs(3481) <= a and not b;
    layer3_outputs(3482) <= not a;
    layer3_outputs(3483) <= a and b;
    layer3_outputs(3484) <= a and b;
    layer3_outputs(3485) <= b;
    layer3_outputs(3486) <= b and not a;
    layer3_outputs(3487) <= not a;
    layer3_outputs(3488) <= not (a xor b);
    layer3_outputs(3489) <= a;
    layer3_outputs(3490) <= a or b;
    layer3_outputs(3491) <= 1'b0;
    layer3_outputs(3492) <= a and not b;
    layer3_outputs(3493) <= b and not a;
    layer3_outputs(3494) <= not (a xor b);
    layer3_outputs(3495) <= a and not b;
    layer3_outputs(3496) <= not a;
    layer3_outputs(3497) <= not a or b;
    layer3_outputs(3498) <= 1'b1;
    layer3_outputs(3499) <= a;
    layer3_outputs(3500) <= a;
    layer3_outputs(3501) <= not (a xor b);
    layer3_outputs(3502) <= a;
    layer3_outputs(3503) <= b and not a;
    layer3_outputs(3504) <= not a or b;
    layer3_outputs(3505) <= not a or b;
    layer3_outputs(3506) <= a xor b;
    layer3_outputs(3507) <= b and not a;
    layer3_outputs(3508) <= a and b;
    layer3_outputs(3509) <= not a or b;
    layer3_outputs(3510) <= not (a or b);
    layer3_outputs(3511) <= 1'b0;
    layer3_outputs(3512) <= 1'b0;
    layer3_outputs(3513) <= not a or b;
    layer3_outputs(3514) <= not (a and b);
    layer3_outputs(3515) <= not a or b;
    layer3_outputs(3516) <= not a;
    layer3_outputs(3517) <= not a;
    layer3_outputs(3518) <= not (a or b);
    layer3_outputs(3519) <= b and not a;
    layer3_outputs(3520) <= not (a and b);
    layer3_outputs(3521) <= a or b;
    layer3_outputs(3522) <= a or b;
    layer3_outputs(3523) <= a and b;
    layer3_outputs(3524) <= a or b;
    layer3_outputs(3525) <= not b;
    layer3_outputs(3526) <= a and not b;
    layer3_outputs(3527) <= not (a and b);
    layer3_outputs(3528) <= not b;
    layer3_outputs(3529) <= not b or a;
    layer3_outputs(3530) <= not b or a;
    layer3_outputs(3531) <= a and b;
    layer3_outputs(3532) <= not b or a;
    layer3_outputs(3533) <= 1'b1;
    layer3_outputs(3534) <= a or b;
    layer3_outputs(3535) <= a and b;
    layer3_outputs(3536) <= a and not b;
    layer3_outputs(3537) <= a xor b;
    layer3_outputs(3538) <= 1'b1;
    layer3_outputs(3539) <= b and not a;
    layer3_outputs(3540) <= 1'b0;
    layer3_outputs(3541) <= a or b;
    layer3_outputs(3542) <= not a or b;
    layer3_outputs(3543) <= not b;
    layer3_outputs(3544) <= not a;
    layer3_outputs(3545) <= a or b;
    layer3_outputs(3546) <= b;
    layer3_outputs(3547) <= a and not b;
    layer3_outputs(3548) <= b and not a;
    layer3_outputs(3549) <= a;
    layer3_outputs(3550) <= not b or a;
    layer3_outputs(3551) <= a and not b;
    layer3_outputs(3552) <= 1'b1;
    layer3_outputs(3553) <= not b;
    layer3_outputs(3554) <= 1'b0;
    layer3_outputs(3555) <= not a or b;
    layer3_outputs(3556) <= a or b;
    layer3_outputs(3557) <= b and not a;
    layer3_outputs(3558) <= a xor b;
    layer3_outputs(3559) <= b;
    layer3_outputs(3560) <= not b or a;
    layer3_outputs(3561) <= b;
    layer3_outputs(3562) <= a;
    layer3_outputs(3563) <= not b;
    layer3_outputs(3564) <= 1'b1;
    layer3_outputs(3565) <= a;
    layer3_outputs(3566) <= b;
    layer3_outputs(3567) <= not (a and b);
    layer3_outputs(3568) <= not (a and b);
    layer3_outputs(3569) <= not (a and b);
    layer3_outputs(3570) <= not a or b;
    layer3_outputs(3571) <= not (a and b);
    layer3_outputs(3572) <= 1'b0;
    layer3_outputs(3573) <= b and not a;
    layer3_outputs(3574) <= 1'b0;
    layer3_outputs(3575) <= not (a xor b);
    layer3_outputs(3576) <= b and not a;
    layer3_outputs(3577) <= a and not b;
    layer3_outputs(3578) <= b and not a;
    layer3_outputs(3579) <= b and not a;
    layer3_outputs(3580) <= a or b;
    layer3_outputs(3581) <= not b;
    layer3_outputs(3582) <= not (a xor b);
    layer3_outputs(3583) <= a or b;
    layer3_outputs(3584) <= not (a and b);
    layer3_outputs(3585) <= a and not b;
    layer3_outputs(3586) <= a or b;
    layer3_outputs(3587) <= not a;
    layer3_outputs(3588) <= b and not a;
    layer3_outputs(3589) <= not a;
    layer3_outputs(3590) <= a and b;
    layer3_outputs(3591) <= b;
    layer3_outputs(3592) <= b and not a;
    layer3_outputs(3593) <= a or b;
    layer3_outputs(3594) <= not (a or b);
    layer3_outputs(3595) <= not a or b;
    layer3_outputs(3596) <= not a or b;
    layer3_outputs(3597) <= a and not b;
    layer3_outputs(3598) <= a;
    layer3_outputs(3599) <= not b;
    layer3_outputs(3600) <= not a;
    layer3_outputs(3601) <= b and not a;
    layer3_outputs(3602) <= not a;
    layer3_outputs(3603) <= a or b;
    layer3_outputs(3604) <= 1'b0;
    layer3_outputs(3605) <= not a or b;
    layer3_outputs(3606) <= b;
    layer3_outputs(3607) <= b and not a;
    layer3_outputs(3608) <= not b;
    layer3_outputs(3609) <= not (a and b);
    layer3_outputs(3610) <= 1'b0;
    layer3_outputs(3611) <= not a;
    layer3_outputs(3612) <= a and not b;
    layer3_outputs(3613) <= not b or a;
    layer3_outputs(3614) <= not a;
    layer3_outputs(3615) <= b;
    layer3_outputs(3616) <= 1'b0;
    layer3_outputs(3617) <= not a;
    layer3_outputs(3618) <= not a;
    layer3_outputs(3619) <= a or b;
    layer3_outputs(3620) <= 1'b0;
    layer3_outputs(3621) <= a xor b;
    layer3_outputs(3622) <= not (a and b);
    layer3_outputs(3623) <= not a;
    layer3_outputs(3624) <= a;
    layer3_outputs(3625) <= not (a and b);
    layer3_outputs(3626) <= not (a or b);
    layer3_outputs(3627) <= not (a or b);
    layer3_outputs(3628) <= not (a and b);
    layer3_outputs(3629) <= a and b;
    layer3_outputs(3630) <= a and not b;
    layer3_outputs(3631) <= not (a and b);
    layer3_outputs(3632) <= a and not b;
    layer3_outputs(3633) <= 1'b1;
    layer3_outputs(3634) <= a or b;
    layer3_outputs(3635) <= not a;
    layer3_outputs(3636) <= not (a or b);
    layer3_outputs(3637) <= a xor b;
    layer3_outputs(3638) <= a and not b;
    layer3_outputs(3639) <= a;
    layer3_outputs(3640) <= a and not b;
    layer3_outputs(3641) <= a;
    layer3_outputs(3642) <= a or b;
    layer3_outputs(3643) <= a or b;
    layer3_outputs(3644) <= not a or b;
    layer3_outputs(3645) <= a and b;
    layer3_outputs(3646) <= not b;
    layer3_outputs(3647) <= not b;
    layer3_outputs(3648) <= not a or b;
    layer3_outputs(3649) <= not a;
    layer3_outputs(3650) <= not a;
    layer3_outputs(3651) <= not (a and b);
    layer3_outputs(3652) <= not a;
    layer3_outputs(3653) <= not (a or b);
    layer3_outputs(3654) <= a;
    layer3_outputs(3655) <= not b;
    layer3_outputs(3656) <= not b;
    layer3_outputs(3657) <= a;
    layer3_outputs(3658) <= 1'b0;
    layer3_outputs(3659) <= not (a or b);
    layer3_outputs(3660) <= not (a or b);
    layer3_outputs(3661) <= a;
    layer3_outputs(3662) <= 1'b1;
    layer3_outputs(3663) <= 1'b0;
    layer3_outputs(3664) <= not a;
    layer3_outputs(3665) <= 1'b0;
    layer3_outputs(3666) <= 1'b0;
    layer3_outputs(3667) <= not b or a;
    layer3_outputs(3668) <= a;
    layer3_outputs(3669) <= a;
    layer3_outputs(3670) <= 1'b1;
    layer3_outputs(3671) <= not b or a;
    layer3_outputs(3672) <= not a or b;
    layer3_outputs(3673) <= not (a xor b);
    layer3_outputs(3674) <= a;
    layer3_outputs(3675) <= not a or b;
    layer3_outputs(3676) <= 1'b0;
    layer3_outputs(3677) <= not a;
    layer3_outputs(3678) <= not (a or b);
    layer3_outputs(3679) <= 1'b1;
    layer3_outputs(3680) <= a and not b;
    layer3_outputs(3681) <= not b or a;
    layer3_outputs(3682) <= a or b;
    layer3_outputs(3683) <= a;
    layer3_outputs(3684) <= not b or a;
    layer3_outputs(3685) <= not (a or b);
    layer3_outputs(3686) <= not a;
    layer3_outputs(3687) <= 1'b1;
    layer3_outputs(3688) <= not (a and b);
    layer3_outputs(3689) <= a and not b;
    layer3_outputs(3690) <= not (a and b);
    layer3_outputs(3691) <= not a or b;
    layer3_outputs(3692) <= not b;
    layer3_outputs(3693) <= not b;
    layer3_outputs(3694) <= a and not b;
    layer3_outputs(3695) <= not b;
    layer3_outputs(3696) <= 1'b1;
    layer3_outputs(3697) <= a and b;
    layer3_outputs(3698) <= not (a or b);
    layer3_outputs(3699) <= not (a and b);
    layer3_outputs(3700) <= a and b;
    layer3_outputs(3701) <= not (a or b);
    layer3_outputs(3702) <= not b;
    layer3_outputs(3703) <= not (a or b);
    layer3_outputs(3704) <= a and not b;
    layer3_outputs(3705) <= b and not a;
    layer3_outputs(3706) <= not a or b;
    layer3_outputs(3707) <= not (a and b);
    layer3_outputs(3708) <= a or b;
    layer3_outputs(3709) <= not (a xor b);
    layer3_outputs(3710) <= not (a or b);
    layer3_outputs(3711) <= b and not a;
    layer3_outputs(3712) <= a;
    layer3_outputs(3713) <= a and not b;
    layer3_outputs(3714) <= not b;
    layer3_outputs(3715) <= a;
    layer3_outputs(3716) <= b;
    layer3_outputs(3717) <= a or b;
    layer3_outputs(3718) <= not b;
    layer3_outputs(3719) <= not a or b;
    layer3_outputs(3720) <= a or b;
    layer3_outputs(3721) <= not (a and b);
    layer3_outputs(3722) <= a;
    layer3_outputs(3723) <= not b or a;
    layer3_outputs(3724) <= not b or a;
    layer3_outputs(3725) <= a or b;
    layer3_outputs(3726) <= not a or b;
    layer3_outputs(3727) <= not b or a;
    layer3_outputs(3728) <= a;
    layer3_outputs(3729) <= not (a or b);
    layer3_outputs(3730) <= b and not a;
    layer3_outputs(3731) <= b;
    layer3_outputs(3732) <= a and not b;
    layer3_outputs(3733) <= not (a and b);
    layer3_outputs(3734) <= a and b;
    layer3_outputs(3735) <= not a or b;
    layer3_outputs(3736) <= not (a or b);
    layer3_outputs(3737) <= b and not a;
    layer3_outputs(3738) <= a and not b;
    layer3_outputs(3739) <= a and not b;
    layer3_outputs(3740) <= 1'b1;
    layer3_outputs(3741) <= 1'b0;
    layer3_outputs(3742) <= a and not b;
    layer3_outputs(3743) <= a and not b;
    layer3_outputs(3744) <= a and b;
    layer3_outputs(3745) <= not b or a;
    layer3_outputs(3746) <= a and not b;
    layer3_outputs(3747) <= b and not a;
    layer3_outputs(3748) <= b and not a;
    layer3_outputs(3749) <= a and b;
    layer3_outputs(3750) <= not a;
    layer3_outputs(3751) <= a;
    layer3_outputs(3752) <= not (a and b);
    layer3_outputs(3753) <= not b;
    layer3_outputs(3754) <= not (a and b);
    layer3_outputs(3755) <= not a or b;
    layer3_outputs(3756) <= not a;
    layer3_outputs(3757) <= 1'b1;
    layer3_outputs(3758) <= a or b;
    layer3_outputs(3759) <= a xor b;
    layer3_outputs(3760) <= not (a and b);
    layer3_outputs(3761) <= not b or a;
    layer3_outputs(3762) <= not (a and b);
    layer3_outputs(3763) <= not (a or b);
    layer3_outputs(3764) <= 1'b1;
    layer3_outputs(3765) <= not b;
    layer3_outputs(3766) <= not (a xor b);
    layer3_outputs(3767) <= not (a and b);
    layer3_outputs(3768) <= not b;
    layer3_outputs(3769) <= a and b;
    layer3_outputs(3770) <= 1'b0;
    layer3_outputs(3771) <= not (a or b);
    layer3_outputs(3772) <= not b;
    layer3_outputs(3773) <= b;
    layer3_outputs(3774) <= not (a or b);
    layer3_outputs(3775) <= not a or b;
    layer3_outputs(3776) <= 1'b0;
    layer3_outputs(3777) <= not (a or b);
    layer3_outputs(3778) <= a and not b;
    layer3_outputs(3779) <= not (a or b);
    layer3_outputs(3780) <= 1'b1;
    layer3_outputs(3781) <= 1'b1;
    layer3_outputs(3782) <= not b;
    layer3_outputs(3783) <= not a;
    layer3_outputs(3784) <= not (a or b);
    layer3_outputs(3785) <= a xor b;
    layer3_outputs(3786) <= b;
    layer3_outputs(3787) <= a or b;
    layer3_outputs(3788) <= not a;
    layer3_outputs(3789) <= not a;
    layer3_outputs(3790) <= a xor b;
    layer3_outputs(3791) <= not a;
    layer3_outputs(3792) <= b;
    layer3_outputs(3793) <= b and not a;
    layer3_outputs(3794) <= not b;
    layer3_outputs(3795) <= b and not a;
    layer3_outputs(3796) <= not b or a;
    layer3_outputs(3797) <= a;
    layer3_outputs(3798) <= not (a and b);
    layer3_outputs(3799) <= a and b;
    layer3_outputs(3800) <= not a;
    layer3_outputs(3801) <= not a;
    layer3_outputs(3802) <= 1'b1;
    layer3_outputs(3803) <= 1'b0;
    layer3_outputs(3804) <= a or b;
    layer3_outputs(3805) <= a;
    layer3_outputs(3806) <= 1'b0;
    layer3_outputs(3807) <= not b or a;
    layer3_outputs(3808) <= not a;
    layer3_outputs(3809) <= not (a and b);
    layer3_outputs(3810) <= b;
    layer3_outputs(3811) <= a and b;
    layer3_outputs(3812) <= a;
    layer3_outputs(3813) <= not a or b;
    layer3_outputs(3814) <= 1'b0;
    layer3_outputs(3815) <= not a or b;
    layer3_outputs(3816) <= a and not b;
    layer3_outputs(3817) <= b and not a;
    layer3_outputs(3818) <= not b or a;
    layer3_outputs(3819) <= not a or b;
    layer3_outputs(3820) <= not a;
    layer3_outputs(3821) <= b;
    layer3_outputs(3822) <= a and b;
    layer3_outputs(3823) <= 1'b1;
    layer3_outputs(3824) <= not (a and b);
    layer3_outputs(3825) <= a or b;
    layer3_outputs(3826) <= not b;
    layer3_outputs(3827) <= not a;
    layer3_outputs(3828) <= a xor b;
    layer3_outputs(3829) <= not (a and b);
    layer3_outputs(3830) <= not (a and b);
    layer3_outputs(3831) <= a or b;
    layer3_outputs(3832) <= not a or b;
    layer3_outputs(3833) <= not a;
    layer3_outputs(3834) <= 1'b1;
    layer3_outputs(3835) <= b and not a;
    layer3_outputs(3836) <= not (a and b);
    layer3_outputs(3837) <= b and not a;
    layer3_outputs(3838) <= a and not b;
    layer3_outputs(3839) <= 1'b1;
    layer3_outputs(3840) <= 1'b0;
    layer3_outputs(3841) <= not (a and b);
    layer3_outputs(3842) <= not a;
    layer3_outputs(3843) <= 1'b1;
    layer3_outputs(3844) <= b;
    layer3_outputs(3845) <= not a;
    layer3_outputs(3846) <= not b;
    layer3_outputs(3847) <= b and not a;
    layer3_outputs(3848) <= not a;
    layer3_outputs(3849) <= a and b;
    layer3_outputs(3850) <= not b;
    layer3_outputs(3851) <= a;
    layer3_outputs(3852) <= not a or b;
    layer3_outputs(3853) <= not a or b;
    layer3_outputs(3854) <= not (a xor b);
    layer3_outputs(3855) <= a;
    layer3_outputs(3856) <= not b;
    layer3_outputs(3857) <= 1'b1;
    layer3_outputs(3858) <= 1'b1;
    layer3_outputs(3859) <= a or b;
    layer3_outputs(3860) <= not a;
    layer3_outputs(3861) <= b;
    layer3_outputs(3862) <= not (a or b);
    layer3_outputs(3863) <= not b or a;
    layer3_outputs(3864) <= not a;
    layer3_outputs(3865) <= 1'b1;
    layer3_outputs(3866) <= not b;
    layer3_outputs(3867) <= b and not a;
    layer3_outputs(3868) <= a and b;
    layer3_outputs(3869) <= not (a and b);
    layer3_outputs(3870) <= not a or b;
    layer3_outputs(3871) <= not (a xor b);
    layer3_outputs(3872) <= not (a and b);
    layer3_outputs(3873) <= 1'b0;
    layer3_outputs(3874) <= a;
    layer3_outputs(3875) <= a and b;
    layer3_outputs(3876) <= not a or b;
    layer3_outputs(3877) <= not a;
    layer3_outputs(3878) <= a xor b;
    layer3_outputs(3879) <= not a;
    layer3_outputs(3880) <= a xor b;
    layer3_outputs(3881) <= a;
    layer3_outputs(3882) <= not (a or b);
    layer3_outputs(3883) <= not (a and b);
    layer3_outputs(3884) <= a and not b;
    layer3_outputs(3885) <= a xor b;
    layer3_outputs(3886) <= a and b;
    layer3_outputs(3887) <= a or b;
    layer3_outputs(3888) <= not a;
    layer3_outputs(3889) <= not a;
    layer3_outputs(3890) <= b and not a;
    layer3_outputs(3891) <= a;
    layer3_outputs(3892) <= not a or b;
    layer3_outputs(3893) <= a and not b;
    layer3_outputs(3894) <= a and not b;
    layer3_outputs(3895) <= a and not b;
    layer3_outputs(3896) <= b;
    layer3_outputs(3897) <= not (a or b);
    layer3_outputs(3898) <= a and b;
    layer3_outputs(3899) <= 1'b0;
    layer3_outputs(3900) <= 1'b0;
    layer3_outputs(3901) <= not b;
    layer3_outputs(3902) <= a;
    layer3_outputs(3903) <= 1'b1;
    layer3_outputs(3904) <= 1'b1;
    layer3_outputs(3905) <= a;
    layer3_outputs(3906) <= a or b;
    layer3_outputs(3907) <= a xor b;
    layer3_outputs(3908) <= not a or b;
    layer3_outputs(3909) <= a or b;
    layer3_outputs(3910) <= not a or b;
    layer3_outputs(3911) <= a and not b;
    layer3_outputs(3912) <= not a or b;
    layer3_outputs(3913) <= not a;
    layer3_outputs(3914) <= b and not a;
    layer3_outputs(3915) <= not (a or b);
    layer3_outputs(3916) <= not (a and b);
    layer3_outputs(3917) <= not b;
    layer3_outputs(3918) <= not a or b;
    layer3_outputs(3919) <= not (a and b);
    layer3_outputs(3920) <= not b or a;
    layer3_outputs(3921) <= b and not a;
    layer3_outputs(3922) <= a and b;
    layer3_outputs(3923) <= not b;
    layer3_outputs(3924) <= 1'b1;
    layer3_outputs(3925) <= b;
    layer3_outputs(3926) <= not a or b;
    layer3_outputs(3927) <= not b or a;
    layer3_outputs(3928) <= a xor b;
    layer3_outputs(3929) <= a or b;
    layer3_outputs(3930) <= not a;
    layer3_outputs(3931) <= a and b;
    layer3_outputs(3932) <= 1'b0;
    layer3_outputs(3933) <= not a;
    layer3_outputs(3934) <= a and b;
    layer3_outputs(3935) <= not (a and b);
    layer3_outputs(3936) <= 1'b1;
    layer3_outputs(3937) <= 1'b1;
    layer3_outputs(3938) <= not (a and b);
    layer3_outputs(3939) <= b and not a;
    layer3_outputs(3940) <= not a or b;
    layer3_outputs(3941) <= 1'b0;
    layer3_outputs(3942) <= a or b;
    layer3_outputs(3943) <= not b;
    layer3_outputs(3944) <= a and not b;
    layer3_outputs(3945) <= not a;
    layer3_outputs(3946) <= a and b;
    layer3_outputs(3947) <= not (a and b);
    layer3_outputs(3948) <= not b or a;
    layer3_outputs(3949) <= a or b;
    layer3_outputs(3950) <= not b;
    layer3_outputs(3951) <= not b;
    layer3_outputs(3952) <= a;
    layer3_outputs(3953) <= 1'b0;
    layer3_outputs(3954) <= 1'b1;
    layer3_outputs(3955) <= a or b;
    layer3_outputs(3956) <= not b;
    layer3_outputs(3957) <= 1'b0;
    layer3_outputs(3958) <= a;
    layer3_outputs(3959) <= a;
    layer3_outputs(3960) <= 1'b1;
    layer3_outputs(3961) <= a;
    layer3_outputs(3962) <= b;
    layer3_outputs(3963) <= a and not b;
    layer3_outputs(3964) <= a;
    layer3_outputs(3965) <= b and not a;
    layer3_outputs(3966) <= b;
    layer3_outputs(3967) <= a and b;
    layer3_outputs(3968) <= 1'b0;
    layer3_outputs(3969) <= not (a or b);
    layer3_outputs(3970) <= not (a and b);
    layer3_outputs(3971) <= not b;
    layer3_outputs(3972) <= not (a or b);
    layer3_outputs(3973) <= not a;
    layer3_outputs(3974) <= a xor b;
    layer3_outputs(3975) <= 1'b1;
    layer3_outputs(3976) <= 1'b1;
    layer3_outputs(3977) <= a or b;
    layer3_outputs(3978) <= not a or b;
    layer3_outputs(3979) <= not a;
    layer3_outputs(3980) <= a and b;
    layer3_outputs(3981) <= a and not b;
    layer3_outputs(3982) <= a or b;
    layer3_outputs(3983) <= 1'b1;
    layer3_outputs(3984) <= a or b;
    layer3_outputs(3985) <= not (a and b);
    layer3_outputs(3986) <= 1'b1;
    layer3_outputs(3987) <= not b or a;
    layer3_outputs(3988) <= a and not b;
    layer3_outputs(3989) <= not a or b;
    layer3_outputs(3990) <= b and not a;
    layer3_outputs(3991) <= not a;
    layer3_outputs(3992) <= a and b;
    layer3_outputs(3993) <= 1'b1;
    layer3_outputs(3994) <= a and b;
    layer3_outputs(3995) <= not a;
    layer3_outputs(3996) <= 1'b1;
    layer3_outputs(3997) <= not (a xor b);
    layer3_outputs(3998) <= a or b;
    layer3_outputs(3999) <= not b;
    layer3_outputs(4000) <= not (a or b);
    layer3_outputs(4001) <= not a or b;
    layer3_outputs(4002) <= not a;
    layer3_outputs(4003) <= b;
    layer3_outputs(4004) <= 1'b0;
    layer3_outputs(4005) <= not (a or b);
    layer3_outputs(4006) <= a xor b;
    layer3_outputs(4007) <= not a;
    layer3_outputs(4008) <= not b or a;
    layer3_outputs(4009) <= a and not b;
    layer3_outputs(4010) <= not b;
    layer3_outputs(4011) <= not (a and b);
    layer3_outputs(4012) <= a or b;
    layer3_outputs(4013) <= not (a or b);
    layer3_outputs(4014) <= a and not b;
    layer3_outputs(4015) <= not b or a;
    layer3_outputs(4016) <= 1'b0;
    layer3_outputs(4017) <= not (a and b);
    layer3_outputs(4018) <= a;
    layer3_outputs(4019) <= b and not a;
    layer3_outputs(4020) <= not (a or b);
    layer3_outputs(4021) <= not (a and b);
    layer3_outputs(4022) <= a and b;
    layer3_outputs(4023) <= b and not a;
    layer3_outputs(4024) <= not (a or b);
    layer3_outputs(4025) <= a;
    layer3_outputs(4026) <= 1'b1;
    layer3_outputs(4027) <= not (a or b);
    layer3_outputs(4028) <= b;
    layer3_outputs(4029) <= not b;
    layer3_outputs(4030) <= not a or b;
    layer3_outputs(4031) <= b and not a;
    layer3_outputs(4032) <= not b;
    layer3_outputs(4033) <= not b;
    layer3_outputs(4034) <= not b;
    layer3_outputs(4035) <= not b;
    layer3_outputs(4036) <= a and not b;
    layer3_outputs(4037) <= a or b;
    layer3_outputs(4038) <= not a or b;
    layer3_outputs(4039) <= b;
    layer3_outputs(4040) <= not a or b;
    layer3_outputs(4041) <= a and not b;
    layer3_outputs(4042) <= b and not a;
    layer3_outputs(4043) <= a or b;
    layer3_outputs(4044) <= 1'b1;
    layer3_outputs(4045) <= 1'b0;
    layer3_outputs(4046) <= b;
    layer3_outputs(4047) <= a xor b;
    layer3_outputs(4048) <= a and b;
    layer3_outputs(4049) <= a and not b;
    layer3_outputs(4050) <= 1'b0;
    layer3_outputs(4051) <= not (a and b);
    layer3_outputs(4052) <= not a;
    layer3_outputs(4053) <= not a;
    layer3_outputs(4054) <= a or b;
    layer3_outputs(4055) <= not (a or b);
    layer3_outputs(4056) <= b and not a;
    layer3_outputs(4057) <= 1'b0;
    layer3_outputs(4058) <= not (a or b);
    layer3_outputs(4059) <= a or b;
    layer3_outputs(4060) <= 1'b0;
    layer3_outputs(4061) <= b;
    layer3_outputs(4062) <= 1'b0;
    layer3_outputs(4063) <= 1'b1;
    layer3_outputs(4064) <= not (a or b);
    layer3_outputs(4065) <= not a or b;
    layer3_outputs(4066) <= 1'b1;
    layer3_outputs(4067) <= a;
    layer3_outputs(4068) <= b;
    layer3_outputs(4069) <= a;
    layer3_outputs(4070) <= b;
    layer3_outputs(4071) <= 1'b0;
    layer3_outputs(4072) <= not b;
    layer3_outputs(4073) <= a and b;
    layer3_outputs(4074) <= a and b;
    layer3_outputs(4075) <= 1'b1;
    layer3_outputs(4076) <= a or b;
    layer3_outputs(4077) <= a xor b;
    layer3_outputs(4078) <= b;
    layer3_outputs(4079) <= b and not a;
    layer3_outputs(4080) <= 1'b1;
    layer3_outputs(4081) <= a and not b;
    layer3_outputs(4082) <= not a or b;
    layer3_outputs(4083) <= a and b;
    layer3_outputs(4084) <= not (a xor b);
    layer3_outputs(4085) <= 1'b0;
    layer3_outputs(4086) <= not b or a;
    layer3_outputs(4087) <= not b or a;
    layer3_outputs(4088) <= b and not a;
    layer3_outputs(4089) <= b;
    layer3_outputs(4090) <= a and b;
    layer3_outputs(4091) <= not (a or b);
    layer3_outputs(4092) <= a and not b;
    layer3_outputs(4093) <= not a or b;
    layer3_outputs(4094) <= not a;
    layer3_outputs(4095) <= b;
    layer3_outputs(4096) <= 1'b1;
    layer3_outputs(4097) <= b and not a;
    layer3_outputs(4098) <= not b;
    layer3_outputs(4099) <= not (a or b);
    layer3_outputs(4100) <= not (a and b);
    layer3_outputs(4101) <= not (a or b);
    layer3_outputs(4102) <= a and not b;
    layer3_outputs(4103) <= not b;
    layer3_outputs(4104) <= not (a xor b);
    layer3_outputs(4105) <= a or b;
    layer3_outputs(4106) <= b;
    layer3_outputs(4107) <= a;
    layer3_outputs(4108) <= b and not a;
    layer3_outputs(4109) <= 1'b0;
    layer3_outputs(4110) <= not b;
    layer3_outputs(4111) <= not (a xor b);
    layer3_outputs(4112) <= b;
    layer3_outputs(4113) <= a and not b;
    layer3_outputs(4114) <= b;
    layer3_outputs(4115) <= a or b;
    layer3_outputs(4116) <= not a;
    layer3_outputs(4117) <= 1'b1;
    layer3_outputs(4118) <= a and b;
    layer3_outputs(4119) <= b and not a;
    layer3_outputs(4120) <= 1'b0;
    layer3_outputs(4121) <= a and b;
    layer3_outputs(4122) <= b;
    layer3_outputs(4123) <= not (a and b);
    layer3_outputs(4124) <= a and not b;
    layer3_outputs(4125) <= b and not a;
    layer3_outputs(4126) <= a and not b;
    layer3_outputs(4127) <= not b or a;
    layer3_outputs(4128) <= 1'b1;
    layer3_outputs(4129) <= b;
    layer3_outputs(4130) <= b and not a;
    layer3_outputs(4131) <= 1'b1;
    layer3_outputs(4132) <= a and b;
    layer3_outputs(4133) <= not (a or b);
    layer3_outputs(4134) <= a;
    layer3_outputs(4135) <= not b;
    layer3_outputs(4136) <= a;
    layer3_outputs(4137) <= 1'b1;
    layer3_outputs(4138) <= a and b;
    layer3_outputs(4139) <= not (a and b);
    layer3_outputs(4140) <= 1'b1;
    layer3_outputs(4141) <= a and not b;
    layer3_outputs(4142) <= not (a or b);
    layer3_outputs(4143) <= a;
    layer3_outputs(4144) <= a or b;
    layer3_outputs(4145) <= 1'b0;
    layer3_outputs(4146) <= not b or a;
    layer3_outputs(4147) <= not b or a;
    layer3_outputs(4148) <= b and not a;
    layer3_outputs(4149) <= 1'b0;
    layer3_outputs(4150) <= 1'b0;
    layer3_outputs(4151) <= b and not a;
    layer3_outputs(4152) <= b and not a;
    layer3_outputs(4153) <= b;
    layer3_outputs(4154) <= 1'b0;
    layer3_outputs(4155) <= not (a or b);
    layer3_outputs(4156) <= not a or b;
    layer3_outputs(4157) <= a and b;
    layer3_outputs(4158) <= a and not b;
    layer3_outputs(4159) <= not a;
    layer3_outputs(4160) <= b;
    layer3_outputs(4161) <= not (a xor b);
    layer3_outputs(4162) <= a and b;
    layer3_outputs(4163) <= b and not a;
    layer3_outputs(4164) <= not a;
    layer3_outputs(4165) <= a;
    layer3_outputs(4166) <= not (a and b);
    layer3_outputs(4167) <= b;
    layer3_outputs(4168) <= a and not b;
    layer3_outputs(4169) <= 1'b0;
    layer3_outputs(4170) <= not (a and b);
    layer3_outputs(4171) <= a and b;
    layer3_outputs(4172) <= 1'b1;
    layer3_outputs(4173) <= 1'b0;
    layer3_outputs(4174) <= not a or b;
    layer3_outputs(4175) <= 1'b0;
    layer3_outputs(4176) <= b and not a;
    layer3_outputs(4177) <= not a;
    layer3_outputs(4178) <= a xor b;
    layer3_outputs(4179) <= a or b;
    layer3_outputs(4180) <= a or b;
    layer3_outputs(4181) <= b and not a;
    layer3_outputs(4182) <= 1'b0;
    layer3_outputs(4183) <= not b;
    layer3_outputs(4184) <= a;
    layer3_outputs(4185) <= a and b;
    layer3_outputs(4186) <= not (a and b);
    layer3_outputs(4187) <= a and not b;
    layer3_outputs(4188) <= not (a and b);
    layer3_outputs(4189) <= a and b;
    layer3_outputs(4190) <= not b;
    layer3_outputs(4191) <= 1'b0;
    layer3_outputs(4192) <= not a;
    layer3_outputs(4193) <= not b;
    layer3_outputs(4194) <= not a or b;
    layer3_outputs(4195) <= not (a or b);
    layer3_outputs(4196) <= not b or a;
    layer3_outputs(4197) <= not (a and b);
    layer3_outputs(4198) <= not a or b;
    layer3_outputs(4199) <= a;
    layer3_outputs(4200) <= not (a or b);
    layer3_outputs(4201) <= b and not a;
    layer3_outputs(4202) <= a and not b;
    layer3_outputs(4203) <= a;
    layer3_outputs(4204) <= a and b;
    layer3_outputs(4205) <= b;
    layer3_outputs(4206) <= not a;
    layer3_outputs(4207) <= 1'b0;
    layer3_outputs(4208) <= not (a and b);
    layer3_outputs(4209) <= not b;
    layer3_outputs(4210) <= not b;
    layer3_outputs(4211) <= a and not b;
    layer3_outputs(4212) <= 1'b0;
    layer3_outputs(4213) <= not b or a;
    layer3_outputs(4214) <= not (a or b);
    layer3_outputs(4215) <= a;
    layer3_outputs(4216) <= not (a or b);
    layer3_outputs(4217) <= a xor b;
    layer3_outputs(4218) <= a;
    layer3_outputs(4219) <= not a or b;
    layer3_outputs(4220) <= not a;
    layer3_outputs(4221) <= not b or a;
    layer3_outputs(4222) <= not (a xor b);
    layer3_outputs(4223) <= a;
    layer3_outputs(4224) <= not (a and b);
    layer3_outputs(4225) <= not a or b;
    layer3_outputs(4226) <= 1'b1;
    layer3_outputs(4227) <= 1'b0;
    layer3_outputs(4228) <= a or b;
    layer3_outputs(4229) <= 1'b0;
    layer3_outputs(4230) <= a and not b;
    layer3_outputs(4231) <= a;
    layer3_outputs(4232) <= a;
    layer3_outputs(4233) <= not b or a;
    layer3_outputs(4234) <= a and not b;
    layer3_outputs(4235) <= not (a and b);
    layer3_outputs(4236) <= not b;
    layer3_outputs(4237) <= not a or b;
    layer3_outputs(4238) <= 1'b1;
    layer3_outputs(4239) <= not b or a;
    layer3_outputs(4240) <= not b or a;
    layer3_outputs(4241) <= not b or a;
    layer3_outputs(4242) <= a and not b;
    layer3_outputs(4243) <= not a;
    layer3_outputs(4244) <= 1'b1;
    layer3_outputs(4245) <= a or b;
    layer3_outputs(4246) <= not (a or b);
    layer3_outputs(4247) <= not b;
    layer3_outputs(4248) <= not (a or b);
    layer3_outputs(4249) <= not a;
    layer3_outputs(4250) <= a;
    layer3_outputs(4251) <= not b or a;
    layer3_outputs(4252) <= not (a or b);
    layer3_outputs(4253) <= a and b;
    layer3_outputs(4254) <= a and not b;
    layer3_outputs(4255) <= not (a and b);
    layer3_outputs(4256) <= a or b;
    layer3_outputs(4257) <= 1'b1;
    layer3_outputs(4258) <= a or b;
    layer3_outputs(4259) <= b;
    layer3_outputs(4260) <= a and not b;
    layer3_outputs(4261) <= 1'b0;
    layer3_outputs(4262) <= not (a and b);
    layer3_outputs(4263) <= 1'b0;
    layer3_outputs(4264) <= b and not a;
    layer3_outputs(4265) <= not b or a;
    layer3_outputs(4266) <= not b or a;
    layer3_outputs(4267) <= 1'b1;
    layer3_outputs(4268) <= not a;
    layer3_outputs(4269) <= 1'b0;
    layer3_outputs(4270) <= a and b;
    layer3_outputs(4271) <= not (a or b);
    layer3_outputs(4272) <= not b;
    layer3_outputs(4273) <= 1'b0;
    layer3_outputs(4274) <= not (a and b);
    layer3_outputs(4275) <= not (a xor b);
    layer3_outputs(4276) <= not b or a;
    layer3_outputs(4277) <= b;
    layer3_outputs(4278) <= not (a and b);
    layer3_outputs(4279) <= b and not a;
    layer3_outputs(4280) <= b;
    layer3_outputs(4281) <= a or b;
    layer3_outputs(4282) <= not b;
    layer3_outputs(4283) <= b and not a;
    layer3_outputs(4284) <= b and not a;
    layer3_outputs(4285) <= not a or b;
    layer3_outputs(4286) <= not b or a;
    layer3_outputs(4287) <= not (a or b);
    layer3_outputs(4288) <= a and b;
    layer3_outputs(4289) <= not (a and b);
    layer3_outputs(4290) <= a and not b;
    layer3_outputs(4291) <= 1'b0;
    layer3_outputs(4292) <= 1'b0;
    layer3_outputs(4293) <= not b;
    layer3_outputs(4294) <= a and not b;
    layer3_outputs(4295) <= a or b;
    layer3_outputs(4296) <= a and not b;
    layer3_outputs(4297) <= not (a and b);
    layer3_outputs(4298) <= b;
    layer3_outputs(4299) <= not (a or b);
    layer3_outputs(4300) <= b;
    layer3_outputs(4301) <= not b or a;
    layer3_outputs(4302) <= a and not b;
    layer3_outputs(4303) <= not (a or b);
    layer3_outputs(4304) <= a and not b;
    layer3_outputs(4305) <= not (a and b);
    layer3_outputs(4306) <= not b;
    layer3_outputs(4307) <= not b or a;
    layer3_outputs(4308) <= not (a and b);
    layer3_outputs(4309) <= not b or a;
    layer3_outputs(4310) <= a or b;
    layer3_outputs(4311) <= not b or a;
    layer3_outputs(4312) <= a or b;
    layer3_outputs(4313) <= not (a or b);
    layer3_outputs(4314) <= b;
    layer3_outputs(4315) <= not a;
    layer3_outputs(4316) <= not b;
    layer3_outputs(4317) <= 1'b1;
    layer3_outputs(4318) <= not (a or b);
    layer3_outputs(4319) <= not (a xor b);
    layer3_outputs(4320) <= not b;
    layer3_outputs(4321) <= a xor b;
    layer3_outputs(4322) <= not (a and b);
    layer3_outputs(4323) <= b;
    layer3_outputs(4324) <= not a or b;
    layer3_outputs(4325) <= b;
    layer3_outputs(4326) <= not a or b;
    layer3_outputs(4327) <= a and b;
    layer3_outputs(4328) <= b;
    layer3_outputs(4329) <= not a or b;
    layer3_outputs(4330) <= a;
    layer3_outputs(4331) <= 1'b1;
    layer3_outputs(4332) <= not (a and b);
    layer3_outputs(4333) <= not a;
    layer3_outputs(4334) <= a and b;
    layer3_outputs(4335) <= not (a and b);
    layer3_outputs(4336) <= not (a or b);
    layer3_outputs(4337) <= a;
    layer3_outputs(4338) <= a and not b;
    layer3_outputs(4339) <= a;
    layer3_outputs(4340) <= b and not a;
    layer3_outputs(4341) <= b;
    layer3_outputs(4342) <= b and not a;
    layer3_outputs(4343) <= b and not a;
    layer3_outputs(4344) <= not b;
    layer3_outputs(4345) <= not (a and b);
    layer3_outputs(4346) <= not (a and b);
    layer3_outputs(4347) <= not (a and b);
    layer3_outputs(4348) <= not (a or b);
    layer3_outputs(4349) <= a or b;
    layer3_outputs(4350) <= a xor b;
    layer3_outputs(4351) <= not (a and b);
    layer3_outputs(4352) <= not (a xor b);
    layer3_outputs(4353) <= a or b;
    layer3_outputs(4354) <= not (a and b);
    layer3_outputs(4355) <= not (a or b);
    layer3_outputs(4356) <= not (a or b);
    layer3_outputs(4357) <= 1'b0;
    layer3_outputs(4358) <= not (a and b);
    layer3_outputs(4359) <= a and b;
    layer3_outputs(4360) <= 1'b0;
    layer3_outputs(4361) <= not b or a;
    layer3_outputs(4362) <= 1'b0;
    layer3_outputs(4363) <= 1'b0;
    layer3_outputs(4364) <= a and not b;
    layer3_outputs(4365) <= a and b;
    layer3_outputs(4366) <= a;
    layer3_outputs(4367) <= 1'b1;
    layer3_outputs(4368) <= not (a and b);
    layer3_outputs(4369) <= a and not b;
    layer3_outputs(4370) <= 1'b1;
    layer3_outputs(4371) <= not b or a;
    layer3_outputs(4372) <= 1'b0;
    layer3_outputs(4373) <= not b or a;
    layer3_outputs(4374) <= 1'b1;
    layer3_outputs(4375) <= 1'b1;
    layer3_outputs(4376) <= a and not b;
    layer3_outputs(4377) <= a and b;
    layer3_outputs(4378) <= a or b;
    layer3_outputs(4379) <= not b;
    layer3_outputs(4380) <= b;
    layer3_outputs(4381) <= not a or b;
    layer3_outputs(4382) <= not (a or b);
    layer3_outputs(4383) <= not a or b;
    layer3_outputs(4384) <= a and not b;
    layer3_outputs(4385) <= 1'b1;
    layer3_outputs(4386) <= b;
    layer3_outputs(4387) <= a or b;
    layer3_outputs(4388) <= b;
    layer3_outputs(4389) <= not b or a;
    layer3_outputs(4390) <= b and not a;
    layer3_outputs(4391) <= not a or b;
    layer3_outputs(4392) <= 1'b0;
    layer3_outputs(4393) <= b and not a;
    layer3_outputs(4394) <= not (a and b);
    layer3_outputs(4395) <= a or b;
    layer3_outputs(4396) <= 1'b1;
    layer3_outputs(4397) <= a;
    layer3_outputs(4398) <= not (a or b);
    layer3_outputs(4399) <= a or b;
    layer3_outputs(4400) <= not b or a;
    layer3_outputs(4401) <= not a or b;
    layer3_outputs(4402) <= not (a or b);
    layer3_outputs(4403) <= 1'b1;
    layer3_outputs(4404) <= a and b;
    layer3_outputs(4405) <= not (a and b);
    layer3_outputs(4406) <= a;
    layer3_outputs(4407) <= not (a or b);
    layer3_outputs(4408) <= 1'b0;
    layer3_outputs(4409) <= a and b;
    layer3_outputs(4410) <= not b;
    layer3_outputs(4411) <= 1'b1;
    layer3_outputs(4412) <= not b or a;
    layer3_outputs(4413) <= a and b;
    layer3_outputs(4414) <= not (a and b);
    layer3_outputs(4415) <= not b;
    layer3_outputs(4416) <= a;
    layer3_outputs(4417) <= a;
    layer3_outputs(4418) <= 1'b0;
    layer3_outputs(4419) <= not b;
    layer3_outputs(4420) <= a and b;
    layer3_outputs(4421) <= not a;
    layer3_outputs(4422) <= a xor b;
    layer3_outputs(4423) <= a and b;
    layer3_outputs(4424) <= b and not a;
    layer3_outputs(4425) <= b;
    layer3_outputs(4426) <= b and not a;
    layer3_outputs(4427) <= b and not a;
    layer3_outputs(4428) <= 1'b1;
    layer3_outputs(4429) <= not (a or b);
    layer3_outputs(4430) <= not (a xor b);
    layer3_outputs(4431) <= not (a xor b);
    layer3_outputs(4432) <= not (a or b);
    layer3_outputs(4433) <= b and not a;
    layer3_outputs(4434) <= a and not b;
    layer3_outputs(4435) <= not (a or b);
    layer3_outputs(4436) <= a or b;
    layer3_outputs(4437) <= a;
    layer3_outputs(4438) <= b;
    layer3_outputs(4439) <= not b;
    layer3_outputs(4440) <= b and not a;
    layer3_outputs(4441) <= not a or b;
    layer3_outputs(4442) <= a;
    layer3_outputs(4443) <= not (a and b);
    layer3_outputs(4444) <= b and not a;
    layer3_outputs(4445) <= not b or a;
    layer3_outputs(4446) <= a and b;
    layer3_outputs(4447) <= a or b;
    layer3_outputs(4448) <= not b;
    layer3_outputs(4449) <= 1'b1;
    layer3_outputs(4450) <= a and b;
    layer3_outputs(4451) <= not (a and b);
    layer3_outputs(4452) <= a and b;
    layer3_outputs(4453) <= b and not a;
    layer3_outputs(4454) <= b;
    layer3_outputs(4455) <= b and not a;
    layer3_outputs(4456) <= not b or a;
    layer3_outputs(4457) <= not a;
    layer3_outputs(4458) <= 1'b0;
    layer3_outputs(4459) <= b;
    layer3_outputs(4460) <= 1'b0;
    layer3_outputs(4461) <= not a or b;
    layer3_outputs(4462) <= not a;
    layer3_outputs(4463) <= a and b;
    layer3_outputs(4464) <= a or b;
    layer3_outputs(4465) <= not b;
    layer3_outputs(4466) <= b and not a;
    layer3_outputs(4467) <= not a;
    layer3_outputs(4468) <= not (a and b);
    layer3_outputs(4469) <= a;
    layer3_outputs(4470) <= a or b;
    layer3_outputs(4471) <= not a;
    layer3_outputs(4472) <= a;
    layer3_outputs(4473) <= not a;
    layer3_outputs(4474) <= a and not b;
    layer3_outputs(4475) <= not b;
    layer3_outputs(4476) <= a;
    layer3_outputs(4477) <= not b;
    layer3_outputs(4478) <= 1'b0;
    layer3_outputs(4479) <= not a or b;
    layer3_outputs(4480) <= 1'b1;
    layer3_outputs(4481) <= not a;
    layer3_outputs(4482) <= a and not b;
    layer3_outputs(4483) <= not (a and b);
    layer3_outputs(4484) <= 1'b0;
    layer3_outputs(4485) <= b and not a;
    layer3_outputs(4486) <= not (a xor b);
    layer3_outputs(4487) <= not b;
    layer3_outputs(4488) <= 1'b0;
    layer3_outputs(4489) <= 1'b1;
    layer3_outputs(4490) <= a or b;
    layer3_outputs(4491) <= a;
    layer3_outputs(4492) <= b and not a;
    layer3_outputs(4493) <= not a;
    layer3_outputs(4494) <= b and not a;
    layer3_outputs(4495) <= b and not a;
    layer3_outputs(4496) <= b and not a;
    layer3_outputs(4497) <= not (a or b);
    layer3_outputs(4498) <= b;
    layer3_outputs(4499) <= not b;
    layer3_outputs(4500) <= 1'b0;
    layer3_outputs(4501) <= a or b;
    layer3_outputs(4502) <= not b;
    layer3_outputs(4503) <= a and b;
    layer3_outputs(4504) <= b and not a;
    layer3_outputs(4505) <= not a;
    layer3_outputs(4506) <= not (a and b);
    layer3_outputs(4507) <= 1'b0;
    layer3_outputs(4508) <= 1'b1;
    layer3_outputs(4509) <= a and b;
    layer3_outputs(4510) <= a;
    layer3_outputs(4511) <= not a;
    layer3_outputs(4512) <= 1'b0;
    layer3_outputs(4513) <= not b;
    layer3_outputs(4514) <= a;
    layer3_outputs(4515) <= 1'b0;
    layer3_outputs(4516) <= not a;
    layer3_outputs(4517) <= a and b;
    layer3_outputs(4518) <= 1'b0;
    layer3_outputs(4519) <= a or b;
    layer3_outputs(4520) <= not a or b;
    layer3_outputs(4521) <= not (a or b);
    layer3_outputs(4522) <= b and not a;
    layer3_outputs(4523) <= a or b;
    layer3_outputs(4524) <= not b or a;
    layer3_outputs(4525) <= not b or a;
    layer3_outputs(4526) <= not b or a;
    layer3_outputs(4527) <= b and not a;
    layer3_outputs(4528) <= not b;
    layer3_outputs(4529) <= not a or b;
    layer3_outputs(4530) <= not (a and b);
    layer3_outputs(4531) <= not b or a;
    layer3_outputs(4532) <= a and b;
    layer3_outputs(4533) <= b;
    layer3_outputs(4534) <= not (a or b);
    layer3_outputs(4535) <= 1'b1;
    layer3_outputs(4536) <= a;
    layer3_outputs(4537) <= 1'b0;
    layer3_outputs(4538) <= not b;
    layer3_outputs(4539) <= a;
    layer3_outputs(4540) <= a and not b;
    layer3_outputs(4541) <= not b;
    layer3_outputs(4542) <= b and not a;
    layer3_outputs(4543) <= 1'b0;
    layer3_outputs(4544) <= not b or a;
    layer3_outputs(4545) <= a or b;
    layer3_outputs(4546) <= a xor b;
    layer3_outputs(4547) <= not b;
    layer3_outputs(4548) <= not a or b;
    layer3_outputs(4549) <= not a or b;
    layer3_outputs(4550) <= not (a or b);
    layer3_outputs(4551) <= not (a or b);
    layer3_outputs(4552) <= not (a and b);
    layer3_outputs(4553) <= a;
    layer3_outputs(4554) <= not b;
    layer3_outputs(4555) <= b;
    layer3_outputs(4556) <= not b;
    layer3_outputs(4557) <= not (a and b);
    layer3_outputs(4558) <= not a;
    layer3_outputs(4559) <= b and not a;
    layer3_outputs(4560) <= 1'b0;
    layer3_outputs(4561) <= a and b;
    layer3_outputs(4562) <= not b or a;
    layer3_outputs(4563) <= not (a or b);
    layer3_outputs(4564) <= not b or a;
    layer3_outputs(4565) <= not a or b;
    layer3_outputs(4566) <= not b or a;
    layer3_outputs(4567) <= not b;
    layer3_outputs(4568) <= b and not a;
    layer3_outputs(4569) <= 1'b1;
    layer3_outputs(4570) <= b and not a;
    layer3_outputs(4571) <= a and b;
    layer3_outputs(4572) <= 1'b0;
    layer3_outputs(4573) <= a or b;
    layer3_outputs(4574) <= b and not a;
    layer3_outputs(4575) <= not b or a;
    layer3_outputs(4576) <= not (a and b);
    layer3_outputs(4577) <= not b or a;
    layer3_outputs(4578) <= not (a and b);
    layer3_outputs(4579) <= not a or b;
    layer3_outputs(4580) <= a;
    layer3_outputs(4581) <= not b;
    layer3_outputs(4582) <= not a or b;
    layer3_outputs(4583) <= not b;
    layer3_outputs(4584) <= not (a and b);
    layer3_outputs(4585) <= a and not b;
    layer3_outputs(4586) <= not b or a;
    layer3_outputs(4587) <= a;
    layer3_outputs(4588) <= b and not a;
    layer3_outputs(4589) <= a and b;
    layer3_outputs(4590) <= not a;
    layer3_outputs(4591) <= not a or b;
    layer3_outputs(4592) <= a or b;
    layer3_outputs(4593) <= 1'b0;
    layer3_outputs(4594) <= a;
    layer3_outputs(4595) <= b and not a;
    layer3_outputs(4596) <= b and not a;
    layer3_outputs(4597) <= not b;
    layer3_outputs(4598) <= not a or b;
    layer3_outputs(4599) <= not b;
    layer3_outputs(4600) <= not (a and b);
    layer3_outputs(4601) <= not a or b;
    layer3_outputs(4602) <= not b or a;
    layer3_outputs(4603) <= not (a and b);
    layer3_outputs(4604) <= a;
    layer3_outputs(4605) <= 1'b0;
    layer3_outputs(4606) <= not (a and b);
    layer3_outputs(4607) <= not b or a;
    layer3_outputs(4608) <= 1'b1;
    layer3_outputs(4609) <= a or b;
    layer3_outputs(4610) <= a and b;
    layer3_outputs(4611) <= 1'b1;
    layer3_outputs(4612) <= not b or a;
    layer3_outputs(4613) <= b and not a;
    layer3_outputs(4614) <= a and not b;
    layer3_outputs(4615) <= not (a or b);
    layer3_outputs(4616) <= not a or b;
    layer3_outputs(4617) <= not a or b;
    layer3_outputs(4618) <= 1'b0;
    layer3_outputs(4619) <= b and not a;
    layer3_outputs(4620) <= 1'b0;
    layer3_outputs(4621) <= 1'b0;
    layer3_outputs(4622) <= not a;
    layer3_outputs(4623) <= not b;
    layer3_outputs(4624) <= 1'b0;
    layer3_outputs(4625) <= a;
    layer3_outputs(4626) <= 1'b0;
    layer3_outputs(4627) <= a and not b;
    layer3_outputs(4628) <= not (a and b);
    layer3_outputs(4629) <= not b or a;
    layer3_outputs(4630) <= a and b;
    layer3_outputs(4631) <= not a or b;
    layer3_outputs(4632) <= not a;
    layer3_outputs(4633) <= not a or b;
    layer3_outputs(4634) <= b;
    layer3_outputs(4635) <= a xor b;
    layer3_outputs(4636) <= not a or b;
    layer3_outputs(4637) <= 1'b1;
    layer3_outputs(4638) <= 1'b1;
    layer3_outputs(4639) <= b;
    layer3_outputs(4640) <= not b or a;
    layer3_outputs(4641) <= not (a or b);
    layer3_outputs(4642) <= b;
    layer3_outputs(4643) <= b and not a;
    layer3_outputs(4644) <= a;
    layer3_outputs(4645) <= 1'b1;
    layer3_outputs(4646) <= not a or b;
    layer3_outputs(4647) <= a and not b;
    layer3_outputs(4648) <= a;
    layer3_outputs(4649) <= not a;
    layer3_outputs(4650) <= not b;
    layer3_outputs(4651) <= a and not b;
    layer3_outputs(4652) <= a and not b;
    layer3_outputs(4653) <= not b;
    layer3_outputs(4654) <= not a or b;
    layer3_outputs(4655) <= not b or a;
    layer3_outputs(4656) <= a;
    layer3_outputs(4657) <= not a;
    layer3_outputs(4658) <= 1'b0;
    layer3_outputs(4659) <= a or b;
    layer3_outputs(4660) <= a;
    layer3_outputs(4661) <= not a or b;
    layer3_outputs(4662) <= a;
    layer3_outputs(4663) <= not b;
    layer3_outputs(4664) <= b and not a;
    layer3_outputs(4665) <= not b;
    layer3_outputs(4666) <= not b;
    layer3_outputs(4667) <= not (a and b);
    layer3_outputs(4668) <= a or b;
    layer3_outputs(4669) <= not b;
    layer3_outputs(4670) <= not (a or b);
    layer3_outputs(4671) <= a and not b;
    layer3_outputs(4672) <= a;
    layer3_outputs(4673) <= a or b;
    layer3_outputs(4674) <= not a or b;
    layer3_outputs(4675) <= not b or a;
    layer3_outputs(4676) <= a or b;
    layer3_outputs(4677) <= not b or a;
    layer3_outputs(4678) <= b and not a;
    layer3_outputs(4679) <= not b;
    layer3_outputs(4680) <= a xor b;
    layer3_outputs(4681) <= not a;
    layer3_outputs(4682) <= b and not a;
    layer3_outputs(4683) <= not (a or b);
    layer3_outputs(4684) <= not (a or b);
    layer3_outputs(4685) <= not a or b;
    layer3_outputs(4686) <= not b;
    layer3_outputs(4687) <= not b;
    layer3_outputs(4688) <= a;
    layer3_outputs(4689) <= not a or b;
    layer3_outputs(4690) <= not a;
    layer3_outputs(4691) <= b and not a;
    layer3_outputs(4692) <= not (a or b);
    layer3_outputs(4693) <= not b;
    layer3_outputs(4694) <= not b;
    layer3_outputs(4695) <= a and b;
    layer3_outputs(4696) <= b;
    layer3_outputs(4697) <= a xor b;
    layer3_outputs(4698) <= 1'b0;
    layer3_outputs(4699) <= a or b;
    layer3_outputs(4700) <= b;
    layer3_outputs(4701) <= 1'b0;
    layer3_outputs(4702) <= a;
    layer3_outputs(4703) <= b;
    layer3_outputs(4704) <= not (a and b);
    layer3_outputs(4705) <= 1'b0;
    layer3_outputs(4706) <= b;
    layer3_outputs(4707) <= not (a or b);
    layer3_outputs(4708) <= 1'b0;
    layer3_outputs(4709) <= not b;
    layer3_outputs(4710) <= not a or b;
    layer3_outputs(4711) <= not a;
    layer3_outputs(4712) <= a;
    layer3_outputs(4713) <= b;
    layer3_outputs(4714) <= not b or a;
    layer3_outputs(4715) <= not (a or b);
    layer3_outputs(4716) <= not (a and b);
    layer3_outputs(4717) <= 1'b1;
    layer3_outputs(4718) <= not a;
    layer3_outputs(4719) <= a or b;
    layer3_outputs(4720) <= b and not a;
    layer3_outputs(4721) <= not a;
    layer3_outputs(4722) <= b;
    layer3_outputs(4723) <= 1'b1;
    layer3_outputs(4724) <= not b;
    layer3_outputs(4725) <= not b;
    layer3_outputs(4726) <= b;
    layer3_outputs(4727) <= a and b;
    layer3_outputs(4728) <= not b or a;
    layer3_outputs(4729) <= not a or b;
    layer3_outputs(4730) <= not (a and b);
    layer3_outputs(4731) <= not (a or b);
    layer3_outputs(4732) <= b;
    layer3_outputs(4733) <= not b or a;
    layer3_outputs(4734) <= not b or a;
    layer3_outputs(4735) <= a or b;
    layer3_outputs(4736) <= a or b;
    layer3_outputs(4737) <= not (a xor b);
    layer3_outputs(4738) <= 1'b1;
    layer3_outputs(4739) <= not (a and b);
    layer3_outputs(4740) <= 1'b0;
    layer3_outputs(4741) <= b;
    layer3_outputs(4742) <= a and not b;
    layer3_outputs(4743) <= not a or b;
    layer3_outputs(4744) <= not b or a;
    layer3_outputs(4745) <= a xor b;
    layer3_outputs(4746) <= 1'b1;
    layer3_outputs(4747) <= not b or a;
    layer3_outputs(4748) <= a and b;
    layer3_outputs(4749) <= b and not a;
    layer3_outputs(4750) <= not b;
    layer3_outputs(4751) <= b and not a;
    layer3_outputs(4752) <= a and b;
    layer3_outputs(4753) <= not (a or b);
    layer3_outputs(4754) <= b and not a;
    layer3_outputs(4755) <= a or b;
    layer3_outputs(4756) <= a;
    layer3_outputs(4757) <= a and b;
    layer3_outputs(4758) <= a xor b;
    layer3_outputs(4759) <= a;
    layer3_outputs(4760) <= not (a or b);
    layer3_outputs(4761) <= a and not b;
    layer3_outputs(4762) <= 1'b0;
    layer3_outputs(4763) <= a;
    layer3_outputs(4764) <= a and b;
    layer3_outputs(4765) <= not (a and b);
    layer3_outputs(4766) <= b;
    layer3_outputs(4767) <= a or b;
    layer3_outputs(4768) <= a and b;
    layer3_outputs(4769) <= 1'b1;
    layer3_outputs(4770) <= 1'b0;
    layer3_outputs(4771) <= b and not a;
    layer3_outputs(4772) <= b;
    layer3_outputs(4773) <= not b;
    layer3_outputs(4774) <= not b;
    layer3_outputs(4775) <= not b;
    layer3_outputs(4776) <= not (a or b);
    layer3_outputs(4777) <= a and b;
    layer3_outputs(4778) <= 1'b1;
    layer3_outputs(4779) <= not b;
    layer3_outputs(4780) <= 1'b0;
    layer3_outputs(4781) <= b;
    layer3_outputs(4782) <= not a or b;
    layer3_outputs(4783) <= 1'b1;
    layer3_outputs(4784) <= not (a xor b);
    layer3_outputs(4785) <= b and not a;
    layer3_outputs(4786) <= not b;
    layer3_outputs(4787) <= not b or a;
    layer3_outputs(4788) <= 1'b1;
    layer3_outputs(4789) <= 1'b0;
    layer3_outputs(4790) <= a;
    layer3_outputs(4791) <= b;
    layer3_outputs(4792) <= not b;
    layer3_outputs(4793) <= 1'b1;
    layer3_outputs(4794) <= 1'b1;
    layer3_outputs(4795) <= 1'b0;
    layer3_outputs(4796) <= b;
    layer3_outputs(4797) <= not b or a;
    layer3_outputs(4798) <= b;
    layer3_outputs(4799) <= b and not a;
    layer3_outputs(4800) <= not b or a;
    layer3_outputs(4801) <= a or b;
    layer3_outputs(4802) <= 1'b1;
    layer3_outputs(4803) <= not (a xor b);
    layer3_outputs(4804) <= not a;
    layer3_outputs(4805) <= not a;
    layer3_outputs(4806) <= a or b;
    layer3_outputs(4807) <= b and not a;
    layer3_outputs(4808) <= 1'b1;
    layer3_outputs(4809) <= a and b;
    layer3_outputs(4810) <= b;
    layer3_outputs(4811) <= a;
    layer3_outputs(4812) <= b;
    layer3_outputs(4813) <= not a;
    layer3_outputs(4814) <= a and b;
    layer3_outputs(4815) <= not b or a;
    layer3_outputs(4816) <= a and b;
    layer3_outputs(4817) <= not (a and b);
    layer3_outputs(4818) <= a;
    layer3_outputs(4819) <= not b or a;
    layer3_outputs(4820) <= a and not b;
    layer3_outputs(4821) <= not b or a;
    layer3_outputs(4822) <= not a or b;
    layer3_outputs(4823) <= a and not b;
    layer3_outputs(4824) <= b and not a;
    layer3_outputs(4825) <= not a;
    layer3_outputs(4826) <= a and b;
    layer3_outputs(4827) <= a and b;
    layer3_outputs(4828) <= b and not a;
    layer3_outputs(4829) <= a and b;
    layer3_outputs(4830) <= not (a or b);
    layer3_outputs(4831) <= not b;
    layer3_outputs(4832) <= 1'b0;
    layer3_outputs(4833) <= 1'b0;
    layer3_outputs(4834) <= b and not a;
    layer3_outputs(4835) <= a;
    layer3_outputs(4836) <= a or b;
    layer3_outputs(4837) <= a and not b;
    layer3_outputs(4838) <= 1'b0;
    layer3_outputs(4839) <= 1'b0;
    layer3_outputs(4840) <= not (a and b);
    layer3_outputs(4841) <= not (a and b);
    layer3_outputs(4842) <= a;
    layer3_outputs(4843) <= a and b;
    layer3_outputs(4844) <= not a or b;
    layer3_outputs(4845) <= not b;
    layer3_outputs(4846) <= not (a or b);
    layer3_outputs(4847) <= a;
    layer3_outputs(4848) <= 1'b1;
    layer3_outputs(4849) <= a or b;
    layer3_outputs(4850) <= a or b;
    layer3_outputs(4851) <= a;
    layer3_outputs(4852) <= 1'b0;
    layer3_outputs(4853) <= not b or a;
    layer3_outputs(4854) <= not b;
    layer3_outputs(4855) <= not a;
    layer3_outputs(4856) <= not (a or b);
    layer3_outputs(4857) <= a;
    layer3_outputs(4858) <= b;
    layer3_outputs(4859) <= not (a or b);
    layer3_outputs(4860) <= not (a or b);
    layer3_outputs(4861) <= b;
    layer3_outputs(4862) <= 1'b0;
    layer3_outputs(4863) <= 1'b0;
    layer3_outputs(4864) <= not b;
    layer3_outputs(4865) <= a and b;
    layer3_outputs(4866) <= b and not a;
    layer3_outputs(4867) <= not a;
    layer3_outputs(4868) <= not (a xor b);
    layer3_outputs(4869) <= not b or a;
    layer3_outputs(4870) <= not (a and b);
    layer3_outputs(4871) <= not b or a;
    layer3_outputs(4872) <= b and not a;
    layer3_outputs(4873) <= a and not b;
    layer3_outputs(4874) <= 1'b1;
    layer3_outputs(4875) <= a and not b;
    layer3_outputs(4876) <= a xor b;
    layer3_outputs(4877) <= not (a or b);
    layer3_outputs(4878) <= 1'b1;
    layer3_outputs(4879) <= a and b;
    layer3_outputs(4880) <= not a;
    layer3_outputs(4881) <= not a;
    layer3_outputs(4882) <= not a;
    layer3_outputs(4883) <= not (a and b);
    layer3_outputs(4884) <= a and not b;
    layer3_outputs(4885) <= b;
    layer3_outputs(4886) <= b;
    layer3_outputs(4887) <= not (a and b);
    layer3_outputs(4888) <= a or b;
    layer3_outputs(4889) <= not b;
    layer3_outputs(4890) <= not a;
    layer3_outputs(4891) <= a or b;
    layer3_outputs(4892) <= 1'b0;
    layer3_outputs(4893) <= b;
    layer3_outputs(4894) <= not b or a;
    layer3_outputs(4895) <= not (a and b);
    layer3_outputs(4896) <= b;
    layer3_outputs(4897) <= not b;
    layer3_outputs(4898) <= not (a and b);
    layer3_outputs(4899) <= a;
    layer3_outputs(4900) <= b and not a;
    layer3_outputs(4901) <= 1'b1;
    layer3_outputs(4902) <= 1'b1;
    layer3_outputs(4903) <= not (a xor b);
    layer3_outputs(4904) <= a or b;
    layer3_outputs(4905) <= not (a xor b);
    layer3_outputs(4906) <= 1'b0;
    layer3_outputs(4907) <= not a;
    layer3_outputs(4908) <= not b or a;
    layer3_outputs(4909) <= a;
    layer3_outputs(4910) <= not b;
    layer3_outputs(4911) <= a and b;
    layer3_outputs(4912) <= not a;
    layer3_outputs(4913) <= 1'b1;
    layer3_outputs(4914) <= b and not a;
    layer3_outputs(4915) <= not b or a;
    layer3_outputs(4916) <= a or b;
    layer3_outputs(4917) <= not a;
    layer3_outputs(4918) <= not b or a;
    layer3_outputs(4919) <= 1'b0;
    layer3_outputs(4920) <= a;
    layer3_outputs(4921) <= a and not b;
    layer3_outputs(4922) <= b;
    layer3_outputs(4923) <= a and b;
    layer3_outputs(4924) <= 1'b1;
    layer3_outputs(4925) <= b;
    layer3_outputs(4926) <= 1'b1;
    layer3_outputs(4927) <= 1'b0;
    layer3_outputs(4928) <= a and b;
    layer3_outputs(4929) <= not b or a;
    layer3_outputs(4930) <= 1'b1;
    layer3_outputs(4931) <= not b or a;
    layer3_outputs(4932) <= a;
    layer3_outputs(4933) <= 1'b0;
    layer3_outputs(4934) <= not a;
    layer3_outputs(4935) <= b;
    layer3_outputs(4936) <= not a;
    layer3_outputs(4937) <= not (a xor b);
    layer3_outputs(4938) <= 1'b0;
    layer3_outputs(4939) <= a and b;
    layer3_outputs(4940) <= b;
    layer3_outputs(4941) <= a or b;
    layer3_outputs(4942) <= a;
    layer3_outputs(4943) <= 1'b1;
    layer3_outputs(4944) <= not (a and b);
    layer3_outputs(4945) <= 1'b1;
    layer3_outputs(4946) <= a;
    layer3_outputs(4947) <= a or b;
    layer3_outputs(4948) <= b and not a;
    layer3_outputs(4949) <= not b or a;
    layer3_outputs(4950) <= 1'b1;
    layer3_outputs(4951) <= not a;
    layer3_outputs(4952) <= 1'b0;
    layer3_outputs(4953) <= b;
    layer3_outputs(4954) <= 1'b0;
    layer3_outputs(4955) <= not a;
    layer3_outputs(4956) <= not b or a;
    layer3_outputs(4957) <= a and b;
    layer3_outputs(4958) <= not (a or b);
    layer3_outputs(4959) <= not b or a;
    layer3_outputs(4960) <= a and b;
    layer3_outputs(4961) <= not (a and b);
    layer3_outputs(4962) <= a;
    layer3_outputs(4963) <= not a;
    layer3_outputs(4964) <= a and not b;
    layer3_outputs(4965) <= a;
    layer3_outputs(4966) <= not a or b;
    layer3_outputs(4967) <= a or b;
    layer3_outputs(4968) <= a and b;
    layer3_outputs(4969) <= not (a or b);
    layer3_outputs(4970) <= b;
    layer3_outputs(4971) <= a and not b;
    layer3_outputs(4972) <= not b or a;
    layer3_outputs(4973) <= b;
    layer3_outputs(4974) <= not a;
    layer3_outputs(4975) <= a xor b;
    layer3_outputs(4976) <= not a;
    layer3_outputs(4977) <= not (a and b);
    layer3_outputs(4978) <= a and not b;
    layer3_outputs(4979) <= not a or b;
    layer3_outputs(4980) <= a;
    layer3_outputs(4981) <= a xor b;
    layer3_outputs(4982) <= b;
    layer3_outputs(4983) <= not b;
    layer3_outputs(4984) <= not a;
    layer3_outputs(4985) <= a;
    layer3_outputs(4986) <= not a;
    layer3_outputs(4987) <= a and b;
    layer3_outputs(4988) <= not b;
    layer3_outputs(4989) <= a and not b;
    layer3_outputs(4990) <= b;
    layer3_outputs(4991) <= 1'b1;
    layer3_outputs(4992) <= not (a and b);
    layer3_outputs(4993) <= not b;
    layer3_outputs(4994) <= not b or a;
    layer3_outputs(4995) <= a and b;
    layer3_outputs(4996) <= not a or b;
    layer3_outputs(4997) <= a;
    layer3_outputs(4998) <= not b;
    layer3_outputs(4999) <= 1'b0;
    layer3_outputs(5000) <= b;
    layer3_outputs(5001) <= 1'b0;
    layer3_outputs(5002) <= 1'b1;
    layer3_outputs(5003) <= not a;
    layer3_outputs(5004) <= 1'b1;
    layer3_outputs(5005) <= not a;
    layer3_outputs(5006) <= not b;
    layer3_outputs(5007) <= not a or b;
    layer3_outputs(5008) <= not (a or b);
    layer3_outputs(5009) <= not b;
    layer3_outputs(5010) <= 1'b0;
    layer3_outputs(5011) <= not b or a;
    layer3_outputs(5012) <= a;
    layer3_outputs(5013) <= not a;
    layer3_outputs(5014) <= a and not b;
    layer3_outputs(5015) <= b;
    layer3_outputs(5016) <= a and b;
    layer3_outputs(5017) <= a and b;
    layer3_outputs(5018) <= a;
    layer3_outputs(5019) <= a or b;
    layer3_outputs(5020) <= b and not a;
    layer3_outputs(5021) <= a xor b;
    layer3_outputs(5022) <= a and not b;
    layer3_outputs(5023) <= not (a or b);
    layer3_outputs(5024) <= b;
    layer3_outputs(5025) <= b;
    layer3_outputs(5026) <= a;
    layer3_outputs(5027) <= a and not b;
    layer3_outputs(5028) <= not a or b;
    layer3_outputs(5029) <= a and not b;
    layer3_outputs(5030) <= 1'b1;
    layer3_outputs(5031) <= not b or a;
    layer3_outputs(5032) <= not a or b;
    layer3_outputs(5033) <= a and b;
    layer3_outputs(5034) <= a or b;
    layer3_outputs(5035) <= not (a and b);
    layer3_outputs(5036) <= a and b;
    layer3_outputs(5037) <= b;
    layer3_outputs(5038) <= 1'b1;
    layer3_outputs(5039) <= not (a or b);
    layer3_outputs(5040) <= not (a and b);
    layer3_outputs(5041) <= not b;
    layer3_outputs(5042) <= a xor b;
    layer3_outputs(5043) <= b and not a;
    layer3_outputs(5044) <= not a;
    layer3_outputs(5045) <= a xor b;
    layer3_outputs(5046) <= 1'b0;
    layer3_outputs(5047) <= a and not b;
    layer3_outputs(5048) <= not (a and b);
    layer3_outputs(5049) <= not (a or b);
    layer3_outputs(5050) <= not b or a;
    layer3_outputs(5051) <= not a or b;
    layer3_outputs(5052) <= 1'b1;
    layer3_outputs(5053) <= a and b;
    layer3_outputs(5054) <= 1'b1;
    layer3_outputs(5055) <= not (a and b);
    layer3_outputs(5056) <= b;
    layer3_outputs(5057) <= b and not a;
    layer3_outputs(5058) <= a or b;
    layer3_outputs(5059) <= 1'b1;
    layer3_outputs(5060) <= a and b;
    layer3_outputs(5061) <= not b or a;
    layer3_outputs(5062) <= not b;
    layer3_outputs(5063) <= not b;
    layer3_outputs(5064) <= b and not a;
    layer3_outputs(5065) <= a or b;
    layer3_outputs(5066) <= 1'b0;
    layer3_outputs(5067) <= b;
    layer3_outputs(5068) <= not a;
    layer3_outputs(5069) <= not (a or b);
    layer3_outputs(5070) <= not b or a;
    layer3_outputs(5071) <= not a or b;
    layer3_outputs(5072) <= a and not b;
    layer3_outputs(5073) <= not (a xor b);
    layer3_outputs(5074) <= not b;
    layer3_outputs(5075) <= b and not a;
    layer3_outputs(5076) <= not (a and b);
    layer3_outputs(5077) <= 1'b0;
    layer3_outputs(5078) <= not b or a;
    layer3_outputs(5079) <= not a;
    layer3_outputs(5080) <= 1'b0;
    layer3_outputs(5081) <= b;
    layer3_outputs(5082) <= not (a and b);
    layer3_outputs(5083) <= not b;
    layer3_outputs(5084) <= a and b;
    layer3_outputs(5085) <= a and not b;
    layer3_outputs(5086) <= not (a or b);
    layer3_outputs(5087) <= not b;
    layer3_outputs(5088) <= a;
    layer3_outputs(5089) <= a xor b;
    layer3_outputs(5090) <= 1'b0;
    layer3_outputs(5091) <= a and not b;
    layer3_outputs(5092) <= not a or b;
    layer3_outputs(5093) <= a or b;
    layer3_outputs(5094) <= 1'b0;
    layer3_outputs(5095) <= not b or a;
    layer3_outputs(5096) <= not a;
    layer3_outputs(5097) <= not (a and b);
    layer3_outputs(5098) <= not (a or b);
    layer3_outputs(5099) <= not b or a;
    layer3_outputs(5100) <= 1'b0;
    layer3_outputs(5101) <= not (a and b);
    layer3_outputs(5102) <= 1'b1;
    layer3_outputs(5103) <= b;
    layer3_outputs(5104) <= b;
    layer3_outputs(5105) <= not (a and b);
    layer3_outputs(5106) <= 1'b1;
    layer3_outputs(5107) <= not a or b;
    layer3_outputs(5108) <= a or b;
    layer3_outputs(5109) <= not b or a;
    layer3_outputs(5110) <= a;
    layer3_outputs(5111) <= a;
    layer3_outputs(5112) <= a or b;
    layer3_outputs(5113) <= 1'b1;
    layer3_outputs(5114) <= a and b;
    layer3_outputs(5115) <= a xor b;
    layer3_outputs(5116) <= not a or b;
    layer3_outputs(5117) <= not a;
    layer3_outputs(5118) <= b and not a;
    layer3_outputs(5119) <= not (a or b);
    layer3_outputs(5120) <= not a or b;
    layer3_outputs(5121) <= not a;
    layer3_outputs(5122) <= not (a and b);
    layer3_outputs(5123) <= not a or b;
    layer3_outputs(5124) <= 1'b0;
    layer3_outputs(5125) <= not a;
    layer3_outputs(5126) <= 1'b1;
    layer3_outputs(5127) <= a and not b;
    layer3_outputs(5128) <= b and not a;
    layer3_outputs(5129) <= not b;
    layer3_outputs(5130) <= b;
    layer3_outputs(5131) <= not (a or b);
    layer3_outputs(5132) <= a and b;
    layer3_outputs(5133) <= 1'b0;
    layer3_outputs(5134) <= a;
    layer3_outputs(5135) <= not b;
    layer3_outputs(5136) <= not a;
    layer3_outputs(5137) <= not (a or b);
    layer3_outputs(5138) <= 1'b1;
    layer3_outputs(5139) <= a or b;
    layer3_outputs(5140) <= 1'b1;
    layer3_outputs(5141) <= a and b;
    layer3_outputs(5142) <= 1'b1;
    layer3_outputs(5143) <= 1'b0;
    layer3_outputs(5144) <= 1'b1;
    layer3_outputs(5145) <= not b or a;
    layer3_outputs(5146) <= a and not b;
    layer3_outputs(5147) <= b and not a;
    layer3_outputs(5148) <= 1'b1;
    layer3_outputs(5149) <= 1'b0;
    layer3_outputs(5150) <= not (a xor b);
    layer3_outputs(5151) <= a and not b;
    layer3_outputs(5152) <= a or b;
    layer3_outputs(5153) <= a and not b;
    layer3_outputs(5154) <= b and not a;
    layer3_outputs(5155) <= not a or b;
    layer3_outputs(5156) <= a;
    layer3_outputs(5157) <= not a;
    layer3_outputs(5158) <= not b or a;
    layer3_outputs(5159) <= a xor b;
    layer3_outputs(5160) <= not (a or b);
    layer3_outputs(5161) <= not b;
    layer3_outputs(5162) <= a or b;
    layer3_outputs(5163) <= 1'b0;
    layer3_outputs(5164) <= b;
    layer3_outputs(5165) <= not a or b;
    layer3_outputs(5166) <= b and not a;
    layer3_outputs(5167) <= a xor b;
    layer3_outputs(5168) <= not a;
    layer3_outputs(5169) <= not a;
    layer3_outputs(5170) <= a;
    layer3_outputs(5171) <= b;
    layer3_outputs(5172) <= not (a or b);
    layer3_outputs(5173) <= 1'b0;
    layer3_outputs(5174) <= not a or b;
    layer3_outputs(5175) <= not (a and b);
    layer3_outputs(5176) <= not b or a;
    layer3_outputs(5177) <= not (a and b);
    layer3_outputs(5178) <= b;
    layer3_outputs(5179) <= 1'b0;
    layer3_outputs(5180) <= 1'b1;
    layer3_outputs(5181) <= b;
    layer3_outputs(5182) <= not a or b;
    layer3_outputs(5183) <= not (a or b);
    layer3_outputs(5184) <= not a;
    layer3_outputs(5185) <= not (a xor b);
    layer3_outputs(5186) <= a or b;
    layer3_outputs(5187) <= 1'b1;
    layer3_outputs(5188) <= a;
    layer3_outputs(5189) <= not a;
    layer3_outputs(5190) <= b and not a;
    layer3_outputs(5191) <= a or b;
    layer3_outputs(5192) <= not b;
    layer3_outputs(5193) <= a and b;
    layer3_outputs(5194) <= not a or b;
    layer3_outputs(5195) <= 1'b0;
    layer3_outputs(5196) <= not a or b;
    layer3_outputs(5197) <= not b or a;
    layer3_outputs(5198) <= not a;
    layer3_outputs(5199) <= a and b;
    layer3_outputs(5200) <= 1'b1;
    layer3_outputs(5201) <= 1'b1;
    layer3_outputs(5202) <= not (a or b);
    layer3_outputs(5203) <= not a;
    layer3_outputs(5204) <= b;
    layer3_outputs(5205) <= b and not a;
    layer3_outputs(5206) <= not (a or b);
    layer3_outputs(5207) <= 1'b0;
    layer3_outputs(5208) <= not (a and b);
    layer3_outputs(5209) <= b;
    layer3_outputs(5210) <= a and b;
    layer3_outputs(5211) <= not (a and b);
    layer3_outputs(5212) <= a and not b;
    layer3_outputs(5213) <= not b;
    layer3_outputs(5214) <= 1'b0;
    layer3_outputs(5215) <= b and not a;
    layer3_outputs(5216) <= a xor b;
    layer3_outputs(5217) <= a and b;
    layer3_outputs(5218) <= a or b;
    layer3_outputs(5219) <= not a or b;
    layer3_outputs(5220) <= 1'b0;
    layer3_outputs(5221) <= b and not a;
    layer3_outputs(5222) <= not b;
    layer3_outputs(5223) <= a or b;
    layer3_outputs(5224) <= b;
    layer3_outputs(5225) <= not b or a;
    layer3_outputs(5226) <= not (a and b);
    layer3_outputs(5227) <= a and not b;
    layer3_outputs(5228) <= b;
    layer3_outputs(5229) <= not (a and b);
    layer3_outputs(5230) <= a or b;
    layer3_outputs(5231) <= 1'b1;
    layer3_outputs(5232) <= a or b;
    layer3_outputs(5233) <= not (a xor b);
    layer3_outputs(5234) <= 1'b1;
    layer3_outputs(5235) <= a and not b;
    layer3_outputs(5236) <= a or b;
    layer3_outputs(5237) <= 1'b1;
    layer3_outputs(5238) <= b and not a;
    layer3_outputs(5239) <= 1'b0;
    layer3_outputs(5240) <= not (a or b);
    layer3_outputs(5241) <= 1'b1;
    layer3_outputs(5242) <= b and not a;
    layer3_outputs(5243) <= not a or b;
    layer3_outputs(5244) <= a and b;
    layer3_outputs(5245) <= 1'b0;
    layer3_outputs(5246) <= a or b;
    layer3_outputs(5247) <= 1'b1;
    layer3_outputs(5248) <= not b;
    layer3_outputs(5249) <= 1'b1;
    layer3_outputs(5250) <= b and not a;
    layer3_outputs(5251) <= b and not a;
    layer3_outputs(5252) <= not a;
    layer3_outputs(5253) <= not a or b;
    layer3_outputs(5254) <= a or b;
    layer3_outputs(5255) <= a and not b;
    layer3_outputs(5256) <= 1'b0;
    layer3_outputs(5257) <= 1'b1;
    layer3_outputs(5258) <= not a or b;
    layer3_outputs(5259) <= not (a or b);
    layer3_outputs(5260) <= not b or a;
    layer3_outputs(5261) <= not (a and b);
    layer3_outputs(5262) <= 1'b0;
    layer3_outputs(5263) <= b and not a;
    layer3_outputs(5264) <= a xor b;
    layer3_outputs(5265) <= not (a and b);
    layer3_outputs(5266) <= not a or b;
    layer3_outputs(5267) <= 1'b1;
    layer3_outputs(5268) <= a and not b;
    layer3_outputs(5269) <= a xor b;
    layer3_outputs(5270) <= 1'b1;
    layer3_outputs(5271) <= not b or a;
    layer3_outputs(5272) <= a xor b;
    layer3_outputs(5273) <= b;
    layer3_outputs(5274) <= 1'b0;
    layer3_outputs(5275) <= 1'b0;
    layer3_outputs(5276) <= a;
    layer3_outputs(5277) <= not (a xor b);
    layer3_outputs(5278) <= not b;
    layer3_outputs(5279) <= not b or a;
    layer3_outputs(5280) <= 1'b1;
    layer3_outputs(5281) <= not a or b;
    layer3_outputs(5282) <= not a or b;
    layer3_outputs(5283) <= a;
    layer3_outputs(5284) <= 1'b1;
    layer3_outputs(5285) <= a and not b;
    layer3_outputs(5286) <= b and not a;
    layer3_outputs(5287) <= a and not b;
    layer3_outputs(5288) <= not a or b;
    layer3_outputs(5289) <= a;
    layer3_outputs(5290) <= not b or a;
    layer3_outputs(5291) <= not a or b;
    layer3_outputs(5292) <= not (a and b);
    layer3_outputs(5293) <= not (a xor b);
    layer3_outputs(5294) <= not (a and b);
    layer3_outputs(5295) <= 1'b0;
    layer3_outputs(5296) <= a and not b;
    layer3_outputs(5297) <= b and not a;
    layer3_outputs(5298) <= a and not b;
    layer3_outputs(5299) <= not (a xor b);
    layer3_outputs(5300) <= a or b;
    layer3_outputs(5301) <= a and b;
    layer3_outputs(5302) <= b and not a;
    layer3_outputs(5303) <= a xor b;
    layer3_outputs(5304) <= not b;
    layer3_outputs(5305) <= 1'b1;
    layer3_outputs(5306) <= b and not a;
    layer3_outputs(5307) <= b;
    layer3_outputs(5308) <= 1'b1;
    layer3_outputs(5309) <= a and b;
    layer3_outputs(5310) <= not (a or b);
    layer3_outputs(5311) <= not b or a;
    layer3_outputs(5312) <= not (a or b);
    layer3_outputs(5313) <= 1'b0;
    layer3_outputs(5314) <= a;
    layer3_outputs(5315) <= a and b;
    layer3_outputs(5316) <= not b or a;
    layer3_outputs(5317) <= not (a or b);
    layer3_outputs(5318) <= a and not b;
    layer3_outputs(5319) <= b and not a;
    layer3_outputs(5320) <= a;
    layer3_outputs(5321) <= not a or b;
    layer3_outputs(5322) <= 1'b1;
    layer3_outputs(5323) <= not (a xor b);
    layer3_outputs(5324) <= a and not b;
    layer3_outputs(5325) <= b;
    layer3_outputs(5326) <= not a;
    layer3_outputs(5327) <= not b;
    layer3_outputs(5328) <= not a;
    layer3_outputs(5329) <= b;
    layer3_outputs(5330) <= not a;
    layer3_outputs(5331) <= not (a and b);
    layer3_outputs(5332) <= not b;
    layer3_outputs(5333) <= not (a and b);
    layer3_outputs(5334) <= 1'b0;
    layer3_outputs(5335) <= a;
    layer3_outputs(5336) <= not (a and b);
    layer3_outputs(5337) <= b;
    layer3_outputs(5338) <= not a;
    layer3_outputs(5339) <= not a;
    layer3_outputs(5340) <= not a or b;
    layer3_outputs(5341) <= not b;
    layer3_outputs(5342) <= 1'b1;
    layer3_outputs(5343) <= 1'b0;
    layer3_outputs(5344) <= a or b;
    layer3_outputs(5345) <= b and not a;
    layer3_outputs(5346) <= a;
    layer3_outputs(5347) <= not b;
    layer3_outputs(5348) <= b;
    layer3_outputs(5349) <= not b;
    layer3_outputs(5350) <= 1'b0;
    layer3_outputs(5351) <= not (a and b);
    layer3_outputs(5352) <= not (a and b);
    layer3_outputs(5353) <= a and not b;
    layer3_outputs(5354) <= not (a and b);
    layer3_outputs(5355) <= a or b;
    layer3_outputs(5356) <= 1'b1;
    layer3_outputs(5357) <= b and not a;
    layer3_outputs(5358) <= not b or a;
    layer3_outputs(5359) <= a;
    layer3_outputs(5360) <= 1'b0;
    layer3_outputs(5361) <= not (a and b);
    layer3_outputs(5362) <= a;
    layer3_outputs(5363) <= a xor b;
    layer3_outputs(5364) <= b and not a;
    layer3_outputs(5365) <= a or b;
    layer3_outputs(5366) <= not (a and b);
    layer3_outputs(5367) <= b and not a;
    layer3_outputs(5368) <= a and b;
    layer3_outputs(5369) <= 1'b1;
    layer3_outputs(5370) <= a and not b;
    layer3_outputs(5371) <= 1'b0;
    layer3_outputs(5372) <= not b;
    layer3_outputs(5373) <= 1'b0;
    layer3_outputs(5374) <= not a or b;
    layer3_outputs(5375) <= not b or a;
    layer3_outputs(5376) <= a or b;
    layer3_outputs(5377) <= 1'b1;
    layer3_outputs(5378) <= 1'b0;
    layer3_outputs(5379) <= not a or b;
    layer3_outputs(5380) <= not (a and b);
    layer3_outputs(5381) <= a or b;
    layer3_outputs(5382) <= not (a and b);
    layer3_outputs(5383) <= not a;
    layer3_outputs(5384) <= not b or a;
    layer3_outputs(5385) <= not a;
    layer3_outputs(5386) <= a;
    layer3_outputs(5387) <= a xor b;
    layer3_outputs(5388) <= 1'b0;
    layer3_outputs(5389) <= not (a and b);
    layer3_outputs(5390) <= b;
    layer3_outputs(5391) <= not (a and b);
    layer3_outputs(5392) <= a;
    layer3_outputs(5393) <= not b or a;
    layer3_outputs(5394) <= a xor b;
    layer3_outputs(5395) <= b;
    layer3_outputs(5396) <= a xor b;
    layer3_outputs(5397) <= not b or a;
    layer3_outputs(5398) <= not b;
    layer3_outputs(5399) <= b and not a;
    layer3_outputs(5400) <= b and not a;
    layer3_outputs(5401) <= not b or a;
    layer3_outputs(5402) <= not (a xor b);
    layer3_outputs(5403) <= a or b;
    layer3_outputs(5404) <= not (a or b);
    layer3_outputs(5405) <= b;
    layer3_outputs(5406) <= not b or a;
    layer3_outputs(5407) <= a and not b;
    layer3_outputs(5408) <= not b;
    layer3_outputs(5409) <= not (a or b);
    layer3_outputs(5410) <= a and b;
    layer3_outputs(5411) <= not b;
    layer3_outputs(5412) <= not (a or b);
    layer3_outputs(5413) <= b;
    layer3_outputs(5414) <= not (a or b);
    layer3_outputs(5415) <= not b;
    layer3_outputs(5416) <= not b or a;
    layer3_outputs(5417) <= b and not a;
    layer3_outputs(5418) <= a or b;
    layer3_outputs(5419) <= b;
    layer3_outputs(5420) <= a and not b;
    layer3_outputs(5421) <= not a;
    layer3_outputs(5422) <= a and b;
    layer3_outputs(5423) <= not (a or b);
    layer3_outputs(5424) <= not b or a;
    layer3_outputs(5425) <= not a or b;
    layer3_outputs(5426) <= 1'b1;
    layer3_outputs(5427) <= not b;
    layer3_outputs(5428) <= not a or b;
    layer3_outputs(5429) <= not a or b;
    layer3_outputs(5430) <= not (a and b);
    layer3_outputs(5431) <= 1'b0;
    layer3_outputs(5432) <= 1'b0;
    layer3_outputs(5433) <= 1'b1;
    layer3_outputs(5434) <= not (a or b);
    layer3_outputs(5435) <= not b;
    layer3_outputs(5436) <= a xor b;
    layer3_outputs(5437) <= not a or b;
    layer3_outputs(5438) <= not a;
    layer3_outputs(5439) <= 1'b0;
    layer3_outputs(5440) <= not (a or b);
    layer3_outputs(5441) <= not b;
    layer3_outputs(5442) <= not a;
    layer3_outputs(5443) <= not b or a;
    layer3_outputs(5444) <= not b;
    layer3_outputs(5445) <= not (a xor b);
    layer3_outputs(5446) <= not a;
    layer3_outputs(5447) <= 1'b0;
    layer3_outputs(5448) <= a;
    layer3_outputs(5449) <= a or b;
    layer3_outputs(5450) <= not (a and b);
    layer3_outputs(5451) <= a and b;
    layer3_outputs(5452) <= a and not b;
    layer3_outputs(5453) <= a xor b;
    layer3_outputs(5454) <= a and not b;
    layer3_outputs(5455) <= a and b;
    layer3_outputs(5456) <= a;
    layer3_outputs(5457) <= not (a xor b);
    layer3_outputs(5458) <= b and not a;
    layer3_outputs(5459) <= b and not a;
    layer3_outputs(5460) <= not a;
    layer3_outputs(5461) <= a and not b;
    layer3_outputs(5462) <= not (a or b);
    layer3_outputs(5463) <= a and not b;
    layer3_outputs(5464) <= not b;
    layer3_outputs(5465) <= a and b;
    layer3_outputs(5466) <= b;
    layer3_outputs(5467) <= not a or b;
    layer3_outputs(5468) <= a or b;
    layer3_outputs(5469) <= a or b;
    layer3_outputs(5470) <= not b;
    layer3_outputs(5471) <= not b or a;
    layer3_outputs(5472) <= not (a or b);
    layer3_outputs(5473) <= 1'b1;
    layer3_outputs(5474) <= 1'b0;
    layer3_outputs(5475) <= not b;
    layer3_outputs(5476) <= not a;
    layer3_outputs(5477) <= 1'b1;
    layer3_outputs(5478) <= not b or a;
    layer3_outputs(5479) <= not a;
    layer3_outputs(5480) <= b and not a;
    layer3_outputs(5481) <= a;
    layer3_outputs(5482) <= a and not b;
    layer3_outputs(5483) <= a and b;
    layer3_outputs(5484) <= a;
    layer3_outputs(5485) <= 1'b1;
    layer3_outputs(5486) <= a or b;
    layer3_outputs(5487) <= 1'b0;
    layer3_outputs(5488) <= 1'b1;
    layer3_outputs(5489) <= not (a xor b);
    layer3_outputs(5490) <= not (a or b);
    layer3_outputs(5491) <= a;
    layer3_outputs(5492) <= not (a and b);
    layer3_outputs(5493) <= a xor b;
    layer3_outputs(5494) <= not (a and b);
    layer3_outputs(5495) <= b;
    layer3_outputs(5496) <= a and b;
    layer3_outputs(5497) <= b and not a;
    layer3_outputs(5498) <= a and b;
    layer3_outputs(5499) <= not a;
    layer3_outputs(5500) <= not b;
    layer3_outputs(5501) <= a xor b;
    layer3_outputs(5502) <= a or b;
    layer3_outputs(5503) <= not b or a;
    layer3_outputs(5504) <= a xor b;
    layer3_outputs(5505) <= not a;
    layer3_outputs(5506) <= not (a or b);
    layer3_outputs(5507) <= b and not a;
    layer3_outputs(5508) <= 1'b1;
    layer3_outputs(5509) <= a and not b;
    layer3_outputs(5510) <= not b or a;
    layer3_outputs(5511) <= 1'b0;
    layer3_outputs(5512) <= b and not a;
    layer3_outputs(5513) <= not a;
    layer3_outputs(5514) <= 1'b1;
    layer3_outputs(5515) <= b;
    layer3_outputs(5516) <= b and not a;
    layer3_outputs(5517) <= not (a xor b);
    layer3_outputs(5518) <= a and b;
    layer3_outputs(5519) <= 1'b0;
    layer3_outputs(5520) <= b and not a;
    layer3_outputs(5521) <= not a or b;
    layer3_outputs(5522) <= not a or b;
    layer3_outputs(5523) <= b and not a;
    layer3_outputs(5524) <= a or b;
    layer3_outputs(5525) <= 1'b1;
    layer3_outputs(5526) <= not a;
    layer3_outputs(5527) <= a or b;
    layer3_outputs(5528) <= not b;
    layer3_outputs(5529) <= not a or b;
    layer3_outputs(5530) <= b and not a;
    layer3_outputs(5531) <= not a or b;
    layer3_outputs(5532) <= a or b;
    layer3_outputs(5533) <= not b;
    layer3_outputs(5534) <= b and not a;
    layer3_outputs(5535) <= 1'b1;
    layer3_outputs(5536) <= not b;
    layer3_outputs(5537) <= not a;
    layer3_outputs(5538) <= b;
    layer3_outputs(5539) <= b;
    layer3_outputs(5540) <= b and not a;
    layer3_outputs(5541) <= 1'b0;
    layer3_outputs(5542) <= a xor b;
    layer3_outputs(5543) <= not (a and b);
    layer3_outputs(5544) <= not (a or b);
    layer3_outputs(5545) <= a and b;
    layer3_outputs(5546) <= a;
    layer3_outputs(5547) <= not (a and b);
    layer3_outputs(5548) <= not (a and b);
    layer3_outputs(5549) <= b and not a;
    layer3_outputs(5550) <= not b;
    layer3_outputs(5551) <= not (a or b);
    layer3_outputs(5552) <= not b;
    layer3_outputs(5553) <= 1'b0;
    layer3_outputs(5554) <= 1'b1;
    layer3_outputs(5555) <= not (a or b);
    layer3_outputs(5556) <= 1'b0;
    layer3_outputs(5557) <= not b;
    layer3_outputs(5558) <= not (a and b);
    layer3_outputs(5559) <= a or b;
    layer3_outputs(5560) <= a;
    layer3_outputs(5561) <= not (a or b);
    layer3_outputs(5562) <= not b or a;
    layer3_outputs(5563) <= a or b;
    layer3_outputs(5564) <= not a;
    layer3_outputs(5565) <= not (a xor b);
    layer3_outputs(5566) <= a or b;
    layer3_outputs(5567) <= b and not a;
    layer3_outputs(5568) <= not (a or b);
    layer3_outputs(5569) <= b;
    layer3_outputs(5570) <= not b;
    layer3_outputs(5571) <= a or b;
    layer3_outputs(5572) <= a;
    layer3_outputs(5573) <= not a or b;
    layer3_outputs(5574) <= a or b;
    layer3_outputs(5575) <= a;
    layer3_outputs(5576) <= a and not b;
    layer3_outputs(5577) <= not b or a;
    layer3_outputs(5578) <= b and not a;
    layer3_outputs(5579) <= not a;
    layer3_outputs(5580) <= a or b;
    layer3_outputs(5581) <= not a;
    layer3_outputs(5582) <= b and not a;
    layer3_outputs(5583) <= not b or a;
    layer3_outputs(5584) <= not b or a;
    layer3_outputs(5585) <= not (a and b);
    layer3_outputs(5586) <= not (a and b);
    layer3_outputs(5587) <= 1'b0;
    layer3_outputs(5588) <= b;
    layer3_outputs(5589) <= not b;
    layer3_outputs(5590) <= 1'b1;
    layer3_outputs(5591) <= not a;
    layer3_outputs(5592) <= not (a or b);
    layer3_outputs(5593) <= a;
    layer3_outputs(5594) <= a and not b;
    layer3_outputs(5595) <= not (a and b);
    layer3_outputs(5596) <= 1'b1;
    layer3_outputs(5597) <= not b;
    layer3_outputs(5598) <= not (a or b);
    layer3_outputs(5599) <= 1'b1;
    layer3_outputs(5600) <= a;
    layer3_outputs(5601) <= a and not b;
    layer3_outputs(5602) <= 1'b0;
    layer3_outputs(5603) <= 1'b0;
    layer3_outputs(5604) <= not b or a;
    layer3_outputs(5605) <= not a;
    layer3_outputs(5606) <= a;
    layer3_outputs(5607) <= not b or a;
    layer3_outputs(5608) <= not b or a;
    layer3_outputs(5609) <= b and not a;
    layer3_outputs(5610) <= a and b;
    layer3_outputs(5611) <= b and not a;
    layer3_outputs(5612) <= not a or b;
    layer3_outputs(5613) <= not a;
    layer3_outputs(5614) <= not (a or b);
    layer3_outputs(5615) <= not (a or b);
    layer3_outputs(5616) <= not a or b;
    layer3_outputs(5617) <= b and not a;
    layer3_outputs(5618) <= not (a and b);
    layer3_outputs(5619) <= a and b;
    layer3_outputs(5620) <= not (a and b);
    layer3_outputs(5621) <= not a;
    layer3_outputs(5622) <= a and b;
    layer3_outputs(5623) <= not a;
    layer3_outputs(5624) <= not a or b;
    layer3_outputs(5625) <= not (a and b);
    layer3_outputs(5626) <= a;
    layer3_outputs(5627) <= a and not b;
    layer3_outputs(5628) <= a and b;
    layer3_outputs(5629) <= a and b;
    layer3_outputs(5630) <= b and not a;
    layer3_outputs(5631) <= not b or a;
    layer3_outputs(5632) <= 1'b0;
    layer3_outputs(5633) <= not a;
    layer3_outputs(5634) <= not (a or b);
    layer3_outputs(5635) <= b and not a;
    layer3_outputs(5636) <= 1'b1;
    layer3_outputs(5637) <= a;
    layer3_outputs(5638) <= not b;
    layer3_outputs(5639) <= a and b;
    layer3_outputs(5640) <= not a or b;
    layer3_outputs(5641) <= not b or a;
    layer3_outputs(5642) <= a or b;
    layer3_outputs(5643) <= not b;
    layer3_outputs(5644) <= a xor b;
    layer3_outputs(5645) <= not (a or b);
    layer3_outputs(5646) <= not a or b;
    layer3_outputs(5647) <= a and not b;
    layer3_outputs(5648) <= not b;
    layer3_outputs(5649) <= not a or b;
    layer3_outputs(5650) <= a and b;
    layer3_outputs(5651) <= not a;
    layer3_outputs(5652) <= not (a and b);
    layer3_outputs(5653) <= not b;
    layer3_outputs(5654) <= 1'b0;
    layer3_outputs(5655) <= not b or a;
    layer3_outputs(5656) <= b;
    layer3_outputs(5657) <= a and not b;
    layer3_outputs(5658) <= 1'b1;
    layer3_outputs(5659) <= not b or a;
    layer3_outputs(5660) <= a xor b;
    layer3_outputs(5661) <= not (a or b);
    layer3_outputs(5662) <= not a or b;
    layer3_outputs(5663) <= a and not b;
    layer3_outputs(5664) <= a and b;
    layer3_outputs(5665) <= not b;
    layer3_outputs(5666) <= b and not a;
    layer3_outputs(5667) <= not b;
    layer3_outputs(5668) <= not (a and b);
    layer3_outputs(5669) <= not b;
    layer3_outputs(5670) <= a and b;
    layer3_outputs(5671) <= a;
    layer3_outputs(5672) <= not (a or b);
    layer3_outputs(5673) <= not a or b;
    layer3_outputs(5674) <= not a or b;
    layer3_outputs(5675) <= 1'b1;
    layer3_outputs(5676) <= not (a and b);
    layer3_outputs(5677) <= not (a or b);
    layer3_outputs(5678) <= not (a or b);
    layer3_outputs(5679) <= not (a or b);
    layer3_outputs(5680) <= b and not a;
    layer3_outputs(5681) <= not a;
    layer3_outputs(5682) <= 1'b0;
    layer3_outputs(5683) <= a or b;
    layer3_outputs(5684) <= a and b;
    layer3_outputs(5685) <= not a;
    layer3_outputs(5686) <= not (a xor b);
    layer3_outputs(5687) <= b;
    layer3_outputs(5688) <= a;
    layer3_outputs(5689) <= b;
    layer3_outputs(5690) <= not b or a;
    layer3_outputs(5691) <= not (a and b);
    layer3_outputs(5692) <= a xor b;
    layer3_outputs(5693) <= not (a or b);
    layer3_outputs(5694) <= not (a or b);
    layer3_outputs(5695) <= a;
    layer3_outputs(5696) <= not b;
    layer3_outputs(5697) <= a or b;
    layer3_outputs(5698) <= not b;
    layer3_outputs(5699) <= a and b;
    layer3_outputs(5700) <= a xor b;
    layer3_outputs(5701) <= not b or a;
    layer3_outputs(5702) <= 1'b1;
    layer3_outputs(5703) <= not b;
    layer3_outputs(5704) <= not b or a;
    layer3_outputs(5705) <= a and not b;
    layer3_outputs(5706) <= not a;
    layer3_outputs(5707) <= not a;
    layer3_outputs(5708) <= not a or b;
    layer3_outputs(5709) <= not a;
    layer3_outputs(5710) <= not (a xor b);
    layer3_outputs(5711) <= 1'b0;
    layer3_outputs(5712) <= 1'b1;
    layer3_outputs(5713) <= a and b;
    layer3_outputs(5714) <= not a or b;
    layer3_outputs(5715) <= not (a and b);
    layer3_outputs(5716) <= not b or a;
    layer3_outputs(5717) <= 1'b1;
    layer3_outputs(5718) <= a and not b;
    layer3_outputs(5719) <= b;
    layer3_outputs(5720) <= a;
    layer3_outputs(5721) <= not b;
    layer3_outputs(5722) <= a or b;
    layer3_outputs(5723) <= 1'b0;
    layer3_outputs(5724) <= a or b;
    layer3_outputs(5725) <= not a or b;
    layer3_outputs(5726) <= a;
    layer3_outputs(5727) <= a and b;
    layer3_outputs(5728) <= not a or b;
    layer3_outputs(5729) <= b;
    layer3_outputs(5730) <= a and b;
    layer3_outputs(5731) <= b and not a;
    layer3_outputs(5732) <= not a;
    layer3_outputs(5733) <= not a or b;
    layer3_outputs(5734) <= a and b;
    layer3_outputs(5735) <= not b or a;
    layer3_outputs(5736) <= a and b;
    layer3_outputs(5737) <= a or b;
    layer3_outputs(5738) <= 1'b1;
    layer3_outputs(5739) <= a;
    layer3_outputs(5740) <= b and not a;
    layer3_outputs(5741) <= a and not b;
    layer3_outputs(5742) <= not b or a;
    layer3_outputs(5743) <= 1'b0;
    layer3_outputs(5744) <= a or b;
    layer3_outputs(5745) <= not (a or b);
    layer3_outputs(5746) <= not (a or b);
    layer3_outputs(5747) <= 1'b1;
    layer3_outputs(5748) <= a;
    layer3_outputs(5749) <= not b or a;
    layer3_outputs(5750) <= not b or a;
    layer3_outputs(5751) <= not b;
    layer3_outputs(5752) <= not b or a;
    layer3_outputs(5753) <= not a or b;
    layer3_outputs(5754) <= a;
    layer3_outputs(5755) <= 1'b0;
    layer3_outputs(5756) <= not (a or b);
    layer3_outputs(5757) <= a and not b;
    layer3_outputs(5758) <= a or b;
    layer3_outputs(5759) <= not a or b;
    layer3_outputs(5760) <= 1'b1;
    layer3_outputs(5761) <= not a or b;
    layer3_outputs(5762) <= 1'b1;
    layer3_outputs(5763) <= not a;
    layer3_outputs(5764) <= not a or b;
    layer3_outputs(5765) <= not b;
    layer3_outputs(5766) <= not b;
    layer3_outputs(5767) <= a and b;
    layer3_outputs(5768) <= not b or a;
    layer3_outputs(5769) <= not a;
    layer3_outputs(5770) <= not (a or b);
    layer3_outputs(5771) <= b and not a;
    layer3_outputs(5772) <= not b;
    layer3_outputs(5773) <= 1'b0;
    layer3_outputs(5774) <= not a or b;
    layer3_outputs(5775) <= b and not a;
    layer3_outputs(5776) <= a or b;
    layer3_outputs(5777) <= not b or a;
    layer3_outputs(5778) <= b and not a;
    layer3_outputs(5779) <= b and not a;
    layer3_outputs(5780) <= 1'b1;
    layer3_outputs(5781) <= not (a xor b);
    layer3_outputs(5782) <= not (a xor b);
    layer3_outputs(5783) <= a and not b;
    layer3_outputs(5784) <= not a;
    layer3_outputs(5785) <= not (a and b);
    layer3_outputs(5786) <= a and not b;
    layer3_outputs(5787) <= 1'b1;
    layer3_outputs(5788) <= a and b;
    layer3_outputs(5789) <= not (a or b);
    layer3_outputs(5790) <= 1'b0;
    layer3_outputs(5791) <= a and b;
    layer3_outputs(5792) <= a or b;
    layer3_outputs(5793) <= a and b;
    layer3_outputs(5794) <= not b;
    layer3_outputs(5795) <= b;
    layer3_outputs(5796) <= a;
    layer3_outputs(5797) <= a and not b;
    layer3_outputs(5798) <= not a;
    layer3_outputs(5799) <= a and b;
    layer3_outputs(5800) <= b;
    layer3_outputs(5801) <= a;
    layer3_outputs(5802) <= b;
    layer3_outputs(5803) <= not a or b;
    layer3_outputs(5804) <= not (a or b);
    layer3_outputs(5805) <= b and not a;
    layer3_outputs(5806) <= b and not a;
    layer3_outputs(5807) <= 1'b0;
    layer3_outputs(5808) <= not (a xor b);
    layer3_outputs(5809) <= a;
    layer3_outputs(5810) <= b;
    layer3_outputs(5811) <= b and not a;
    layer3_outputs(5812) <= not b;
    layer3_outputs(5813) <= not b or a;
    layer3_outputs(5814) <= not (a xor b);
    layer3_outputs(5815) <= not a or b;
    layer3_outputs(5816) <= not b or a;
    layer3_outputs(5817) <= a and b;
    layer3_outputs(5818) <= a and b;
    layer3_outputs(5819) <= a or b;
    layer3_outputs(5820) <= 1'b0;
    layer3_outputs(5821) <= a or b;
    layer3_outputs(5822) <= not a;
    layer3_outputs(5823) <= b and not a;
    layer3_outputs(5824) <= a;
    layer3_outputs(5825) <= b;
    layer3_outputs(5826) <= b and not a;
    layer3_outputs(5827) <= a or b;
    layer3_outputs(5828) <= a;
    layer3_outputs(5829) <= b and not a;
    layer3_outputs(5830) <= a;
    layer3_outputs(5831) <= a and b;
    layer3_outputs(5832) <= b;
    layer3_outputs(5833) <= b and not a;
    layer3_outputs(5834) <= not b;
    layer3_outputs(5835) <= a;
    layer3_outputs(5836) <= a;
    layer3_outputs(5837) <= not b;
    layer3_outputs(5838) <= a;
    layer3_outputs(5839) <= a or b;
    layer3_outputs(5840) <= b;
    layer3_outputs(5841) <= a or b;
    layer3_outputs(5842) <= not (a or b);
    layer3_outputs(5843) <= b and not a;
    layer3_outputs(5844) <= a and b;
    layer3_outputs(5845) <= b;
    layer3_outputs(5846) <= not a;
    layer3_outputs(5847) <= not (a xor b);
    layer3_outputs(5848) <= b and not a;
    layer3_outputs(5849) <= a xor b;
    layer3_outputs(5850) <= not (a or b);
    layer3_outputs(5851) <= not (a or b);
    layer3_outputs(5852) <= not a or b;
    layer3_outputs(5853) <= a;
    layer3_outputs(5854) <= 1'b1;
    layer3_outputs(5855) <= 1'b0;
    layer3_outputs(5856) <= a;
    layer3_outputs(5857) <= not b;
    layer3_outputs(5858) <= not a;
    layer3_outputs(5859) <= b;
    layer3_outputs(5860) <= b and not a;
    layer3_outputs(5861) <= b;
    layer3_outputs(5862) <= not (a or b);
    layer3_outputs(5863) <= not a or b;
    layer3_outputs(5864) <= a and b;
    layer3_outputs(5865) <= a or b;
    layer3_outputs(5866) <= a and not b;
    layer3_outputs(5867) <= b and not a;
    layer3_outputs(5868) <= b;
    layer3_outputs(5869) <= a or b;
    layer3_outputs(5870) <= a and not b;
    layer3_outputs(5871) <= a;
    layer3_outputs(5872) <= not a or b;
    layer3_outputs(5873) <= a and not b;
    layer3_outputs(5874) <= not a or b;
    layer3_outputs(5875) <= a or b;
    layer3_outputs(5876) <= a or b;
    layer3_outputs(5877) <= not (a xor b);
    layer3_outputs(5878) <= a or b;
    layer3_outputs(5879) <= not b or a;
    layer3_outputs(5880) <= a and b;
    layer3_outputs(5881) <= not b or a;
    layer3_outputs(5882) <= not (a and b);
    layer3_outputs(5883) <= not b or a;
    layer3_outputs(5884) <= a and b;
    layer3_outputs(5885) <= b and not a;
    layer3_outputs(5886) <= a or b;
    layer3_outputs(5887) <= b and not a;
    layer3_outputs(5888) <= a;
    layer3_outputs(5889) <= not b or a;
    layer3_outputs(5890) <= not a or b;
    layer3_outputs(5891) <= not (a xor b);
    layer3_outputs(5892) <= a and b;
    layer3_outputs(5893) <= not a;
    layer3_outputs(5894) <= not (a and b);
    layer3_outputs(5895) <= b;
    layer3_outputs(5896) <= not a or b;
    layer3_outputs(5897) <= 1'b1;
    layer3_outputs(5898) <= not a or b;
    layer3_outputs(5899) <= a and not b;
    layer3_outputs(5900) <= a xor b;
    layer3_outputs(5901) <= 1'b1;
    layer3_outputs(5902) <= 1'b0;
    layer3_outputs(5903) <= not a or b;
    layer3_outputs(5904) <= 1'b1;
    layer3_outputs(5905) <= not a or b;
    layer3_outputs(5906) <= a or b;
    layer3_outputs(5907) <= not a;
    layer3_outputs(5908) <= a or b;
    layer3_outputs(5909) <= 1'b0;
    layer3_outputs(5910) <= not a;
    layer3_outputs(5911) <= not (a or b);
    layer3_outputs(5912) <= 1'b1;
    layer3_outputs(5913) <= not a or b;
    layer3_outputs(5914) <= not b;
    layer3_outputs(5915) <= not (a or b);
    layer3_outputs(5916) <= 1'b1;
    layer3_outputs(5917) <= b;
    layer3_outputs(5918) <= b;
    layer3_outputs(5919) <= not a;
    layer3_outputs(5920) <= b;
    layer3_outputs(5921) <= a xor b;
    layer3_outputs(5922) <= not (a or b);
    layer3_outputs(5923) <= b;
    layer3_outputs(5924) <= a or b;
    layer3_outputs(5925) <= b and not a;
    layer3_outputs(5926) <= not (a or b);
    layer3_outputs(5927) <= a and not b;
    layer3_outputs(5928) <= a;
    layer3_outputs(5929) <= a;
    layer3_outputs(5930) <= not (a and b);
    layer3_outputs(5931) <= not a;
    layer3_outputs(5932) <= not a;
    layer3_outputs(5933) <= not a or b;
    layer3_outputs(5934) <= not (a or b);
    layer3_outputs(5935) <= 1'b1;
    layer3_outputs(5936) <= not a;
    layer3_outputs(5937) <= b;
    layer3_outputs(5938) <= a or b;
    layer3_outputs(5939) <= not b or a;
    layer3_outputs(5940) <= a and b;
    layer3_outputs(5941) <= a or b;
    layer3_outputs(5942) <= 1'b0;
    layer3_outputs(5943) <= not (a and b);
    layer3_outputs(5944) <= not a;
    layer3_outputs(5945) <= not a or b;
    layer3_outputs(5946) <= a or b;
    layer3_outputs(5947) <= not (a and b);
    layer3_outputs(5948) <= not a;
    layer3_outputs(5949) <= a;
    layer3_outputs(5950) <= not (a and b);
    layer3_outputs(5951) <= a and b;
    layer3_outputs(5952) <= not a or b;
    layer3_outputs(5953) <= b;
    layer3_outputs(5954) <= a and b;
    layer3_outputs(5955) <= not a or b;
    layer3_outputs(5956) <= 1'b1;
    layer3_outputs(5957) <= 1'b1;
    layer3_outputs(5958) <= b;
    layer3_outputs(5959) <= 1'b0;
    layer3_outputs(5960) <= b and not a;
    layer3_outputs(5961) <= not a or b;
    layer3_outputs(5962) <= a and b;
    layer3_outputs(5963) <= not b or a;
    layer3_outputs(5964) <= a;
    layer3_outputs(5965) <= not a or b;
    layer3_outputs(5966) <= not a;
    layer3_outputs(5967) <= 1'b1;
    layer3_outputs(5968) <= a;
    layer3_outputs(5969) <= not (a or b);
    layer3_outputs(5970) <= not (a or b);
    layer3_outputs(5971) <= 1'b0;
    layer3_outputs(5972) <= not a;
    layer3_outputs(5973) <= not (a and b);
    layer3_outputs(5974) <= a or b;
    layer3_outputs(5975) <= not (a xor b);
    layer3_outputs(5976) <= not b or a;
    layer3_outputs(5977) <= not b or a;
    layer3_outputs(5978) <= not (a or b);
    layer3_outputs(5979) <= a;
    layer3_outputs(5980) <= not (a and b);
    layer3_outputs(5981) <= b;
    layer3_outputs(5982) <= not b or a;
    layer3_outputs(5983) <= not b;
    layer3_outputs(5984) <= b and not a;
    layer3_outputs(5985) <= a and b;
    layer3_outputs(5986) <= not a or b;
    layer3_outputs(5987) <= a and not b;
    layer3_outputs(5988) <= not (a or b);
    layer3_outputs(5989) <= a xor b;
    layer3_outputs(5990) <= b and not a;
    layer3_outputs(5991) <= b and not a;
    layer3_outputs(5992) <= a and b;
    layer3_outputs(5993) <= 1'b1;
    layer3_outputs(5994) <= not (a and b);
    layer3_outputs(5995) <= not a;
    layer3_outputs(5996) <= not a or b;
    layer3_outputs(5997) <= not (a and b);
    layer3_outputs(5998) <= not (a and b);
    layer3_outputs(5999) <= b and not a;
    layer3_outputs(6000) <= not (a xor b);
    layer3_outputs(6001) <= not (a or b);
    layer3_outputs(6002) <= not a;
    layer3_outputs(6003) <= not b or a;
    layer3_outputs(6004) <= not b;
    layer3_outputs(6005) <= 1'b0;
    layer3_outputs(6006) <= not (a and b);
    layer3_outputs(6007) <= a;
    layer3_outputs(6008) <= not a;
    layer3_outputs(6009) <= b and not a;
    layer3_outputs(6010) <= b and not a;
    layer3_outputs(6011) <= 1'b1;
    layer3_outputs(6012) <= not a or b;
    layer3_outputs(6013) <= a or b;
    layer3_outputs(6014) <= not b;
    layer3_outputs(6015) <= a and not b;
    layer3_outputs(6016) <= not (a or b);
    layer3_outputs(6017) <= not b or a;
    layer3_outputs(6018) <= a xor b;
    layer3_outputs(6019) <= not (a and b);
    layer3_outputs(6020) <= not b;
    layer3_outputs(6021) <= not b or a;
    layer3_outputs(6022) <= b and not a;
    layer3_outputs(6023) <= b and not a;
    layer3_outputs(6024) <= a and b;
    layer3_outputs(6025) <= not b or a;
    layer3_outputs(6026) <= b and not a;
    layer3_outputs(6027) <= a and b;
    layer3_outputs(6028) <= b;
    layer3_outputs(6029) <= b;
    layer3_outputs(6030) <= a or b;
    layer3_outputs(6031) <= b and not a;
    layer3_outputs(6032) <= a;
    layer3_outputs(6033) <= a;
    layer3_outputs(6034) <= a and not b;
    layer3_outputs(6035) <= not b or a;
    layer3_outputs(6036) <= not (a and b);
    layer3_outputs(6037) <= a and not b;
    layer3_outputs(6038) <= a or b;
    layer3_outputs(6039) <= not a or b;
    layer3_outputs(6040) <= a and not b;
    layer3_outputs(6041) <= b;
    layer3_outputs(6042) <= not b;
    layer3_outputs(6043) <= a xor b;
    layer3_outputs(6044) <= 1'b0;
    layer3_outputs(6045) <= not (a or b);
    layer3_outputs(6046) <= not b;
    layer3_outputs(6047) <= a and b;
    layer3_outputs(6048) <= a and b;
    layer3_outputs(6049) <= b and not a;
    layer3_outputs(6050) <= not b or a;
    layer3_outputs(6051) <= a and b;
    layer3_outputs(6052) <= b;
    layer3_outputs(6053) <= 1'b1;
    layer3_outputs(6054) <= b and not a;
    layer3_outputs(6055) <= not b or a;
    layer3_outputs(6056) <= not b;
    layer3_outputs(6057) <= not (a and b);
    layer3_outputs(6058) <= a;
    layer3_outputs(6059) <= not a;
    layer3_outputs(6060) <= not (a or b);
    layer3_outputs(6061) <= not a;
    layer3_outputs(6062) <= 1'b1;
    layer3_outputs(6063) <= a or b;
    layer3_outputs(6064) <= not (a or b);
    layer3_outputs(6065) <= not a;
    layer3_outputs(6066) <= b and not a;
    layer3_outputs(6067) <= not a or b;
    layer3_outputs(6068) <= a or b;
    layer3_outputs(6069) <= a and b;
    layer3_outputs(6070) <= not a;
    layer3_outputs(6071) <= a or b;
    layer3_outputs(6072) <= not b or a;
    layer3_outputs(6073) <= b;
    layer3_outputs(6074) <= not b or a;
    layer3_outputs(6075) <= a or b;
    layer3_outputs(6076) <= a and not b;
    layer3_outputs(6077) <= a or b;
    layer3_outputs(6078) <= not (a or b);
    layer3_outputs(6079) <= not b;
    layer3_outputs(6080) <= not a;
    layer3_outputs(6081) <= a;
    layer3_outputs(6082) <= a and b;
    layer3_outputs(6083) <= not a or b;
    layer3_outputs(6084) <= b and not a;
    layer3_outputs(6085) <= b;
    layer3_outputs(6086) <= 1'b0;
    layer3_outputs(6087) <= not a;
    layer3_outputs(6088) <= a and not b;
    layer3_outputs(6089) <= not a or b;
    layer3_outputs(6090) <= 1'b0;
    layer3_outputs(6091) <= 1'b0;
    layer3_outputs(6092) <= a and b;
    layer3_outputs(6093) <= 1'b0;
    layer3_outputs(6094) <= 1'b0;
    layer3_outputs(6095) <= a;
    layer3_outputs(6096) <= a;
    layer3_outputs(6097) <= not a;
    layer3_outputs(6098) <= a or b;
    layer3_outputs(6099) <= not a;
    layer3_outputs(6100) <= b;
    layer3_outputs(6101) <= b and not a;
    layer3_outputs(6102) <= not b or a;
    layer3_outputs(6103) <= a and b;
    layer3_outputs(6104) <= not (a and b);
    layer3_outputs(6105) <= a;
    layer3_outputs(6106) <= not b;
    layer3_outputs(6107) <= not b or a;
    layer3_outputs(6108) <= not b or a;
    layer3_outputs(6109) <= b;
    layer3_outputs(6110) <= b;
    layer3_outputs(6111) <= 1'b0;
    layer3_outputs(6112) <= 1'b1;
    layer3_outputs(6113) <= not (a and b);
    layer3_outputs(6114) <= not a or b;
    layer3_outputs(6115) <= 1'b1;
    layer3_outputs(6116) <= a and b;
    layer3_outputs(6117) <= 1'b1;
    layer3_outputs(6118) <= b;
    layer3_outputs(6119) <= b and not a;
    layer3_outputs(6120) <= b;
    layer3_outputs(6121) <= 1'b1;
    layer3_outputs(6122) <= not (a xor b);
    layer3_outputs(6123) <= a and not b;
    layer3_outputs(6124) <= a or b;
    layer3_outputs(6125) <= b and not a;
    layer3_outputs(6126) <= b and not a;
    layer3_outputs(6127) <= a and not b;
    layer3_outputs(6128) <= a or b;
    layer3_outputs(6129) <= a or b;
    layer3_outputs(6130) <= not (a and b);
    layer3_outputs(6131) <= a and not b;
    layer3_outputs(6132) <= not b or a;
    layer3_outputs(6133) <= a;
    layer3_outputs(6134) <= a and not b;
    layer3_outputs(6135) <= b;
    layer3_outputs(6136) <= not b;
    layer3_outputs(6137) <= a and not b;
    layer3_outputs(6138) <= a or b;
    layer3_outputs(6139) <= not (a and b);
    layer3_outputs(6140) <= a and b;
    layer3_outputs(6141) <= 1'b0;
    layer3_outputs(6142) <= 1'b1;
    layer3_outputs(6143) <= not a or b;
    layer3_outputs(6144) <= a;
    layer3_outputs(6145) <= not a;
    layer3_outputs(6146) <= a and b;
    layer3_outputs(6147) <= a or b;
    layer3_outputs(6148) <= 1'b0;
    layer3_outputs(6149) <= a and b;
    layer3_outputs(6150) <= 1'b1;
    layer3_outputs(6151) <= not b;
    layer3_outputs(6152) <= a and not b;
    layer3_outputs(6153) <= b;
    layer3_outputs(6154) <= 1'b1;
    layer3_outputs(6155) <= a or b;
    layer3_outputs(6156) <= a and not b;
    layer3_outputs(6157) <= 1'b0;
    layer3_outputs(6158) <= a and not b;
    layer3_outputs(6159) <= not a or b;
    layer3_outputs(6160) <= 1'b0;
    layer3_outputs(6161) <= 1'b1;
    layer3_outputs(6162) <= not b or a;
    layer3_outputs(6163) <= a and not b;
    layer3_outputs(6164) <= not b or a;
    layer3_outputs(6165) <= not (a and b);
    layer3_outputs(6166) <= 1'b1;
    layer3_outputs(6167) <= not b;
    layer3_outputs(6168) <= not a or b;
    layer3_outputs(6169) <= 1'b0;
    layer3_outputs(6170) <= not a or b;
    layer3_outputs(6171) <= b and not a;
    layer3_outputs(6172) <= 1'b1;
    layer3_outputs(6173) <= a and b;
    layer3_outputs(6174) <= a or b;
    layer3_outputs(6175) <= not a or b;
    layer3_outputs(6176) <= b;
    layer3_outputs(6177) <= not b;
    layer3_outputs(6178) <= a and not b;
    layer3_outputs(6179) <= a or b;
    layer3_outputs(6180) <= a and not b;
    layer3_outputs(6181) <= not b;
    layer3_outputs(6182) <= a and not b;
    layer3_outputs(6183) <= 1'b1;
    layer3_outputs(6184) <= a and b;
    layer3_outputs(6185) <= a and not b;
    layer3_outputs(6186) <= not (a or b);
    layer3_outputs(6187) <= 1'b1;
    layer3_outputs(6188) <= not (a and b);
    layer3_outputs(6189) <= not (a or b);
    layer3_outputs(6190) <= 1'b1;
    layer3_outputs(6191) <= not (a or b);
    layer3_outputs(6192) <= not b or a;
    layer3_outputs(6193) <= not a;
    layer3_outputs(6194) <= a;
    layer3_outputs(6195) <= not a;
    layer3_outputs(6196) <= 1'b1;
    layer3_outputs(6197) <= not a or b;
    layer3_outputs(6198) <= not b;
    layer3_outputs(6199) <= 1'b0;
    layer3_outputs(6200) <= b;
    layer3_outputs(6201) <= a;
    layer3_outputs(6202) <= 1'b1;
    layer3_outputs(6203) <= a;
    layer3_outputs(6204) <= not b;
    layer3_outputs(6205) <= a and not b;
    layer3_outputs(6206) <= not a or b;
    layer3_outputs(6207) <= b and not a;
    layer3_outputs(6208) <= a;
    layer3_outputs(6209) <= 1'b1;
    layer3_outputs(6210) <= a;
    layer3_outputs(6211) <= not b;
    layer3_outputs(6212) <= not b;
    layer3_outputs(6213) <= a or b;
    layer3_outputs(6214) <= a and not b;
    layer3_outputs(6215) <= 1'b0;
    layer3_outputs(6216) <= 1'b0;
    layer3_outputs(6217) <= a or b;
    layer3_outputs(6218) <= b and not a;
    layer3_outputs(6219) <= a and not b;
    layer3_outputs(6220) <= not a or b;
    layer3_outputs(6221) <= 1'b1;
    layer3_outputs(6222) <= not b;
    layer3_outputs(6223) <= not a or b;
    layer3_outputs(6224) <= not b;
    layer3_outputs(6225) <= not a or b;
    layer3_outputs(6226) <= not a or b;
    layer3_outputs(6227) <= b;
    layer3_outputs(6228) <= a or b;
    layer3_outputs(6229) <= not a;
    layer3_outputs(6230) <= not b;
    layer3_outputs(6231) <= not b;
    layer3_outputs(6232) <= not b or a;
    layer3_outputs(6233) <= a;
    layer3_outputs(6234) <= b and not a;
    layer3_outputs(6235) <= a and not b;
    layer3_outputs(6236) <= not a;
    layer3_outputs(6237) <= not a;
    layer3_outputs(6238) <= a or b;
    layer3_outputs(6239) <= a or b;
    layer3_outputs(6240) <= 1'b0;
    layer3_outputs(6241) <= b;
    layer3_outputs(6242) <= a or b;
    layer3_outputs(6243) <= 1'b0;
    layer3_outputs(6244) <= a;
    layer3_outputs(6245) <= not b or a;
    layer3_outputs(6246) <= not a or b;
    layer3_outputs(6247) <= b;
    layer3_outputs(6248) <= not (a and b);
    layer3_outputs(6249) <= 1'b1;
    layer3_outputs(6250) <= 1'b0;
    layer3_outputs(6251) <= not a or b;
    layer3_outputs(6252) <= not b;
    layer3_outputs(6253) <= not (a and b);
    layer3_outputs(6254) <= not b or a;
    layer3_outputs(6255) <= a and not b;
    layer3_outputs(6256) <= b and not a;
    layer3_outputs(6257) <= not b or a;
    layer3_outputs(6258) <= not b or a;
    layer3_outputs(6259) <= not (a or b);
    layer3_outputs(6260) <= a and not b;
    layer3_outputs(6261) <= b and not a;
    layer3_outputs(6262) <= b and not a;
    layer3_outputs(6263) <= not (a xor b);
    layer3_outputs(6264) <= not b;
    layer3_outputs(6265) <= not (a or b);
    layer3_outputs(6266) <= not (a and b);
    layer3_outputs(6267) <= a or b;
    layer3_outputs(6268) <= a and not b;
    layer3_outputs(6269) <= a xor b;
    layer3_outputs(6270) <= b and not a;
    layer3_outputs(6271) <= not b;
    layer3_outputs(6272) <= a and b;
    layer3_outputs(6273) <= not (a or b);
    layer3_outputs(6274) <= 1'b1;
    layer3_outputs(6275) <= not (a and b);
    layer3_outputs(6276) <= b;
    layer3_outputs(6277) <= not b;
    layer3_outputs(6278) <= not b;
    layer3_outputs(6279) <= not b or a;
    layer3_outputs(6280) <= 1'b1;
    layer3_outputs(6281) <= 1'b1;
    layer3_outputs(6282) <= b;
    layer3_outputs(6283) <= not (a xor b);
    layer3_outputs(6284) <= a xor b;
    layer3_outputs(6285) <= not (a xor b);
    layer3_outputs(6286) <= b and not a;
    layer3_outputs(6287) <= not (a xor b);
    layer3_outputs(6288) <= not b;
    layer3_outputs(6289) <= b and not a;
    layer3_outputs(6290) <= b and not a;
    layer3_outputs(6291) <= not a;
    layer3_outputs(6292) <= not a;
    layer3_outputs(6293) <= a and b;
    layer3_outputs(6294) <= not b or a;
    layer3_outputs(6295) <= b and not a;
    layer3_outputs(6296) <= 1'b1;
    layer3_outputs(6297) <= 1'b1;
    layer3_outputs(6298) <= b;
    layer3_outputs(6299) <= not (a or b);
    layer3_outputs(6300) <= not b;
    layer3_outputs(6301) <= 1'b0;
    layer3_outputs(6302) <= b and not a;
    layer3_outputs(6303) <= not (a or b);
    layer3_outputs(6304) <= a and not b;
    layer3_outputs(6305) <= a and b;
    layer3_outputs(6306) <= a or b;
    layer3_outputs(6307) <= a or b;
    layer3_outputs(6308) <= not b;
    layer3_outputs(6309) <= 1'b0;
    layer3_outputs(6310) <= not b;
    layer3_outputs(6311) <= 1'b0;
    layer3_outputs(6312) <= a or b;
    layer3_outputs(6313) <= 1'b0;
    layer3_outputs(6314) <= a and not b;
    layer3_outputs(6315) <= not (a and b);
    layer3_outputs(6316) <= not (a and b);
    layer3_outputs(6317) <= 1'b1;
    layer3_outputs(6318) <= a or b;
    layer3_outputs(6319) <= 1'b0;
    layer3_outputs(6320) <= not (a xor b);
    layer3_outputs(6321) <= a and not b;
    layer3_outputs(6322) <= not b or a;
    layer3_outputs(6323) <= b and not a;
    layer3_outputs(6324) <= not (a or b);
    layer3_outputs(6325) <= not (a xor b);
    layer3_outputs(6326) <= a;
    layer3_outputs(6327) <= a or b;
    layer3_outputs(6328) <= not (a and b);
    layer3_outputs(6329) <= a;
    layer3_outputs(6330) <= 1'b0;
    layer3_outputs(6331) <= b and not a;
    layer3_outputs(6332) <= a or b;
    layer3_outputs(6333) <= not (a or b);
    layer3_outputs(6334) <= a and b;
    layer3_outputs(6335) <= not a or b;
    layer3_outputs(6336) <= not (a or b);
    layer3_outputs(6337) <= a or b;
    layer3_outputs(6338) <= not (a and b);
    layer3_outputs(6339) <= a;
    layer3_outputs(6340) <= not a;
    layer3_outputs(6341) <= a;
    layer3_outputs(6342) <= a and not b;
    layer3_outputs(6343) <= not b or a;
    layer3_outputs(6344) <= a;
    layer3_outputs(6345) <= not (a and b);
    layer3_outputs(6346) <= b and not a;
    layer3_outputs(6347) <= a or b;
    layer3_outputs(6348) <= a and not b;
    layer3_outputs(6349) <= not b;
    layer3_outputs(6350) <= not a or b;
    layer3_outputs(6351) <= a;
    layer3_outputs(6352) <= not a or b;
    layer3_outputs(6353) <= not a;
    layer3_outputs(6354) <= not (a and b);
    layer3_outputs(6355) <= not (a or b);
    layer3_outputs(6356) <= 1'b1;
    layer3_outputs(6357) <= a;
    layer3_outputs(6358) <= 1'b0;
    layer3_outputs(6359) <= not a or b;
    layer3_outputs(6360) <= b;
    layer3_outputs(6361) <= a and b;
    layer3_outputs(6362) <= not (a or b);
    layer3_outputs(6363) <= 1'b0;
    layer3_outputs(6364) <= a xor b;
    layer3_outputs(6365) <= 1'b0;
    layer3_outputs(6366) <= 1'b0;
    layer3_outputs(6367) <= a and b;
    layer3_outputs(6368) <= a or b;
    layer3_outputs(6369) <= a and not b;
    layer3_outputs(6370) <= not a or b;
    layer3_outputs(6371) <= b and not a;
    layer3_outputs(6372) <= not b;
    layer3_outputs(6373) <= not b or a;
    layer3_outputs(6374) <= a or b;
    layer3_outputs(6375) <= not b;
    layer3_outputs(6376) <= not b or a;
    layer3_outputs(6377) <= not a;
    layer3_outputs(6378) <= b and not a;
    layer3_outputs(6379) <= not (a and b);
    layer3_outputs(6380) <= b;
    layer3_outputs(6381) <= not (a or b);
    layer3_outputs(6382) <= a and not b;
    layer3_outputs(6383) <= a or b;
    layer3_outputs(6384) <= not (a or b);
    layer3_outputs(6385) <= not (a and b);
    layer3_outputs(6386) <= not b;
    layer3_outputs(6387) <= 1'b0;
    layer3_outputs(6388) <= 1'b1;
    layer3_outputs(6389) <= 1'b1;
    layer3_outputs(6390) <= not b or a;
    layer3_outputs(6391) <= not a;
    layer3_outputs(6392) <= a and not b;
    layer3_outputs(6393) <= 1'b0;
    layer3_outputs(6394) <= a and b;
    layer3_outputs(6395) <= not b;
    layer3_outputs(6396) <= not a;
    layer3_outputs(6397) <= not a or b;
    layer3_outputs(6398) <= b and not a;
    layer3_outputs(6399) <= not (a or b);
    layer3_outputs(6400) <= a or b;
    layer3_outputs(6401) <= a;
    layer3_outputs(6402) <= b;
    layer3_outputs(6403) <= a and b;
    layer3_outputs(6404) <= a xor b;
    layer3_outputs(6405) <= a and b;
    layer3_outputs(6406) <= b and not a;
    layer3_outputs(6407) <= a and not b;
    layer3_outputs(6408) <= not a or b;
    layer3_outputs(6409) <= not (a or b);
    layer3_outputs(6410) <= a;
    layer3_outputs(6411) <= a;
    layer3_outputs(6412) <= a;
    layer3_outputs(6413) <= not b;
    layer3_outputs(6414) <= b and not a;
    layer3_outputs(6415) <= not b or a;
    layer3_outputs(6416) <= b;
    layer3_outputs(6417) <= not a or b;
    layer3_outputs(6418) <= a and not b;
    layer3_outputs(6419) <= b and not a;
    layer3_outputs(6420) <= a and b;
    layer3_outputs(6421) <= not a or b;
    layer3_outputs(6422) <= not b or a;
    layer3_outputs(6423) <= a and b;
    layer3_outputs(6424) <= a;
    layer3_outputs(6425) <= a and b;
    layer3_outputs(6426) <= a or b;
    layer3_outputs(6427) <= not (a and b);
    layer3_outputs(6428) <= not (a or b);
    layer3_outputs(6429) <= a and not b;
    layer3_outputs(6430) <= a and not b;
    layer3_outputs(6431) <= a and b;
    layer3_outputs(6432) <= not a or b;
    layer3_outputs(6433) <= not a or b;
    layer3_outputs(6434) <= a and b;
    layer3_outputs(6435) <= not b;
    layer3_outputs(6436) <= 1'b1;
    layer3_outputs(6437) <= a;
    layer3_outputs(6438) <= a and not b;
    layer3_outputs(6439) <= a and b;
    layer3_outputs(6440) <= not b or a;
    layer3_outputs(6441) <= 1'b1;
    layer3_outputs(6442) <= 1'b0;
    layer3_outputs(6443) <= not b;
    layer3_outputs(6444) <= not a;
    layer3_outputs(6445) <= b;
    layer3_outputs(6446) <= a xor b;
    layer3_outputs(6447) <= not a or b;
    layer3_outputs(6448) <= b and not a;
    layer3_outputs(6449) <= 1'b1;
    layer3_outputs(6450) <= not (a and b);
    layer3_outputs(6451) <= not a or b;
    layer3_outputs(6452) <= not a;
    layer3_outputs(6453) <= a;
    layer3_outputs(6454) <= a or b;
    layer3_outputs(6455) <= not a or b;
    layer3_outputs(6456) <= not a;
    layer3_outputs(6457) <= not (a and b);
    layer3_outputs(6458) <= not (a or b);
    layer3_outputs(6459) <= a and b;
    layer3_outputs(6460) <= not a;
    layer3_outputs(6461) <= not b;
    layer3_outputs(6462) <= 1'b0;
    layer3_outputs(6463) <= a or b;
    layer3_outputs(6464) <= 1'b0;
    layer3_outputs(6465) <= a and b;
    layer3_outputs(6466) <= not (a and b);
    layer3_outputs(6467) <= b and not a;
    layer3_outputs(6468) <= a and not b;
    layer3_outputs(6469) <= b and not a;
    layer3_outputs(6470) <= not (a xor b);
    layer3_outputs(6471) <= not (a or b);
    layer3_outputs(6472) <= not a;
    layer3_outputs(6473) <= not a;
    layer3_outputs(6474) <= a and b;
    layer3_outputs(6475) <= not a;
    layer3_outputs(6476) <= a or b;
    layer3_outputs(6477) <= not (a xor b);
    layer3_outputs(6478) <= b;
    layer3_outputs(6479) <= a;
    layer3_outputs(6480) <= not a;
    layer3_outputs(6481) <= b and not a;
    layer3_outputs(6482) <= not (a and b);
    layer3_outputs(6483) <= not b;
    layer3_outputs(6484) <= not (a xor b);
    layer3_outputs(6485) <= not b;
    layer3_outputs(6486) <= 1'b1;
    layer3_outputs(6487) <= not a;
    layer3_outputs(6488) <= not a;
    layer3_outputs(6489) <= not b or a;
    layer3_outputs(6490) <= not b;
    layer3_outputs(6491) <= not (a xor b);
    layer3_outputs(6492) <= not (a and b);
    layer3_outputs(6493) <= a and b;
    layer3_outputs(6494) <= a;
    layer3_outputs(6495) <= not b or a;
    layer3_outputs(6496) <= a and not b;
    layer3_outputs(6497) <= not b or a;
    layer3_outputs(6498) <= not a or b;
    layer3_outputs(6499) <= not (a or b);
    layer3_outputs(6500) <= not (a xor b);
    layer3_outputs(6501) <= not a;
    layer3_outputs(6502) <= a or b;
    layer3_outputs(6503) <= 1'b1;
    layer3_outputs(6504) <= a and b;
    layer3_outputs(6505) <= a and b;
    layer3_outputs(6506) <= a and not b;
    layer3_outputs(6507) <= b and not a;
    layer3_outputs(6508) <= b;
    layer3_outputs(6509) <= not (a xor b);
    layer3_outputs(6510) <= a and not b;
    layer3_outputs(6511) <= a xor b;
    layer3_outputs(6512) <= 1'b1;
    layer3_outputs(6513) <= b and not a;
    layer3_outputs(6514) <= not b;
    layer3_outputs(6515) <= a or b;
    layer3_outputs(6516) <= a;
    layer3_outputs(6517) <= not b;
    layer3_outputs(6518) <= 1'b1;
    layer3_outputs(6519) <= not b or a;
    layer3_outputs(6520) <= not (a and b);
    layer3_outputs(6521) <= not a;
    layer3_outputs(6522) <= not b or a;
    layer3_outputs(6523) <= a and b;
    layer3_outputs(6524) <= 1'b1;
    layer3_outputs(6525) <= not a;
    layer3_outputs(6526) <= a;
    layer3_outputs(6527) <= a or b;
    layer3_outputs(6528) <= a and b;
    layer3_outputs(6529) <= a;
    layer3_outputs(6530) <= a and b;
    layer3_outputs(6531) <= 1'b0;
    layer3_outputs(6532) <= a;
    layer3_outputs(6533) <= a or b;
    layer3_outputs(6534) <= a and not b;
    layer3_outputs(6535) <= not (a xor b);
    layer3_outputs(6536) <= not b or a;
    layer3_outputs(6537) <= a or b;
    layer3_outputs(6538) <= a and not b;
    layer3_outputs(6539) <= a;
    layer3_outputs(6540) <= a and not b;
    layer3_outputs(6541) <= 1'b1;
    layer3_outputs(6542) <= b;
    layer3_outputs(6543) <= a and not b;
    layer3_outputs(6544) <= not (a and b);
    layer3_outputs(6545) <= b and not a;
    layer3_outputs(6546) <= not (a and b);
    layer3_outputs(6547) <= a;
    layer3_outputs(6548) <= a and b;
    layer3_outputs(6549) <= 1'b0;
    layer3_outputs(6550) <= 1'b1;
    layer3_outputs(6551) <= not (a and b);
    layer3_outputs(6552) <= not (a and b);
    layer3_outputs(6553) <= not (a xor b);
    layer3_outputs(6554) <= not a;
    layer3_outputs(6555) <= 1'b1;
    layer3_outputs(6556) <= 1'b0;
    layer3_outputs(6557) <= not a;
    layer3_outputs(6558) <= not (a and b);
    layer3_outputs(6559) <= 1'b0;
    layer3_outputs(6560) <= a and b;
    layer3_outputs(6561) <= 1'b1;
    layer3_outputs(6562) <= a and b;
    layer3_outputs(6563) <= a xor b;
    layer3_outputs(6564) <= b and not a;
    layer3_outputs(6565) <= a and b;
    layer3_outputs(6566) <= a or b;
    layer3_outputs(6567) <= not b or a;
    layer3_outputs(6568) <= not a;
    layer3_outputs(6569) <= a xor b;
    layer3_outputs(6570) <= a;
    layer3_outputs(6571) <= not (a or b);
    layer3_outputs(6572) <= b and not a;
    layer3_outputs(6573) <= not (a or b);
    layer3_outputs(6574) <= a and b;
    layer3_outputs(6575) <= not (a or b);
    layer3_outputs(6576) <= not a;
    layer3_outputs(6577) <= b and not a;
    layer3_outputs(6578) <= a or b;
    layer3_outputs(6579) <= a or b;
    layer3_outputs(6580) <= not b;
    layer3_outputs(6581) <= b;
    layer3_outputs(6582) <= not a or b;
    layer3_outputs(6583) <= not a;
    layer3_outputs(6584) <= a or b;
    layer3_outputs(6585) <= not (a or b);
    layer3_outputs(6586) <= not (a or b);
    layer3_outputs(6587) <= b and not a;
    layer3_outputs(6588) <= a or b;
    layer3_outputs(6589) <= not b or a;
    layer3_outputs(6590) <= a or b;
    layer3_outputs(6591) <= a or b;
    layer3_outputs(6592) <= a and b;
    layer3_outputs(6593) <= b;
    layer3_outputs(6594) <= not b;
    layer3_outputs(6595) <= not (a and b);
    layer3_outputs(6596) <= 1'b1;
    layer3_outputs(6597) <= a;
    layer3_outputs(6598) <= not a or b;
    layer3_outputs(6599) <= b and not a;
    layer3_outputs(6600) <= not b;
    layer3_outputs(6601) <= a and not b;
    layer3_outputs(6602) <= not (a and b);
    layer3_outputs(6603) <= 1'b1;
    layer3_outputs(6604) <= b and not a;
    layer3_outputs(6605) <= not (a and b);
    layer3_outputs(6606) <= b and not a;
    layer3_outputs(6607) <= not (a and b);
    layer3_outputs(6608) <= not (a or b);
    layer3_outputs(6609) <= a;
    layer3_outputs(6610) <= a and not b;
    layer3_outputs(6611) <= not (a or b);
    layer3_outputs(6612) <= a and b;
    layer3_outputs(6613) <= a or b;
    layer3_outputs(6614) <= b;
    layer3_outputs(6615) <= b and not a;
    layer3_outputs(6616) <= not b or a;
    layer3_outputs(6617) <= not b;
    layer3_outputs(6618) <= 1'b1;
    layer3_outputs(6619) <= not (a and b);
    layer3_outputs(6620) <= a or b;
    layer3_outputs(6621) <= a and not b;
    layer3_outputs(6622) <= b;
    layer3_outputs(6623) <= a;
    layer3_outputs(6624) <= not (a and b);
    layer3_outputs(6625) <= not (a and b);
    layer3_outputs(6626) <= a and b;
    layer3_outputs(6627) <= 1'b0;
    layer3_outputs(6628) <= not a;
    layer3_outputs(6629) <= not b or a;
    layer3_outputs(6630) <= a and b;
    layer3_outputs(6631) <= not b;
    layer3_outputs(6632) <= a;
    layer3_outputs(6633) <= a and b;
    layer3_outputs(6634) <= not b;
    layer3_outputs(6635) <= not b or a;
    layer3_outputs(6636) <= not (a xor b);
    layer3_outputs(6637) <= a;
    layer3_outputs(6638) <= b and not a;
    layer3_outputs(6639) <= b and not a;
    layer3_outputs(6640) <= not b or a;
    layer3_outputs(6641) <= b and not a;
    layer3_outputs(6642) <= not a or b;
    layer3_outputs(6643) <= not (a or b);
    layer3_outputs(6644) <= b;
    layer3_outputs(6645) <= 1'b0;
    layer3_outputs(6646) <= a and not b;
    layer3_outputs(6647) <= a and b;
    layer3_outputs(6648) <= 1'b1;
    layer3_outputs(6649) <= b;
    layer3_outputs(6650) <= 1'b0;
    layer3_outputs(6651) <= 1'b1;
    layer3_outputs(6652) <= a and not b;
    layer3_outputs(6653) <= 1'b1;
    layer3_outputs(6654) <= a and b;
    layer3_outputs(6655) <= a and b;
    layer3_outputs(6656) <= not a or b;
    layer3_outputs(6657) <= 1'b0;
    layer3_outputs(6658) <= not a or b;
    layer3_outputs(6659) <= b and not a;
    layer3_outputs(6660) <= a and b;
    layer3_outputs(6661) <= 1'b0;
    layer3_outputs(6662) <= a or b;
    layer3_outputs(6663) <= a xor b;
    layer3_outputs(6664) <= 1'b1;
    layer3_outputs(6665) <= not b or a;
    layer3_outputs(6666) <= not (a or b);
    layer3_outputs(6667) <= a and b;
    layer3_outputs(6668) <= not b or a;
    layer3_outputs(6669) <= 1'b0;
    layer3_outputs(6670) <= b;
    layer3_outputs(6671) <= a;
    layer3_outputs(6672) <= not (a xor b);
    layer3_outputs(6673) <= 1'b0;
    layer3_outputs(6674) <= 1'b1;
    layer3_outputs(6675) <= not a;
    layer3_outputs(6676) <= b;
    layer3_outputs(6677) <= 1'b1;
    layer3_outputs(6678) <= not (a and b);
    layer3_outputs(6679) <= b and not a;
    layer3_outputs(6680) <= 1'b1;
    layer3_outputs(6681) <= a xor b;
    layer3_outputs(6682) <= a and not b;
    layer3_outputs(6683) <= a and not b;
    layer3_outputs(6684) <= b and not a;
    layer3_outputs(6685) <= not a;
    layer3_outputs(6686) <= b;
    layer3_outputs(6687) <= not a;
    layer3_outputs(6688) <= not a or b;
    layer3_outputs(6689) <= a and not b;
    layer3_outputs(6690) <= not b;
    layer3_outputs(6691) <= not (a or b);
    layer3_outputs(6692) <= a;
    layer3_outputs(6693) <= a or b;
    layer3_outputs(6694) <= 1'b0;
    layer3_outputs(6695) <= a or b;
    layer3_outputs(6696) <= a xor b;
    layer3_outputs(6697) <= 1'b1;
    layer3_outputs(6698) <= a and not b;
    layer3_outputs(6699) <= a and b;
    layer3_outputs(6700) <= a xor b;
    layer3_outputs(6701) <= a and b;
    layer3_outputs(6702) <= a and not b;
    layer3_outputs(6703) <= 1'b1;
    layer3_outputs(6704) <= 1'b1;
    layer3_outputs(6705) <= b;
    layer3_outputs(6706) <= b and not a;
    layer3_outputs(6707) <= b;
    layer3_outputs(6708) <= 1'b0;
    layer3_outputs(6709) <= not (a and b);
    layer3_outputs(6710) <= b and not a;
    layer3_outputs(6711) <= a and not b;
    layer3_outputs(6712) <= not (a or b);
    layer3_outputs(6713) <= a or b;
    layer3_outputs(6714) <= not a or b;
    layer3_outputs(6715) <= a or b;
    layer3_outputs(6716) <= 1'b0;
    layer3_outputs(6717) <= not a or b;
    layer3_outputs(6718) <= 1'b1;
    layer3_outputs(6719) <= 1'b1;
    layer3_outputs(6720) <= b and not a;
    layer3_outputs(6721) <= a xor b;
    layer3_outputs(6722) <= not b or a;
    layer3_outputs(6723) <= not a;
    layer3_outputs(6724) <= a and not b;
    layer3_outputs(6725) <= not (a and b);
    layer3_outputs(6726) <= not b;
    layer3_outputs(6727) <= 1'b1;
    layer3_outputs(6728) <= 1'b0;
    layer3_outputs(6729) <= not b;
    layer3_outputs(6730) <= not b or a;
    layer3_outputs(6731) <= a and not b;
    layer3_outputs(6732) <= not a;
    layer3_outputs(6733) <= not b;
    layer3_outputs(6734) <= not b;
    layer3_outputs(6735) <= a;
    layer3_outputs(6736) <= a and b;
    layer3_outputs(6737) <= a and b;
    layer3_outputs(6738) <= 1'b1;
    layer3_outputs(6739) <= a or b;
    layer3_outputs(6740) <= not (a and b);
    layer3_outputs(6741) <= not b;
    layer3_outputs(6742) <= a and b;
    layer3_outputs(6743) <= a xor b;
    layer3_outputs(6744) <= not (a and b);
    layer3_outputs(6745) <= not a;
    layer3_outputs(6746) <= a or b;
    layer3_outputs(6747) <= a and not b;
    layer3_outputs(6748) <= a and not b;
    layer3_outputs(6749) <= b and not a;
    layer3_outputs(6750) <= a and b;
    layer3_outputs(6751) <= a;
    layer3_outputs(6752) <= not (a and b);
    layer3_outputs(6753) <= a and b;
    layer3_outputs(6754) <= b;
    layer3_outputs(6755) <= not a;
    layer3_outputs(6756) <= 1'b1;
    layer3_outputs(6757) <= not (a xor b);
    layer3_outputs(6758) <= not (a or b);
    layer3_outputs(6759) <= a and not b;
    layer3_outputs(6760) <= not (a or b);
    layer3_outputs(6761) <= 1'b0;
    layer3_outputs(6762) <= not a;
    layer3_outputs(6763) <= not (a and b);
    layer3_outputs(6764) <= 1'b1;
    layer3_outputs(6765) <= 1'b0;
    layer3_outputs(6766) <= b;
    layer3_outputs(6767) <= a;
    layer3_outputs(6768) <= 1'b0;
    layer3_outputs(6769) <= not b;
    layer3_outputs(6770) <= not a or b;
    layer3_outputs(6771) <= not (a and b);
    layer3_outputs(6772) <= not (a or b);
    layer3_outputs(6773) <= not b;
    layer3_outputs(6774) <= 1'b1;
    layer3_outputs(6775) <= a or b;
    layer3_outputs(6776) <= b;
    layer3_outputs(6777) <= not (a and b);
    layer3_outputs(6778) <= 1'b0;
    layer3_outputs(6779) <= 1'b0;
    layer3_outputs(6780) <= not b or a;
    layer3_outputs(6781) <= not (a or b);
    layer3_outputs(6782) <= a;
    layer3_outputs(6783) <= not a;
    layer3_outputs(6784) <= not b or a;
    layer3_outputs(6785) <= not a;
    layer3_outputs(6786) <= 1'b1;
    layer3_outputs(6787) <= not b or a;
    layer3_outputs(6788) <= a;
    layer3_outputs(6789) <= 1'b1;
    layer3_outputs(6790) <= not a;
    layer3_outputs(6791) <= 1'b1;
    layer3_outputs(6792) <= a or b;
    layer3_outputs(6793) <= a and not b;
    layer3_outputs(6794) <= not (a and b);
    layer3_outputs(6795) <= not b or a;
    layer3_outputs(6796) <= b;
    layer3_outputs(6797) <= not (a or b);
    layer3_outputs(6798) <= not (a and b);
    layer3_outputs(6799) <= 1'b1;
    layer3_outputs(6800) <= b and not a;
    layer3_outputs(6801) <= 1'b1;
    layer3_outputs(6802) <= a xor b;
    layer3_outputs(6803) <= not (a or b);
    layer3_outputs(6804) <= not b;
    layer3_outputs(6805) <= a;
    layer3_outputs(6806) <= 1'b1;
    layer3_outputs(6807) <= not (a or b);
    layer3_outputs(6808) <= a;
    layer3_outputs(6809) <= not (a xor b);
    layer3_outputs(6810) <= a and not b;
    layer3_outputs(6811) <= 1'b0;
    layer3_outputs(6812) <= a and not b;
    layer3_outputs(6813) <= a and b;
    layer3_outputs(6814) <= b;
    layer3_outputs(6815) <= 1'b0;
    layer3_outputs(6816) <= a;
    layer3_outputs(6817) <= a xor b;
    layer3_outputs(6818) <= not b;
    layer3_outputs(6819) <= a;
    layer3_outputs(6820) <= not (a and b);
    layer3_outputs(6821) <= not (a or b);
    layer3_outputs(6822) <= a and b;
    layer3_outputs(6823) <= not b or a;
    layer3_outputs(6824) <= not b or a;
    layer3_outputs(6825) <= not a or b;
    layer3_outputs(6826) <= not a;
    layer3_outputs(6827) <= 1'b0;
    layer3_outputs(6828) <= 1'b1;
    layer3_outputs(6829) <= not a;
    layer3_outputs(6830) <= not (a or b);
    layer3_outputs(6831) <= not a;
    layer3_outputs(6832) <= a and b;
    layer3_outputs(6833) <= not a or b;
    layer3_outputs(6834) <= not b;
    layer3_outputs(6835) <= not a or b;
    layer3_outputs(6836) <= b and not a;
    layer3_outputs(6837) <= a and not b;
    layer3_outputs(6838) <= a or b;
    layer3_outputs(6839) <= not b;
    layer3_outputs(6840) <= not b;
    layer3_outputs(6841) <= not (a and b);
    layer3_outputs(6842) <= not a;
    layer3_outputs(6843) <= a or b;
    layer3_outputs(6844) <= 1'b1;
    layer3_outputs(6845) <= a or b;
    layer3_outputs(6846) <= a;
    layer3_outputs(6847) <= a and b;
    layer3_outputs(6848) <= not (a or b);
    layer3_outputs(6849) <= not (a or b);
    layer3_outputs(6850) <= not (a or b);
    layer3_outputs(6851) <= 1'b0;
    layer3_outputs(6852) <= not (a or b);
    layer3_outputs(6853) <= 1'b1;
    layer3_outputs(6854) <= not a or b;
    layer3_outputs(6855) <= a;
    layer3_outputs(6856) <= a and b;
    layer3_outputs(6857) <= b and not a;
    layer3_outputs(6858) <= not (a and b);
    layer3_outputs(6859) <= 1'b1;
    layer3_outputs(6860) <= a;
    layer3_outputs(6861) <= not b;
    layer3_outputs(6862) <= a or b;
    layer3_outputs(6863) <= 1'b0;
    layer3_outputs(6864) <= b;
    layer3_outputs(6865) <= b and not a;
    layer3_outputs(6866) <= not b;
    layer3_outputs(6867) <= not b or a;
    layer3_outputs(6868) <= not (a and b);
    layer3_outputs(6869) <= not a or b;
    layer3_outputs(6870) <= 1'b0;
    layer3_outputs(6871) <= a or b;
    layer3_outputs(6872) <= b and not a;
    layer3_outputs(6873) <= not b;
    layer3_outputs(6874) <= not a or b;
    layer3_outputs(6875) <= not a;
    layer3_outputs(6876) <= b and not a;
    layer3_outputs(6877) <= not (a and b);
    layer3_outputs(6878) <= not b or a;
    layer3_outputs(6879) <= not b;
    layer3_outputs(6880) <= not a;
    layer3_outputs(6881) <= not a;
    layer3_outputs(6882) <= not (a and b);
    layer3_outputs(6883) <= not b or a;
    layer3_outputs(6884) <= a and b;
    layer3_outputs(6885) <= 1'b1;
    layer3_outputs(6886) <= b;
    layer3_outputs(6887) <= not b;
    layer3_outputs(6888) <= a and b;
    layer3_outputs(6889) <= a or b;
    layer3_outputs(6890) <= not (a or b);
    layer3_outputs(6891) <= not a;
    layer3_outputs(6892) <= a;
    layer3_outputs(6893) <= not (a xor b);
    layer3_outputs(6894) <= b and not a;
    layer3_outputs(6895) <= b and not a;
    layer3_outputs(6896) <= 1'b0;
    layer3_outputs(6897) <= not a;
    layer3_outputs(6898) <= a and b;
    layer3_outputs(6899) <= b;
    layer3_outputs(6900) <= 1'b1;
    layer3_outputs(6901) <= a xor b;
    layer3_outputs(6902) <= not a;
    layer3_outputs(6903) <= 1'b1;
    layer3_outputs(6904) <= a or b;
    layer3_outputs(6905) <= not b;
    layer3_outputs(6906) <= not (a xor b);
    layer3_outputs(6907) <= not a or b;
    layer3_outputs(6908) <= a;
    layer3_outputs(6909) <= 1'b1;
    layer3_outputs(6910) <= not a or b;
    layer3_outputs(6911) <= b;
    layer3_outputs(6912) <= b;
    layer3_outputs(6913) <= b;
    layer3_outputs(6914) <= a or b;
    layer3_outputs(6915) <= not b or a;
    layer3_outputs(6916) <= not (a or b);
    layer3_outputs(6917) <= 1'b0;
    layer3_outputs(6918) <= not a;
    layer3_outputs(6919) <= not a;
    layer3_outputs(6920) <= 1'b1;
    layer3_outputs(6921) <= a and b;
    layer3_outputs(6922) <= not (a and b);
    layer3_outputs(6923) <= not (a or b);
    layer3_outputs(6924) <= not a or b;
    layer3_outputs(6925) <= a;
    layer3_outputs(6926) <= b;
    layer3_outputs(6927) <= b;
    layer3_outputs(6928) <= b;
    layer3_outputs(6929) <= a and not b;
    layer3_outputs(6930) <= b;
    layer3_outputs(6931) <= 1'b1;
    layer3_outputs(6932) <= 1'b0;
    layer3_outputs(6933) <= a and not b;
    layer3_outputs(6934) <= b and not a;
    layer3_outputs(6935) <= 1'b1;
    layer3_outputs(6936) <= not (a xor b);
    layer3_outputs(6937) <= not (a and b);
    layer3_outputs(6938) <= not a or b;
    layer3_outputs(6939) <= not a or b;
    layer3_outputs(6940) <= 1'b0;
    layer3_outputs(6941) <= a and not b;
    layer3_outputs(6942) <= not a or b;
    layer3_outputs(6943) <= 1'b1;
    layer3_outputs(6944) <= 1'b1;
    layer3_outputs(6945) <= not (a or b);
    layer3_outputs(6946) <= a;
    layer3_outputs(6947) <= 1'b0;
    layer3_outputs(6948) <= b;
    layer3_outputs(6949) <= a;
    layer3_outputs(6950) <= a and b;
    layer3_outputs(6951) <= b and not a;
    layer3_outputs(6952) <= b and not a;
    layer3_outputs(6953) <= a and b;
    layer3_outputs(6954) <= not b;
    layer3_outputs(6955) <= a and not b;
    layer3_outputs(6956) <= not b or a;
    layer3_outputs(6957) <= not b or a;
    layer3_outputs(6958) <= b and not a;
    layer3_outputs(6959) <= 1'b1;
    layer3_outputs(6960) <= b and not a;
    layer3_outputs(6961) <= a and not b;
    layer3_outputs(6962) <= a or b;
    layer3_outputs(6963) <= a;
    layer3_outputs(6964) <= not a or b;
    layer3_outputs(6965) <= not b;
    layer3_outputs(6966) <= not a or b;
    layer3_outputs(6967) <= 1'b1;
    layer3_outputs(6968) <= not a or b;
    layer3_outputs(6969) <= a;
    layer3_outputs(6970) <= not a or b;
    layer3_outputs(6971) <= a or b;
    layer3_outputs(6972) <= not (a or b);
    layer3_outputs(6973) <= b and not a;
    layer3_outputs(6974) <= 1'b1;
    layer3_outputs(6975) <= not a or b;
    layer3_outputs(6976) <= b and not a;
    layer3_outputs(6977) <= 1'b1;
    layer3_outputs(6978) <= b;
    layer3_outputs(6979) <= not (a or b);
    layer3_outputs(6980) <= a or b;
    layer3_outputs(6981) <= b;
    layer3_outputs(6982) <= b;
    layer3_outputs(6983) <= not (a and b);
    layer3_outputs(6984) <= not (a xor b);
    layer3_outputs(6985) <= a;
    layer3_outputs(6986) <= a and b;
    layer3_outputs(6987) <= a and not b;
    layer3_outputs(6988) <= a;
    layer3_outputs(6989) <= a and b;
    layer3_outputs(6990) <= a and not b;
    layer3_outputs(6991) <= a and not b;
    layer3_outputs(6992) <= 1'b1;
    layer3_outputs(6993) <= b;
    layer3_outputs(6994) <= a and not b;
    layer3_outputs(6995) <= a and not b;
    layer3_outputs(6996) <= 1'b1;
    layer3_outputs(6997) <= a or b;
    layer3_outputs(6998) <= b;
    layer3_outputs(6999) <= a and not b;
    layer3_outputs(7000) <= a or b;
    layer3_outputs(7001) <= a and b;
    layer3_outputs(7002) <= not (a or b);
    layer3_outputs(7003) <= not b;
    layer3_outputs(7004) <= b;
    layer3_outputs(7005) <= 1'b1;
    layer3_outputs(7006) <= not a;
    layer3_outputs(7007) <= a and not b;
    layer3_outputs(7008) <= 1'b0;
    layer3_outputs(7009) <= not (a and b);
    layer3_outputs(7010) <= 1'b1;
    layer3_outputs(7011) <= not a;
    layer3_outputs(7012) <= a and not b;
    layer3_outputs(7013) <= a;
    layer3_outputs(7014) <= a or b;
    layer3_outputs(7015) <= a and not b;
    layer3_outputs(7016) <= a and not b;
    layer3_outputs(7017) <= a or b;
    layer3_outputs(7018) <= 1'b0;
    layer3_outputs(7019) <= 1'b0;
    layer3_outputs(7020) <= b and not a;
    layer3_outputs(7021) <= not (a or b);
    layer3_outputs(7022) <= not a;
    layer3_outputs(7023) <= not a;
    layer3_outputs(7024) <= b;
    layer3_outputs(7025) <= not a or b;
    layer3_outputs(7026) <= 1'b0;
    layer3_outputs(7027) <= a;
    layer3_outputs(7028) <= 1'b1;
    layer3_outputs(7029) <= a and b;
    layer3_outputs(7030) <= 1'b1;
    layer3_outputs(7031) <= a and not b;
    layer3_outputs(7032) <= a or b;
    layer3_outputs(7033) <= a and b;
    layer3_outputs(7034) <= b and not a;
    layer3_outputs(7035) <= not b;
    layer3_outputs(7036) <= 1'b0;
    layer3_outputs(7037) <= 1'b1;
    layer3_outputs(7038) <= a and not b;
    layer3_outputs(7039) <= b;
    layer3_outputs(7040) <= not (a and b);
    layer3_outputs(7041) <= not a or b;
    layer3_outputs(7042) <= 1'b0;
    layer3_outputs(7043) <= b;
    layer3_outputs(7044) <= not (a and b);
    layer3_outputs(7045) <= 1'b0;
    layer3_outputs(7046) <= b and not a;
    layer3_outputs(7047) <= not (a or b);
    layer3_outputs(7048) <= b and not a;
    layer3_outputs(7049) <= a and b;
    layer3_outputs(7050) <= not a;
    layer3_outputs(7051) <= not b;
    layer3_outputs(7052) <= a and b;
    layer3_outputs(7053) <= b;
    layer3_outputs(7054) <= 1'b0;
    layer3_outputs(7055) <= b and not a;
    layer3_outputs(7056) <= b and not a;
    layer3_outputs(7057) <= not a;
    layer3_outputs(7058) <= a and not b;
    layer3_outputs(7059) <= not b;
    layer3_outputs(7060) <= b;
    layer3_outputs(7061) <= a;
    layer3_outputs(7062) <= not b;
    layer3_outputs(7063) <= not a or b;
    layer3_outputs(7064) <= a;
    layer3_outputs(7065) <= not (a and b);
    layer3_outputs(7066) <= a or b;
    layer3_outputs(7067) <= 1'b1;
    layer3_outputs(7068) <= b;
    layer3_outputs(7069) <= not a;
    layer3_outputs(7070) <= a and not b;
    layer3_outputs(7071) <= not b or a;
    layer3_outputs(7072) <= a and b;
    layer3_outputs(7073) <= a xor b;
    layer3_outputs(7074) <= not b or a;
    layer3_outputs(7075) <= 1'b0;
    layer3_outputs(7076) <= b;
    layer3_outputs(7077) <= not (a and b);
    layer3_outputs(7078) <= b;
    layer3_outputs(7079) <= a or b;
    layer3_outputs(7080) <= 1'b1;
    layer3_outputs(7081) <= b and not a;
    layer3_outputs(7082) <= 1'b0;
    layer3_outputs(7083) <= a;
    layer3_outputs(7084) <= not a or b;
    layer3_outputs(7085) <= not b or a;
    layer3_outputs(7086) <= 1'b0;
    layer3_outputs(7087) <= 1'b0;
    layer3_outputs(7088) <= not a;
    layer3_outputs(7089) <= a and b;
    layer3_outputs(7090) <= not a;
    layer3_outputs(7091) <= 1'b1;
    layer3_outputs(7092) <= 1'b0;
    layer3_outputs(7093) <= b and not a;
    layer3_outputs(7094) <= not a or b;
    layer3_outputs(7095) <= not a or b;
    layer3_outputs(7096) <= not a;
    layer3_outputs(7097) <= a;
    layer3_outputs(7098) <= a xor b;
    layer3_outputs(7099) <= a;
    layer3_outputs(7100) <= a;
    layer3_outputs(7101) <= 1'b1;
    layer3_outputs(7102) <= not (a and b);
    layer3_outputs(7103) <= not b or a;
    layer3_outputs(7104) <= a and not b;
    layer3_outputs(7105) <= 1'b0;
    layer3_outputs(7106) <= a;
    layer3_outputs(7107) <= not (a and b);
    layer3_outputs(7108) <= not b or a;
    layer3_outputs(7109) <= not a or b;
    layer3_outputs(7110) <= not (a or b);
    layer3_outputs(7111) <= not (a xor b);
    layer3_outputs(7112) <= not b or a;
    layer3_outputs(7113) <= a and not b;
    layer3_outputs(7114) <= a or b;
    layer3_outputs(7115) <= not (a or b);
    layer3_outputs(7116) <= a and b;
    layer3_outputs(7117) <= b and not a;
    layer3_outputs(7118) <= a and not b;
    layer3_outputs(7119) <= 1'b0;
    layer3_outputs(7120) <= b and not a;
    layer3_outputs(7121) <= a and b;
    layer3_outputs(7122) <= a and b;
    layer3_outputs(7123) <= b;
    layer3_outputs(7124) <= a or b;
    layer3_outputs(7125) <= b;
    layer3_outputs(7126) <= not a or b;
    layer3_outputs(7127) <= a;
    layer3_outputs(7128) <= not (a or b);
    layer3_outputs(7129) <= not (a or b);
    layer3_outputs(7130) <= not a;
    layer3_outputs(7131) <= not b;
    layer3_outputs(7132) <= b;
    layer3_outputs(7133) <= a or b;
    layer3_outputs(7134) <= b and not a;
    layer3_outputs(7135) <= 1'b1;
    layer3_outputs(7136) <= not b;
    layer3_outputs(7137) <= a and b;
    layer3_outputs(7138) <= 1'b1;
    layer3_outputs(7139) <= 1'b1;
    layer3_outputs(7140) <= b;
    layer3_outputs(7141) <= b and not a;
    layer3_outputs(7142) <= not a or b;
    layer3_outputs(7143) <= not a or b;
    layer3_outputs(7144) <= a and b;
    layer3_outputs(7145) <= not a or b;
    layer3_outputs(7146) <= not b;
    layer3_outputs(7147) <= a;
    layer3_outputs(7148) <= not b or a;
    layer3_outputs(7149) <= not a or b;
    layer3_outputs(7150) <= not (a and b);
    layer3_outputs(7151) <= 1'b1;
    layer3_outputs(7152) <= not (a and b);
    layer3_outputs(7153) <= not b or a;
    layer3_outputs(7154) <= b and not a;
    layer3_outputs(7155) <= a;
    layer3_outputs(7156) <= b and not a;
    layer3_outputs(7157) <= a and b;
    layer3_outputs(7158) <= 1'b1;
    layer3_outputs(7159) <= not a or b;
    layer3_outputs(7160) <= a;
    layer3_outputs(7161) <= a xor b;
    layer3_outputs(7162) <= a and not b;
    layer3_outputs(7163) <= a and not b;
    layer3_outputs(7164) <= not a or b;
    layer3_outputs(7165) <= not (a xor b);
    layer3_outputs(7166) <= not (a or b);
    layer3_outputs(7167) <= not a or b;
    layer3_outputs(7168) <= a or b;
    layer3_outputs(7169) <= b;
    layer3_outputs(7170) <= not a;
    layer3_outputs(7171) <= a and not b;
    layer3_outputs(7172) <= a and not b;
    layer3_outputs(7173) <= a and b;
    layer3_outputs(7174) <= not b or a;
    layer3_outputs(7175) <= not b or a;
    layer3_outputs(7176) <= 1'b0;
    layer3_outputs(7177) <= a and not b;
    layer3_outputs(7178) <= a and b;
    layer3_outputs(7179) <= b and not a;
    layer3_outputs(7180) <= a or b;
    layer3_outputs(7181) <= a and not b;
    layer3_outputs(7182) <= not b;
    layer3_outputs(7183) <= a or b;
    layer3_outputs(7184) <= 1'b0;
    layer3_outputs(7185) <= not a;
    layer3_outputs(7186) <= not (a and b);
    layer3_outputs(7187) <= 1'b1;
    layer3_outputs(7188) <= 1'b1;
    layer3_outputs(7189) <= a xor b;
    layer3_outputs(7190) <= a;
    layer3_outputs(7191) <= b and not a;
    layer3_outputs(7192) <= a and b;
    layer3_outputs(7193) <= not b or a;
    layer3_outputs(7194) <= 1'b0;
    layer3_outputs(7195) <= not a;
    layer3_outputs(7196) <= not a;
    layer3_outputs(7197) <= a or b;
    layer3_outputs(7198) <= a;
    layer3_outputs(7199) <= not a or b;
    layer3_outputs(7200) <= 1'b1;
    layer3_outputs(7201) <= not a or b;
    layer3_outputs(7202) <= not a or b;
    layer3_outputs(7203) <= b and not a;
    layer3_outputs(7204) <= a or b;
    layer3_outputs(7205) <= not (a or b);
    layer3_outputs(7206) <= b and not a;
    layer3_outputs(7207) <= a;
    layer3_outputs(7208) <= not b or a;
    layer3_outputs(7209) <= 1'b1;
    layer3_outputs(7210) <= 1'b0;
    layer3_outputs(7211) <= a;
    layer3_outputs(7212) <= a;
    layer3_outputs(7213) <= a and not b;
    layer3_outputs(7214) <= b;
    layer3_outputs(7215) <= a;
    layer3_outputs(7216) <= not (a and b);
    layer3_outputs(7217) <= b;
    layer3_outputs(7218) <= not (a and b);
    layer3_outputs(7219) <= a xor b;
    layer3_outputs(7220) <= not b;
    layer3_outputs(7221) <= 1'b1;
    layer3_outputs(7222) <= b;
    layer3_outputs(7223) <= a;
    layer3_outputs(7224) <= not a;
    layer3_outputs(7225) <= not (a and b);
    layer3_outputs(7226) <= b;
    layer3_outputs(7227) <= not (a or b);
    layer3_outputs(7228) <= a;
    layer3_outputs(7229) <= b;
    layer3_outputs(7230) <= a and not b;
    layer3_outputs(7231) <= a;
    layer3_outputs(7232) <= b;
    layer3_outputs(7233) <= a and not b;
    layer3_outputs(7234) <= not (a or b);
    layer3_outputs(7235) <= not (a and b);
    layer3_outputs(7236) <= not (a and b);
    layer3_outputs(7237) <= a or b;
    layer3_outputs(7238) <= not b or a;
    layer3_outputs(7239) <= a and not b;
    layer3_outputs(7240) <= 1'b0;
    layer3_outputs(7241) <= not b or a;
    layer3_outputs(7242) <= 1'b0;
    layer3_outputs(7243) <= a;
    layer3_outputs(7244) <= 1'b1;
    layer3_outputs(7245) <= not (a and b);
    layer3_outputs(7246) <= not b or a;
    layer3_outputs(7247) <= a;
    layer3_outputs(7248) <= 1'b1;
    layer3_outputs(7249) <= a and not b;
    layer3_outputs(7250) <= not (a or b);
    layer3_outputs(7251) <= a and b;
    layer3_outputs(7252) <= 1'b1;
    layer3_outputs(7253) <= a and b;
    layer3_outputs(7254) <= not a;
    layer3_outputs(7255) <= not (a xor b);
    layer3_outputs(7256) <= not b;
    layer3_outputs(7257) <= a and b;
    layer3_outputs(7258) <= not a or b;
    layer3_outputs(7259) <= not (a and b);
    layer3_outputs(7260) <= not a;
    layer3_outputs(7261) <= 1'b0;
    layer3_outputs(7262) <= not (a or b);
    layer3_outputs(7263) <= 1'b0;
    layer3_outputs(7264) <= 1'b1;
    layer3_outputs(7265) <= not (a and b);
    layer3_outputs(7266) <= b;
    layer3_outputs(7267) <= a or b;
    layer3_outputs(7268) <= not a or b;
    layer3_outputs(7269) <= not (a and b);
    layer3_outputs(7270) <= 1'b1;
    layer3_outputs(7271) <= not b or a;
    layer3_outputs(7272) <= 1'b1;
    layer3_outputs(7273) <= b;
    layer3_outputs(7274) <= not b;
    layer3_outputs(7275) <= a or b;
    layer3_outputs(7276) <= not (a and b);
    layer3_outputs(7277) <= 1'b0;
    layer3_outputs(7278) <= not a or b;
    layer3_outputs(7279) <= a;
    layer3_outputs(7280) <= b;
    layer3_outputs(7281) <= not (a or b);
    layer3_outputs(7282) <= not b or a;
    layer3_outputs(7283) <= 1'b0;
    layer3_outputs(7284) <= not (a or b);
    layer3_outputs(7285) <= not (a xor b);
    layer3_outputs(7286) <= 1'b1;
    layer3_outputs(7287) <= not a;
    layer3_outputs(7288) <= not a or b;
    layer3_outputs(7289) <= not b;
    layer3_outputs(7290) <= not (a and b);
    layer3_outputs(7291) <= 1'b1;
    layer3_outputs(7292) <= 1'b0;
    layer3_outputs(7293) <= not (a or b);
    layer3_outputs(7294) <= not b or a;
    layer3_outputs(7295) <= b;
    layer3_outputs(7296) <= b and not a;
    layer3_outputs(7297) <= a or b;
    layer3_outputs(7298) <= not (a and b);
    layer3_outputs(7299) <= b;
    layer3_outputs(7300) <= a and b;
    layer3_outputs(7301) <= a;
    layer3_outputs(7302) <= not (a and b);
    layer3_outputs(7303) <= a;
    layer3_outputs(7304) <= 1'b1;
    layer3_outputs(7305) <= a xor b;
    layer3_outputs(7306) <= a or b;
    layer3_outputs(7307) <= not (a and b);
    layer3_outputs(7308) <= not b or a;
    layer3_outputs(7309) <= a and not b;
    layer3_outputs(7310) <= not (a or b);
    layer3_outputs(7311) <= not a;
    layer3_outputs(7312) <= not (a or b);
    layer3_outputs(7313) <= b;
    layer3_outputs(7314) <= a and not b;
    layer3_outputs(7315) <= b;
    layer3_outputs(7316) <= not (a or b);
    layer3_outputs(7317) <= not a;
    layer3_outputs(7318) <= a or b;
    layer3_outputs(7319) <= not b;
    layer3_outputs(7320) <= not b;
    layer3_outputs(7321) <= not b;
    layer3_outputs(7322) <= b;
    layer3_outputs(7323) <= not (a and b);
    layer3_outputs(7324) <= b and not a;
    layer3_outputs(7325) <= a and b;
    layer3_outputs(7326) <= 1'b0;
    layer3_outputs(7327) <= not b or a;
    layer3_outputs(7328) <= not b;
    layer3_outputs(7329) <= a;
    layer3_outputs(7330) <= not (a or b);
    layer3_outputs(7331) <= b and not a;
    layer3_outputs(7332) <= b and not a;
    layer3_outputs(7333) <= a or b;
    layer3_outputs(7334) <= a and not b;
    layer3_outputs(7335) <= a and not b;
    layer3_outputs(7336) <= not b;
    layer3_outputs(7337) <= b;
    layer3_outputs(7338) <= not a;
    layer3_outputs(7339) <= a xor b;
    layer3_outputs(7340) <= not b or a;
    layer3_outputs(7341) <= a and not b;
    layer3_outputs(7342) <= not b;
    layer3_outputs(7343) <= 1'b0;
    layer3_outputs(7344) <= not a or b;
    layer3_outputs(7345) <= not (a and b);
    layer3_outputs(7346) <= not (a and b);
    layer3_outputs(7347) <= not b;
    layer3_outputs(7348) <= 1'b0;
    layer3_outputs(7349) <= a;
    layer3_outputs(7350) <= a and b;
    layer3_outputs(7351) <= a or b;
    layer3_outputs(7352) <= 1'b1;
    layer3_outputs(7353) <= not a;
    layer3_outputs(7354) <= not b;
    layer3_outputs(7355) <= not a or b;
    layer3_outputs(7356) <= not (a and b);
    layer3_outputs(7357) <= 1'b0;
    layer3_outputs(7358) <= not b;
    layer3_outputs(7359) <= not b;
    layer3_outputs(7360) <= not b;
    layer3_outputs(7361) <= not a or b;
    layer3_outputs(7362) <= not (a or b);
    layer3_outputs(7363) <= b;
    layer3_outputs(7364) <= 1'b0;
    layer3_outputs(7365) <= not (a xor b);
    layer3_outputs(7366) <= not a or b;
    layer3_outputs(7367) <= not b;
    layer3_outputs(7368) <= not b;
    layer3_outputs(7369) <= not (a or b);
    layer3_outputs(7370) <= not (a and b);
    layer3_outputs(7371) <= a and not b;
    layer3_outputs(7372) <= not (a or b);
    layer3_outputs(7373) <= not b;
    layer3_outputs(7374) <= a and not b;
    layer3_outputs(7375) <= not a or b;
    layer3_outputs(7376) <= not b;
    layer3_outputs(7377) <= 1'b0;
    layer3_outputs(7378) <= a and b;
    layer3_outputs(7379) <= not (a and b);
    layer3_outputs(7380) <= not b;
    layer3_outputs(7381) <= not a or b;
    layer3_outputs(7382) <= not b;
    layer3_outputs(7383) <= not a or b;
    layer3_outputs(7384) <= b and not a;
    layer3_outputs(7385) <= a;
    layer3_outputs(7386) <= not (a or b);
    layer3_outputs(7387) <= 1'b1;
    layer3_outputs(7388) <= a or b;
    layer3_outputs(7389) <= not a;
    layer3_outputs(7390) <= not (a or b);
    layer3_outputs(7391) <= a;
    layer3_outputs(7392) <= b;
    layer3_outputs(7393) <= not a;
    layer3_outputs(7394) <= not b or a;
    layer3_outputs(7395) <= not (a or b);
    layer3_outputs(7396) <= 1'b0;
    layer3_outputs(7397) <= b;
    layer3_outputs(7398) <= a or b;
    layer3_outputs(7399) <= a or b;
    layer3_outputs(7400) <= not (a and b);
    layer3_outputs(7401) <= 1'b0;
    layer3_outputs(7402) <= 1'b1;
    layer3_outputs(7403) <= not b;
    layer3_outputs(7404) <= b;
    layer3_outputs(7405) <= a and b;
    layer3_outputs(7406) <= a;
    layer3_outputs(7407) <= a;
    layer3_outputs(7408) <= not a;
    layer3_outputs(7409) <= not a or b;
    layer3_outputs(7410) <= a or b;
    layer3_outputs(7411) <= b;
    layer3_outputs(7412) <= not (a or b);
    layer3_outputs(7413) <= a and not b;
    layer3_outputs(7414) <= b;
    layer3_outputs(7415) <= not b;
    layer3_outputs(7416) <= not (a or b);
    layer3_outputs(7417) <= not a;
    layer3_outputs(7418) <= not (a or b);
    layer3_outputs(7419) <= not a or b;
    layer3_outputs(7420) <= a;
    layer3_outputs(7421) <= a and not b;
    layer3_outputs(7422) <= 1'b0;
    layer3_outputs(7423) <= a and not b;
    layer3_outputs(7424) <= b and not a;
    layer3_outputs(7425) <= 1'b0;
    layer3_outputs(7426) <= a or b;
    layer3_outputs(7427) <= a and b;
    layer3_outputs(7428) <= not b;
    layer3_outputs(7429) <= 1'b1;
    layer3_outputs(7430) <= a or b;
    layer3_outputs(7431) <= b and not a;
    layer3_outputs(7432) <= a and not b;
    layer3_outputs(7433) <= not (a or b);
    layer3_outputs(7434) <= not (a or b);
    layer3_outputs(7435) <= a or b;
    layer3_outputs(7436) <= a or b;
    layer3_outputs(7437) <= not (a and b);
    layer3_outputs(7438) <= not (a and b);
    layer3_outputs(7439) <= b and not a;
    layer3_outputs(7440) <= a or b;
    layer3_outputs(7441) <= a and b;
    layer3_outputs(7442) <= a and not b;
    layer3_outputs(7443) <= 1'b0;
    layer3_outputs(7444) <= not (a or b);
    layer3_outputs(7445) <= not (a xor b);
    layer3_outputs(7446) <= not b;
    layer3_outputs(7447) <= b;
    layer3_outputs(7448) <= not (a xor b);
    layer3_outputs(7449) <= not a or b;
    layer3_outputs(7450) <= not (a or b);
    layer3_outputs(7451) <= not (a and b);
    layer3_outputs(7452) <= 1'b0;
    layer3_outputs(7453) <= not (a or b);
    layer3_outputs(7454) <= not a;
    layer3_outputs(7455) <= b and not a;
    layer3_outputs(7456) <= not (a and b);
    layer3_outputs(7457) <= a and not b;
    layer3_outputs(7458) <= a;
    layer3_outputs(7459) <= b and not a;
    layer3_outputs(7460) <= not (a xor b);
    layer3_outputs(7461) <= a and b;
    layer3_outputs(7462) <= b and not a;
    layer3_outputs(7463) <= not b;
    layer3_outputs(7464) <= 1'b0;
    layer3_outputs(7465) <= not a;
    layer3_outputs(7466) <= b;
    layer3_outputs(7467) <= a;
    layer3_outputs(7468) <= a;
    layer3_outputs(7469) <= not b or a;
    layer3_outputs(7470) <= not a or b;
    layer3_outputs(7471) <= a and b;
    layer3_outputs(7472) <= a xor b;
    layer3_outputs(7473) <= not b or a;
    layer3_outputs(7474) <= not b;
    layer3_outputs(7475) <= not a;
    layer3_outputs(7476) <= a or b;
    layer3_outputs(7477) <= 1'b1;
    layer3_outputs(7478) <= not b;
    layer3_outputs(7479) <= not b or a;
    layer3_outputs(7480) <= not b or a;
    layer3_outputs(7481) <= 1'b0;
    layer3_outputs(7482) <= b;
    layer3_outputs(7483) <= not (a or b);
    layer3_outputs(7484) <= a;
    layer3_outputs(7485) <= a and b;
    layer3_outputs(7486) <= a and not b;
    layer3_outputs(7487) <= a;
    layer3_outputs(7488) <= a and not b;
    layer3_outputs(7489) <= not (a or b);
    layer3_outputs(7490) <= not (a or b);
    layer3_outputs(7491) <= b;
    layer3_outputs(7492) <= not a;
    layer3_outputs(7493) <= not b;
    layer3_outputs(7494) <= 1'b0;
    layer3_outputs(7495) <= a or b;
    layer3_outputs(7496) <= not b;
    layer3_outputs(7497) <= not (a or b);
    layer3_outputs(7498) <= not (a xor b);
    layer3_outputs(7499) <= 1'b0;
    layer3_outputs(7500) <= a and b;
    layer3_outputs(7501) <= a or b;
    layer3_outputs(7502) <= not b;
    layer3_outputs(7503) <= a or b;
    layer3_outputs(7504) <= 1'b0;
    layer3_outputs(7505) <= b and not a;
    layer3_outputs(7506) <= 1'b1;
    layer3_outputs(7507) <= not b or a;
    layer3_outputs(7508) <= not a or b;
    layer3_outputs(7509) <= not (a xor b);
    layer3_outputs(7510) <= not (a and b);
    layer3_outputs(7511) <= a;
    layer3_outputs(7512) <= a and not b;
    layer3_outputs(7513) <= a;
    layer3_outputs(7514) <= a and not b;
    layer3_outputs(7515) <= b and not a;
    layer3_outputs(7516) <= not b;
    layer3_outputs(7517) <= b and not a;
    layer3_outputs(7518) <= a and b;
    layer3_outputs(7519) <= not a or b;
    layer3_outputs(7520) <= not a;
    layer3_outputs(7521) <= 1'b0;
    layer3_outputs(7522) <= not a or b;
    layer3_outputs(7523) <= not b or a;
    layer3_outputs(7524) <= not (a and b);
    layer3_outputs(7525) <= not (a xor b);
    layer3_outputs(7526) <= not b or a;
    layer3_outputs(7527) <= 1'b0;
    layer3_outputs(7528) <= b and not a;
    layer3_outputs(7529) <= not b;
    layer3_outputs(7530) <= b;
    layer3_outputs(7531) <= not (a or b);
    layer3_outputs(7532) <= b and not a;
    layer3_outputs(7533) <= not a;
    layer3_outputs(7534) <= 1'b1;
    layer3_outputs(7535) <= a and b;
    layer3_outputs(7536) <= not (a or b);
    layer3_outputs(7537) <= not (a and b);
    layer3_outputs(7538) <= not b;
    layer3_outputs(7539) <= a xor b;
    layer3_outputs(7540) <= not a or b;
    layer3_outputs(7541) <= 1'b1;
    layer3_outputs(7542) <= a;
    layer3_outputs(7543) <= not (a or b);
    layer3_outputs(7544) <= not b or a;
    layer3_outputs(7545) <= a and b;
    layer3_outputs(7546) <= not a;
    layer3_outputs(7547) <= not b;
    layer3_outputs(7548) <= a or b;
    layer3_outputs(7549) <= not a;
    layer3_outputs(7550) <= a;
    layer3_outputs(7551) <= not a or b;
    layer3_outputs(7552) <= 1'b1;
    layer3_outputs(7553) <= b;
    layer3_outputs(7554) <= b;
    layer3_outputs(7555) <= not b or a;
    layer3_outputs(7556) <= not (a or b);
    layer3_outputs(7557) <= not (a xor b);
    layer3_outputs(7558) <= not (a or b);
    layer3_outputs(7559) <= b and not a;
    layer3_outputs(7560) <= 1'b1;
    layer3_outputs(7561) <= not a;
    layer3_outputs(7562) <= a;
    layer3_outputs(7563) <= a and b;
    layer3_outputs(7564) <= b and not a;
    layer3_outputs(7565) <= a or b;
    layer3_outputs(7566) <= 1'b0;
    layer3_outputs(7567) <= not (a or b);
    layer3_outputs(7568) <= b;
    layer3_outputs(7569) <= a and b;
    layer3_outputs(7570) <= not b;
    layer3_outputs(7571) <= not (a and b);
    layer3_outputs(7572) <= not b or a;
    layer3_outputs(7573) <= a and not b;
    layer3_outputs(7574) <= a;
    layer3_outputs(7575) <= a;
    layer3_outputs(7576) <= b;
    layer3_outputs(7577) <= not b;
    layer3_outputs(7578) <= not a or b;
    layer3_outputs(7579) <= not b;
    layer3_outputs(7580) <= not b or a;
    layer3_outputs(7581) <= not (a or b);
    layer3_outputs(7582) <= 1'b1;
    layer3_outputs(7583) <= a or b;
    layer3_outputs(7584) <= 1'b0;
    layer3_outputs(7585) <= not (a or b);
    layer3_outputs(7586) <= a and not b;
    layer3_outputs(7587) <= not b or a;
    layer3_outputs(7588) <= 1'b0;
    layer3_outputs(7589) <= not (a and b);
    layer3_outputs(7590) <= a or b;
    layer3_outputs(7591) <= not a or b;
    layer3_outputs(7592) <= a;
    layer3_outputs(7593) <= a;
    layer3_outputs(7594) <= b;
    layer3_outputs(7595) <= a;
    layer3_outputs(7596) <= not (a and b);
    layer3_outputs(7597) <= 1'b1;
    layer3_outputs(7598) <= not (a or b);
    layer3_outputs(7599) <= a or b;
    layer3_outputs(7600) <= not b;
    layer3_outputs(7601) <= not (a xor b);
    layer3_outputs(7602) <= a and not b;
    layer3_outputs(7603) <= not (a or b);
    layer3_outputs(7604) <= b;
    layer3_outputs(7605) <= a;
    layer3_outputs(7606) <= not b or a;
    layer3_outputs(7607) <= not (a xor b);
    layer3_outputs(7608) <= b and not a;
    layer3_outputs(7609) <= b;
    layer3_outputs(7610) <= not b;
    layer3_outputs(7611) <= 1'b1;
    layer3_outputs(7612) <= not b;
    layer3_outputs(7613) <= a;
    layer3_outputs(7614) <= not (a or b);
    layer3_outputs(7615) <= not b or a;
    layer3_outputs(7616) <= a or b;
    layer3_outputs(7617) <= 1'b1;
    layer3_outputs(7618) <= 1'b0;
    layer3_outputs(7619) <= 1'b0;
    layer3_outputs(7620) <= 1'b0;
    layer3_outputs(7621) <= 1'b0;
    layer3_outputs(7622) <= 1'b0;
    layer3_outputs(7623) <= not a or b;
    layer3_outputs(7624) <= b and not a;
    layer3_outputs(7625) <= b;
    layer3_outputs(7626) <= not (a and b);
    layer3_outputs(7627) <= a and not b;
    layer3_outputs(7628) <= b and not a;
    layer3_outputs(7629) <= not b;
    layer3_outputs(7630) <= a or b;
    layer3_outputs(7631) <= not b;
    layer3_outputs(7632) <= 1'b0;
    layer3_outputs(7633) <= not b or a;
    layer3_outputs(7634) <= not (a or b);
    layer3_outputs(7635) <= b;
    layer3_outputs(7636) <= not b or a;
    layer3_outputs(7637) <= a;
    layer3_outputs(7638) <= a xor b;
    layer3_outputs(7639) <= a;
    layer3_outputs(7640) <= not b or a;
    layer3_outputs(7641) <= a and b;
    layer3_outputs(7642) <= 1'b1;
    layer3_outputs(7643) <= not (a or b);
    layer3_outputs(7644) <= a or b;
    layer3_outputs(7645) <= 1'b1;
    layer3_outputs(7646) <= a or b;
    layer3_outputs(7647) <= a and not b;
    layer3_outputs(7648) <= not b or a;
    layer3_outputs(7649) <= a and b;
    layer3_outputs(7650) <= not (a xor b);
    layer3_outputs(7651) <= not b or a;
    layer3_outputs(7652) <= not b;
    layer3_outputs(7653) <= not a or b;
    layer3_outputs(7654) <= 1'b1;
    layer3_outputs(7655) <= a and not b;
    layer3_outputs(7656) <= a or b;
    layer3_outputs(7657) <= 1'b1;
    layer3_outputs(7658) <= b;
    layer3_outputs(7659) <= a or b;
    layer3_outputs(7660) <= a or b;
    layer3_outputs(7661) <= not (a or b);
    layer3_outputs(7662) <= not b;
    layer3_outputs(7663) <= a;
    layer3_outputs(7664) <= not b;
    layer3_outputs(7665) <= not a;
    layer3_outputs(7666) <= a and not b;
    layer3_outputs(7667) <= 1'b0;
    layer3_outputs(7668) <= a and not b;
    layer3_outputs(7669) <= a;
    layer3_outputs(7670) <= a and b;
    layer3_outputs(7671) <= b;
    layer3_outputs(7672) <= 1'b1;
    layer3_outputs(7673) <= a and not b;
    layer3_outputs(7674) <= b;
    layer3_outputs(7675) <= not (a or b);
    layer3_outputs(7676) <= 1'b0;
    layer3_outputs(7677) <= not b;
    layer3_outputs(7678) <= a and not b;
    layer3_outputs(7679) <= not (a and b);
    layer3_outputs(7680) <= a and b;
    layer3_outputs(7681) <= not (a or b);
    layer3_outputs(7682) <= a;
    layer3_outputs(7683) <= not a;
    layer3_outputs(7684) <= b and not a;
    layer3_outputs(7685) <= a and not b;
    layer3_outputs(7686) <= a;
    layer3_outputs(7687) <= 1'b0;
    layer3_outputs(7688) <= a and b;
    layer3_outputs(7689) <= not a or b;
    layer3_outputs(7690) <= not (a and b);
    layer3_outputs(7691) <= not a;
    layer3_outputs(7692) <= a;
    layer3_outputs(7693) <= not (a or b);
    layer3_outputs(7694) <= 1'b1;
    layer3_outputs(7695) <= not a or b;
    layer3_outputs(7696) <= 1'b0;
    layer3_outputs(7697) <= not b;
    layer3_outputs(7698) <= not (a or b);
    layer3_outputs(7699) <= not b or a;
    layer3_outputs(7700) <= not (a and b);
    layer3_outputs(7701) <= a and b;
    layer3_outputs(7702) <= 1'b0;
    layer3_outputs(7703) <= a and b;
    layer3_outputs(7704) <= 1'b0;
    layer3_outputs(7705) <= a xor b;
    layer3_outputs(7706) <= b and not a;
    layer3_outputs(7707) <= not b or a;
    layer3_outputs(7708) <= a and b;
    layer3_outputs(7709) <= a or b;
    layer3_outputs(7710) <= not a or b;
    layer3_outputs(7711) <= 1'b1;
    layer3_outputs(7712) <= not (a or b);
    layer3_outputs(7713) <= not (a xor b);
    layer3_outputs(7714) <= not (a and b);
    layer3_outputs(7715) <= not a;
    layer3_outputs(7716) <= b;
    layer3_outputs(7717) <= 1'b1;
    layer3_outputs(7718) <= not (a or b);
    layer3_outputs(7719) <= a and b;
    layer3_outputs(7720) <= b;
    layer3_outputs(7721) <= b;
    layer3_outputs(7722) <= not (a or b);
    layer3_outputs(7723) <= b;
    layer3_outputs(7724) <= not b;
    layer3_outputs(7725) <= b;
    layer3_outputs(7726) <= not a;
    layer3_outputs(7727) <= b;
    layer3_outputs(7728) <= not b or a;
    layer3_outputs(7729) <= b;
    layer3_outputs(7730) <= a and b;
    layer3_outputs(7731) <= not (a and b);
    layer3_outputs(7732) <= not b;
    layer3_outputs(7733) <= a;
    layer3_outputs(7734) <= b and not a;
    layer3_outputs(7735) <= 1'b0;
    layer3_outputs(7736) <= not (a and b);
    layer3_outputs(7737) <= not (a and b);
    layer3_outputs(7738) <= a and b;
    layer3_outputs(7739) <= a or b;
    layer3_outputs(7740) <= a;
    layer3_outputs(7741) <= a and not b;
    layer3_outputs(7742) <= not a;
    layer3_outputs(7743) <= not a or b;
    layer3_outputs(7744) <= a and b;
    layer3_outputs(7745) <= a and not b;
    layer3_outputs(7746) <= not a;
    layer3_outputs(7747) <= b;
    layer3_outputs(7748) <= 1'b0;
    layer3_outputs(7749) <= not a;
    layer3_outputs(7750) <= not b or a;
    layer3_outputs(7751) <= b and not a;
    layer3_outputs(7752) <= a xor b;
    layer3_outputs(7753) <= a or b;
    layer3_outputs(7754) <= not a;
    layer3_outputs(7755) <= b and not a;
    layer3_outputs(7756) <= a xor b;
    layer3_outputs(7757) <= 1'b1;
    layer3_outputs(7758) <= not b;
    layer3_outputs(7759) <= b;
    layer3_outputs(7760) <= a and not b;
    layer3_outputs(7761) <= not b;
    layer3_outputs(7762) <= a and not b;
    layer3_outputs(7763) <= a and not b;
    layer3_outputs(7764) <= b and not a;
    layer3_outputs(7765) <= not b or a;
    layer3_outputs(7766) <= b;
    layer3_outputs(7767) <= a xor b;
    layer3_outputs(7768) <= not b;
    layer3_outputs(7769) <= a or b;
    layer3_outputs(7770) <= 1'b1;
    layer3_outputs(7771) <= a;
    layer3_outputs(7772) <= b;
    layer3_outputs(7773) <= not a or b;
    layer3_outputs(7774) <= not (a and b);
    layer3_outputs(7775) <= not (a xor b);
    layer3_outputs(7776) <= a;
    layer3_outputs(7777) <= a or b;
    layer3_outputs(7778) <= not a;
    layer3_outputs(7779) <= b;
    layer3_outputs(7780) <= b and not a;
    layer3_outputs(7781) <= 1'b1;
    layer3_outputs(7782) <= not a;
    layer3_outputs(7783) <= not (a and b);
    layer3_outputs(7784) <= a and not b;
    layer3_outputs(7785) <= 1'b1;
    layer3_outputs(7786) <= a xor b;
    layer3_outputs(7787) <= b and not a;
    layer3_outputs(7788) <= not a;
    layer3_outputs(7789) <= 1'b0;
    layer3_outputs(7790) <= a;
    layer3_outputs(7791) <= not (a and b);
    layer3_outputs(7792) <= not b;
    layer3_outputs(7793) <= 1'b0;
    layer3_outputs(7794) <= not a or b;
    layer3_outputs(7795) <= a;
    layer3_outputs(7796) <= 1'b1;
    layer3_outputs(7797) <= not (a or b);
    layer3_outputs(7798) <= a and not b;
    layer3_outputs(7799) <= not b or a;
    layer3_outputs(7800) <= a and b;
    layer3_outputs(7801) <= a or b;
    layer3_outputs(7802) <= not a or b;
    layer3_outputs(7803) <= a or b;
    layer3_outputs(7804) <= not b;
    layer3_outputs(7805) <= a;
    layer3_outputs(7806) <= a and b;
    layer3_outputs(7807) <= not a or b;
    layer3_outputs(7808) <= a and not b;
    layer3_outputs(7809) <= b;
    layer3_outputs(7810) <= not a;
    layer3_outputs(7811) <= not a;
    layer3_outputs(7812) <= a and not b;
    layer3_outputs(7813) <= not b or a;
    layer3_outputs(7814) <= not b or a;
    layer3_outputs(7815) <= 1'b0;
    layer3_outputs(7816) <= not (a and b);
    layer3_outputs(7817) <= not (a and b);
    layer3_outputs(7818) <= not b or a;
    layer3_outputs(7819) <= b and not a;
    layer3_outputs(7820) <= not a;
    layer3_outputs(7821) <= b;
    layer3_outputs(7822) <= b;
    layer3_outputs(7823) <= 1'b0;
    layer3_outputs(7824) <= not (a or b);
    layer3_outputs(7825) <= 1'b1;
    layer3_outputs(7826) <= not (a and b);
    layer3_outputs(7827) <= not b;
    layer3_outputs(7828) <= not (a and b);
    layer3_outputs(7829) <= a;
    layer3_outputs(7830) <= a;
    layer3_outputs(7831) <= 1'b0;
    layer3_outputs(7832) <= not (a and b);
    layer3_outputs(7833) <= not a;
    layer3_outputs(7834) <= a and b;
    layer3_outputs(7835) <= a and not b;
    layer3_outputs(7836) <= b;
    layer3_outputs(7837) <= a and not b;
    layer3_outputs(7838) <= a and b;
    layer3_outputs(7839) <= 1'b0;
    layer3_outputs(7840) <= a and b;
    layer3_outputs(7841) <= a and not b;
    layer3_outputs(7842) <= 1'b1;
    layer3_outputs(7843) <= a and b;
    layer3_outputs(7844) <= a;
    layer3_outputs(7845) <= a and not b;
    layer3_outputs(7846) <= a and b;
    layer3_outputs(7847) <= 1'b1;
    layer3_outputs(7848) <= not b;
    layer3_outputs(7849) <= b;
    layer3_outputs(7850) <= a and not b;
    layer3_outputs(7851) <= not (a or b);
    layer3_outputs(7852) <= not b or a;
    layer3_outputs(7853) <= a and b;
    layer3_outputs(7854) <= not a or b;
    layer3_outputs(7855) <= a xor b;
    layer3_outputs(7856) <= b and not a;
    layer3_outputs(7857) <= not a;
    layer3_outputs(7858) <= not a;
    layer3_outputs(7859) <= not (a and b);
    layer3_outputs(7860) <= a;
    layer3_outputs(7861) <= a and not b;
    layer3_outputs(7862) <= a;
    layer3_outputs(7863) <= not (a or b);
    layer3_outputs(7864) <= 1'b0;
    layer3_outputs(7865) <= a and not b;
    layer3_outputs(7866) <= not a;
    layer3_outputs(7867) <= a;
    layer3_outputs(7868) <= not a or b;
    layer3_outputs(7869) <= not b or a;
    layer3_outputs(7870) <= a and not b;
    layer3_outputs(7871) <= 1'b0;
    layer3_outputs(7872) <= 1'b0;
    layer3_outputs(7873) <= a or b;
    layer3_outputs(7874) <= b;
    layer3_outputs(7875) <= a and not b;
    layer3_outputs(7876) <= 1'b1;
    layer3_outputs(7877) <= not (a or b);
    layer3_outputs(7878) <= a;
    layer3_outputs(7879) <= a or b;
    layer3_outputs(7880) <= a and b;
    layer3_outputs(7881) <= 1'b0;
    layer3_outputs(7882) <= b;
    layer3_outputs(7883) <= b and not a;
    layer3_outputs(7884) <= b and not a;
    layer3_outputs(7885) <= a and b;
    layer3_outputs(7886) <= not (a or b);
    layer3_outputs(7887) <= a and b;
    layer3_outputs(7888) <= not a or b;
    layer3_outputs(7889) <= not a;
    layer3_outputs(7890) <= 1'b0;
    layer3_outputs(7891) <= not (a and b);
    layer3_outputs(7892) <= b;
    layer3_outputs(7893) <= a and not b;
    layer3_outputs(7894) <= a;
    layer3_outputs(7895) <= a;
    layer3_outputs(7896) <= not b;
    layer3_outputs(7897) <= a and not b;
    layer3_outputs(7898) <= not (a and b);
    layer3_outputs(7899) <= not a;
    layer3_outputs(7900) <= a;
    layer3_outputs(7901) <= a and not b;
    layer3_outputs(7902) <= not a;
    layer3_outputs(7903) <= 1'b0;
    layer3_outputs(7904) <= a;
    layer3_outputs(7905) <= b;
    layer3_outputs(7906) <= not b or a;
    layer3_outputs(7907) <= 1'b1;
    layer3_outputs(7908) <= not (a and b);
    layer3_outputs(7909) <= not a;
    layer3_outputs(7910) <= not (a or b);
    layer3_outputs(7911) <= 1'b1;
    layer3_outputs(7912) <= b;
    layer3_outputs(7913) <= b and not a;
    layer3_outputs(7914) <= a;
    layer3_outputs(7915) <= not (a and b);
    layer3_outputs(7916) <= a and not b;
    layer3_outputs(7917) <= a xor b;
    layer3_outputs(7918) <= not a;
    layer3_outputs(7919) <= not (a and b);
    layer3_outputs(7920) <= not a or b;
    layer3_outputs(7921) <= a and b;
    layer3_outputs(7922) <= a;
    layer3_outputs(7923) <= a or b;
    layer3_outputs(7924) <= a or b;
    layer3_outputs(7925) <= not a;
    layer3_outputs(7926) <= not a or b;
    layer3_outputs(7927) <= not b or a;
    layer3_outputs(7928) <= b;
    layer3_outputs(7929) <= a xor b;
    layer3_outputs(7930) <= a or b;
    layer3_outputs(7931) <= a and not b;
    layer3_outputs(7932) <= 1'b1;
    layer3_outputs(7933) <= not (a and b);
    layer3_outputs(7934) <= a or b;
    layer3_outputs(7935) <= not (a xor b);
    layer3_outputs(7936) <= a and b;
    layer3_outputs(7937) <= a;
    layer3_outputs(7938) <= a and not b;
    layer3_outputs(7939) <= 1'b0;
    layer3_outputs(7940) <= b and not a;
    layer3_outputs(7941) <= 1'b1;
    layer3_outputs(7942) <= b and not a;
    layer3_outputs(7943) <= b and not a;
    layer3_outputs(7944) <= 1'b0;
    layer3_outputs(7945) <= a and b;
    layer3_outputs(7946) <= 1'b0;
    layer3_outputs(7947) <= b;
    layer3_outputs(7948) <= not (a or b);
    layer3_outputs(7949) <= not a or b;
    layer3_outputs(7950) <= not (a and b);
    layer3_outputs(7951) <= 1'b0;
    layer3_outputs(7952) <= not (a or b);
    layer3_outputs(7953) <= 1'b0;
    layer3_outputs(7954) <= not b;
    layer3_outputs(7955) <= not b;
    layer3_outputs(7956) <= 1'b1;
    layer3_outputs(7957) <= a and not b;
    layer3_outputs(7958) <= 1'b1;
    layer3_outputs(7959) <= 1'b0;
    layer3_outputs(7960) <= 1'b0;
    layer3_outputs(7961) <= not (a and b);
    layer3_outputs(7962) <= not (a or b);
    layer3_outputs(7963) <= not a or b;
    layer3_outputs(7964) <= a and not b;
    layer3_outputs(7965) <= 1'b1;
    layer3_outputs(7966) <= not a or b;
    layer3_outputs(7967) <= not a or b;
    layer3_outputs(7968) <= not b or a;
    layer3_outputs(7969) <= 1'b1;
    layer3_outputs(7970) <= not a;
    layer3_outputs(7971) <= not (a and b);
    layer3_outputs(7972) <= a and not b;
    layer3_outputs(7973) <= not a or b;
    layer3_outputs(7974) <= a and b;
    layer3_outputs(7975) <= not (a or b);
    layer3_outputs(7976) <= not (a and b);
    layer3_outputs(7977) <= not b or a;
    layer3_outputs(7978) <= a and not b;
    layer3_outputs(7979) <= not (a and b);
    layer3_outputs(7980) <= not (a and b);
    layer3_outputs(7981) <= 1'b1;
    layer3_outputs(7982) <= a or b;
    layer3_outputs(7983) <= not b or a;
    layer3_outputs(7984) <= b;
    layer3_outputs(7985) <= 1'b0;
    layer3_outputs(7986) <= not a;
    layer3_outputs(7987) <= a;
    layer3_outputs(7988) <= b;
    layer3_outputs(7989) <= not (a and b);
    layer3_outputs(7990) <= b and not a;
    layer3_outputs(7991) <= not (a or b);
    layer3_outputs(7992) <= not (a or b);
    layer3_outputs(7993) <= not (a or b);
    layer3_outputs(7994) <= not b or a;
    layer3_outputs(7995) <= 1'b0;
    layer3_outputs(7996) <= 1'b0;
    layer3_outputs(7997) <= not a;
    layer3_outputs(7998) <= not b;
    layer3_outputs(7999) <= a;
    layer3_outputs(8000) <= not a;
    layer3_outputs(8001) <= 1'b0;
    layer3_outputs(8002) <= a and not b;
    layer3_outputs(8003) <= a;
    layer3_outputs(8004) <= a or b;
    layer3_outputs(8005) <= a;
    layer3_outputs(8006) <= not (a and b);
    layer3_outputs(8007) <= not b;
    layer3_outputs(8008) <= 1'b0;
    layer3_outputs(8009) <= not (a or b);
    layer3_outputs(8010) <= not a or b;
    layer3_outputs(8011) <= not a or b;
    layer3_outputs(8012) <= not (a and b);
    layer3_outputs(8013) <= not b or a;
    layer3_outputs(8014) <= b;
    layer3_outputs(8015) <= not b or a;
    layer3_outputs(8016) <= not a or b;
    layer3_outputs(8017) <= a or b;
    layer3_outputs(8018) <= b;
    layer3_outputs(8019) <= a and not b;
    layer3_outputs(8020) <= 1'b1;
    layer3_outputs(8021) <= not (a or b);
    layer3_outputs(8022) <= not (a or b);
    layer3_outputs(8023) <= b;
    layer3_outputs(8024) <= a;
    layer3_outputs(8025) <= not (a or b);
    layer3_outputs(8026) <= not (a or b);
    layer3_outputs(8027) <= not b or a;
    layer3_outputs(8028) <= not (a and b);
    layer3_outputs(8029) <= a or b;
    layer3_outputs(8030) <= a or b;
    layer3_outputs(8031) <= not b;
    layer3_outputs(8032) <= a;
    layer3_outputs(8033) <= a or b;
    layer3_outputs(8034) <= not b or a;
    layer3_outputs(8035) <= not b or a;
    layer3_outputs(8036) <= not a or b;
    layer3_outputs(8037) <= a or b;
    layer3_outputs(8038) <= b;
    layer3_outputs(8039) <= not b or a;
    layer3_outputs(8040) <= 1'b0;
    layer3_outputs(8041) <= b and not a;
    layer3_outputs(8042) <= not (a xor b);
    layer3_outputs(8043) <= 1'b0;
    layer3_outputs(8044) <= not b or a;
    layer3_outputs(8045) <= not (a and b);
    layer3_outputs(8046) <= not (a and b);
    layer3_outputs(8047) <= 1'b1;
    layer3_outputs(8048) <= a and b;
    layer3_outputs(8049) <= a;
    layer3_outputs(8050) <= b and not a;
    layer3_outputs(8051) <= a and not b;
    layer3_outputs(8052) <= not b or a;
    layer3_outputs(8053) <= a and not b;
    layer3_outputs(8054) <= a;
    layer3_outputs(8055) <= not a;
    layer3_outputs(8056) <= not b or a;
    layer3_outputs(8057) <= 1'b0;
    layer3_outputs(8058) <= b and not a;
    layer3_outputs(8059) <= not (a or b);
    layer3_outputs(8060) <= not b;
    layer3_outputs(8061) <= a and not b;
    layer3_outputs(8062) <= 1'b0;
    layer3_outputs(8063) <= 1'b1;
    layer3_outputs(8064) <= 1'b0;
    layer3_outputs(8065) <= a and not b;
    layer3_outputs(8066) <= not b or a;
    layer3_outputs(8067) <= a and not b;
    layer3_outputs(8068) <= b;
    layer3_outputs(8069) <= 1'b1;
    layer3_outputs(8070) <= 1'b1;
    layer3_outputs(8071) <= not a;
    layer3_outputs(8072) <= not (a xor b);
    layer3_outputs(8073) <= 1'b0;
    layer3_outputs(8074) <= b;
    layer3_outputs(8075) <= not (a or b);
    layer3_outputs(8076) <= a;
    layer3_outputs(8077) <= a;
    layer3_outputs(8078) <= a and not b;
    layer3_outputs(8079) <= b;
    layer3_outputs(8080) <= not (a or b);
    layer3_outputs(8081) <= a and not b;
    layer3_outputs(8082) <= a and not b;
    layer3_outputs(8083) <= 1'b1;
    layer3_outputs(8084) <= not (a xor b);
    layer3_outputs(8085) <= a or b;
    layer3_outputs(8086) <= not a or b;
    layer3_outputs(8087) <= not b or a;
    layer3_outputs(8088) <= not (a or b);
    layer3_outputs(8089) <= not (a and b);
    layer3_outputs(8090) <= not (a or b);
    layer3_outputs(8091) <= b and not a;
    layer3_outputs(8092) <= 1'b0;
    layer3_outputs(8093) <= not b or a;
    layer3_outputs(8094) <= a and b;
    layer3_outputs(8095) <= not a;
    layer3_outputs(8096) <= not (a or b);
    layer3_outputs(8097) <= 1'b1;
    layer3_outputs(8098) <= not a;
    layer3_outputs(8099) <= 1'b1;
    layer3_outputs(8100) <= not b;
    layer3_outputs(8101) <= b;
    layer3_outputs(8102) <= not b;
    layer3_outputs(8103) <= a;
    layer3_outputs(8104) <= a xor b;
    layer3_outputs(8105) <= a and not b;
    layer3_outputs(8106) <= 1'b0;
    layer3_outputs(8107) <= 1'b0;
    layer3_outputs(8108) <= not b;
    layer3_outputs(8109) <= b;
    layer3_outputs(8110) <= not (a xor b);
    layer3_outputs(8111) <= a or b;
    layer3_outputs(8112) <= not b or a;
    layer3_outputs(8113) <= not b;
    layer3_outputs(8114) <= not b;
    layer3_outputs(8115) <= not a;
    layer3_outputs(8116) <= a and not b;
    layer3_outputs(8117) <= not b or a;
    layer3_outputs(8118) <= 1'b1;
    layer3_outputs(8119) <= a;
    layer3_outputs(8120) <= 1'b1;
    layer3_outputs(8121) <= not b or a;
    layer3_outputs(8122) <= a and not b;
    layer3_outputs(8123) <= a and not b;
    layer3_outputs(8124) <= not (a and b);
    layer3_outputs(8125) <= not a;
    layer3_outputs(8126) <= 1'b0;
    layer3_outputs(8127) <= a or b;
    layer3_outputs(8128) <= not b or a;
    layer3_outputs(8129) <= a;
    layer3_outputs(8130) <= not (a and b);
    layer3_outputs(8131) <= b;
    layer3_outputs(8132) <= b;
    layer3_outputs(8133) <= b;
    layer3_outputs(8134) <= not (a or b);
    layer3_outputs(8135) <= a and not b;
    layer3_outputs(8136) <= not a;
    layer3_outputs(8137) <= not (a or b);
    layer3_outputs(8138) <= a and b;
    layer3_outputs(8139) <= b;
    layer3_outputs(8140) <= 1'b1;
    layer3_outputs(8141) <= not (a or b);
    layer3_outputs(8142) <= b and not a;
    layer3_outputs(8143) <= not b or a;
    layer3_outputs(8144) <= not (a or b);
    layer3_outputs(8145) <= not (a and b);
    layer3_outputs(8146) <= 1'b0;
    layer3_outputs(8147) <= a and b;
    layer3_outputs(8148) <= 1'b0;
    layer3_outputs(8149) <= b and not a;
    layer3_outputs(8150) <= b;
    layer3_outputs(8151) <= not b;
    layer3_outputs(8152) <= not (a and b);
    layer3_outputs(8153) <= not (a or b);
    layer3_outputs(8154) <= not a;
    layer3_outputs(8155) <= not b or a;
    layer3_outputs(8156) <= 1'b0;
    layer3_outputs(8157) <= not b or a;
    layer3_outputs(8158) <= a;
    layer3_outputs(8159) <= not a or b;
    layer3_outputs(8160) <= a and not b;
    layer3_outputs(8161) <= not (a xor b);
    layer3_outputs(8162) <= not a;
    layer3_outputs(8163) <= not b;
    layer3_outputs(8164) <= 1'b1;
    layer3_outputs(8165) <= not (a and b);
    layer3_outputs(8166) <= not (a or b);
    layer3_outputs(8167) <= not b;
    layer3_outputs(8168) <= 1'b0;
    layer3_outputs(8169) <= a;
    layer3_outputs(8170) <= a and not b;
    layer3_outputs(8171) <= a and not b;
    layer3_outputs(8172) <= not (a xor b);
    layer3_outputs(8173) <= a or b;
    layer3_outputs(8174) <= not b or a;
    layer3_outputs(8175) <= 1'b0;
    layer3_outputs(8176) <= a and b;
    layer3_outputs(8177) <= not b;
    layer3_outputs(8178) <= 1'b0;
    layer3_outputs(8179) <= not (a and b);
    layer3_outputs(8180) <= not a;
    layer3_outputs(8181) <= a;
    layer3_outputs(8182) <= a and not b;
    layer3_outputs(8183) <= not b or a;
    layer3_outputs(8184) <= a or b;
    layer3_outputs(8185) <= not a or b;
    layer3_outputs(8186) <= not (a and b);
    layer3_outputs(8187) <= 1'b0;
    layer3_outputs(8188) <= not b or a;
    layer3_outputs(8189) <= a and b;
    layer3_outputs(8190) <= 1'b1;
    layer3_outputs(8191) <= not b or a;
    layer3_outputs(8192) <= not a or b;
    layer3_outputs(8193) <= a and not b;
    layer3_outputs(8194) <= not a or b;
    layer3_outputs(8195) <= not b;
    layer3_outputs(8196) <= not a;
    layer3_outputs(8197) <= b;
    layer3_outputs(8198) <= b and not a;
    layer3_outputs(8199) <= a and b;
    layer3_outputs(8200) <= a or b;
    layer3_outputs(8201) <= a and b;
    layer3_outputs(8202) <= a and not b;
    layer3_outputs(8203) <= 1'b1;
    layer3_outputs(8204) <= not a or b;
    layer3_outputs(8205) <= not b;
    layer3_outputs(8206) <= b and not a;
    layer3_outputs(8207) <= not (a or b);
    layer3_outputs(8208) <= not b;
    layer3_outputs(8209) <= 1'b1;
    layer3_outputs(8210) <= not a;
    layer3_outputs(8211) <= 1'b1;
    layer3_outputs(8212) <= 1'b1;
    layer3_outputs(8213) <= not a or b;
    layer3_outputs(8214) <= a and not b;
    layer3_outputs(8215) <= not a;
    layer3_outputs(8216) <= a and b;
    layer3_outputs(8217) <= b;
    layer3_outputs(8218) <= b;
    layer3_outputs(8219) <= 1'b0;
    layer3_outputs(8220) <= b;
    layer3_outputs(8221) <= not b;
    layer3_outputs(8222) <= not (a xor b);
    layer3_outputs(8223) <= a and not b;
    layer3_outputs(8224) <= b;
    layer3_outputs(8225) <= not (a or b);
    layer3_outputs(8226) <= not (a or b);
    layer3_outputs(8227) <= 1'b0;
    layer3_outputs(8228) <= not a;
    layer3_outputs(8229) <= b;
    layer3_outputs(8230) <= not a;
    layer3_outputs(8231) <= not a or b;
    layer3_outputs(8232) <= not a or b;
    layer3_outputs(8233) <= a or b;
    layer3_outputs(8234) <= a xor b;
    layer3_outputs(8235) <= a and not b;
    layer3_outputs(8236) <= not (a or b);
    layer3_outputs(8237) <= b;
    layer3_outputs(8238) <= b and not a;
    layer3_outputs(8239) <= not (a or b);
    layer3_outputs(8240) <= a and b;
    layer3_outputs(8241) <= not (a xor b);
    layer3_outputs(8242) <= a and b;
    layer3_outputs(8243) <= a;
    layer3_outputs(8244) <= 1'b1;
    layer3_outputs(8245) <= a;
    layer3_outputs(8246) <= not (a xor b);
    layer3_outputs(8247) <= b;
    layer3_outputs(8248) <= 1'b0;
    layer3_outputs(8249) <= not (a xor b);
    layer3_outputs(8250) <= a and b;
    layer3_outputs(8251) <= not a;
    layer3_outputs(8252) <= a or b;
    layer3_outputs(8253) <= not b;
    layer3_outputs(8254) <= a and not b;
    layer3_outputs(8255) <= not (a and b);
    layer3_outputs(8256) <= not a or b;
    layer3_outputs(8257) <= not b;
    layer3_outputs(8258) <= not a or b;
    layer3_outputs(8259) <= a and not b;
    layer3_outputs(8260) <= not b;
    layer3_outputs(8261) <= a and b;
    layer3_outputs(8262) <= not b or a;
    layer3_outputs(8263) <= b and not a;
    layer3_outputs(8264) <= not (a and b);
    layer3_outputs(8265) <= not (a and b);
    layer3_outputs(8266) <= a and b;
    layer3_outputs(8267) <= not a;
    layer3_outputs(8268) <= a and b;
    layer3_outputs(8269) <= 1'b1;
    layer3_outputs(8270) <= not b or a;
    layer3_outputs(8271) <= not a;
    layer3_outputs(8272) <= not (a or b);
    layer3_outputs(8273) <= not (a or b);
    layer3_outputs(8274) <= not (a or b);
    layer3_outputs(8275) <= a xor b;
    layer3_outputs(8276) <= a;
    layer3_outputs(8277) <= not a;
    layer3_outputs(8278) <= b and not a;
    layer3_outputs(8279) <= a or b;
    layer3_outputs(8280) <= 1'b0;
    layer3_outputs(8281) <= a;
    layer3_outputs(8282) <= 1'b1;
    layer3_outputs(8283) <= a;
    layer3_outputs(8284) <= not a;
    layer3_outputs(8285) <= not b or a;
    layer3_outputs(8286) <= a and not b;
    layer3_outputs(8287) <= not b or a;
    layer3_outputs(8288) <= 1'b1;
    layer3_outputs(8289) <= not a;
    layer3_outputs(8290) <= a and b;
    layer3_outputs(8291) <= b and not a;
    layer3_outputs(8292) <= not a or b;
    layer3_outputs(8293) <= a and b;
    layer3_outputs(8294) <= not (a or b);
    layer3_outputs(8295) <= 1'b0;
    layer3_outputs(8296) <= b and not a;
    layer3_outputs(8297) <= b and not a;
    layer3_outputs(8298) <= b;
    layer3_outputs(8299) <= not (a or b);
    layer3_outputs(8300) <= not a;
    layer3_outputs(8301) <= not (a and b);
    layer3_outputs(8302) <= not a;
    layer3_outputs(8303) <= 1'b0;
    layer3_outputs(8304) <= not (a or b);
    layer3_outputs(8305) <= b and not a;
    layer3_outputs(8306) <= not (a or b);
    layer3_outputs(8307) <= b;
    layer3_outputs(8308) <= b;
    layer3_outputs(8309) <= not (a and b);
    layer3_outputs(8310) <= not b or a;
    layer3_outputs(8311) <= a;
    layer3_outputs(8312) <= 1'b0;
    layer3_outputs(8313) <= not (a xor b);
    layer3_outputs(8314) <= a and not b;
    layer3_outputs(8315) <= 1'b1;
    layer3_outputs(8316) <= not a;
    layer3_outputs(8317) <= 1'b0;
    layer3_outputs(8318) <= a and b;
    layer3_outputs(8319) <= not a or b;
    layer3_outputs(8320) <= 1'b1;
    layer3_outputs(8321) <= 1'b0;
    layer3_outputs(8322) <= not b or a;
    layer3_outputs(8323) <= not (a and b);
    layer3_outputs(8324) <= 1'b0;
    layer3_outputs(8325) <= not a or b;
    layer3_outputs(8326) <= not b;
    layer3_outputs(8327) <= a and not b;
    layer3_outputs(8328) <= 1'b0;
    layer3_outputs(8329) <= b;
    layer3_outputs(8330) <= a;
    layer3_outputs(8331) <= a;
    layer3_outputs(8332) <= not b;
    layer3_outputs(8333) <= not a or b;
    layer3_outputs(8334) <= not b or a;
    layer3_outputs(8335) <= a and b;
    layer3_outputs(8336) <= a or b;
    layer3_outputs(8337) <= not (a and b);
    layer3_outputs(8338) <= a xor b;
    layer3_outputs(8339) <= not b;
    layer3_outputs(8340) <= a and not b;
    layer3_outputs(8341) <= a or b;
    layer3_outputs(8342) <= a;
    layer3_outputs(8343) <= a and b;
    layer3_outputs(8344) <= a and b;
    layer3_outputs(8345) <= not b;
    layer3_outputs(8346) <= 1'b1;
    layer3_outputs(8347) <= not a;
    layer3_outputs(8348) <= b;
    layer3_outputs(8349) <= a or b;
    layer3_outputs(8350) <= b;
    layer3_outputs(8351) <= a and not b;
    layer3_outputs(8352) <= not (a xor b);
    layer3_outputs(8353) <= 1'b1;
    layer3_outputs(8354) <= not (a or b);
    layer3_outputs(8355) <= not (a and b);
    layer3_outputs(8356) <= b;
    layer3_outputs(8357) <= b and not a;
    layer3_outputs(8358) <= not b;
    layer3_outputs(8359) <= a and not b;
    layer3_outputs(8360) <= a and not b;
    layer3_outputs(8361) <= b;
    layer3_outputs(8362) <= not a or b;
    layer3_outputs(8363) <= a or b;
    layer3_outputs(8364) <= a or b;
    layer3_outputs(8365) <= b and not a;
    layer3_outputs(8366) <= b;
    layer3_outputs(8367) <= 1'b1;
    layer3_outputs(8368) <= not (a or b);
    layer3_outputs(8369) <= b and not a;
    layer3_outputs(8370) <= 1'b0;
    layer3_outputs(8371) <= not (a and b);
    layer3_outputs(8372) <= not (a and b);
    layer3_outputs(8373) <= a xor b;
    layer3_outputs(8374) <= not b or a;
    layer3_outputs(8375) <= 1'b0;
    layer3_outputs(8376) <= a and not b;
    layer3_outputs(8377) <= a and b;
    layer3_outputs(8378) <= a and b;
    layer3_outputs(8379) <= not b;
    layer3_outputs(8380) <= 1'b0;
    layer3_outputs(8381) <= 1'b0;
    layer3_outputs(8382) <= not (a or b);
    layer3_outputs(8383) <= b and not a;
    layer3_outputs(8384) <= not b or a;
    layer3_outputs(8385) <= not (a or b);
    layer3_outputs(8386) <= not (a or b);
    layer3_outputs(8387) <= a and b;
    layer3_outputs(8388) <= b;
    layer3_outputs(8389) <= 1'b0;
    layer3_outputs(8390) <= not b or a;
    layer3_outputs(8391) <= 1'b1;
    layer3_outputs(8392) <= a and not b;
    layer3_outputs(8393) <= 1'b1;
    layer3_outputs(8394) <= 1'b1;
    layer3_outputs(8395) <= b;
    layer3_outputs(8396) <= a and b;
    layer3_outputs(8397) <= not b;
    layer3_outputs(8398) <= not a;
    layer3_outputs(8399) <= not (a or b);
    layer3_outputs(8400) <= b and not a;
    layer3_outputs(8401) <= not (a or b);
    layer3_outputs(8402) <= 1'b1;
    layer3_outputs(8403) <= not b;
    layer3_outputs(8404) <= not a or b;
    layer3_outputs(8405) <= a;
    layer3_outputs(8406) <= not (a or b);
    layer3_outputs(8407) <= not (a or b);
    layer3_outputs(8408) <= a or b;
    layer3_outputs(8409) <= 1'b1;
    layer3_outputs(8410) <= 1'b0;
    layer3_outputs(8411) <= a or b;
    layer3_outputs(8412) <= b;
    layer3_outputs(8413) <= a and not b;
    layer3_outputs(8414) <= 1'b0;
    layer3_outputs(8415) <= 1'b0;
    layer3_outputs(8416) <= a and b;
    layer3_outputs(8417) <= not a;
    layer3_outputs(8418) <= not (a and b);
    layer3_outputs(8419) <= not a;
    layer3_outputs(8420) <= not a or b;
    layer3_outputs(8421) <= b;
    layer3_outputs(8422) <= 1'b0;
    layer3_outputs(8423) <= not (a and b);
    layer3_outputs(8424) <= 1'b0;
    layer3_outputs(8425) <= not (a or b);
    layer3_outputs(8426) <= b;
    layer3_outputs(8427) <= b;
    layer3_outputs(8428) <= b and not a;
    layer3_outputs(8429) <= 1'b1;
    layer3_outputs(8430) <= 1'b0;
    layer3_outputs(8431) <= b;
    layer3_outputs(8432) <= a;
    layer3_outputs(8433) <= 1'b0;
    layer3_outputs(8434) <= not b;
    layer3_outputs(8435) <= b;
    layer3_outputs(8436) <= 1'b0;
    layer3_outputs(8437) <= a;
    layer3_outputs(8438) <= not b;
    layer3_outputs(8439) <= not (a and b);
    layer3_outputs(8440) <= not (a or b);
    layer3_outputs(8441) <= not a or b;
    layer3_outputs(8442) <= a;
    layer3_outputs(8443) <= not a or b;
    layer3_outputs(8444) <= not a;
    layer3_outputs(8445) <= not a or b;
    layer3_outputs(8446) <= a and not b;
    layer3_outputs(8447) <= 1'b1;
    layer3_outputs(8448) <= 1'b0;
    layer3_outputs(8449) <= a;
    layer3_outputs(8450) <= a or b;
    layer3_outputs(8451) <= not (a or b);
    layer3_outputs(8452) <= not (a and b);
    layer3_outputs(8453) <= not b;
    layer3_outputs(8454) <= not a;
    layer3_outputs(8455) <= b and not a;
    layer3_outputs(8456) <= a and not b;
    layer3_outputs(8457) <= 1'b0;
    layer3_outputs(8458) <= b;
    layer3_outputs(8459) <= 1'b1;
    layer3_outputs(8460) <= b and not a;
    layer3_outputs(8461) <= not b or a;
    layer3_outputs(8462) <= not a or b;
    layer3_outputs(8463) <= b and not a;
    layer3_outputs(8464) <= a and not b;
    layer3_outputs(8465) <= not (a or b);
    layer3_outputs(8466) <= a and b;
    layer3_outputs(8467) <= a;
    layer3_outputs(8468) <= 1'b1;
    layer3_outputs(8469) <= b;
    layer3_outputs(8470) <= a;
    layer3_outputs(8471) <= b;
    layer3_outputs(8472) <= not (a or b);
    layer3_outputs(8473) <= a and not b;
    layer3_outputs(8474) <= 1'b1;
    layer3_outputs(8475) <= 1'b0;
    layer3_outputs(8476) <= b and not a;
    layer3_outputs(8477) <= a or b;
    layer3_outputs(8478) <= a and b;
    layer3_outputs(8479) <= b and not a;
    layer3_outputs(8480) <= 1'b0;
    layer3_outputs(8481) <= not a;
    layer3_outputs(8482) <= not a;
    layer3_outputs(8483) <= not b;
    layer3_outputs(8484) <= not a or b;
    layer3_outputs(8485) <= 1'b0;
    layer3_outputs(8486) <= 1'b1;
    layer3_outputs(8487) <= b and not a;
    layer3_outputs(8488) <= not (a and b);
    layer3_outputs(8489) <= a or b;
    layer3_outputs(8490) <= not a or b;
    layer3_outputs(8491) <= not a or b;
    layer3_outputs(8492) <= a and b;
    layer3_outputs(8493) <= a or b;
    layer3_outputs(8494) <= not a or b;
    layer3_outputs(8495) <= a or b;
    layer3_outputs(8496) <= a and b;
    layer3_outputs(8497) <= not b or a;
    layer3_outputs(8498) <= a and b;
    layer3_outputs(8499) <= not b;
    layer3_outputs(8500) <= b and not a;
    layer3_outputs(8501) <= a;
    layer3_outputs(8502) <= a and b;
    layer3_outputs(8503) <= a and not b;
    layer3_outputs(8504) <= not a or b;
    layer3_outputs(8505) <= not (a xor b);
    layer3_outputs(8506) <= not (a xor b);
    layer3_outputs(8507) <= b and not a;
    layer3_outputs(8508) <= a or b;
    layer3_outputs(8509) <= a and not b;
    layer3_outputs(8510) <= not (a or b);
    layer3_outputs(8511) <= 1'b1;
    layer3_outputs(8512) <= not b or a;
    layer3_outputs(8513) <= not (a and b);
    layer3_outputs(8514) <= a xor b;
    layer3_outputs(8515) <= a and b;
    layer3_outputs(8516) <= 1'b1;
    layer3_outputs(8517) <= a and not b;
    layer3_outputs(8518) <= a or b;
    layer3_outputs(8519) <= b and not a;
    layer3_outputs(8520) <= a and b;
    layer3_outputs(8521) <= not b;
    layer3_outputs(8522) <= not (a xor b);
    layer3_outputs(8523) <= 1'b1;
    layer3_outputs(8524) <= not b;
    layer3_outputs(8525) <= not b or a;
    layer3_outputs(8526) <= a xor b;
    layer3_outputs(8527) <= not b or a;
    layer3_outputs(8528) <= not (a xor b);
    layer3_outputs(8529) <= a or b;
    layer3_outputs(8530) <= not b or a;
    layer3_outputs(8531) <= a or b;
    layer3_outputs(8532) <= 1'b0;
    layer3_outputs(8533) <= not a;
    layer3_outputs(8534) <= not (a xor b);
    layer3_outputs(8535) <= not (a or b);
    layer3_outputs(8536) <= b;
    layer3_outputs(8537) <= a;
    layer3_outputs(8538) <= 1'b0;
    layer3_outputs(8539) <= a and b;
    layer3_outputs(8540) <= b;
    layer3_outputs(8541) <= not b or a;
    layer3_outputs(8542) <= not b or a;
    layer3_outputs(8543) <= 1'b1;
    layer3_outputs(8544) <= 1'b0;
    layer3_outputs(8545) <= not (a or b);
    layer3_outputs(8546) <= not (a and b);
    layer3_outputs(8547) <= a and b;
    layer3_outputs(8548) <= not a or b;
    layer3_outputs(8549) <= not b or a;
    layer3_outputs(8550) <= a and b;
    layer3_outputs(8551) <= a and not b;
    layer3_outputs(8552) <= not b or a;
    layer3_outputs(8553) <= not b;
    layer3_outputs(8554) <= not b or a;
    layer3_outputs(8555) <= b and not a;
    layer3_outputs(8556) <= not (a and b);
    layer3_outputs(8557) <= not (a or b);
    layer3_outputs(8558) <= not a or b;
    layer3_outputs(8559) <= b;
    layer3_outputs(8560) <= not (a xor b);
    layer3_outputs(8561) <= a or b;
    layer3_outputs(8562) <= b;
    layer3_outputs(8563) <= not b;
    layer3_outputs(8564) <= not (a xor b);
    layer3_outputs(8565) <= a;
    layer3_outputs(8566) <= not a;
    layer3_outputs(8567) <= not a or b;
    layer3_outputs(8568) <= a and not b;
    layer3_outputs(8569) <= a and b;
    layer3_outputs(8570) <= b;
    layer3_outputs(8571) <= b and not a;
    layer3_outputs(8572) <= not a or b;
    layer3_outputs(8573) <= not (a or b);
    layer3_outputs(8574) <= not b or a;
    layer3_outputs(8575) <= a xor b;
    layer3_outputs(8576) <= 1'b1;
    layer3_outputs(8577) <= a or b;
    layer3_outputs(8578) <= a and not b;
    layer3_outputs(8579) <= 1'b0;
    layer3_outputs(8580) <= not b;
    layer3_outputs(8581) <= a and b;
    layer3_outputs(8582) <= 1'b0;
    layer3_outputs(8583) <= not (a xor b);
    layer3_outputs(8584) <= not (a or b);
    layer3_outputs(8585) <= a and b;
    layer3_outputs(8586) <= not b;
    layer3_outputs(8587) <= 1'b0;
    layer3_outputs(8588) <= not (a and b);
    layer3_outputs(8589) <= b;
    layer3_outputs(8590) <= not (a or b);
    layer3_outputs(8591) <= not (a or b);
    layer3_outputs(8592) <= not a;
    layer3_outputs(8593) <= 1'b1;
    layer3_outputs(8594) <= not (a or b);
    layer3_outputs(8595) <= not (a and b);
    layer3_outputs(8596) <= not (a and b);
    layer3_outputs(8597) <= a;
    layer3_outputs(8598) <= not a;
    layer3_outputs(8599) <= a or b;
    layer3_outputs(8600) <= not a;
    layer3_outputs(8601) <= a and b;
    layer3_outputs(8602) <= not (a xor b);
    layer3_outputs(8603) <= a and b;
    layer3_outputs(8604) <= 1'b1;
    layer3_outputs(8605) <= not a;
    layer3_outputs(8606) <= 1'b0;
    layer3_outputs(8607) <= 1'b1;
    layer3_outputs(8608) <= a and not b;
    layer3_outputs(8609) <= b and not a;
    layer3_outputs(8610) <= 1'b1;
    layer3_outputs(8611) <= 1'b0;
    layer3_outputs(8612) <= 1'b1;
    layer3_outputs(8613) <= not a or b;
    layer3_outputs(8614) <= a or b;
    layer3_outputs(8615) <= a and b;
    layer3_outputs(8616) <= a;
    layer3_outputs(8617) <= b;
    layer3_outputs(8618) <= a or b;
    layer3_outputs(8619) <= b and not a;
    layer3_outputs(8620) <= a;
    layer3_outputs(8621) <= not a or b;
    layer3_outputs(8622) <= a xor b;
    layer3_outputs(8623) <= not (a or b);
    layer3_outputs(8624) <= not a;
    layer3_outputs(8625) <= b and not a;
    layer3_outputs(8626) <= not (a xor b);
    layer3_outputs(8627) <= not (a or b);
    layer3_outputs(8628) <= not b or a;
    layer3_outputs(8629) <= not b;
    layer3_outputs(8630) <= a and b;
    layer3_outputs(8631) <= 1'b1;
    layer3_outputs(8632) <= a and b;
    layer3_outputs(8633) <= not b;
    layer3_outputs(8634) <= not (a or b);
    layer3_outputs(8635) <= not a;
    layer3_outputs(8636) <= a or b;
    layer3_outputs(8637) <= 1'b1;
    layer3_outputs(8638) <= a or b;
    layer3_outputs(8639) <= a;
    layer3_outputs(8640) <= 1'b0;
    layer3_outputs(8641) <= not b or a;
    layer3_outputs(8642) <= not a;
    layer3_outputs(8643) <= b;
    layer3_outputs(8644) <= 1'b1;
    layer3_outputs(8645) <= not b;
    layer3_outputs(8646) <= a or b;
    layer3_outputs(8647) <= a and not b;
    layer3_outputs(8648) <= not (a or b);
    layer3_outputs(8649) <= not a or b;
    layer3_outputs(8650) <= not (a xor b);
    layer3_outputs(8651) <= b and not a;
    layer3_outputs(8652) <= a and not b;
    layer3_outputs(8653) <= b;
    layer3_outputs(8654) <= a;
    layer3_outputs(8655) <= a or b;
    layer3_outputs(8656) <= b and not a;
    layer3_outputs(8657) <= not a or b;
    layer3_outputs(8658) <= not b;
    layer3_outputs(8659) <= b and not a;
    layer3_outputs(8660) <= 1'b1;
    layer3_outputs(8661) <= not (a or b);
    layer3_outputs(8662) <= not b or a;
    layer3_outputs(8663) <= not a;
    layer3_outputs(8664) <= not a or b;
    layer3_outputs(8665) <= not b;
    layer3_outputs(8666) <= 1'b1;
    layer3_outputs(8667) <= b;
    layer3_outputs(8668) <= a or b;
    layer3_outputs(8669) <= a and b;
    layer3_outputs(8670) <= a and b;
    layer3_outputs(8671) <= a and b;
    layer3_outputs(8672) <= not (a or b);
    layer3_outputs(8673) <= a and not b;
    layer3_outputs(8674) <= 1'b0;
    layer3_outputs(8675) <= a xor b;
    layer3_outputs(8676) <= 1'b1;
    layer3_outputs(8677) <= b;
    layer3_outputs(8678) <= not a or b;
    layer3_outputs(8679) <= a or b;
    layer3_outputs(8680) <= b and not a;
    layer3_outputs(8681) <= not a;
    layer3_outputs(8682) <= a;
    layer3_outputs(8683) <= not (a or b);
    layer3_outputs(8684) <= b and not a;
    layer3_outputs(8685) <= a and not b;
    layer3_outputs(8686) <= a and b;
    layer3_outputs(8687) <= not (a or b);
    layer3_outputs(8688) <= b and not a;
    layer3_outputs(8689) <= not a;
    layer3_outputs(8690) <= not b or a;
    layer3_outputs(8691) <= not b or a;
    layer3_outputs(8692) <= not (a or b);
    layer3_outputs(8693) <= not b or a;
    layer3_outputs(8694) <= a and b;
    layer3_outputs(8695) <= b;
    layer3_outputs(8696) <= 1'b1;
    layer3_outputs(8697) <= not a or b;
    layer3_outputs(8698) <= 1'b1;
    layer3_outputs(8699) <= a;
    layer3_outputs(8700) <= 1'b0;
    layer3_outputs(8701) <= a and b;
    layer3_outputs(8702) <= a and b;
    layer3_outputs(8703) <= a and b;
    layer3_outputs(8704) <= b;
    layer3_outputs(8705) <= not (a and b);
    layer3_outputs(8706) <= 1'b1;
    layer3_outputs(8707) <= not (a and b);
    layer3_outputs(8708) <= not a;
    layer3_outputs(8709) <= b;
    layer3_outputs(8710) <= 1'b0;
    layer3_outputs(8711) <= a and not b;
    layer3_outputs(8712) <= b and not a;
    layer3_outputs(8713) <= not a;
    layer3_outputs(8714) <= a;
    layer3_outputs(8715) <= b and not a;
    layer3_outputs(8716) <= not b;
    layer3_outputs(8717) <= a or b;
    layer3_outputs(8718) <= not b or a;
    layer3_outputs(8719) <= not (a and b);
    layer3_outputs(8720) <= not (a and b);
    layer3_outputs(8721) <= b;
    layer3_outputs(8722) <= 1'b1;
    layer3_outputs(8723) <= not (a xor b);
    layer3_outputs(8724) <= 1'b1;
    layer3_outputs(8725) <= not b;
    layer3_outputs(8726) <= a and not b;
    layer3_outputs(8727) <= not (a or b);
    layer3_outputs(8728) <= a xor b;
    layer3_outputs(8729) <= not b or a;
    layer3_outputs(8730) <= 1'b0;
    layer3_outputs(8731) <= not b;
    layer3_outputs(8732) <= not b;
    layer3_outputs(8733) <= b and not a;
    layer3_outputs(8734) <= not b or a;
    layer3_outputs(8735) <= a and b;
    layer3_outputs(8736) <= not b;
    layer3_outputs(8737) <= 1'b1;
    layer3_outputs(8738) <= not a;
    layer3_outputs(8739) <= not b;
    layer3_outputs(8740) <= 1'b1;
    layer3_outputs(8741) <= not (a and b);
    layer3_outputs(8742) <= b and not a;
    layer3_outputs(8743) <= 1'b0;
    layer3_outputs(8744) <= not (a and b);
    layer3_outputs(8745) <= a and not b;
    layer3_outputs(8746) <= a or b;
    layer3_outputs(8747) <= not (a and b);
    layer3_outputs(8748) <= a xor b;
    layer3_outputs(8749) <= b and not a;
    layer3_outputs(8750) <= a and not b;
    layer3_outputs(8751) <= not (a and b);
    layer3_outputs(8752) <= 1'b0;
    layer3_outputs(8753) <= a;
    layer3_outputs(8754) <= not a;
    layer3_outputs(8755) <= not a or b;
    layer3_outputs(8756) <= a xor b;
    layer3_outputs(8757) <= 1'b1;
    layer3_outputs(8758) <= b;
    layer3_outputs(8759) <= a;
    layer3_outputs(8760) <= not a or b;
    layer3_outputs(8761) <= a and not b;
    layer3_outputs(8762) <= a and b;
    layer3_outputs(8763) <= not a or b;
    layer3_outputs(8764) <= a xor b;
    layer3_outputs(8765) <= a or b;
    layer3_outputs(8766) <= a or b;
    layer3_outputs(8767) <= not a or b;
    layer3_outputs(8768) <= 1'b1;
    layer3_outputs(8769) <= a and b;
    layer3_outputs(8770) <= not a;
    layer3_outputs(8771) <= 1'b1;
    layer3_outputs(8772) <= b and not a;
    layer3_outputs(8773) <= b;
    layer3_outputs(8774) <= b and not a;
    layer3_outputs(8775) <= 1'b1;
    layer3_outputs(8776) <= not (a or b);
    layer3_outputs(8777) <= 1'b1;
    layer3_outputs(8778) <= not b;
    layer3_outputs(8779) <= not (a xor b);
    layer3_outputs(8780) <= not (a or b);
    layer3_outputs(8781) <= not b or a;
    layer3_outputs(8782) <= not (a and b);
    layer3_outputs(8783) <= 1'b1;
    layer3_outputs(8784) <= b;
    layer3_outputs(8785) <= not b;
    layer3_outputs(8786) <= not b;
    layer3_outputs(8787) <= not (a or b);
    layer3_outputs(8788) <= b;
    layer3_outputs(8789) <= not b or a;
    layer3_outputs(8790) <= not b or a;
    layer3_outputs(8791) <= not (a or b);
    layer3_outputs(8792) <= a and not b;
    layer3_outputs(8793) <= b;
    layer3_outputs(8794) <= a;
    layer3_outputs(8795) <= not (a xor b);
    layer3_outputs(8796) <= not b or a;
    layer3_outputs(8797) <= b;
    layer3_outputs(8798) <= not a;
    layer3_outputs(8799) <= 1'b0;
    layer3_outputs(8800) <= 1'b0;
    layer3_outputs(8801) <= 1'b1;
    layer3_outputs(8802) <= not b;
    layer3_outputs(8803) <= not (a or b);
    layer3_outputs(8804) <= b and not a;
    layer3_outputs(8805) <= not b or a;
    layer3_outputs(8806) <= not b;
    layer3_outputs(8807) <= not a or b;
    layer3_outputs(8808) <= not (a or b);
    layer3_outputs(8809) <= b;
    layer3_outputs(8810) <= a or b;
    layer3_outputs(8811) <= not a;
    layer3_outputs(8812) <= a and b;
    layer3_outputs(8813) <= 1'b1;
    layer3_outputs(8814) <= a and b;
    layer3_outputs(8815) <= 1'b1;
    layer3_outputs(8816) <= b and not a;
    layer3_outputs(8817) <= not a or b;
    layer3_outputs(8818) <= not b or a;
    layer3_outputs(8819) <= not a;
    layer3_outputs(8820) <= a;
    layer3_outputs(8821) <= b and not a;
    layer3_outputs(8822) <= not (a xor b);
    layer3_outputs(8823) <= not b;
    layer3_outputs(8824) <= 1'b0;
    layer3_outputs(8825) <= a or b;
    layer3_outputs(8826) <= b;
    layer3_outputs(8827) <= a and b;
    layer3_outputs(8828) <= b and not a;
    layer3_outputs(8829) <= 1'b1;
    layer3_outputs(8830) <= not a;
    layer3_outputs(8831) <= 1'b0;
    layer3_outputs(8832) <= 1'b1;
    layer3_outputs(8833) <= not (a and b);
    layer3_outputs(8834) <= a and b;
    layer3_outputs(8835) <= not b;
    layer3_outputs(8836) <= a and b;
    layer3_outputs(8837) <= 1'b1;
    layer3_outputs(8838) <= a and b;
    layer3_outputs(8839) <= not b or a;
    layer3_outputs(8840) <= not b or a;
    layer3_outputs(8841) <= b and not a;
    layer3_outputs(8842) <= not (a and b);
    layer3_outputs(8843) <= not b or a;
    layer3_outputs(8844) <= not b;
    layer3_outputs(8845) <= a or b;
    layer3_outputs(8846) <= b;
    layer3_outputs(8847) <= a and b;
    layer3_outputs(8848) <= not b or a;
    layer3_outputs(8849) <= not b;
    layer3_outputs(8850) <= not (a or b);
    layer3_outputs(8851) <= not a or b;
    layer3_outputs(8852) <= a;
    layer3_outputs(8853) <= not b;
    layer3_outputs(8854) <= not b or a;
    layer3_outputs(8855) <= a xor b;
    layer3_outputs(8856) <= a or b;
    layer3_outputs(8857) <= not b or a;
    layer3_outputs(8858) <= b;
    layer3_outputs(8859) <= a or b;
    layer3_outputs(8860) <= not a or b;
    layer3_outputs(8861) <= a and b;
    layer3_outputs(8862) <= a and not b;
    layer3_outputs(8863) <= b;
    layer3_outputs(8864) <= not a;
    layer3_outputs(8865) <= a and not b;
    layer3_outputs(8866) <= not a;
    layer3_outputs(8867) <= not b or a;
    layer3_outputs(8868) <= not b;
    layer3_outputs(8869) <= not (a or b);
    layer3_outputs(8870) <= not a;
    layer3_outputs(8871) <= 1'b0;
    layer3_outputs(8872) <= a and b;
    layer3_outputs(8873) <= not (a or b);
    layer3_outputs(8874) <= 1'b0;
    layer3_outputs(8875) <= a and not b;
    layer3_outputs(8876) <= a or b;
    layer3_outputs(8877) <= not b;
    layer3_outputs(8878) <= not (a xor b);
    layer3_outputs(8879) <= b;
    layer3_outputs(8880) <= not a;
    layer3_outputs(8881) <= b and not a;
    layer3_outputs(8882) <= a;
    layer3_outputs(8883) <= a or b;
    layer3_outputs(8884) <= not a;
    layer3_outputs(8885) <= a or b;
    layer3_outputs(8886) <= a xor b;
    layer3_outputs(8887) <= not (a or b);
    layer3_outputs(8888) <= a or b;
    layer3_outputs(8889) <= not (a and b);
    layer3_outputs(8890) <= 1'b1;
    layer3_outputs(8891) <= b;
    layer3_outputs(8892) <= b;
    layer3_outputs(8893) <= a and b;
    layer3_outputs(8894) <= not a or b;
    layer3_outputs(8895) <= 1'b1;
    layer3_outputs(8896) <= not b or a;
    layer3_outputs(8897) <= a;
    layer3_outputs(8898) <= not b or a;
    layer3_outputs(8899) <= not (a and b);
    layer3_outputs(8900) <= a and not b;
    layer3_outputs(8901) <= a;
    layer3_outputs(8902) <= 1'b1;
    layer3_outputs(8903) <= b;
    layer3_outputs(8904) <= 1'b0;
    layer3_outputs(8905) <= a and not b;
    layer3_outputs(8906) <= a;
    layer3_outputs(8907) <= b;
    layer3_outputs(8908) <= b and not a;
    layer3_outputs(8909) <= 1'b0;
    layer3_outputs(8910) <= not a;
    layer3_outputs(8911) <= b and not a;
    layer3_outputs(8912) <= a and not b;
    layer3_outputs(8913) <= b;
    layer3_outputs(8914) <= not a;
    layer3_outputs(8915) <= a and b;
    layer3_outputs(8916) <= not (a or b);
    layer3_outputs(8917) <= 1'b1;
    layer3_outputs(8918) <= b and not a;
    layer3_outputs(8919) <= b and not a;
    layer3_outputs(8920) <= not b;
    layer3_outputs(8921) <= not a or b;
    layer3_outputs(8922) <= a and not b;
    layer3_outputs(8923) <= 1'b0;
    layer3_outputs(8924) <= b;
    layer3_outputs(8925) <= a or b;
    layer3_outputs(8926) <= not b or a;
    layer3_outputs(8927) <= 1'b0;
    layer3_outputs(8928) <= a and not b;
    layer3_outputs(8929) <= 1'b1;
    layer3_outputs(8930) <= not a;
    layer3_outputs(8931) <= a and b;
    layer3_outputs(8932) <= a or b;
    layer3_outputs(8933) <= not b or a;
    layer3_outputs(8934) <= not a;
    layer3_outputs(8935) <= 1'b0;
    layer3_outputs(8936) <= not a or b;
    layer3_outputs(8937) <= not a or b;
    layer3_outputs(8938) <= a;
    layer3_outputs(8939) <= a;
    layer3_outputs(8940) <= 1'b0;
    layer3_outputs(8941) <= not b;
    layer3_outputs(8942) <= b;
    layer3_outputs(8943) <= 1'b0;
    layer3_outputs(8944) <= 1'b1;
    layer3_outputs(8945) <= not b or a;
    layer3_outputs(8946) <= not a or b;
    layer3_outputs(8947) <= a and not b;
    layer3_outputs(8948) <= b and not a;
    layer3_outputs(8949) <= not a;
    layer3_outputs(8950) <= not a or b;
    layer3_outputs(8951) <= not b;
    layer3_outputs(8952) <= 1'b0;
    layer3_outputs(8953) <= a and not b;
    layer3_outputs(8954) <= not a;
    layer3_outputs(8955) <= not b;
    layer3_outputs(8956) <= 1'b0;
    layer3_outputs(8957) <= a and b;
    layer3_outputs(8958) <= not a;
    layer3_outputs(8959) <= b;
    layer3_outputs(8960) <= not a or b;
    layer3_outputs(8961) <= a and not b;
    layer3_outputs(8962) <= not b or a;
    layer3_outputs(8963) <= not (a or b);
    layer3_outputs(8964) <= not (a or b);
    layer3_outputs(8965) <= not b or a;
    layer3_outputs(8966) <= not (a and b);
    layer3_outputs(8967) <= a or b;
    layer3_outputs(8968) <= a and b;
    layer3_outputs(8969) <= a or b;
    layer3_outputs(8970) <= a;
    layer3_outputs(8971) <= 1'b0;
    layer3_outputs(8972) <= a and not b;
    layer3_outputs(8973) <= a or b;
    layer3_outputs(8974) <= not (a or b);
    layer3_outputs(8975) <= not (a and b);
    layer3_outputs(8976) <= 1'b0;
    layer3_outputs(8977) <= not b or a;
    layer3_outputs(8978) <= b and not a;
    layer3_outputs(8979) <= 1'b1;
    layer3_outputs(8980) <= a and not b;
    layer3_outputs(8981) <= not a or b;
    layer3_outputs(8982) <= a or b;
    layer3_outputs(8983) <= b;
    layer3_outputs(8984) <= not a;
    layer3_outputs(8985) <= not a or b;
    layer3_outputs(8986) <= not (a and b);
    layer3_outputs(8987) <= not b;
    layer3_outputs(8988) <= b;
    layer3_outputs(8989) <= b and not a;
    layer3_outputs(8990) <= 1'b0;
    layer3_outputs(8991) <= a and not b;
    layer3_outputs(8992) <= not b;
    layer3_outputs(8993) <= b and not a;
    layer3_outputs(8994) <= a;
    layer3_outputs(8995) <= b and not a;
    layer3_outputs(8996) <= 1'b0;
    layer3_outputs(8997) <= a and not b;
    layer3_outputs(8998) <= not a or b;
    layer3_outputs(8999) <= a and not b;
    layer3_outputs(9000) <= not b or a;
    layer3_outputs(9001) <= a and b;
    layer3_outputs(9002) <= a or b;
    layer3_outputs(9003) <= 1'b0;
    layer3_outputs(9004) <= not a or b;
    layer3_outputs(9005) <= not b or a;
    layer3_outputs(9006) <= not (a or b);
    layer3_outputs(9007) <= 1'b1;
    layer3_outputs(9008) <= a and b;
    layer3_outputs(9009) <= 1'b1;
    layer3_outputs(9010) <= b;
    layer3_outputs(9011) <= a and not b;
    layer3_outputs(9012) <= b;
    layer3_outputs(9013) <= not b or a;
    layer3_outputs(9014) <= not (a or b);
    layer3_outputs(9015) <= not (a and b);
    layer3_outputs(9016) <= 1'b0;
    layer3_outputs(9017) <= 1'b0;
    layer3_outputs(9018) <= not (a xor b);
    layer3_outputs(9019) <= not a or b;
    layer3_outputs(9020) <= not (a and b);
    layer3_outputs(9021) <= not (a or b);
    layer3_outputs(9022) <= a xor b;
    layer3_outputs(9023) <= 1'b0;
    layer3_outputs(9024) <= not a;
    layer3_outputs(9025) <= not (a xor b);
    layer3_outputs(9026) <= 1'b1;
    layer3_outputs(9027) <= b;
    layer3_outputs(9028) <= a and not b;
    layer3_outputs(9029) <= not (a and b);
    layer3_outputs(9030) <= not (a or b);
    layer3_outputs(9031) <= a and b;
    layer3_outputs(9032) <= a and b;
    layer3_outputs(9033) <= a and b;
    layer3_outputs(9034) <= not a;
    layer3_outputs(9035) <= not (a and b);
    layer3_outputs(9036) <= not b;
    layer3_outputs(9037) <= not (a xor b);
    layer3_outputs(9038) <= a;
    layer3_outputs(9039) <= 1'b0;
    layer3_outputs(9040) <= a xor b;
    layer3_outputs(9041) <= a;
    layer3_outputs(9042) <= a or b;
    layer3_outputs(9043) <= a and not b;
    layer3_outputs(9044) <= b and not a;
    layer3_outputs(9045) <= a and b;
    layer3_outputs(9046) <= not (a or b);
    layer3_outputs(9047) <= not a;
    layer3_outputs(9048) <= not (a xor b);
    layer3_outputs(9049) <= not b;
    layer3_outputs(9050) <= 1'b1;
    layer3_outputs(9051) <= 1'b1;
    layer3_outputs(9052) <= a and not b;
    layer3_outputs(9053) <= not a;
    layer3_outputs(9054) <= a or b;
    layer3_outputs(9055) <= not b;
    layer3_outputs(9056) <= not (a and b);
    layer3_outputs(9057) <= a xor b;
    layer3_outputs(9058) <= 1'b0;
    layer3_outputs(9059) <= not a;
    layer3_outputs(9060) <= a and b;
    layer3_outputs(9061) <= a and not b;
    layer3_outputs(9062) <= a and b;
    layer3_outputs(9063) <= b;
    layer3_outputs(9064) <= not (a or b);
    layer3_outputs(9065) <= not (a and b);
    layer3_outputs(9066) <= a xor b;
    layer3_outputs(9067) <= 1'b1;
    layer3_outputs(9068) <= not b;
    layer3_outputs(9069) <= 1'b0;
    layer3_outputs(9070) <= 1'b0;
    layer3_outputs(9071) <= b and not a;
    layer3_outputs(9072) <= a;
    layer3_outputs(9073) <= not (a or b);
    layer3_outputs(9074) <= not b;
    layer3_outputs(9075) <= b;
    layer3_outputs(9076) <= 1'b1;
    layer3_outputs(9077) <= not a;
    layer3_outputs(9078) <= a;
    layer3_outputs(9079) <= a;
    layer3_outputs(9080) <= not b or a;
    layer3_outputs(9081) <= a or b;
    layer3_outputs(9082) <= not (a and b);
    layer3_outputs(9083) <= a xor b;
    layer3_outputs(9084) <= b and not a;
    layer3_outputs(9085) <= a or b;
    layer3_outputs(9086) <= not b;
    layer3_outputs(9087) <= 1'b1;
    layer3_outputs(9088) <= a;
    layer3_outputs(9089) <= 1'b0;
    layer3_outputs(9090) <= 1'b0;
    layer3_outputs(9091) <= not b or a;
    layer3_outputs(9092) <= a and b;
    layer3_outputs(9093) <= 1'b1;
    layer3_outputs(9094) <= a and b;
    layer3_outputs(9095) <= 1'b0;
    layer3_outputs(9096) <= b and not a;
    layer3_outputs(9097) <= 1'b1;
    layer3_outputs(9098) <= 1'b0;
    layer3_outputs(9099) <= a;
    layer3_outputs(9100) <= a;
    layer3_outputs(9101) <= not (a and b);
    layer3_outputs(9102) <= b and not a;
    layer3_outputs(9103) <= a and b;
    layer3_outputs(9104) <= not a or b;
    layer3_outputs(9105) <= a and not b;
    layer3_outputs(9106) <= a;
    layer3_outputs(9107) <= not b;
    layer3_outputs(9108) <= a xor b;
    layer3_outputs(9109) <= not a or b;
    layer3_outputs(9110) <= a and not b;
    layer3_outputs(9111) <= not (a xor b);
    layer3_outputs(9112) <= b and not a;
    layer3_outputs(9113) <= a and b;
    layer3_outputs(9114) <= 1'b1;
    layer3_outputs(9115) <= a and not b;
    layer3_outputs(9116) <= not b or a;
    layer3_outputs(9117) <= b;
    layer3_outputs(9118) <= a xor b;
    layer3_outputs(9119) <= not a or b;
    layer3_outputs(9120) <= 1'b0;
    layer3_outputs(9121) <= not b or a;
    layer3_outputs(9122) <= a or b;
    layer3_outputs(9123) <= not (a or b);
    layer3_outputs(9124) <= a and b;
    layer3_outputs(9125) <= 1'b1;
    layer3_outputs(9126) <= not a;
    layer3_outputs(9127) <= not a;
    layer3_outputs(9128) <= a or b;
    layer3_outputs(9129) <= a or b;
    layer3_outputs(9130) <= not a or b;
    layer3_outputs(9131) <= not b;
    layer3_outputs(9132) <= not a;
    layer3_outputs(9133) <= not (a and b);
    layer3_outputs(9134) <= 1'b0;
    layer3_outputs(9135) <= b and not a;
    layer3_outputs(9136) <= b and not a;
    layer3_outputs(9137) <= a;
    layer3_outputs(9138) <= a xor b;
    layer3_outputs(9139) <= a;
    layer3_outputs(9140) <= b and not a;
    layer3_outputs(9141) <= a;
    layer3_outputs(9142) <= not (a or b);
    layer3_outputs(9143) <= a or b;
    layer3_outputs(9144) <= a and b;
    layer3_outputs(9145) <= 1'b0;
    layer3_outputs(9146) <= a and b;
    layer3_outputs(9147) <= not b;
    layer3_outputs(9148) <= not (a or b);
    layer3_outputs(9149) <= 1'b0;
    layer3_outputs(9150) <= not b;
    layer3_outputs(9151) <= 1'b1;
    layer3_outputs(9152) <= not b;
    layer3_outputs(9153) <= a and not b;
    layer3_outputs(9154) <= not (a or b);
    layer3_outputs(9155) <= b and not a;
    layer3_outputs(9156) <= b;
    layer3_outputs(9157) <= b and not a;
    layer3_outputs(9158) <= 1'b0;
    layer3_outputs(9159) <= not (a and b);
    layer3_outputs(9160) <= a and b;
    layer3_outputs(9161) <= a or b;
    layer3_outputs(9162) <= not b or a;
    layer3_outputs(9163) <= a xor b;
    layer3_outputs(9164) <= not a or b;
    layer3_outputs(9165) <= not (a and b);
    layer3_outputs(9166) <= not b;
    layer3_outputs(9167) <= a and not b;
    layer3_outputs(9168) <= 1'b1;
    layer3_outputs(9169) <= b and not a;
    layer3_outputs(9170) <= not b or a;
    layer3_outputs(9171) <= a and b;
    layer3_outputs(9172) <= not a;
    layer3_outputs(9173) <= not (a or b);
    layer3_outputs(9174) <= b;
    layer3_outputs(9175) <= a and not b;
    layer3_outputs(9176) <= not a;
    layer3_outputs(9177) <= a;
    layer3_outputs(9178) <= b;
    layer3_outputs(9179) <= 1'b1;
    layer3_outputs(9180) <= not a or b;
    layer3_outputs(9181) <= not (a or b);
    layer3_outputs(9182) <= not a or b;
    layer3_outputs(9183) <= a xor b;
    layer3_outputs(9184) <= a and b;
    layer3_outputs(9185) <= not a or b;
    layer3_outputs(9186) <= a or b;
    layer3_outputs(9187) <= a and not b;
    layer3_outputs(9188) <= a and b;
    layer3_outputs(9189) <= not a;
    layer3_outputs(9190) <= not b;
    layer3_outputs(9191) <= not (a or b);
    layer3_outputs(9192) <= not b or a;
    layer3_outputs(9193) <= a and not b;
    layer3_outputs(9194) <= not b;
    layer3_outputs(9195) <= not (a xor b);
    layer3_outputs(9196) <= not b or a;
    layer3_outputs(9197) <= not a or b;
    layer3_outputs(9198) <= a or b;
    layer3_outputs(9199) <= 1'b1;
    layer3_outputs(9200) <= 1'b1;
    layer3_outputs(9201) <= 1'b0;
    layer3_outputs(9202) <= a or b;
    layer3_outputs(9203) <= a;
    layer3_outputs(9204) <= not a or b;
    layer3_outputs(9205) <= 1'b0;
    layer3_outputs(9206) <= b;
    layer3_outputs(9207) <= not (a and b);
    layer3_outputs(9208) <= a or b;
    layer3_outputs(9209) <= b and not a;
    layer3_outputs(9210) <= not b;
    layer3_outputs(9211) <= b and not a;
    layer3_outputs(9212) <= a;
    layer3_outputs(9213) <= not a;
    layer3_outputs(9214) <= b and not a;
    layer3_outputs(9215) <= not (a or b);
    layer3_outputs(9216) <= not (a or b);
    layer3_outputs(9217) <= 1'b0;
    layer3_outputs(9218) <= not (a or b);
    layer3_outputs(9219) <= a xor b;
    layer3_outputs(9220) <= 1'b1;
    layer3_outputs(9221) <= 1'b1;
    layer3_outputs(9222) <= not a;
    layer3_outputs(9223) <= not (a or b);
    layer3_outputs(9224) <= not b;
    layer3_outputs(9225) <= b;
    layer3_outputs(9226) <= a and not b;
    layer3_outputs(9227) <= not a or b;
    layer3_outputs(9228) <= a and not b;
    layer3_outputs(9229) <= b;
    layer3_outputs(9230) <= a and b;
    layer3_outputs(9231) <= a;
    layer3_outputs(9232) <= a and b;
    layer3_outputs(9233) <= 1'b0;
    layer3_outputs(9234) <= 1'b0;
    layer3_outputs(9235) <= not b;
    layer3_outputs(9236) <= a;
    layer3_outputs(9237) <= 1'b0;
    layer3_outputs(9238) <= b and not a;
    layer3_outputs(9239) <= a xor b;
    layer3_outputs(9240) <= a and b;
    layer3_outputs(9241) <= 1'b0;
    layer3_outputs(9242) <= not b;
    layer3_outputs(9243) <= a and not b;
    layer3_outputs(9244) <= not a;
    layer3_outputs(9245) <= a and b;
    layer3_outputs(9246) <= a or b;
    layer3_outputs(9247) <= a;
    layer3_outputs(9248) <= b and not a;
    layer3_outputs(9249) <= not (a and b);
    layer3_outputs(9250) <= not (a xor b);
    layer3_outputs(9251) <= a and b;
    layer3_outputs(9252) <= a xor b;
    layer3_outputs(9253) <= b;
    layer3_outputs(9254) <= 1'b0;
    layer3_outputs(9255) <= b and not a;
    layer3_outputs(9256) <= a and not b;
    layer3_outputs(9257) <= not a;
    layer3_outputs(9258) <= a or b;
    layer3_outputs(9259) <= 1'b0;
    layer3_outputs(9260) <= not a;
    layer3_outputs(9261) <= not (a or b);
    layer3_outputs(9262) <= not b or a;
    layer3_outputs(9263) <= a and b;
    layer3_outputs(9264) <= not b or a;
    layer3_outputs(9265) <= a;
    layer3_outputs(9266) <= not a or b;
    layer3_outputs(9267) <= b;
    layer3_outputs(9268) <= a;
    layer3_outputs(9269) <= not b or a;
    layer3_outputs(9270) <= a and b;
    layer3_outputs(9271) <= 1'b1;
    layer3_outputs(9272) <= b;
    layer3_outputs(9273) <= 1'b0;
    layer3_outputs(9274) <= a and not b;
    layer3_outputs(9275) <= not a;
    layer3_outputs(9276) <= not a;
    layer3_outputs(9277) <= b and not a;
    layer3_outputs(9278) <= not b or a;
    layer3_outputs(9279) <= a or b;
    layer3_outputs(9280) <= not (a and b);
    layer3_outputs(9281) <= not b or a;
    layer3_outputs(9282) <= a;
    layer3_outputs(9283) <= a and b;
    layer3_outputs(9284) <= 1'b0;
    layer3_outputs(9285) <= a;
    layer3_outputs(9286) <= not b or a;
    layer3_outputs(9287) <= not (a or b);
    layer3_outputs(9288) <= a;
    layer3_outputs(9289) <= not (a and b);
    layer3_outputs(9290) <= b and not a;
    layer3_outputs(9291) <= 1'b0;
    layer3_outputs(9292) <= a or b;
    layer3_outputs(9293) <= 1'b1;
    layer3_outputs(9294) <= not b or a;
    layer3_outputs(9295) <= b;
    layer3_outputs(9296) <= a and not b;
    layer3_outputs(9297) <= a and b;
    layer3_outputs(9298) <= not a or b;
    layer3_outputs(9299) <= a xor b;
    layer3_outputs(9300) <= not b or a;
    layer3_outputs(9301) <= not (a and b);
    layer3_outputs(9302) <= a;
    layer3_outputs(9303) <= 1'b1;
    layer3_outputs(9304) <= a or b;
    layer3_outputs(9305) <= b and not a;
    layer3_outputs(9306) <= not a or b;
    layer3_outputs(9307) <= a xor b;
    layer3_outputs(9308) <= 1'b0;
    layer3_outputs(9309) <= not b;
    layer3_outputs(9310) <= b;
    layer3_outputs(9311) <= not (a or b);
    layer3_outputs(9312) <= not b;
    layer3_outputs(9313) <= b and not a;
    layer3_outputs(9314) <= a;
    layer3_outputs(9315) <= a or b;
    layer3_outputs(9316) <= 1'b0;
    layer3_outputs(9317) <= a;
    layer3_outputs(9318) <= not b or a;
    layer3_outputs(9319) <= a and not b;
    layer3_outputs(9320) <= not a;
    layer3_outputs(9321) <= not (a or b);
    layer3_outputs(9322) <= 1'b1;
    layer3_outputs(9323) <= 1'b1;
    layer3_outputs(9324) <= not b or a;
    layer3_outputs(9325) <= not b;
    layer3_outputs(9326) <= a and not b;
    layer3_outputs(9327) <= a and not b;
    layer3_outputs(9328) <= not a;
    layer3_outputs(9329) <= a and b;
    layer3_outputs(9330) <= not a or b;
    layer3_outputs(9331) <= 1'b0;
    layer3_outputs(9332) <= 1'b0;
    layer3_outputs(9333) <= not (a or b);
    layer3_outputs(9334) <= b and not a;
    layer3_outputs(9335) <= a and b;
    layer3_outputs(9336) <= a and not b;
    layer3_outputs(9337) <= not b;
    layer3_outputs(9338) <= a;
    layer3_outputs(9339) <= a xor b;
    layer3_outputs(9340) <= b and not a;
    layer3_outputs(9341) <= not a;
    layer3_outputs(9342) <= b and not a;
    layer3_outputs(9343) <= b;
    layer3_outputs(9344) <= a or b;
    layer3_outputs(9345) <= 1'b1;
    layer3_outputs(9346) <= 1'b1;
    layer3_outputs(9347) <= a or b;
    layer3_outputs(9348) <= not (a xor b);
    layer3_outputs(9349) <= a and b;
    layer3_outputs(9350) <= a and not b;
    layer3_outputs(9351) <= not a or b;
    layer3_outputs(9352) <= 1'b1;
    layer3_outputs(9353) <= a or b;
    layer3_outputs(9354) <= a or b;
    layer3_outputs(9355) <= not b;
    layer3_outputs(9356) <= a or b;
    layer3_outputs(9357) <= a or b;
    layer3_outputs(9358) <= not (a and b);
    layer3_outputs(9359) <= not a;
    layer3_outputs(9360) <= a;
    layer3_outputs(9361) <= a and not b;
    layer3_outputs(9362) <= 1'b1;
    layer3_outputs(9363) <= a and b;
    layer3_outputs(9364) <= not b or a;
    layer3_outputs(9365) <= not a;
    layer3_outputs(9366) <= a and not b;
    layer3_outputs(9367) <= not a;
    layer3_outputs(9368) <= a and b;
    layer3_outputs(9369) <= a and b;
    layer3_outputs(9370) <= not a;
    layer3_outputs(9371) <= a and b;
    layer3_outputs(9372) <= a;
    layer3_outputs(9373) <= a or b;
    layer3_outputs(9374) <= not (a xor b);
    layer3_outputs(9375) <= not a or b;
    layer3_outputs(9376) <= a and b;
    layer3_outputs(9377) <= b and not a;
    layer3_outputs(9378) <= not a or b;
    layer3_outputs(9379) <= b;
    layer3_outputs(9380) <= not (a xor b);
    layer3_outputs(9381) <= a or b;
    layer3_outputs(9382) <= a xor b;
    layer3_outputs(9383) <= not (a xor b);
    layer3_outputs(9384) <= a or b;
    layer3_outputs(9385) <= a or b;
    layer3_outputs(9386) <= a or b;
    layer3_outputs(9387) <= not a or b;
    layer3_outputs(9388) <= a and not b;
    layer3_outputs(9389) <= a and not b;
    layer3_outputs(9390) <= 1'b0;
    layer3_outputs(9391) <= not a or b;
    layer3_outputs(9392) <= a and not b;
    layer3_outputs(9393) <= not (a xor b);
    layer3_outputs(9394) <= 1'b1;
    layer3_outputs(9395) <= a and not b;
    layer3_outputs(9396) <= a xor b;
    layer3_outputs(9397) <= not (a xor b);
    layer3_outputs(9398) <= not a or b;
    layer3_outputs(9399) <= a and not b;
    layer3_outputs(9400) <= 1'b1;
    layer3_outputs(9401) <= a;
    layer3_outputs(9402) <= 1'b0;
    layer3_outputs(9403) <= 1'b1;
    layer3_outputs(9404) <= a;
    layer3_outputs(9405) <= 1'b1;
    layer3_outputs(9406) <= not (a xor b);
    layer3_outputs(9407) <= a xor b;
    layer3_outputs(9408) <= a and not b;
    layer3_outputs(9409) <= not a;
    layer3_outputs(9410) <= 1'b0;
    layer3_outputs(9411) <= not (a or b);
    layer3_outputs(9412) <= not b or a;
    layer3_outputs(9413) <= a or b;
    layer3_outputs(9414) <= b;
    layer3_outputs(9415) <= b;
    layer3_outputs(9416) <= not b;
    layer3_outputs(9417) <= a and not b;
    layer3_outputs(9418) <= not a or b;
    layer3_outputs(9419) <= b and not a;
    layer3_outputs(9420) <= b and not a;
    layer3_outputs(9421) <= b;
    layer3_outputs(9422) <= 1'b1;
    layer3_outputs(9423) <= not a;
    layer3_outputs(9424) <= a;
    layer3_outputs(9425) <= not (a xor b);
    layer3_outputs(9426) <= a;
    layer3_outputs(9427) <= not a or b;
    layer3_outputs(9428) <= a or b;
    layer3_outputs(9429) <= a or b;
    layer3_outputs(9430) <= a or b;
    layer3_outputs(9431) <= b;
    layer3_outputs(9432) <= a;
    layer3_outputs(9433) <= not (a or b);
    layer3_outputs(9434) <= a and not b;
    layer3_outputs(9435) <= 1'b0;
    layer3_outputs(9436) <= a;
    layer3_outputs(9437) <= not a;
    layer3_outputs(9438) <= a;
    layer3_outputs(9439) <= a and b;
    layer3_outputs(9440) <= a;
    layer3_outputs(9441) <= not b;
    layer3_outputs(9442) <= not (a or b);
    layer3_outputs(9443) <= a;
    layer3_outputs(9444) <= not b;
    layer3_outputs(9445) <= a and not b;
    layer3_outputs(9446) <= not b or a;
    layer3_outputs(9447) <= not (a and b);
    layer3_outputs(9448) <= b;
    layer3_outputs(9449) <= b;
    layer3_outputs(9450) <= a xor b;
    layer3_outputs(9451) <= a and not b;
    layer3_outputs(9452) <= 1'b0;
    layer3_outputs(9453) <= not b or a;
    layer3_outputs(9454) <= a and not b;
    layer3_outputs(9455) <= not a;
    layer3_outputs(9456) <= not a or b;
    layer3_outputs(9457) <= 1'b0;
    layer3_outputs(9458) <= not (a and b);
    layer3_outputs(9459) <= b and not a;
    layer3_outputs(9460) <= a or b;
    layer3_outputs(9461) <= not a or b;
    layer3_outputs(9462) <= a and b;
    layer3_outputs(9463) <= not b;
    layer3_outputs(9464) <= 1'b1;
    layer3_outputs(9465) <= not a or b;
    layer3_outputs(9466) <= a xor b;
    layer3_outputs(9467) <= not b;
    layer3_outputs(9468) <= not (a and b);
    layer3_outputs(9469) <= not b;
    layer3_outputs(9470) <= 1'b1;
    layer3_outputs(9471) <= b;
    layer3_outputs(9472) <= a and b;
    layer3_outputs(9473) <= not a;
    layer3_outputs(9474) <= a;
    layer3_outputs(9475) <= 1'b1;
    layer3_outputs(9476) <= not a or b;
    layer3_outputs(9477) <= not (a xor b);
    layer3_outputs(9478) <= b and not a;
    layer3_outputs(9479) <= b and not a;
    layer3_outputs(9480) <= not b or a;
    layer3_outputs(9481) <= not b or a;
    layer3_outputs(9482) <= a and not b;
    layer3_outputs(9483) <= not a;
    layer3_outputs(9484) <= a;
    layer3_outputs(9485) <= not a or b;
    layer3_outputs(9486) <= 1'b0;
    layer3_outputs(9487) <= not (a or b);
    layer3_outputs(9488) <= b and not a;
    layer3_outputs(9489) <= not (a and b);
    layer3_outputs(9490) <= not b or a;
    layer3_outputs(9491) <= not b or a;
    layer3_outputs(9492) <= a and b;
    layer3_outputs(9493) <= 1'b0;
    layer3_outputs(9494) <= b and not a;
    layer3_outputs(9495) <= a or b;
    layer3_outputs(9496) <= 1'b1;
    layer3_outputs(9497) <= not (a and b);
    layer3_outputs(9498) <= not a;
    layer3_outputs(9499) <= not b or a;
    layer3_outputs(9500) <= 1'b0;
    layer3_outputs(9501) <= not a or b;
    layer3_outputs(9502) <= not b;
    layer3_outputs(9503) <= a;
    layer3_outputs(9504) <= b;
    layer3_outputs(9505) <= a and not b;
    layer3_outputs(9506) <= a and not b;
    layer3_outputs(9507) <= a;
    layer3_outputs(9508) <= not b or a;
    layer3_outputs(9509) <= 1'b0;
    layer3_outputs(9510) <= a or b;
    layer3_outputs(9511) <= not (a or b);
    layer3_outputs(9512) <= b;
    layer3_outputs(9513) <= not b;
    layer3_outputs(9514) <= a or b;
    layer3_outputs(9515) <= b and not a;
    layer3_outputs(9516) <= not a;
    layer3_outputs(9517) <= not (a and b);
    layer3_outputs(9518) <= a;
    layer3_outputs(9519) <= b and not a;
    layer3_outputs(9520) <= a or b;
    layer3_outputs(9521) <= 1'b1;
    layer3_outputs(9522) <= not a;
    layer3_outputs(9523) <= a and not b;
    layer3_outputs(9524) <= a and not b;
    layer3_outputs(9525) <= a and not b;
    layer3_outputs(9526) <= not b or a;
    layer3_outputs(9527) <= not (a and b);
    layer3_outputs(9528) <= 1'b1;
    layer3_outputs(9529) <= a and not b;
    layer3_outputs(9530) <= a xor b;
    layer3_outputs(9531) <= b;
    layer3_outputs(9532) <= a xor b;
    layer3_outputs(9533) <= a and b;
    layer3_outputs(9534) <= a;
    layer3_outputs(9535) <= b and not a;
    layer3_outputs(9536) <= b and not a;
    layer3_outputs(9537) <= 1'b1;
    layer3_outputs(9538) <= a and not b;
    layer3_outputs(9539) <= a and b;
    layer3_outputs(9540) <= 1'b1;
    layer3_outputs(9541) <= a or b;
    layer3_outputs(9542) <= a;
    layer3_outputs(9543) <= not b or a;
    layer3_outputs(9544) <= b and not a;
    layer3_outputs(9545) <= a and not b;
    layer3_outputs(9546) <= not b;
    layer3_outputs(9547) <= b;
    layer3_outputs(9548) <= not a or b;
    layer3_outputs(9549) <= not (a xor b);
    layer3_outputs(9550) <= not a or b;
    layer3_outputs(9551) <= 1'b1;
    layer3_outputs(9552) <= not (a and b);
    layer3_outputs(9553) <= not b;
    layer3_outputs(9554) <= not (a or b);
    layer3_outputs(9555) <= a and b;
    layer3_outputs(9556) <= a and not b;
    layer3_outputs(9557) <= not a or b;
    layer3_outputs(9558) <= not (a or b);
    layer3_outputs(9559) <= a;
    layer3_outputs(9560) <= not a;
    layer3_outputs(9561) <= a or b;
    layer3_outputs(9562) <= 1'b0;
    layer3_outputs(9563) <= a and b;
    layer3_outputs(9564) <= a;
    layer3_outputs(9565) <= not (a or b);
    layer3_outputs(9566) <= 1'b1;
    layer3_outputs(9567) <= 1'b0;
    layer3_outputs(9568) <= not (a or b);
    layer3_outputs(9569) <= not b;
    layer3_outputs(9570) <= not (a xor b);
    layer3_outputs(9571) <= not (a or b);
    layer3_outputs(9572) <= not a;
    layer3_outputs(9573) <= not a;
    layer3_outputs(9574) <= a and b;
    layer3_outputs(9575) <= not b or a;
    layer3_outputs(9576) <= a;
    layer3_outputs(9577) <= a and b;
    layer3_outputs(9578) <= not b or a;
    layer3_outputs(9579) <= not (a and b);
    layer3_outputs(9580) <= a and b;
    layer3_outputs(9581) <= b and not a;
    layer3_outputs(9582) <= a;
    layer3_outputs(9583) <= a;
    layer3_outputs(9584) <= not a;
    layer3_outputs(9585) <= a and not b;
    layer3_outputs(9586) <= b and not a;
    layer3_outputs(9587) <= a or b;
    layer3_outputs(9588) <= not (a or b);
    layer3_outputs(9589) <= b;
    layer3_outputs(9590) <= b and not a;
    layer3_outputs(9591) <= b;
    layer3_outputs(9592) <= a xor b;
    layer3_outputs(9593) <= a;
    layer3_outputs(9594) <= a or b;
    layer3_outputs(9595) <= not b or a;
    layer3_outputs(9596) <= not (a and b);
    layer3_outputs(9597) <= a and not b;
    layer3_outputs(9598) <= b and not a;
    layer3_outputs(9599) <= b;
    layer3_outputs(9600) <= not a or b;
    layer3_outputs(9601) <= not a or b;
    layer3_outputs(9602) <= not b or a;
    layer3_outputs(9603) <= a and not b;
    layer3_outputs(9604) <= a;
    layer3_outputs(9605) <= not (a xor b);
    layer3_outputs(9606) <= a or b;
    layer3_outputs(9607) <= 1'b1;
    layer3_outputs(9608) <= 1'b1;
    layer3_outputs(9609) <= a and not b;
    layer3_outputs(9610) <= not b;
    layer3_outputs(9611) <= not (a xor b);
    layer3_outputs(9612) <= not (a and b);
    layer3_outputs(9613) <= not a or b;
    layer3_outputs(9614) <= a xor b;
    layer3_outputs(9615) <= a and not b;
    layer3_outputs(9616) <= 1'b1;
    layer3_outputs(9617) <= a and b;
    layer3_outputs(9618) <= 1'b0;
    layer3_outputs(9619) <= not a;
    layer3_outputs(9620) <= a and not b;
    layer3_outputs(9621) <= 1'b0;
    layer3_outputs(9622) <= a;
    layer3_outputs(9623) <= not (a and b);
    layer3_outputs(9624) <= 1'b1;
    layer3_outputs(9625) <= a and b;
    layer3_outputs(9626) <= a;
    layer3_outputs(9627) <= not b or a;
    layer3_outputs(9628) <= a or b;
    layer3_outputs(9629) <= a or b;
    layer3_outputs(9630) <= not (a and b);
    layer3_outputs(9631) <= 1'b0;
    layer3_outputs(9632) <= b;
    layer3_outputs(9633) <= a and not b;
    layer3_outputs(9634) <= b;
    layer3_outputs(9635) <= not (a and b);
    layer3_outputs(9636) <= a;
    layer3_outputs(9637) <= a xor b;
    layer3_outputs(9638) <= a and b;
    layer3_outputs(9639) <= not b;
    layer3_outputs(9640) <= 1'b1;
    layer3_outputs(9641) <= a xor b;
    layer3_outputs(9642) <= not b;
    layer3_outputs(9643) <= not b or a;
    layer3_outputs(9644) <= not b;
    layer3_outputs(9645) <= a;
    layer3_outputs(9646) <= a and b;
    layer3_outputs(9647) <= b;
    layer3_outputs(9648) <= b and not a;
    layer3_outputs(9649) <= not b;
    layer3_outputs(9650) <= b;
    layer3_outputs(9651) <= not (a or b);
    layer3_outputs(9652) <= 1'b1;
    layer3_outputs(9653) <= not a;
    layer3_outputs(9654) <= b;
    layer3_outputs(9655) <= a or b;
    layer3_outputs(9656) <= a and not b;
    layer3_outputs(9657) <= a and b;
    layer3_outputs(9658) <= not (a and b);
    layer3_outputs(9659) <= not (a or b);
    layer3_outputs(9660) <= not b or a;
    layer3_outputs(9661) <= b and not a;
    layer3_outputs(9662) <= not (a and b);
    layer3_outputs(9663) <= not a;
    layer3_outputs(9664) <= b and not a;
    layer3_outputs(9665) <= a and b;
    layer3_outputs(9666) <= not a or b;
    layer3_outputs(9667) <= not a or b;
    layer3_outputs(9668) <= a and b;
    layer3_outputs(9669) <= b;
    layer3_outputs(9670) <= not (a and b);
    layer3_outputs(9671) <= not a;
    layer3_outputs(9672) <= 1'b1;
    layer3_outputs(9673) <= not (a and b);
    layer3_outputs(9674) <= not (a and b);
    layer3_outputs(9675) <= a or b;
    layer3_outputs(9676) <= b;
    layer3_outputs(9677) <= 1'b1;
    layer3_outputs(9678) <= not b;
    layer3_outputs(9679) <= a;
    layer3_outputs(9680) <= 1'b0;
    layer3_outputs(9681) <= b;
    layer3_outputs(9682) <= a and not b;
    layer3_outputs(9683) <= a and b;
    layer3_outputs(9684) <= b and not a;
    layer3_outputs(9685) <= b and not a;
    layer3_outputs(9686) <= 1'b0;
    layer3_outputs(9687) <= a xor b;
    layer3_outputs(9688) <= not b;
    layer3_outputs(9689) <= a and not b;
    layer3_outputs(9690) <= 1'b0;
    layer3_outputs(9691) <= a xor b;
    layer3_outputs(9692) <= a and not b;
    layer3_outputs(9693) <= a or b;
    layer3_outputs(9694) <= a and b;
    layer3_outputs(9695) <= a;
    layer3_outputs(9696) <= not b;
    layer3_outputs(9697) <= b;
    layer3_outputs(9698) <= not b;
    layer3_outputs(9699) <= a;
    layer3_outputs(9700) <= not b or a;
    layer3_outputs(9701) <= a and not b;
    layer3_outputs(9702) <= a and not b;
    layer3_outputs(9703) <= a and b;
    layer3_outputs(9704) <= a;
    layer3_outputs(9705) <= not (a and b);
    layer3_outputs(9706) <= 1'b1;
    layer3_outputs(9707) <= a;
    layer3_outputs(9708) <= a;
    layer3_outputs(9709) <= a and not b;
    layer3_outputs(9710) <= not a or b;
    layer3_outputs(9711) <= 1'b0;
    layer3_outputs(9712) <= not (a or b);
    layer3_outputs(9713) <= not (a xor b);
    layer3_outputs(9714) <= not b or a;
    layer3_outputs(9715) <= a;
    layer3_outputs(9716) <= a and b;
    layer3_outputs(9717) <= not a or b;
    layer3_outputs(9718) <= b;
    layer3_outputs(9719) <= a or b;
    layer3_outputs(9720) <= not (a and b);
    layer3_outputs(9721) <= a;
    layer3_outputs(9722) <= not (a xor b);
    layer3_outputs(9723) <= a and b;
    layer3_outputs(9724) <= a or b;
    layer3_outputs(9725) <= a xor b;
    layer3_outputs(9726) <= 1'b1;
    layer3_outputs(9727) <= a and b;
    layer3_outputs(9728) <= a and b;
    layer3_outputs(9729) <= 1'b1;
    layer3_outputs(9730) <= a or b;
    layer3_outputs(9731) <= a;
    layer3_outputs(9732) <= not (a or b);
    layer3_outputs(9733) <= b;
    layer3_outputs(9734) <= not (a or b);
    layer3_outputs(9735) <= not (a or b);
    layer3_outputs(9736) <= not (a and b);
    layer3_outputs(9737) <= not a;
    layer3_outputs(9738) <= b;
    layer3_outputs(9739) <= not (a or b);
    layer3_outputs(9740) <= a;
    layer3_outputs(9741) <= not b or a;
    layer3_outputs(9742) <= b and not a;
    layer3_outputs(9743) <= not a;
    layer3_outputs(9744) <= not b or a;
    layer3_outputs(9745) <= not b;
    layer3_outputs(9746) <= a or b;
    layer3_outputs(9747) <= b and not a;
    layer3_outputs(9748) <= not a;
    layer3_outputs(9749) <= not b;
    layer3_outputs(9750) <= not a or b;
    layer3_outputs(9751) <= b and not a;
    layer3_outputs(9752) <= not b;
    layer3_outputs(9753) <= b;
    layer3_outputs(9754) <= a;
    layer3_outputs(9755) <= not (a xor b);
    layer3_outputs(9756) <= not a;
    layer3_outputs(9757) <= a and b;
    layer3_outputs(9758) <= not a;
    layer3_outputs(9759) <= a and b;
    layer3_outputs(9760) <= not a;
    layer3_outputs(9761) <= a or b;
    layer3_outputs(9762) <= a and b;
    layer3_outputs(9763) <= a or b;
    layer3_outputs(9764) <= not a or b;
    layer3_outputs(9765) <= 1'b1;
    layer3_outputs(9766) <= not a or b;
    layer3_outputs(9767) <= b and not a;
    layer3_outputs(9768) <= 1'b0;
    layer3_outputs(9769) <= not b or a;
    layer3_outputs(9770) <= not (a or b);
    layer3_outputs(9771) <= 1'b0;
    layer3_outputs(9772) <= not b;
    layer3_outputs(9773) <= 1'b0;
    layer3_outputs(9774) <= not (a and b);
    layer3_outputs(9775) <= 1'b0;
    layer3_outputs(9776) <= not a or b;
    layer3_outputs(9777) <= not b;
    layer3_outputs(9778) <= b and not a;
    layer3_outputs(9779) <= a or b;
    layer3_outputs(9780) <= 1'b0;
    layer3_outputs(9781) <= 1'b1;
    layer3_outputs(9782) <= 1'b0;
    layer3_outputs(9783) <= not (a xor b);
    layer3_outputs(9784) <= b and not a;
    layer3_outputs(9785) <= not b;
    layer3_outputs(9786) <= b;
    layer3_outputs(9787) <= not (a or b);
    layer3_outputs(9788) <= b and not a;
    layer3_outputs(9789) <= not (a and b);
    layer3_outputs(9790) <= a or b;
    layer3_outputs(9791) <= a and b;
    layer3_outputs(9792) <= b and not a;
    layer3_outputs(9793) <= b;
    layer3_outputs(9794) <= not b or a;
    layer3_outputs(9795) <= 1'b0;
    layer3_outputs(9796) <= b and not a;
    layer3_outputs(9797) <= a and b;
    layer3_outputs(9798) <= a and b;
    layer3_outputs(9799) <= a and b;
    layer3_outputs(9800) <= a;
    layer3_outputs(9801) <= b and not a;
    layer3_outputs(9802) <= a xor b;
    layer3_outputs(9803) <= a;
    layer3_outputs(9804) <= a or b;
    layer3_outputs(9805) <= a and not b;
    layer3_outputs(9806) <= a or b;
    layer3_outputs(9807) <= a and not b;
    layer3_outputs(9808) <= not (a and b);
    layer3_outputs(9809) <= not a or b;
    layer3_outputs(9810) <= 1'b0;
    layer3_outputs(9811) <= not b or a;
    layer3_outputs(9812) <= 1'b0;
    layer3_outputs(9813) <= a and not b;
    layer3_outputs(9814) <= not (a and b);
    layer3_outputs(9815) <= not b or a;
    layer3_outputs(9816) <= not (a or b);
    layer3_outputs(9817) <= b;
    layer3_outputs(9818) <= not a;
    layer3_outputs(9819) <= a or b;
    layer3_outputs(9820) <= a xor b;
    layer3_outputs(9821) <= not (a and b);
    layer3_outputs(9822) <= a and not b;
    layer3_outputs(9823) <= not a or b;
    layer3_outputs(9824) <= a and b;
    layer3_outputs(9825) <= 1'b1;
    layer3_outputs(9826) <= b;
    layer3_outputs(9827) <= not (a and b);
    layer3_outputs(9828) <= not b;
    layer3_outputs(9829) <= a and b;
    layer3_outputs(9830) <= not b or a;
    layer3_outputs(9831) <= 1'b0;
    layer3_outputs(9832) <= 1'b0;
    layer3_outputs(9833) <= a or b;
    layer3_outputs(9834) <= a and not b;
    layer3_outputs(9835) <= a;
    layer3_outputs(9836) <= not a;
    layer3_outputs(9837) <= 1'b1;
    layer3_outputs(9838) <= 1'b0;
    layer3_outputs(9839) <= a and b;
    layer3_outputs(9840) <= a and not b;
    layer3_outputs(9841) <= a and b;
    layer3_outputs(9842) <= a and b;
    layer3_outputs(9843) <= a xor b;
    layer3_outputs(9844) <= not (a and b);
    layer3_outputs(9845) <= a;
    layer3_outputs(9846) <= not a or b;
    layer3_outputs(9847) <= 1'b1;
    layer3_outputs(9848) <= a;
    layer3_outputs(9849) <= not (a or b);
    layer3_outputs(9850) <= not a or b;
    layer3_outputs(9851) <= a and b;
    layer3_outputs(9852) <= not b;
    layer3_outputs(9853) <= not a;
    layer3_outputs(9854) <= not a;
    layer3_outputs(9855) <= not b;
    layer3_outputs(9856) <= not (a or b);
    layer3_outputs(9857) <= not b or a;
    layer3_outputs(9858) <= not a or b;
    layer3_outputs(9859) <= not (a or b);
    layer3_outputs(9860) <= b and not a;
    layer3_outputs(9861) <= b;
    layer3_outputs(9862) <= a and b;
    layer3_outputs(9863) <= a and b;
    layer3_outputs(9864) <= a and not b;
    layer3_outputs(9865) <= b;
    layer3_outputs(9866) <= a;
    layer3_outputs(9867) <= not b;
    layer3_outputs(9868) <= a and b;
    layer3_outputs(9869) <= not a or b;
    layer3_outputs(9870) <= 1'b0;
    layer3_outputs(9871) <= not a or b;
    layer3_outputs(9872) <= b;
    layer3_outputs(9873) <= a and not b;
    layer3_outputs(9874) <= a or b;
    layer3_outputs(9875) <= a and b;
    layer3_outputs(9876) <= b;
    layer3_outputs(9877) <= 1'b1;
    layer3_outputs(9878) <= 1'b1;
    layer3_outputs(9879) <= a;
    layer3_outputs(9880) <= a xor b;
    layer3_outputs(9881) <= a and b;
    layer3_outputs(9882) <= not (a xor b);
    layer3_outputs(9883) <= 1'b1;
    layer3_outputs(9884) <= not (a xor b);
    layer3_outputs(9885) <= a;
    layer3_outputs(9886) <= b and not a;
    layer3_outputs(9887) <= 1'b0;
    layer3_outputs(9888) <= not b or a;
    layer3_outputs(9889) <= not a or b;
    layer3_outputs(9890) <= not a;
    layer3_outputs(9891) <= 1'b0;
    layer3_outputs(9892) <= not b;
    layer3_outputs(9893) <= not b;
    layer3_outputs(9894) <= 1'b0;
    layer3_outputs(9895) <= b;
    layer3_outputs(9896) <= b;
    layer3_outputs(9897) <= b;
    layer3_outputs(9898) <= a and not b;
    layer3_outputs(9899) <= not b or a;
    layer3_outputs(9900) <= not a;
    layer3_outputs(9901) <= a and not b;
    layer3_outputs(9902) <= a and not b;
    layer3_outputs(9903) <= a or b;
    layer3_outputs(9904) <= b and not a;
    layer3_outputs(9905) <= a and b;
    layer3_outputs(9906) <= not a or b;
    layer3_outputs(9907) <= not (a or b);
    layer3_outputs(9908) <= a or b;
    layer3_outputs(9909) <= not (a and b);
    layer3_outputs(9910) <= not (a xor b);
    layer3_outputs(9911) <= b and not a;
    layer3_outputs(9912) <= 1'b1;
    layer3_outputs(9913) <= not b;
    layer3_outputs(9914) <= not (a or b);
    layer3_outputs(9915) <= not b;
    layer3_outputs(9916) <= not b;
    layer3_outputs(9917) <= 1'b1;
    layer3_outputs(9918) <= a or b;
    layer3_outputs(9919) <= 1'b0;
    layer3_outputs(9920) <= not (a and b);
    layer3_outputs(9921) <= b and not a;
    layer3_outputs(9922) <= b and not a;
    layer3_outputs(9923) <= a;
    layer3_outputs(9924) <= not b or a;
    layer3_outputs(9925) <= a and b;
    layer3_outputs(9926) <= not a;
    layer3_outputs(9927) <= not a;
    layer3_outputs(9928) <= a;
    layer3_outputs(9929) <= 1'b0;
    layer3_outputs(9930) <= not b or a;
    layer3_outputs(9931) <= not (a and b);
    layer3_outputs(9932) <= 1'b1;
    layer3_outputs(9933) <= b and not a;
    layer3_outputs(9934) <= not a;
    layer3_outputs(9935) <= b;
    layer3_outputs(9936) <= not b;
    layer3_outputs(9937) <= a and not b;
    layer3_outputs(9938) <= not a;
    layer3_outputs(9939) <= not (a and b);
    layer3_outputs(9940) <= 1'b0;
    layer3_outputs(9941) <= 1'b0;
    layer3_outputs(9942) <= b and not a;
    layer3_outputs(9943) <= a;
    layer3_outputs(9944) <= not (a or b);
    layer3_outputs(9945) <= not (a or b);
    layer3_outputs(9946) <= not (a and b);
    layer3_outputs(9947) <= a and b;
    layer3_outputs(9948) <= b and not a;
    layer3_outputs(9949) <= 1'b1;
    layer3_outputs(9950) <= not a;
    layer3_outputs(9951) <= not (a or b);
    layer3_outputs(9952) <= not (a and b);
    layer3_outputs(9953) <= not a or b;
    layer3_outputs(9954) <= 1'b1;
    layer3_outputs(9955) <= not (a and b);
    layer3_outputs(9956) <= 1'b0;
    layer3_outputs(9957) <= 1'b1;
    layer3_outputs(9958) <= not a;
    layer3_outputs(9959) <= 1'b1;
    layer3_outputs(9960) <= a or b;
    layer3_outputs(9961) <= not b or a;
    layer3_outputs(9962) <= not a;
    layer3_outputs(9963) <= a;
    layer3_outputs(9964) <= not (a and b);
    layer3_outputs(9965) <= b and not a;
    layer3_outputs(9966) <= not (a or b);
    layer3_outputs(9967) <= 1'b0;
    layer3_outputs(9968) <= a and b;
    layer3_outputs(9969) <= not (a or b);
    layer3_outputs(9970) <= 1'b1;
    layer3_outputs(9971) <= not a;
    layer3_outputs(9972) <= b;
    layer3_outputs(9973) <= a and b;
    layer3_outputs(9974) <= not (a and b);
    layer3_outputs(9975) <= not a;
    layer3_outputs(9976) <= not b;
    layer3_outputs(9977) <= a;
    layer3_outputs(9978) <= not a or b;
    layer3_outputs(9979) <= a or b;
    layer3_outputs(9980) <= b;
    layer3_outputs(9981) <= a and not b;
    layer3_outputs(9982) <= a and b;
    layer3_outputs(9983) <= 1'b0;
    layer3_outputs(9984) <= a;
    layer3_outputs(9985) <= b;
    layer3_outputs(9986) <= not a or b;
    layer3_outputs(9987) <= not b or a;
    layer3_outputs(9988) <= not a;
    layer3_outputs(9989) <= not a;
    layer3_outputs(9990) <= b;
    layer3_outputs(9991) <= a or b;
    layer3_outputs(9992) <= not (a and b);
    layer3_outputs(9993) <= not (a or b);
    layer3_outputs(9994) <= not b or a;
    layer3_outputs(9995) <= not a or b;
    layer3_outputs(9996) <= a or b;
    layer3_outputs(9997) <= not a;
    layer3_outputs(9998) <= a or b;
    layer3_outputs(9999) <= not a;
    layer3_outputs(10000) <= b;
    layer3_outputs(10001) <= not (a and b);
    layer3_outputs(10002) <= a and b;
    layer3_outputs(10003) <= not (a or b);
    layer3_outputs(10004) <= b;
    layer3_outputs(10005) <= 1'b1;
    layer3_outputs(10006) <= b;
    layer3_outputs(10007) <= 1'b1;
    layer3_outputs(10008) <= not a;
    layer3_outputs(10009) <= a and not b;
    layer3_outputs(10010) <= not (a and b);
    layer3_outputs(10011) <= b and not a;
    layer3_outputs(10012) <= a and not b;
    layer3_outputs(10013) <= 1'b0;
    layer3_outputs(10014) <= 1'b0;
    layer3_outputs(10015) <= a or b;
    layer3_outputs(10016) <= a and not b;
    layer3_outputs(10017) <= 1'b0;
    layer3_outputs(10018) <= not (a or b);
    layer3_outputs(10019) <= not (a and b);
    layer3_outputs(10020) <= not a;
    layer3_outputs(10021) <= not b or a;
    layer3_outputs(10022) <= not (a and b);
    layer3_outputs(10023) <= b;
    layer3_outputs(10024) <= a or b;
    layer3_outputs(10025) <= 1'b1;
    layer3_outputs(10026) <= 1'b0;
    layer3_outputs(10027) <= not b or a;
    layer3_outputs(10028) <= 1'b0;
    layer3_outputs(10029) <= a;
    layer3_outputs(10030) <= a;
    layer3_outputs(10031) <= 1'b1;
    layer3_outputs(10032) <= a and not b;
    layer3_outputs(10033) <= not (a and b);
    layer3_outputs(10034) <= b and not a;
    layer3_outputs(10035) <= b;
    layer3_outputs(10036) <= b and not a;
    layer3_outputs(10037) <= a and b;
    layer3_outputs(10038) <= a or b;
    layer3_outputs(10039) <= b and not a;
    layer3_outputs(10040) <= 1'b0;
    layer3_outputs(10041) <= 1'b0;
    layer3_outputs(10042) <= 1'b1;
    layer3_outputs(10043) <= 1'b0;
    layer3_outputs(10044) <= b;
    layer3_outputs(10045) <= b;
    layer3_outputs(10046) <= a;
    layer3_outputs(10047) <= not a or b;
    layer3_outputs(10048) <= not (a or b);
    layer3_outputs(10049) <= 1'b0;
    layer3_outputs(10050) <= b;
    layer3_outputs(10051) <= a or b;
    layer3_outputs(10052) <= not a;
    layer3_outputs(10053) <= not b;
    layer3_outputs(10054) <= 1'b0;
    layer3_outputs(10055) <= not (a or b);
    layer3_outputs(10056) <= b;
    layer3_outputs(10057) <= not (a and b);
    layer3_outputs(10058) <= a and not b;
    layer3_outputs(10059) <= a and not b;
    layer3_outputs(10060) <= not a;
    layer3_outputs(10061) <= b;
    layer3_outputs(10062) <= not (a or b);
    layer3_outputs(10063) <= not a;
    layer3_outputs(10064) <= b;
    layer3_outputs(10065) <= not (a and b);
    layer3_outputs(10066) <= b and not a;
    layer3_outputs(10067) <= not (a and b);
    layer3_outputs(10068) <= 1'b1;
    layer3_outputs(10069) <= a xor b;
    layer3_outputs(10070) <= not a or b;
    layer3_outputs(10071) <= b;
    layer3_outputs(10072) <= not (a xor b);
    layer3_outputs(10073) <= a;
    layer3_outputs(10074) <= a and not b;
    layer3_outputs(10075) <= not a;
    layer3_outputs(10076) <= 1'b0;
    layer3_outputs(10077) <= a xor b;
    layer3_outputs(10078) <= not (a and b);
    layer3_outputs(10079) <= not b;
    layer3_outputs(10080) <= not a or b;
    layer3_outputs(10081) <= not a;
    layer3_outputs(10082) <= not a or b;
    layer3_outputs(10083) <= not b;
    layer3_outputs(10084) <= a and not b;
    layer3_outputs(10085) <= a xor b;
    layer3_outputs(10086) <= a and b;
    layer3_outputs(10087) <= 1'b1;
    layer3_outputs(10088) <= not (a and b);
    layer3_outputs(10089) <= b;
    layer3_outputs(10090) <= not b;
    layer3_outputs(10091) <= not b;
    layer3_outputs(10092) <= b;
    layer3_outputs(10093) <= not b or a;
    layer3_outputs(10094) <= 1'b1;
    layer3_outputs(10095) <= 1'b1;
    layer3_outputs(10096) <= not b;
    layer3_outputs(10097) <= not (a or b);
    layer3_outputs(10098) <= b and not a;
    layer3_outputs(10099) <= not (a or b);
    layer3_outputs(10100) <= a xor b;
    layer3_outputs(10101) <= not b;
    layer3_outputs(10102) <= b and not a;
    layer3_outputs(10103) <= not b;
    layer3_outputs(10104) <= not b;
    layer3_outputs(10105) <= b and not a;
    layer3_outputs(10106) <= not b;
    layer3_outputs(10107) <= b;
    layer3_outputs(10108) <= b and not a;
    layer3_outputs(10109) <= a or b;
    layer3_outputs(10110) <= b;
    layer3_outputs(10111) <= a and not b;
    layer3_outputs(10112) <= b and not a;
    layer3_outputs(10113) <= not (a and b);
    layer3_outputs(10114) <= a xor b;
    layer3_outputs(10115) <= 1'b1;
    layer3_outputs(10116) <= 1'b1;
    layer3_outputs(10117) <= not (a and b);
    layer3_outputs(10118) <= not (a or b);
    layer3_outputs(10119) <= b and not a;
    layer3_outputs(10120) <= b and not a;
    layer3_outputs(10121) <= not b;
    layer3_outputs(10122) <= 1'b0;
    layer3_outputs(10123) <= 1'b0;
    layer3_outputs(10124) <= not b or a;
    layer3_outputs(10125) <= 1'b0;
    layer3_outputs(10126) <= a or b;
    layer3_outputs(10127) <= b and not a;
    layer3_outputs(10128) <= a and b;
    layer3_outputs(10129) <= not a or b;
    layer3_outputs(10130) <= not b or a;
    layer3_outputs(10131) <= a;
    layer3_outputs(10132) <= a and not b;
    layer3_outputs(10133) <= not (a and b);
    layer3_outputs(10134) <= 1'b1;
    layer3_outputs(10135) <= 1'b1;
    layer3_outputs(10136) <= 1'b1;
    layer3_outputs(10137) <= a and b;
    layer3_outputs(10138) <= not a or b;
    layer3_outputs(10139) <= not a;
    layer3_outputs(10140) <= not b or a;
    layer3_outputs(10141) <= 1'b1;
    layer3_outputs(10142) <= a;
    layer3_outputs(10143) <= a and not b;
    layer3_outputs(10144) <= 1'b0;
    layer3_outputs(10145) <= not (a or b);
    layer3_outputs(10146) <= a or b;
    layer3_outputs(10147) <= a and b;
    layer3_outputs(10148) <= not a;
    layer3_outputs(10149) <= 1'b0;
    layer3_outputs(10150) <= not a;
    layer3_outputs(10151) <= not (a and b);
    layer3_outputs(10152) <= not (a or b);
    layer3_outputs(10153) <= not a or b;
    layer3_outputs(10154) <= b;
    layer3_outputs(10155) <= b;
    layer3_outputs(10156) <= a or b;
    layer3_outputs(10157) <= b and not a;
    layer3_outputs(10158) <= not b or a;
    layer3_outputs(10159) <= a xor b;
    layer3_outputs(10160) <= 1'b0;
    layer3_outputs(10161) <= a and b;
    layer3_outputs(10162) <= b;
    layer3_outputs(10163) <= b;
    layer3_outputs(10164) <= b;
    layer3_outputs(10165) <= not b;
    layer3_outputs(10166) <= a and b;
    layer3_outputs(10167) <= a xor b;
    layer3_outputs(10168) <= b;
    layer3_outputs(10169) <= a and b;
    layer3_outputs(10170) <= not (a and b);
    layer3_outputs(10171) <= a and b;
    layer3_outputs(10172) <= not a;
    layer3_outputs(10173) <= not (a and b);
    layer3_outputs(10174) <= 1'b1;
    layer3_outputs(10175) <= not (a or b);
    layer3_outputs(10176) <= not (a and b);
    layer3_outputs(10177) <= not (a and b);
    layer3_outputs(10178) <= not a;
    layer3_outputs(10179) <= 1'b0;
    layer3_outputs(10180) <= a and b;
    layer3_outputs(10181) <= a;
    layer3_outputs(10182) <= not b or a;
    layer3_outputs(10183) <= not b or a;
    layer3_outputs(10184) <= 1'b0;
    layer3_outputs(10185) <= a and not b;
    layer3_outputs(10186) <= not (a or b);
    layer3_outputs(10187) <= not (a and b);
    layer3_outputs(10188) <= a xor b;
    layer3_outputs(10189) <= not (a xor b);
    layer3_outputs(10190) <= not (a or b);
    layer3_outputs(10191) <= not (a or b);
    layer3_outputs(10192) <= not (a and b);
    layer3_outputs(10193) <= not b or a;
    layer3_outputs(10194) <= a or b;
    layer3_outputs(10195) <= a;
    layer3_outputs(10196) <= not a;
    layer3_outputs(10197) <= b;
    layer3_outputs(10198) <= not a or b;
    layer3_outputs(10199) <= not b or a;
    layer3_outputs(10200) <= not a or b;
    layer3_outputs(10201) <= b;
    layer3_outputs(10202) <= not b or a;
    layer3_outputs(10203) <= not a;
    layer3_outputs(10204) <= not b;
    layer3_outputs(10205) <= not (a and b);
    layer3_outputs(10206) <= not (a and b);
    layer3_outputs(10207) <= not a;
    layer3_outputs(10208) <= not (a and b);
    layer3_outputs(10209) <= b;
    layer3_outputs(10210) <= not b or a;
    layer3_outputs(10211) <= 1'b0;
    layer3_outputs(10212) <= 1'b0;
    layer3_outputs(10213) <= a and b;
    layer3_outputs(10214) <= not (a and b);
    layer3_outputs(10215) <= a;
    layer3_outputs(10216) <= 1'b0;
    layer3_outputs(10217) <= a and b;
    layer3_outputs(10218) <= a xor b;
    layer3_outputs(10219) <= 1'b0;
    layer3_outputs(10220) <= a and b;
    layer3_outputs(10221) <= a and b;
    layer3_outputs(10222) <= b;
    layer3_outputs(10223) <= not a or b;
    layer3_outputs(10224) <= not b or a;
    layer3_outputs(10225) <= a;
    layer3_outputs(10226) <= not (a and b);
    layer3_outputs(10227) <= not a;
    layer3_outputs(10228) <= a;
    layer3_outputs(10229) <= b and not a;
    layer3_outputs(10230) <= a;
    layer3_outputs(10231) <= b and not a;
    layer3_outputs(10232) <= a or b;
    layer3_outputs(10233) <= a xor b;
    layer3_outputs(10234) <= 1'b0;
    layer3_outputs(10235) <= 1'b1;
    layer3_outputs(10236) <= 1'b1;
    layer3_outputs(10237) <= b and not a;
    layer3_outputs(10238) <= not a or b;
    layer3_outputs(10239) <= 1'b1;
    layer4_outputs(0) <= a or b;
    layer4_outputs(1) <= not b or a;
    layer4_outputs(2) <= 1'b0;
    layer4_outputs(3) <= a xor b;
    layer4_outputs(4) <= a and b;
    layer4_outputs(5) <= not (a or b);
    layer4_outputs(6) <= not a or b;
    layer4_outputs(7) <= 1'b1;
    layer4_outputs(8) <= 1'b1;
    layer4_outputs(9) <= b;
    layer4_outputs(10) <= not (a or b);
    layer4_outputs(11) <= not b;
    layer4_outputs(12) <= a and b;
    layer4_outputs(13) <= a;
    layer4_outputs(14) <= not a;
    layer4_outputs(15) <= not a or b;
    layer4_outputs(16) <= a xor b;
    layer4_outputs(17) <= 1'b1;
    layer4_outputs(18) <= a and not b;
    layer4_outputs(19) <= a;
    layer4_outputs(20) <= not a or b;
    layer4_outputs(21) <= not (a or b);
    layer4_outputs(22) <= not (a and b);
    layer4_outputs(23) <= not (a or b);
    layer4_outputs(24) <= not a;
    layer4_outputs(25) <= b;
    layer4_outputs(26) <= not (a and b);
    layer4_outputs(27) <= 1'b0;
    layer4_outputs(28) <= 1'b1;
    layer4_outputs(29) <= a and not b;
    layer4_outputs(30) <= not (a xor b);
    layer4_outputs(31) <= not (a and b);
    layer4_outputs(32) <= a or b;
    layer4_outputs(33) <= not a;
    layer4_outputs(34) <= a or b;
    layer4_outputs(35) <= b;
    layer4_outputs(36) <= a;
    layer4_outputs(37) <= not b or a;
    layer4_outputs(38) <= a and b;
    layer4_outputs(39) <= a and not b;
    layer4_outputs(40) <= a and b;
    layer4_outputs(41) <= not b;
    layer4_outputs(42) <= not b;
    layer4_outputs(43) <= not (a xor b);
    layer4_outputs(44) <= not (a or b);
    layer4_outputs(45) <= b;
    layer4_outputs(46) <= 1'b1;
    layer4_outputs(47) <= not b or a;
    layer4_outputs(48) <= not (a xor b);
    layer4_outputs(49) <= b;
    layer4_outputs(50) <= a and not b;
    layer4_outputs(51) <= b and not a;
    layer4_outputs(52) <= a and b;
    layer4_outputs(53) <= a and b;
    layer4_outputs(54) <= not a;
    layer4_outputs(55) <= not b or a;
    layer4_outputs(56) <= a and not b;
    layer4_outputs(57) <= a and b;
    layer4_outputs(58) <= b;
    layer4_outputs(59) <= not (a xor b);
    layer4_outputs(60) <= 1'b1;
    layer4_outputs(61) <= not (a or b);
    layer4_outputs(62) <= a and not b;
    layer4_outputs(63) <= a and not b;
    layer4_outputs(64) <= a and not b;
    layer4_outputs(65) <= not a;
    layer4_outputs(66) <= not a or b;
    layer4_outputs(67) <= a and not b;
    layer4_outputs(68) <= not (a or b);
    layer4_outputs(69) <= not (a or b);
    layer4_outputs(70) <= not (a or b);
    layer4_outputs(71) <= not a;
    layer4_outputs(72) <= a and not b;
    layer4_outputs(73) <= not (a and b);
    layer4_outputs(74) <= 1'b1;
    layer4_outputs(75) <= b and not a;
    layer4_outputs(76) <= not b;
    layer4_outputs(77) <= not b or a;
    layer4_outputs(78) <= not (a and b);
    layer4_outputs(79) <= a;
    layer4_outputs(80) <= not (a or b);
    layer4_outputs(81) <= not a;
    layer4_outputs(82) <= not (a or b);
    layer4_outputs(83) <= a and b;
    layer4_outputs(84) <= not (a or b);
    layer4_outputs(85) <= a xor b;
    layer4_outputs(86) <= a and b;
    layer4_outputs(87) <= not b or a;
    layer4_outputs(88) <= a and not b;
    layer4_outputs(89) <= b and not a;
    layer4_outputs(90) <= not b or a;
    layer4_outputs(91) <= b;
    layer4_outputs(92) <= a or b;
    layer4_outputs(93) <= not b;
    layer4_outputs(94) <= a xor b;
    layer4_outputs(95) <= a xor b;
    layer4_outputs(96) <= not a;
    layer4_outputs(97) <= not a;
    layer4_outputs(98) <= not a;
    layer4_outputs(99) <= 1'b1;
    layer4_outputs(100) <= b and not a;
    layer4_outputs(101) <= b and not a;
    layer4_outputs(102) <= not (a xor b);
    layer4_outputs(103) <= not a;
    layer4_outputs(104) <= not (a or b);
    layer4_outputs(105) <= a;
    layer4_outputs(106) <= not b;
    layer4_outputs(107) <= b;
    layer4_outputs(108) <= not b;
    layer4_outputs(109) <= not (a or b);
    layer4_outputs(110) <= b and not a;
    layer4_outputs(111) <= a and b;
    layer4_outputs(112) <= not a or b;
    layer4_outputs(113) <= not (a and b);
    layer4_outputs(114) <= b and not a;
    layer4_outputs(115) <= a and b;
    layer4_outputs(116) <= not b;
    layer4_outputs(117) <= not b;
    layer4_outputs(118) <= a;
    layer4_outputs(119) <= a or b;
    layer4_outputs(120) <= not a or b;
    layer4_outputs(121) <= b;
    layer4_outputs(122) <= b and not a;
    layer4_outputs(123) <= a;
    layer4_outputs(124) <= 1'b0;
    layer4_outputs(125) <= a or b;
    layer4_outputs(126) <= a;
    layer4_outputs(127) <= 1'b0;
    layer4_outputs(128) <= not (a or b);
    layer4_outputs(129) <= not a or b;
    layer4_outputs(130) <= not (a or b);
    layer4_outputs(131) <= b and not a;
    layer4_outputs(132) <= not a;
    layer4_outputs(133) <= b and not a;
    layer4_outputs(134) <= a xor b;
    layer4_outputs(135) <= a;
    layer4_outputs(136) <= a and not b;
    layer4_outputs(137) <= b;
    layer4_outputs(138) <= a and b;
    layer4_outputs(139) <= b;
    layer4_outputs(140) <= 1'b1;
    layer4_outputs(141) <= a or b;
    layer4_outputs(142) <= not b or a;
    layer4_outputs(143) <= 1'b0;
    layer4_outputs(144) <= b;
    layer4_outputs(145) <= a and b;
    layer4_outputs(146) <= not (a and b);
    layer4_outputs(147) <= not a or b;
    layer4_outputs(148) <= not (a and b);
    layer4_outputs(149) <= not b or a;
    layer4_outputs(150) <= not (a and b);
    layer4_outputs(151) <= not (a or b);
    layer4_outputs(152) <= 1'b0;
    layer4_outputs(153) <= a or b;
    layer4_outputs(154) <= a xor b;
    layer4_outputs(155) <= not (a and b);
    layer4_outputs(156) <= a or b;
    layer4_outputs(157) <= not a or b;
    layer4_outputs(158) <= not (a xor b);
    layer4_outputs(159) <= not (a and b);
    layer4_outputs(160) <= a and b;
    layer4_outputs(161) <= not (a or b);
    layer4_outputs(162) <= a xor b;
    layer4_outputs(163) <= b;
    layer4_outputs(164) <= 1'b0;
    layer4_outputs(165) <= not (a and b);
    layer4_outputs(166) <= not (a and b);
    layer4_outputs(167) <= not a;
    layer4_outputs(168) <= b and not a;
    layer4_outputs(169) <= b;
    layer4_outputs(170) <= not a or b;
    layer4_outputs(171) <= a and not b;
    layer4_outputs(172) <= 1'b0;
    layer4_outputs(173) <= a xor b;
    layer4_outputs(174) <= b and not a;
    layer4_outputs(175) <= not b;
    layer4_outputs(176) <= 1'b0;
    layer4_outputs(177) <= not a or b;
    layer4_outputs(178) <= not (a or b);
    layer4_outputs(179) <= not b;
    layer4_outputs(180) <= not (a or b);
    layer4_outputs(181) <= not b or a;
    layer4_outputs(182) <= not (a and b);
    layer4_outputs(183) <= a and b;
    layer4_outputs(184) <= not (a and b);
    layer4_outputs(185) <= not a or b;
    layer4_outputs(186) <= not (a and b);
    layer4_outputs(187) <= not b or a;
    layer4_outputs(188) <= not (a and b);
    layer4_outputs(189) <= not b;
    layer4_outputs(190) <= not b or a;
    layer4_outputs(191) <= a and not b;
    layer4_outputs(192) <= not (a and b);
    layer4_outputs(193) <= not b;
    layer4_outputs(194) <= a or b;
    layer4_outputs(195) <= not (a xor b);
    layer4_outputs(196) <= a and not b;
    layer4_outputs(197) <= b and not a;
    layer4_outputs(198) <= a;
    layer4_outputs(199) <= a;
    layer4_outputs(200) <= not (a and b);
    layer4_outputs(201) <= not (a xor b);
    layer4_outputs(202) <= not a or b;
    layer4_outputs(203) <= 1'b1;
    layer4_outputs(204) <= 1'b0;
    layer4_outputs(205) <= not (a or b);
    layer4_outputs(206) <= a xor b;
    layer4_outputs(207) <= not (a or b);
    layer4_outputs(208) <= not b or a;
    layer4_outputs(209) <= 1'b0;
    layer4_outputs(210) <= 1'b1;
    layer4_outputs(211) <= 1'b1;
    layer4_outputs(212) <= not a or b;
    layer4_outputs(213) <= a;
    layer4_outputs(214) <= a and not b;
    layer4_outputs(215) <= not a;
    layer4_outputs(216) <= b;
    layer4_outputs(217) <= a;
    layer4_outputs(218) <= not (a or b);
    layer4_outputs(219) <= a or b;
    layer4_outputs(220) <= a or b;
    layer4_outputs(221) <= a and not b;
    layer4_outputs(222) <= not (a and b);
    layer4_outputs(223) <= a or b;
    layer4_outputs(224) <= not (a and b);
    layer4_outputs(225) <= not a or b;
    layer4_outputs(226) <= a or b;
    layer4_outputs(227) <= not (a xor b);
    layer4_outputs(228) <= 1'b1;
    layer4_outputs(229) <= a and not b;
    layer4_outputs(230) <= not a;
    layer4_outputs(231) <= not a;
    layer4_outputs(232) <= b;
    layer4_outputs(233) <= not a;
    layer4_outputs(234) <= not (a and b);
    layer4_outputs(235) <= b and not a;
    layer4_outputs(236) <= b;
    layer4_outputs(237) <= a and not b;
    layer4_outputs(238) <= a or b;
    layer4_outputs(239) <= a;
    layer4_outputs(240) <= a or b;
    layer4_outputs(241) <= a and b;
    layer4_outputs(242) <= not a;
    layer4_outputs(243) <= a xor b;
    layer4_outputs(244) <= not b or a;
    layer4_outputs(245) <= not (a and b);
    layer4_outputs(246) <= a and not b;
    layer4_outputs(247) <= a xor b;
    layer4_outputs(248) <= not a;
    layer4_outputs(249) <= not (a xor b);
    layer4_outputs(250) <= not a;
    layer4_outputs(251) <= not a or b;
    layer4_outputs(252) <= a and not b;
    layer4_outputs(253) <= a and not b;
    layer4_outputs(254) <= a and b;
    layer4_outputs(255) <= a;
    layer4_outputs(256) <= b;
    layer4_outputs(257) <= b and not a;
    layer4_outputs(258) <= b and not a;
    layer4_outputs(259) <= a;
    layer4_outputs(260) <= 1'b0;
    layer4_outputs(261) <= not (a and b);
    layer4_outputs(262) <= a or b;
    layer4_outputs(263) <= b and not a;
    layer4_outputs(264) <= not b or a;
    layer4_outputs(265) <= a and b;
    layer4_outputs(266) <= not b or a;
    layer4_outputs(267) <= not b or a;
    layer4_outputs(268) <= b and not a;
    layer4_outputs(269) <= b and not a;
    layer4_outputs(270) <= not a or b;
    layer4_outputs(271) <= a and not b;
    layer4_outputs(272) <= not b;
    layer4_outputs(273) <= not b;
    layer4_outputs(274) <= not (a or b);
    layer4_outputs(275) <= 1'b1;
    layer4_outputs(276) <= not (a and b);
    layer4_outputs(277) <= a;
    layer4_outputs(278) <= not (a and b);
    layer4_outputs(279) <= a;
    layer4_outputs(280) <= 1'b0;
    layer4_outputs(281) <= b;
    layer4_outputs(282) <= not (a or b);
    layer4_outputs(283) <= not a;
    layer4_outputs(284) <= not b;
    layer4_outputs(285) <= not b or a;
    layer4_outputs(286) <= a;
    layer4_outputs(287) <= a and not b;
    layer4_outputs(288) <= a and b;
    layer4_outputs(289) <= a;
    layer4_outputs(290) <= 1'b0;
    layer4_outputs(291) <= a or b;
    layer4_outputs(292) <= not b or a;
    layer4_outputs(293) <= a and not b;
    layer4_outputs(294) <= not b;
    layer4_outputs(295) <= 1'b0;
    layer4_outputs(296) <= a and not b;
    layer4_outputs(297) <= b;
    layer4_outputs(298) <= not (a or b);
    layer4_outputs(299) <= not (a or b);
    layer4_outputs(300) <= not (a or b);
    layer4_outputs(301) <= 1'b0;
    layer4_outputs(302) <= not b;
    layer4_outputs(303) <= not a;
    layer4_outputs(304) <= 1'b0;
    layer4_outputs(305) <= not (a and b);
    layer4_outputs(306) <= b;
    layer4_outputs(307) <= not a or b;
    layer4_outputs(308) <= 1'b0;
    layer4_outputs(309) <= 1'b0;
    layer4_outputs(310) <= a and b;
    layer4_outputs(311) <= not (a xor b);
    layer4_outputs(312) <= b and not a;
    layer4_outputs(313) <= not b;
    layer4_outputs(314) <= not (a or b);
    layer4_outputs(315) <= not a or b;
    layer4_outputs(316) <= not a;
    layer4_outputs(317) <= not (a or b);
    layer4_outputs(318) <= a and b;
    layer4_outputs(319) <= a;
    layer4_outputs(320) <= b and not a;
    layer4_outputs(321) <= b and not a;
    layer4_outputs(322) <= not b or a;
    layer4_outputs(323) <= a;
    layer4_outputs(324) <= not b;
    layer4_outputs(325) <= not a or b;
    layer4_outputs(326) <= not b or a;
    layer4_outputs(327) <= not (a and b);
    layer4_outputs(328) <= b and not a;
    layer4_outputs(329) <= not b;
    layer4_outputs(330) <= 1'b0;
    layer4_outputs(331) <= not (a and b);
    layer4_outputs(332) <= 1'b1;
    layer4_outputs(333) <= not (a and b);
    layer4_outputs(334) <= not (a or b);
    layer4_outputs(335) <= not b or a;
    layer4_outputs(336) <= a or b;
    layer4_outputs(337) <= not (a and b);
    layer4_outputs(338) <= 1'b0;
    layer4_outputs(339) <= a and b;
    layer4_outputs(340) <= b;
    layer4_outputs(341) <= 1'b0;
    layer4_outputs(342) <= b and not a;
    layer4_outputs(343) <= not a;
    layer4_outputs(344) <= a xor b;
    layer4_outputs(345) <= a or b;
    layer4_outputs(346) <= not b or a;
    layer4_outputs(347) <= 1'b1;
    layer4_outputs(348) <= not a;
    layer4_outputs(349) <= not a or b;
    layer4_outputs(350) <= a and not b;
    layer4_outputs(351) <= not a;
    layer4_outputs(352) <= not (a or b);
    layer4_outputs(353) <= a and b;
    layer4_outputs(354) <= not a or b;
    layer4_outputs(355) <= not (a or b);
    layer4_outputs(356) <= a or b;
    layer4_outputs(357) <= 1'b1;
    layer4_outputs(358) <= not (a and b);
    layer4_outputs(359) <= not b;
    layer4_outputs(360) <= b;
    layer4_outputs(361) <= b and not a;
    layer4_outputs(362) <= not (a and b);
    layer4_outputs(363) <= not a;
    layer4_outputs(364) <= a and b;
    layer4_outputs(365) <= 1'b1;
    layer4_outputs(366) <= b and not a;
    layer4_outputs(367) <= not (a xor b);
    layer4_outputs(368) <= a or b;
    layer4_outputs(369) <= a;
    layer4_outputs(370) <= not b;
    layer4_outputs(371) <= b and not a;
    layer4_outputs(372) <= a and b;
    layer4_outputs(373) <= not (a xor b);
    layer4_outputs(374) <= a and b;
    layer4_outputs(375) <= a and not b;
    layer4_outputs(376) <= a or b;
    layer4_outputs(377) <= not a;
    layer4_outputs(378) <= not b or a;
    layer4_outputs(379) <= 1'b0;
    layer4_outputs(380) <= not b or a;
    layer4_outputs(381) <= a;
    layer4_outputs(382) <= a or b;
    layer4_outputs(383) <= a and b;
    layer4_outputs(384) <= a;
    layer4_outputs(385) <= a or b;
    layer4_outputs(386) <= a and not b;
    layer4_outputs(387) <= not (a or b);
    layer4_outputs(388) <= not (a and b);
    layer4_outputs(389) <= not b;
    layer4_outputs(390) <= not a or b;
    layer4_outputs(391) <= a and not b;
    layer4_outputs(392) <= not b or a;
    layer4_outputs(393) <= a;
    layer4_outputs(394) <= not a or b;
    layer4_outputs(395) <= a xor b;
    layer4_outputs(396) <= not (a xor b);
    layer4_outputs(397) <= not a or b;
    layer4_outputs(398) <= not (a or b);
    layer4_outputs(399) <= not a or b;
    layer4_outputs(400) <= not a or b;
    layer4_outputs(401) <= not (a or b);
    layer4_outputs(402) <= not b or a;
    layer4_outputs(403) <= a;
    layer4_outputs(404) <= a;
    layer4_outputs(405) <= 1'b1;
    layer4_outputs(406) <= not b;
    layer4_outputs(407) <= a;
    layer4_outputs(408) <= not b or a;
    layer4_outputs(409) <= not (a and b);
    layer4_outputs(410) <= not b;
    layer4_outputs(411) <= not a;
    layer4_outputs(412) <= a or b;
    layer4_outputs(413) <= not a or b;
    layer4_outputs(414) <= a and b;
    layer4_outputs(415) <= a or b;
    layer4_outputs(416) <= 1'b0;
    layer4_outputs(417) <= not (a and b);
    layer4_outputs(418) <= not (a or b);
    layer4_outputs(419) <= not (a xor b);
    layer4_outputs(420) <= a;
    layer4_outputs(421) <= not (a or b);
    layer4_outputs(422) <= not (a and b);
    layer4_outputs(423) <= not (a and b);
    layer4_outputs(424) <= a and b;
    layer4_outputs(425) <= a xor b;
    layer4_outputs(426) <= a or b;
    layer4_outputs(427) <= not a or b;
    layer4_outputs(428) <= a and not b;
    layer4_outputs(429) <= a or b;
    layer4_outputs(430) <= not (a and b);
    layer4_outputs(431) <= a;
    layer4_outputs(432) <= a or b;
    layer4_outputs(433) <= a or b;
    layer4_outputs(434) <= not a or b;
    layer4_outputs(435) <= b and not a;
    layer4_outputs(436) <= not (a xor b);
    layer4_outputs(437) <= b and not a;
    layer4_outputs(438) <= not a or b;
    layer4_outputs(439) <= 1'b1;
    layer4_outputs(440) <= a and b;
    layer4_outputs(441) <= a and b;
    layer4_outputs(442) <= a;
    layer4_outputs(443) <= not (a and b);
    layer4_outputs(444) <= not a;
    layer4_outputs(445) <= a or b;
    layer4_outputs(446) <= a and not b;
    layer4_outputs(447) <= b;
    layer4_outputs(448) <= a and not b;
    layer4_outputs(449) <= not b;
    layer4_outputs(450) <= not a;
    layer4_outputs(451) <= not (a and b);
    layer4_outputs(452) <= a or b;
    layer4_outputs(453) <= not a or b;
    layer4_outputs(454) <= b and not a;
    layer4_outputs(455) <= 1'b1;
    layer4_outputs(456) <= not (a xor b);
    layer4_outputs(457) <= a and not b;
    layer4_outputs(458) <= not a or b;
    layer4_outputs(459) <= a or b;
    layer4_outputs(460) <= b and not a;
    layer4_outputs(461) <= b;
    layer4_outputs(462) <= not (a and b);
    layer4_outputs(463) <= b;
    layer4_outputs(464) <= not (a xor b);
    layer4_outputs(465) <= a;
    layer4_outputs(466) <= not (a and b);
    layer4_outputs(467) <= not a;
    layer4_outputs(468) <= b and not a;
    layer4_outputs(469) <= a or b;
    layer4_outputs(470) <= 1'b1;
    layer4_outputs(471) <= b and not a;
    layer4_outputs(472) <= 1'b0;
    layer4_outputs(473) <= not b or a;
    layer4_outputs(474) <= not (a or b);
    layer4_outputs(475) <= 1'b1;
    layer4_outputs(476) <= not b or a;
    layer4_outputs(477) <= not b;
    layer4_outputs(478) <= not a;
    layer4_outputs(479) <= not (a or b);
    layer4_outputs(480) <= not b or a;
    layer4_outputs(481) <= b;
    layer4_outputs(482) <= not a;
    layer4_outputs(483) <= a and b;
    layer4_outputs(484) <= not a or b;
    layer4_outputs(485) <= not b;
    layer4_outputs(486) <= not a;
    layer4_outputs(487) <= b and not a;
    layer4_outputs(488) <= b;
    layer4_outputs(489) <= a and not b;
    layer4_outputs(490) <= a or b;
    layer4_outputs(491) <= not a or b;
    layer4_outputs(492) <= not a or b;
    layer4_outputs(493) <= not b;
    layer4_outputs(494) <= not b;
    layer4_outputs(495) <= a or b;
    layer4_outputs(496) <= a xor b;
    layer4_outputs(497) <= a;
    layer4_outputs(498) <= a xor b;
    layer4_outputs(499) <= not a or b;
    layer4_outputs(500) <= b and not a;
    layer4_outputs(501) <= 1'b0;
    layer4_outputs(502) <= a and b;
    layer4_outputs(503) <= not b or a;
    layer4_outputs(504) <= not b or a;
    layer4_outputs(505) <= 1'b0;
    layer4_outputs(506) <= not (a and b);
    layer4_outputs(507) <= a and b;
    layer4_outputs(508) <= not (a or b);
    layer4_outputs(509) <= not a or b;
    layer4_outputs(510) <= a and not b;
    layer4_outputs(511) <= b and not a;
    layer4_outputs(512) <= a and not b;
    layer4_outputs(513) <= a and not b;
    layer4_outputs(514) <= not (a or b);
    layer4_outputs(515) <= not b;
    layer4_outputs(516) <= a;
    layer4_outputs(517) <= a;
    layer4_outputs(518) <= not a or b;
    layer4_outputs(519) <= a and b;
    layer4_outputs(520) <= a and b;
    layer4_outputs(521) <= not (a xor b);
    layer4_outputs(522) <= not b or a;
    layer4_outputs(523) <= a;
    layer4_outputs(524) <= not (a and b);
    layer4_outputs(525) <= not b;
    layer4_outputs(526) <= not (a or b);
    layer4_outputs(527) <= a and not b;
    layer4_outputs(528) <= a or b;
    layer4_outputs(529) <= not (a xor b);
    layer4_outputs(530) <= b and not a;
    layer4_outputs(531) <= b and not a;
    layer4_outputs(532) <= 1'b0;
    layer4_outputs(533) <= a and not b;
    layer4_outputs(534) <= b;
    layer4_outputs(535) <= not a;
    layer4_outputs(536) <= not a;
    layer4_outputs(537) <= not (a or b);
    layer4_outputs(538) <= 1'b1;
    layer4_outputs(539) <= a xor b;
    layer4_outputs(540) <= a and b;
    layer4_outputs(541) <= 1'b0;
    layer4_outputs(542) <= not b or a;
    layer4_outputs(543) <= not (a or b);
    layer4_outputs(544) <= b;
    layer4_outputs(545) <= a and not b;
    layer4_outputs(546) <= not b;
    layer4_outputs(547) <= not b;
    layer4_outputs(548) <= a and b;
    layer4_outputs(549) <= not a;
    layer4_outputs(550) <= not a or b;
    layer4_outputs(551) <= b and not a;
    layer4_outputs(552) <= a xor b;
    layer4_outputs(553) <= a;
    layer4_outputs(554) <= b and not a;
    layer4_outputs(555) <= b;
    layer4_outputs(556) <= 1'b0;
    layer4_outputs(557) <= not a or b;
    layer4_outputs(558) <= a and not b;
    layer4_outputs(559) <= not (a xor b);
    layer4_outputs(560) <= not b;
    layer4_outputs(561) <= b and not a;
    layer4_outputs(562) <= a xor b;
    layer4_outputs(563) <= a and not b;
    layer4_outputs(564) <= a xor b;
    layer4_outputs(565) <= not a;
    layer4_outputs(566) <= not a or b;
    layer4_outputs(567) <= not (a and b);
    layer4_outputs(568) <= b and not a;
    layer4_outputs(569) <= a xor b;
    layer4_outputs(570) <= not a;
    layer4_outputs(571) <= not a;
    layer4_outputs(572) <= a and not b;
    layer4_outputs(573) <= 1'b1;
    layer4_outputs(574) <= not (a or b);
    layer4_outputs(575) <= a or b;
    layer4_outputs(576) <= not a;
    layer4_outputs(577) <= not a or b;
    layer4_outputs(578) <= not a;
    layer4_outputs(579) <= not b or a;
    layer4_outputs(580) <= b;
    layer4_outputs(581) <= not (a or b);
    layer4_outputs(582) <= not (a and b);
    layer4_outputs(583) <= b and not a;
    layer4_outputs(584) <= not a or b;
    layer4_outputs(585) <= a;
    layer4_outputs(586) <= a or b;
    layer4_outputs(587) <= 1'b1;
    layer4_outputs(588) <= b;
    layer4_outputs(589) <= not a or b;
    layer4_outputs(590) <= a and b;
    layer4_outputs(591) <= a and not b;
    layer4_outputs(592) <= b and not a;
    layer4_outputs(593) <= 1'b0;
    layer4_outputs(594) <= not b or a;
    layer4_outputs(595) <= b;
    layer4_outputs(596) <= not a or b;
    layer4_outputs(597) <= a;
    layer4_outputs(598) <= 1'b0;
    layer4_outputs(599) <= b and not a;
    layer4_outputs(600) <= not (a and b);
    layer4_outputs(601) <= 1'b0;
    layer4_outputs(602) <= a and not b;
    layer4_outputs(603) <= a or b;
    layer4_outputs(604) <= not b or a;
    layer4_outputs(605) <= not (a or b);
    layer4_outputs(606) <= not b;
    layer4_outputs(607) <= not (a and b);
    layer4_outputs(608) <= 1'b0;
    layer4_outputs(609) <= a and not b;
    layer4_outputs(610) <= not (a xor b);
    layer4_outputs(611) <= a and b;
    layer4_outputs(612) <= a and not b;
    layer4_outputs(613) <= not a or b;
    layer4_outputs(614) <= a and b;
    layer4_outputs(615) <= not (a or b);
    layer4_outputs(616) <= a;
    layer4_outputs(617) <= 1'b1;
    layer4_outputs(618) <= not b;
    layer4_outputs(619) <= a and b;
    layer4_outputs(620) <= not (a and b);
    layer4_outputs(621) <= a xor b;
    layer4_outputs(622) <= a and not b;
    layer4_outputs(623) <= 1'b0;
    layer4_outputs(624) <= not b or a;
    layer4_outputs(625) <= a or b;
    layer4_outputs(626) <= not b;
    layer4_outputs(627) <= a;
    layer4_outputs(628) <= not (a and b);
    layer4_outputs(629) <= not b;
    layer4_outputs(630) <= a;
    layer4_outputs(631) <= 1'b1;
    layer4_outputs(632) <= 1'b1;
    layer4_outputs(633) <= a and not b;
    layer4_outputs(634) <= b and not a;
    layer4_outputs(635) <= not a or b;
    layer4_outputs(636) <= not (a or b);
    layer4_outputs(637) <= not a;
    layer4_outputs(638) <= not (a or b);
    layer4_outputs(639) <= not b;
    layer4_outputs(640) <= b;
    layer4_outputs(641) <= not b;
    layer4_outputs(642) <= a and b;
    layer4_outputs(643) <= a;
    layer4_outputs(644) <= a and not b;
    layer4_outputs(645) <= 1'b0;
    layer4_outputs(646) <= not b;
    layer4_outputs(647) <= not (a xor b);
    layer4_outputs(648) <= not (a and b);
    layer4_outputs(649) <= b;
    layer4_outputs(650) <= not (a or b);
    layer4_outputs(651) <= b and not a;
    layer4_outputs(652) <= not b or a;
    layer4_outputs(653) <= not a;
    layer4_outputs(654) <= 1'b1;
    layer4_outputs(655) <= not a or b;
    layer4_outputs(656) <= not b or a;
    layer4_outputs(657) <= not a;
    layer4_outputs(658) <= 1'b0;
    layer4_outputs(659) <= b;
    layer4_outputs(660) <= not b or a;
    layer4_outputs(661) <= not (a and b);
    layer4_outputs(662) <= a and b;
    layer4_outputs(663) <= not b or a;
    layer4_outputs(664) <= not a or b;
    layer4_outputs(665) <= b;
    layer4_outputs(666) <= 1'b1;
    layer4_outputs(667) <= 1'b1;
    layer4_outputs(668) <= not (a or b);
    layer4_outputs(669) <= not a;
    layer4_outputs(670) <= a and not b;
    layer4_outputs(671) <= not (a or b);
    layer4_outputs(672) <= not b or a;
    layer4_outputs(673) <= not a;
    layer4_outputs(674) <= not b;
    layer4_outputs(675) <= not (a and b);
    layer4_outputs(676) <= a xor b;
    layer4_outputs(677) <= a;
    layer4_outputs(678) <= not (a or b);
    layer4_outputs(679) <= not b;
    layer4_outputs(680) <= 1'b0;
    layer4_outputs(681) <= not a;
    layer4_outputs(682) <= a;
    layer4_outputs(683) <= not b;
    layer4_outputs(684) <= not a or b;
    layer4_outputs(685) <= a xor b;
    layer4_outputs(686) <= not (a or b);
    layer4_outputs(687) <= 1'b1;
    layer4_outputs(688) <= a;
    layer4_outputs(689) <= not a or b;
    layer4_outputs(690) <= not (a or b);
    layer4_outputs(691) <= a and not b;
    layer4_outputs(692) <= 1'b0;
    layer4_outputs(693) <= a xor b;
    layer4_outputs(694) <= a and not b;
    layer4_outputs(695) <= a and not b;
    layer4_outputs(696) <= a and not b;
    layer4_outputs(697) <= not a;
    layer4_outputs(698) <= a xor b;
    layer4_outputs(699) <= not b;
    layer4_outputs(700) <= not a;
    layer4_outputs(701) <= 1'b0;
    layer4_outputs(702) <= not b or a;
    layer4_outputs(703) <= not a;
    layer4_outputs(704) <= 1'b0;
    layer4_outputs(705) <= b and not a;
    layer4_outputs(706) <= b;
    layer4_outputs(707) <= a and b;
    layer4_outputs(708) <= not b or a;
    layer4_outputs(709) <= b;
    layer4_outputs(710) <= a and not b;
    layer4_outputs(711) <= not b;
    layer4_outputs(712) <= not (a xor b);
    layer4_outputs(713) <= a or b;
    layer4_outputs(714) <= b and not a;
    layer4_outputs(715) <= not b or a;
    layer4_outputs(716) <= 1'b0;
    layer4_outputs(717) <= a;
    layer4_outputs(718) <= a and b;
    layer4_outputs(719) <= not a;
    layer4_outputs(720) <= a or b;
    layer4_outputs(721) <= a or b;
    layer4_outputs(722) <= not a or b;
    layer4_outputs(723) <= 1'b1;
    layer4_outputs(724) <= a;
    layer4_outputs(725) <= a or b;
    layer4_outputs(726) <= a xor b;
    layer4_outputs(727) <= 1'b0;
    layer4_outputs(728) <= not (a xor b);
    layer4_outputs(729) <= a or b;
    layer4_outputs(730) <= not b;
    layer4_outputs(731) <= 1'b1;
    layer4_outputs(732) <= 1'b1;
    layer4_outputs(733) <= 1'b0;
    layer4_outputs(734) <= not a or b;
    layer4_outputs(735) <= not (a or b);
    layer4_outputs(736) <= b;
    layer4_outputs(737) <= b and not a;
    layer4_outputs(738) <= not a;
    layer4_outputs(739) <= 1'b0;
    layer4_outputs(740) <= not (a or b);
    layer4_outputs(741) <= b and not a;
    layer4_outputs(742) <= not (a or b);
    layer4_outputs(743) <= b and not a;
    layer4_outputs(744) <= not b or a;
    layer4_outputs(745) <= a and not b;
    layer4_outputs(746) <= a;
    layer4_outputs(747) <= a and b;
    layer4_outputs(748) <= a or b;
    layer4_outputs(749) <= not b;
    layer4_outputs(750) <= a and b;
    layer4_outputs(751) <= a;
    layer4_outputs(752) <= not b or a;
    layer4_outputs(753) <= not (a and b);
    layer4_outputs(754) <= not b;
    layer4_outputs(755) <= a and b;
    layer4_outputs(756) <= not b;
    layer4_outputs(757) <= b;
    layer4_outputs(758) <= a or b;
    layer4_outputs(759) <= not b or a;
    layer4_outputs(760) <= 1'b0;
    layer4_outputs(761) <= not b;
    layer4_outputs(762) <= a and b;
    layer4_outputs(763) <= b and not a;
    layer4_outputs(764) <= not (a or b);
    layer4_outputs(765) <= 1'b0;
    layer4_outputs(766) <= not (a and b);
    layer4_outputs(767) <= 1'b0;
    layer4_outputs(768) <= b;
    layer4_outputs(769) <= a;
    layer4_outputs(770) <= not (a or b);
    layer4_outputs(771) <= not a;
    layer4_outputs(772) <= not b;
    layer4_outputs(773) <= a and b;
    layer4_outputs(774) <= a and b;
    layer4_outputs(775) <= b and not a;
    layer4_outputs(776) <= not (a and b);
    layer4_outputs(777) <= b;
    layer4_outputs(778) <= not b or a;
    layer4_outputs(779) <= a;
    layer4_outputs(780) <= not (a and b);
    layer4_outputs(781) <= a;
    layer4_outputs(782) <= b;
    layer4_outputs(783) <= a and b;
    layer4_outputs(784) <= 1'b0;
    layer4_outputs(785) <= not b;
    layer4_outputs(786) <= 1'b1;
    layer4_outputs(787) <= not b or a;
    layer4_outputs(788) <= not (a or b);
    layer4_outputs(789) <= b and not a;
    layer4_outputs(790) <= not (a xor b);
    layer4_outputs(791) <= a or b;
    layer4_outputs(792) <= b;
    layer4_outputs(793) <= not (a and b);
    layer4_outputs(794) <= a;
    layer4_outputs(795) <= not b;
    layer4_outputs(796) <= a and not b;
    layer4_outputs(797) <= not a or b;
    layer4_outputs(798) <= not b or a;
    layer4_outputs(799) <= not a or b;
    layer4_outputs(800) <= a;
    layer4_outputs(801) <= 1'b1;
    layer4_outputs(802) <= not a;
    layer4_outputs(803) <= not (a or b);
    layer4_outputs(804) <= not (a or b);
    layer4_outputs(805) <= not a;
    layer4_outputs(806) <= a and b;
    layer4_outputs(807) <= not b;
    layer4_outputs(808) <= not a or b;
    layer4_outputs(809) <= a xor b;
    layer4_outputs(810) <= not b;
    layer4_outputs(811) <= not (a or b);
    layer4_outputs(812) <= b;
    layer4_outputs(813) <= not b;
    layer4_outputs(814) <= a;
    layer4_outputs(815) <= a and not b;
    layer4_outputs(816) <= 1'b1;
    layer4_outputs(817) <= not a;
    layer4_outputs(818) <= a or b;
    layer4_outputs(819) <= not b or a;
    layer4_outputs(820) <= not b;
    layer4_outputs(821) <= a or b;
    layer4_outputs(822) <= not a;
    layer4_outputs(823) <= 1'b1;
    layer4_outputs(824) <= not a;
    layer4_outputs(825) <= not a;
    layer4_outputs(826) <= not a;
    layer4_outputs(827) <= a;
    layer4_outputs(828) <= 1'b0;
    layer4_outputs(829) <= not a;
    layer4_outputs(830) <= not a or b;
    layer4_outputs(831) <= 1'b0;
    layer4_outputs(832) <= not a or b;
    layer4_outputs(833) <= not (a and b);
    layer4_outputs(834) <= 1'b0;
    layer4_outputs(835) <= a;
    layer4_outputs(836) <= 1'b1;
    layer4_outputs(837) <= not b;
    layer4_outputs(838) <= a;
    layer4_outputs(839) <= b;
    layer4_outputs(840) <= not b;
    layer4_outputs(841) <= not a;
    layer4_outputs(842) <= not (a and b);
    layer4_outputs(843) <= a;
    layer4_outputs(844) <= not (a or b);
    layer4_outputs(845) <= a or b;
    layer4_outputs(846) <= not (a and b);
    layer4_outputs(847) <= not (a and b);
    layer4_outputs(848) <= not a or b;
    layer4_outputs(849) <= 1'b0;
    layer4_outputs(850) <= not (a or b);
    layer4_outputs(851) <= a and not b;
    layer4_outputs(852) <= a or b;
    layer4_outputs(853) <= 1'b0;
    layer4_outputs(854) <= a or b;
    layer4_outputs(855) <= a or b;
    layer4_outputs(856) <= 1'b0;
    layer4_outputs(857) <= not a;
    layer4_outputs(858) <= not a or b;
    layer4_outputs(859) <= b;
    layer4_outputs(860) <= not b;
    layer4_outputs(861) <= not (a and b);
    layer4_outputs(862) <= b;
    layer4_outputs(863) <= b and not a;
    layer4_outputs(864) <= a and b;
    layer4_outputs(865) <= a xor b;
    layer4_outputs(866) <= not (a or b);
    layer4_outputs(867) <= a;
    layer4_outputs(868) <= 1'b1;
    layer4_outputs(869) <= 1'b1;
    layer4_outputs(870) <= not b or a;
    layer4_outputs(871) <= b and not a;
    layer4_outputs(872) <= a;
    layer4_outputs(873) <= b and not a;
    layer4_outputs(874) <= 1'b1;
    layer4_outputs(875) <= b and not a;
    layer4_outputs(876) <= a and b;
    layer4_outputs(877) <= 1'b1;
    layer4_outputs(878) <= 1'b1;
    layer4_outputs(879) <= a or b;
    layer4_outputs(880) <= a;
    layer4_outputs(881) <= b;
    layer4_outputs(882) <= not a or b;
    layer4_outputs(883) <= not a;
    layer4_outputs(884) <= not (a or b);
    layer4_outputs(885) <= 1'b0;
    layer4_outputs(886) <= not (a and b);
    layer4_outputs(887) <= a or b;
    layer4_outputs(888) <= a and not b;
    layer4_outputs(889) <= a and not b;
    layer4_outputs(890) <= a;
    layer4_outputs(891) <= not b;
    layer4_outputs(892) <= not (a and b);
    layer4_outputs(893) <= a or b;
    layer4_outputs(894) <= 1'b1;
    layer4_outputs(895) <= a and not b;
    layer4_outputs(896) <= 1'b0;
    layer4_outputs(897) <= not b;
    layer4_outputs(898) <= 1'b1;
    layer4_outputs(899) <= 1'b1;
    layer4_outputs(900) <= not b;
    layer4_outputs(901) <= b;
    layer4_outputs(902) <= not a;
    layer4_outputs(903) <= a or b;
    layer4_outputs(904) <= not a;
    layer4_outputs(905) <= not (a xor b);
    layer4_outputs(906) <= not (a and b);
    layer4_outputs(907) <= not (a or b);
    layer4_outputs(908) <= not (a or b);
    layer4_outputs(909) <= a;
    layer4_outputs(910) <= not b;
    layer4_outputs(911) <= b and not a;
    layer4_outputs(912) <= a and b;
    layer4_outputs(913) <= not a;
    layer4_outputs(914) <= b and not a;
    layer4_outputs(915) <= 1'b0;
    layer4_outputs(916) <= not b or a;
    layer4_outputs(917) <= not (a and b);
    layer4_outputs(918) <= a;
    layer4_outputs(919) <= a or b;
    layer4_outputs(920) <= not a or b;
    layer4_outputs(921) <= not a;
    layer4_outputs(922) <= not b;
    layer4_outputs(923) <= not (a xor b);
    layer4_outputs(924) <= a or b;
    layer4_outputs(925) <= a and b;
    layer4_outputs(926) <= a xor b;
    layer4_outputs(927) <= a and b;
    layer4_outputs(928) <= not b;
    layer4_outputs(929) <= b;
    layer4_outputs(930) <= a or b;
    layer4_outputs(931) <= b;
    layer4_outputs(932) <= b and not a;
    layer4_outputs(933) <= 1'b1;
    layer4_outputs(934) <= not (a and b);
    layer4_outputs(935) <= a and not b;
    layer4_outputs(936) <= not a or b;
    layer4_outputs(937) <= b and not a;
    layer4_outputs(938) <= a and b;
    layer4_outputs(939) <= not a;
    layer4_outputs(940) <= not (a or b);
    layer4_outputs(941) <= 1'b1;
    layer4_outputs(942) <= not a;
    layer4_outputs(943) <= not b;
    layer4_outputs(944) <= a and b;
    layer4_outputs(945) <= not (a and b);
    layer4_outputs(946) <= not (a and b);
    layer4_outputs(947) <= b;
    layer4_outputs(948) <= a and b;
    layer4_outputs(949) <= b;
    layer4_outputs(950) <= b and not a;
    layer4_outputs(951) <= a and not b;
    layer4_outputs(952) <= a and not b;
    layer4_outputs(953) <= not (a or b);
    layer4_outputs(954) <= not b;
    layer4_outputs(955) <= not b;
    layer4_outputs(956) <= 1'b1;
    layer4_outputs(957) <= 1'b0;
    layer4_outputs(958) <= not b;
    layer4_outputs(959) <= a or b;
    layer4_outputs(960) <= not a or b;
    layer4_outputs(961) <= not b or a;
    layer4_outputs(962) <= b;
    layer4_outputs(963) <= not a;
    layer4_outputs(964) <= a and b;
    layer4_outputs(965) <= not b or a;
    layer4_outputs(966) <= not a;
    layer4_outputs(967) <= not a or b;
    layer4_outputs(968) <= a and not b;
    layer4_outputs(969) <= a;
    layer4_outputs(970) <= 1'b1;
    layer4_outputs(971) <= not a or b;
    layer4_outputs(972) <= a and not b;
    layer4_outputs(973) <= a or b;
    layer4_outputs(974) <= not (a and b);
    layer4_outputs(975) <= 1'b1;
    layer4_outputs(976) <= 1'b1;
    layer4_outputs(977) <= not b;
    layer4_outputs(978) <= 1'b1;
    layer4_outputs(979) <= not a;
    layer4_outputs(980) <= not b;
    layer4_outputs(981) <= b and not a;
    layer4_outputs(982) <= not (a and b);
    layer4_outputs(983) <= a;
    layer4_outputs(984) <= a and not b;
    layer4_outputs(985) <= not (a and b);
    layer4_outputs(986) <= 1'b0;
    layer4_outputs(987) <= a and not b;
    layer4_outputs(988) <= not b;
    layer4_outputs(989) <= b and not a;
    layer4_outputs(990) <= b;
    layer4_outputs(991) <= not (a and b);
    layer4_outputs(992) <= b;
    layer4_outputs(993) <= 1'b1;
    layer4_outputs(994) <= not a or b;
    layer4_outputs(995) <= not (a xor b);
    layer4_outputs(996) <= not a;
    layer4_outputs(997) <= a and not b;
    layer4_outputs(998) <= 1'b0;
    layer4_outputs(999) <= a and b;
    layer4_outputs(1000) <= b;
    layer4_outputs(1001) <= not a or b;
    layer4_outputs(1002) <= not b;
    layer4_outputs(1003) <= a or b;
    layer4_outputs(1004) <= not b;
    layer4_outputs(1005) <= not b or a;
    layer4_outputs(1006) <= not (a and b);
    layer4_outputs(1007) <= not b or a;
    layer4_outputs(1008) <= not a or b;
    layer4_outputs(1009) <= not a or b;
    layer4_outputs(1010) <= not a or b;
    layer4_outputs(1011) <= not a or b;
    layer4_outputs(1012) <= 1'b0;
    layer4_outputs(1013) <= not a;
    layer4_outputs(1014) <= a and not b;
    layer4_outputs(1015) <= a;
    layer4_outputs(1016) <= 1'b1;
    layer4_outputs(1017) <= not b or a;
    layer4_outputs(1018) <= 1'b1;
    layer4_outputs(1019) <= not a;
    layer4_outputs(1020) <= not b or a;
    layer4_outputs(1021) <= b;
    layer4_outputs(1022) <= not (a or b);
    layer4_outputs(1023) <= not (a or b);
    layer4_outputs(1024) <= not b or a;
    layer4_outputs(1025) <= b and not a;
    layer4_outputs(1026) <= not (a and b);
    layer4_outputs(1027) <= b;
    layer4_outputs(1028) <= not b;
    layer4_outputs(1029) <= 1'b1;
    layer4_outputs(1030) <= 1'b0;
    layer4_outputs(1031) <= 1'b1;
    layer4_outputs(1032) <= a;
    layer4_outputs(1033) <= not b;
    layer4_outputs(1034) <= not (a or b);
    layer4_outputs(1035) <= a;
    layer4_outputs(1036) <= a or b;
    layer4_outputs(1037) <= b;
    layer4_outputs(1038) <= not (a or b);
    layer4_outputs(1039) <= not a;
    layer4_outputs(1040) <= a and not b;
    layer4_outputs(1041) <= a and not b;
    layer4_outputs(1042) <= not b;
    layer4_outputs(1043) <= not (a and b);
    layer4_outputs(1044) <= 1'b1;
    layer4_outputs(1045) <= a and not b;
    layer4_outputs(1046) <= a and b;
    layer4_outputs(1047) <= a xor b;
    layer4_outputs(1048) <= b;
    layer4_outputs(1049) <= 1'b1;
    layer4_outputs(1050) <= a or b;
    layer4_outputs(1051) <= not (a or b);
    layer4_outputs(1052) <= a and not b;
    layer4_outputs(1053) <= a and not b;
    layer4_outputs(1054) <= a;
    layer4_outputs(1055) <= a xor b;
    layer4_outputs(1056) <= not b;
    layer4_outputs(1057) <= not a;
    layer4_outputs(1058) <= a or b;
    layer4_outputs(1059) <= b and not a;
    layer4_outputs(1060) <= b and not a;
    layer4_outputs(1061) <= a and not b;
    layer4_outputs(1062) <= a or b;
    layer4_outputs(1063) <= a or b;
    layer4_outputs(1064) <= b;
    layer4_outputs(1065) <= b;
    layer4_outputs(1066) <= a;
    layer4_outputs(1067) <= b;
    layer4_outputs(1068) <= not a;
    layer4_outputs(1069) <= not (a and b);
    layer4_outputs(1070) <= a and b;
    layer4_outputs(1071) <= a and b;
    layer4_outputs(1072) <= a and not b;
    layer4_outputs(1073) <= 1'b1;
    layer4_outputs(1074) <= not (a or b);
    layer4_outputs(1075) <= b and not a;
    layer4_outputs(1076) <= 1'b1;
    layer4_outputs(1077) <= b;
    layer4_outputs(1078) <= 1'b1;
    layer4_outputs(1079) <= not (a or b);
    layer4_outputs(1080) <= a and b;
    layer4_outputs(1081) <= a and not b;
    layer4_outputs(1082) <= b and not a;
    layer4_outputs(1083) <= a or b;
    layer4_outputs(1084) <= b;
    layer4_outputs(1085) <= a and b;
    layer4_outputs(1086) <= b;
    layer4_outputs(1087) <= b;
    layer4_outputs(1088) <= not a;
    layer4_outputs(1089) <= not b;
    layer4_outputs(1090) <= 1'b1;
    layer4_outputs(1091) <= a xor b;
    layer4_outputs(1092) <= b and not a;
    layer4_outputs(1093) <= 1'b1;
    layer4_outputs(1094) <= not a;
    layer4_outputs(1095) <= not (a and b);
    layer4_outputs(1096) <= not (a or b);
    layer4_outputs(1097) <= a and b;
    layer4_outputs(1098) <= 1'b1;
    layer4_outputs(1099) <= not b;
    layer4_outputs(1100) <= not b;
    layer4_outputs(1101) <= b and not a;
    layer4_outputs(1102) <= not a or b;
    layer4_outputs(1103) <= not (a xor b);
    layer4_outputs(1104) <= not (a xor b);
    layer4_outputs(1105) <= a;
    layer4_outputs(1106) <= a;
    layer4_outputs(1107) <= a;
    layer4_outputs(1108) <= not (a and b);
    layer4_outputs(1109) <= 1'b1;
    layer4_outputs(1110) <= not b or a;
    layer4_outputs(1111) <= not b or a;
    layer4_outputs(1112) <= not (a or b);
    layer4_outputs(1113) <= a and not b;
    layer4_outputs(1114) <= b and not a;
    layer4_outputs(1115) <= a and b;
    layer4_outputs(1116) <= a or b;
    layer4_outputs(1117) <= 1'b1;
    layer4_outputs(1118) <= a;
    layer4_outputs(1119) <= b and not a;
    layer4_outputs(1120) <= b and not a;
    layer4_outputs(1121) <= not (a xor b);
    layer4_outputs(1122) <= not b or a;
    layer4_outputs(1123) <= not (a or b);
    layer4_outputs(1124) <= not (a and b);
    layer4_outputs(1125) <= 1'b0;
    layer4_outputs(1126) <= not (a and b);
    layer4_outputs(1127) <= a xor b;
    layer4_outputs(1128) <= not b;
    layer4_outputs(1129) <= not (a or b);
    layer4_outputs(1130) <= a and b;
    layer4_outputs(1131) <= not a or b;
    layer4_outputs(1132) <= 1'b1;
    layer4_outputs(1133) <= a;
    layer4_outputs(1134) <= a and not b;
    layer4_outputs(1135) <= not b or a;
    layer4_outputs(1136) <= not (a xor b);
    layer4_outputs(1137) <= a and b;
    layer4_outputs(1138) <= a or b;
    layer4_outputs(1139) <= a and b;
    layer4_outputs(1140) <= a and b;
    layer4_outputs(1141) <= a or b;
    layer4_outputs(1142) <= a;
    layer4_outputs(1143) <= a;
    layer4_outputs(1144) <= b;
    layer4_outputs(1145) <= not b or a;
    layer4_outputs(1146) <= a or b;
    layer4_outputs(1147) <= not (a and b);
    layer4_outputs(1148) <= not (a and b);
    layer4_outputs(1149) <= a and not b;
    layer4_outputs(1150) <= not b or a;
    layer4_outputs(1151) <= a and b;
    layer4_outputs(1152) <= b;
    layer4_outputs(1153) <= a and b;
    layer4_outputs(1154) <= a;
    layer4_outputs(1155) <= 1'b0;
    layer4_outputs(1156) <= b;
    layer4_outputs(1157) <= b and not a;
    layer4_outputs(1158) <= not b;
    layer4_outputs(1159) <= a;
    layer4_outputs(1160) <= not a or b;
    layer4_outputs(1161) <= a and b;
    layer4_outputs(1162) <= 1'b0;
    layer4_outputs(1163) <= not b;
    layer4_outputs(1164) <= b and not a;
    layer4_outputs(1165) <= not a;
    layer4_outputs(1166) <= not (a or b);
    layer4_outputs(1167) <= b and not a;
    layer4_outputs(1168) <= not b;
    layer4_outputs(1169) <= not a or b;
    layer4_outputs(1170) <= not b;
    layer4_outputs(1171) <= not (a and b);
    layer4_outputs(1172) <= a xor b;
    layer4_outputs(1173) <= not a;
    layer4_outputs(1174) <= not (a xor b);
    layer4_outputs(1175) <= not a;
    layer4_outputs(1176) <= 1'b1;
    layer4_outputs(1177) <= a xor b;
    layer4_outputs(1178) <= not a or b;
    layer4_outputs(1179) <= a and b;
    layer4_outputs(1180) <= not b;
    layer4_outputs(1181) <= not (a and b);
    layer4_outputs(1182) <= 1'b0;
    layer4_outputs(1183) <= not (a and b);
    layer4_outputs(1184) <= a;
    layer4_outputs(1185) <= b and not a;
    layer4_outputs(1186) <= b;
    layer4_outputs(1187) <= b;
    layer4_outputs(1188) <= not (a and b);
    layer4_outputs(1189) <= a and b;
    layer4_outputs(1190) <= 1'b1;
    layer4_outputs(1191) <= not b or a;
    layer4_outputs(1192) <= a or b;
    layer4_outputs(1193) <= not (a and b);
    layer4_outputs(1194) <= not (a and b);
    layer4_outputs(1195) <= not a;
    layer4_outputs(1196) <= b;
    layer4_outputs(1197) <= 1'b1;
    layer4_outputs(1198) <= a and b;
    layer4_outputs(1199) <= a;
    layer4_outputs(1200) <= 1'b1;
    layer4_outputs(1201) <= a;
    layer4_outputs(1202) <= not (a and b);
    layer4_outputs(1203) <= not b or a;
    layer4_outputs(1204) <= 1'b0;
    layer4_outputs(1205) <= not a or b;
    layer4_outputs(1206) <= not (a xor b);
    layer4_outputs(1207) <= a xor b;
    layer4_outputs(1208) <= not (a xor b);
    layer4_outputs(1209) <= b;
    layer4_outputs(1210) <= not b or a;
    layer4_outputs(1211) <= 1'b1;
    layer4_outputs(1212) <= a and b;
    layer4_outputs(1213) <= b;
    layer4_outputs(1214) <= not b or a;
    layer4_outputs(1215) <= 1'b0;
    layer4_outputs(1216) <= not a;
    layer4_outputs(1217) <= b and not a;
    layer4_outputs(1218) <= b;
    layer4_outputs(1219) <= b and not a;
    layer4_outputs(1220) <= not (a or b);
    layer4_outputs(1221) <= a or b;
    layer4_outputs(1222) <= a and not b;
    layer4_outputs(1223) <= b;
    layer4_outputs(1224) <= not b or a;
    layer4_outputs(1225) <= not a;
    layer4_outputs(1226) <= not a or b;
    layer4_outputs(1227) <= not b;
    layer4_outputs(1228) <= not b or a;
    layer4_outputs(1229) <= b;
    layer4_outputs(1230) <= not (a or b);
    layer4_outputs(1231) <= a and b;
    layer4_outputs(1232) <= a xor b;
    layer4_outputs(1233) <= not (a or b);
    layer4_outputs(1234) <= not b;
    layer4_outputs(1235) <= not (a and b);
    layer4_outputs(1236) <= a;
    layer4_outputs(1237) <= not b or a;
    layer4_outputs(1238) <= not (a or b);
    layer4_outputs(1239) <= not b;
    layer4_outputs(1240) <= not (a xor b);
    layer4_outputs(1241) <= not b or a;
    layer4_outputs(1242) <= not b or a;
    layer4_outputs(1243) <= 1'b1;
    layer4_outputs(1244) <= not (a and b);
    layer4_outputs(1245) <= b and not a;
    layer4_outputs(1246) <= a;
    layer4_outputs(1247) <= a;
    layer4_outputs(1248) <= b;
    layer4_outputs(1249) <= a;
    layer4_outputs(1250) <= b;
    layer4_outputs(1251) <= not b;
    layer4_outputs(1252) <= a and b;
    layer4_outputs(1253) <= 1'b0;
    layer4_outputs(1254) <= not b or a;
    layer4_outputs(1255) <= a or b;
    layer4_outputs(1256) <= not a or b;
    layer4_outputs(1257) <= b and not a;
    layer4_outputs(1258) <= a;
    layer4_outputs(1259) <= b and not a;
    layer4_outputs(1260) <= 1'b1;
    layer4_outputs(1261) <= a;
    layer4_outputs(1262) <= 1'b1;
    layer4_outputs(1263) <= not (a or b);
    layer4_outputs(1264) <= not b;
    layer4_outputs(1265) <= b;
    layer4_outputs(1266) <= 1'b0;
    layer4_outputs(1267) <= not b;
    layer4_outputs(1268) <= a and b;
    layer4_outputs(1269) <= a or b;
    layer4_outputs(1270) <= a;
    layer4_outputs(1271) <= a;
    layer4_outputs(1272) <= not (a and b);
    layer4_outputs(1273) <= not (a and b);
    layer4_outputs(1274) <= not (a and b);
    layer4_outputs(1275) <= a;
    layer4_outputs(1276) <= not b;
    layer4_outputs(1277) <= not (a and b);
    layer4_outputs(1278) <= not (a and b);
    layer4_outputs(1279) <= a or b;
    layer4_outputs(1280) <= a and b;
    layer4_outputs(1281) <= not b or a;
    layer4_outputs(1282) <= not (a and b);
    layer4_outputs(1283) <= 1'b1;
    layer4_outputs(1284) <= 1'b0;
    layer4_outputs(1285) <= not b or a;
    layer4_outputs(1286) <= not a or b;
    layer4_outputs(1287) <= a and not b;
    layer4_outputs(1288) <= a and b;
    layer4_outputs(1289) <= a;
    layer4_outputs(1290) <= a or b;
    layer4_outputs(1291) <= a xor b;
    layer4_outputs(1292) <= 1'b0;
    layer4_outputs(1293) <= not a;
    layer4_outputs(1294) <= not (a xor b);
    layer4_outputs(1295) <= a and b;
    layer4_outputs(1296) <= a or b;
    layer4_outputs(1297) <= not (a xor b);
    layer4_outputs(1298) <= not (a and b);
    layer4_outputs(1299) <= not a or b;
    layer4_outputs(1300) <= not (a and b);
    layer4_outputs(1301) <= b;
    layer4_outputs(1302) <= not (a or b);
    layer4_outputs(1303) <= not b or a;
    layer4_outputs(1304) <= not b;
    layer4_outputs(1305) <= a or b;
    layer4_outputs(1306) <= not (a or b);
    layer4_outputs(1307) <= not a or b;
    layer4_outputs(1308) <= not b or a;
    layer4_outputs(1309) <= b;
    layer4_outputs(1310) <= a;
    layer4_outputs(1311) <= not b or a;
    layer4_outputs(1312) <= b;
    layer4_outputs(1313) <= b and not a;
    layer4_outputs(1314) <= not (a and b);
    layer4_outputs(1315) <= a;
    layer4_outputs(1316) <= a and b;
    layer4_outputs(1317) <= a or b;
    layer4_outputs(1318) <= not b;
    layer4_outputs(1319) <= b;
    layer4_outputs(1320) <= not (a or b);
    layer4_outputs(1321) <= a;
    layer4_outputs(1322) <= 1'b1;
    layer4_outputs(1323) <= not b or a;
    layer4_outputs(1324) <= a;
    layer4_outputs(1325) <= b;
    layer4_outputs(1326) <= not (a or b);
    layer4_outputs(1327) <= not a or b;
    layer4_outputs(1328) <= a and b;
    layer4_outputs(1329) <= a and not b;
    layer4_outputs(1330) <= not a or b;
    layer4_outputs(1331) <= a or b;
    layer4_outputs(1332) <= b;
    layer4_outputs(1333) <= not (a or b);
    layer4_outputs(1334) <= a;
    layer4_outputs(1335) <= not b;
    layer4_outputs(1336) <= b;
    layer4_outputs(1337) <= 1'b1;
    layer4_outputs(1338) <= a xor b;
    layer4_outputs(1339) <= a or b;
    layer4_outputs(1340) <= not (a xor b);
    layer4_outputs(1341) <= not a or b;
    layer4_outputs(1342) <= 1'b0;
    layer4_outputs(1343) <= not a;
    layer4_outputs(1344) <= a or b;
    layer4_outputs(1345) <= a;
    layer4_outputs(1346) <= not (a and b);
    layer4_outputs(1347) <= not (a xor b);
    layer4_outputs(1348) <= not b;
    layer4_outputs(1349) <= not b;
    layer4_outputs(1350) <= b;
    layer4_outputs(1351) <= a xor b;
    layer4_outputs(1352) <= not (a xor b);
    layer4_outputs(1353) <= a and not b;
    layer4_outputs(1354) <= not a;
    layer4_outputs(1355) <= not b;
    layer4_outputs(1356) <= not (a or b);
    layer4_outputs(1357) <= a;
    layer4_outputs(1358) <= not b;
    layer4_outputs(1359) <= a or b;
    layer4_outputs(1360) <= not (a or b);
    layer4_outputs(1361) <= not a;
    layer4_outputs(1362) <= 1'b0;
    layer4_outputs(1363) <= 1'b1;
    layer4_outputs(1364) <= not a or b;
    layer4_outputs(1365) <= a or b;
    layer4_outputs(1366) <= a or b;
    layer4_outputs(1367) <= b and not a;
    layer4_outputs(1368) <= b;
    layer4_outputs(1369) <= a and b;
    layer4_outputs(1370) <= 1'b0;
    layer4_outputs(1371) <= not (a and b);
    layer4_outputs(1372) <= a and not b;
    layer4_outputs(1373) <= not b;
    layer4_outputs(1374) <= 1'b0;
    layer4_outputs(1375) <= b and not a;
    layer4_outputs(1376) <= b;
    layer4_outputs(1377) <= 1'b1;
    layer4_outputs(1378) <= not (a and b);
    layer4_outputs(1379) <= not b;
    layer4_outputs(1380) <= not b;
    layer4_outputs(1381) <= not (a and b);
    layer4_outputs(1382) <= 1'b1;
    layer4_outputs(1383) <= not b or a;
    layer4_outputs(1384) <= a and not b;
    layer4_outputs(1385) <= a or b;
    layer4_outputs(1386) <= a and b;
    layer4_outputs(1387) <= a and b;
    layer4_outputs(1388) <= 1'b1;
    layer4_outputs(1389) <= a and not b;
    layer4_outputs(1390) <= 1'b1;
    layer4_outputs(1391) <= a and b;
    layer4_outputs(1392) <= not (a and b);
    layer4_outputs(1393) <= a or b;
    layer4_outputs(1394) <= 1'b1;
    layer4_outputs(1395) <= not (a xor b);
    layer4_outputs(1396) <= 1'b1;
    layer4_outputs(1397) <= not b;
    layer4_outputs(1398) <= 1'b0;
    layer4_outputs(1399) <= not b or a;
    layer4_outputs(1400) <= a and not b;
    layer4_outputs(1401) <= b;
    layer4_outputs(1402) <= a or b;
    layer4_outputs(1403) <= not b;
    layer4_outputs(1404) <= b and not a;
    layer4_outputs(1405) <= not (a or b);
    layer4_outputs(1406) <= not a or b;
    layer4_outputs(1407) <= a;
    layer4_outputs(1408) <= a;
    layer4_outputs(1409) <= a and b;
    layer4_outputs(1410) <= not a;
    layer4_outputs(1411) <= 1'b0;
    layer4_outputs(1412) <= b;
    layer4_outputs(1413) <= not a;
    layer4_outputs(1414) <= a and not b;
    layer4_outputs(1415) <= b;
    layer4_outputs(1416) <= b;
    layer4_outputs(1417) <= not a;
    layer4_outputs(1418) <= 1'b0;
    layer4_outputs(1419) <= not a;
    layer4_outputs(1420) <= not b or a;
    layer4_outputs(1421) <= not (a and b);
    layer4_outputs(1422) <= not a;
    layer4_outputs(1423) <= not (a xor b);
    layer4_outputs(1424) <= not b;
    layer4_outputs(1425) <= b;
    layer4_outputs(1426) <= b;
    layer4_outputs(1427) <= not a;
    layer4_outputs(1428) <= b and not a;
    layer4_outputs(1429) <= a or b;
    layer4_outputs(1430) <= not a;
    layer4_outputs(1431) <= a;
    layer4_outputs(1432) <= b;
    layer4_outputs(1433) <= not b;
    layer4_outputs(1434) <= a and b;
    layer4_outputs(1435) <= a;
    layer4_outputs(1436) <= a and b;
    layer4_outputs(1437) <= not b or a;
    layer4_outputs(1438) <= b;
    layer4_outputs(1439) <= a;
    layer4_outputs(1440) <= a and not b;
    layer4_outputs(1441) <= 1'b0;
    layer4_outputs(1442) <= a or b;
    layer4_outputs(1443) <= 1'b1;
    layer4_outputs(1444) <= not b;
    layer4_outputs(1445) <= 1'b1;
    layer4_outputs(1446) <= a or b;
    layer4_outputs(1447) <= not (a and b);
    layer4_outputs(1448) <= a and not b;
    layer4_outputs(1449) <= a xor b;
    layer4_outputs(1450) <= not a or b;
    layer4_outputs(1451) <= a and b;
    layer4_outputs(1452) <= not a or b;
    layer4_outputs(1453) <= not b;
    layer4_outputs(1454) <= not (a or b);
    layer4_outputs(1455) <= not (a or b);
    layer4_outputs(1456) <= not (a and b);
    layer4_outputs(1457) <= a and not b;
    layer4_outputs(1458) <= not b or a;
    layer4_outputs(1459) <= not a;
    layer4_outputs(1460) <= not (a or b);
    layer4_outputs(1461) <= a xor b;
    layer4_outputs(1462) <= not a;
    layer4_outputs(1463) <= a and not b;
    layer4_outputs(1464) <= not (a xor b);
    layer4_outputs(1465) <= a;
    layer4_outputs(1466) <= not b or a;
    layer4_outputs(1467) <= not b;
    layer4_outputs(1468) <= not a;
    layer4_outputs(1469) <= b;
    layer4_outputs(1470) <= not a;
    layer4_outputs(1471) <= not a;
    layer4_outputs(1472) <= not (a and b);
    layer4_outputs(1473) <= a and b;
    layer4_outputs(1474) <= a and not b;
    layer4_outputs(1475) <= not b or a;
    layer4_outputs(1476) <= b and not a;
    layer4_outputs(1477) <= not a;
    layer4_outputs(1478) <= not a or b;
    layer4_outputs(1479) <= b and not a;
    layer4_outputs(1480) <= 1'b1;
    layer4_outputs(1481) <= not a or b;
    layer4_outputs(1482) <= not b;
    layer4_outputs(1483) <= not b or a;
    layer4_outputs(1484) <= a or b;
    layer4_outputs(1485) <= not a;
    layer4_outputs(1486) <= a xor b;
    layer4_outputs(1487) <= a and b;
    layer4_outputs(1488) <= not b or a;
    layer4_outputs(1489) <= b;
    layer4_outputs(1490) <= a;
    layer4_outputs(1491) <= not (a xor b);
    layer4_outputs(1492) <= not a or b;
    layer4_outputs(1493) <= not b or a;
    layer4_outputs(1494) <= 1'b1;
    layer4_outputs(1495) <= 1'b0;
    layer4_outputs(1496) <= not a or b;
    layer4_outputs(1497) <= a and b;
    layer4_outputs(1498) <= not b;
    layer4_outputs(1499) <= a xor b;
    layer4_outputs(1500) <= not b or a;
    layer4_outputs(1501) <= not b or a;
    layer4_outputs(1502) <= not (a or b);
    layer4_outputs(1503) <= 1'b1;
    layer4_outputs(1504) <= not a or b;
    layer4_outputs(1505) <= b and not a;
    layer4_outputs(1506) <= a and b;
    layer4_outputs(1507) <= a and not b;
    layer4_outputs(1508) <= not (a or b);
    layer4_outputs(1509) <= b and not a;
    layer4_outputs(1510) <= not b;
    layer4_outputs(1511) <= a;
    layer4_outputs(1512) <= not a or b;
    layer4_outputs(1513) <= a or b;
    layer4_outputs(1514) <= not b or a;
    layer4_outputs(1515) <= 1'b0;
    layer4_outputs(1516) <= not (a xor b);
    layer4_outputs(1517) <= a or b;
    layer4_outputs(1518) <= not (a and b);
    layer4_outputs(1519) <= b;
    layer4_outputs(1520) <= 1'b1;
    layer4_outputs(1521) <= b and not a;
    layer4_outputs(1522) <= not b;
    layer4_outputs(1523) <= not b;
    layer4_outputs(1524) <= not a;
    layer4_outputs(1525) <= 1'b1;
    layer4_outputs(1526) <= a or b;
    layer4_outputs(1527) <= not a;
    layer4_outputs(1528) <= not (a xor b);
    layer4_outputs(1529) <= not (a and b);
    layer4_outputs(1530) <= a or b;
    layer4_outputs(1531) <= not a;
    layer4_outputs(1532) <= not (a and b);
    layer4_outputs(1533) <= 1'b1;
    layer4_outputs(1534) <= a xor b;
    layer4_outputs(1535) <= a xor b;
    layer4_outputs(1536) <= a or b;
    layer4_outputs(1537) <= not b or a;
    layer4_outputs(1538) <= a and b;
    layer4_outputs(1539) <= a;
    layer4_outputs(1540) <= not (a xor b);
    layer4_outputs(1541) <= not b;
    layer4_outputs(1542) <= a or b;
    layer4_outputs(1543) <= not a or b;
    layer4_outputs(1544) <= a;
    layer4_outputs(1545) <= not (a xor b);
    layer4_outputs(1546) <= b;
    layer4_outputs(1547) <= not (a and b);
    layer4_outputs(1548) <= not a or b;
    layer4_outputs(1549) <= a and not b;
    layer4_outputs(1550) <= not b or a;
    layer4_outputs(1551) <= a and not b;
    layer4_outputs(1552) <= not a;
    layer4_outputs(1553) <= b and not a;
    layer4_outputs(1554) <= not b;
    layer4_outputs(1555) <= a and not b;
    layer4_outputs(1556) <= a;
    layer4_outputs(1557) <= not (a or b);
    layer4_outputs(1558) <= b;
    layer4_outputs(1559) <= not a;
    layer4_outputs(1560) <= not (a and b);
    layer4_outputs(1561) <= not a or b;
    layer4_outputs(1562) <= not a or b;
    layer4_outputs(1563) <= a and not b;
    layer4_outputs(1564) <= b and not a;
    layer4_outputs(1565) <= not b or a;
    layer4_outputs(1566) <= 1'b1;
    layer4_outputs(1567) <= a and not b;
    layer4_outputs(1568) <= a;
    layer4_outputs(1569) <= a or b;
    layer4_outputs(1570) <= a;
    layer4_outputs(1571) <= b and not a;
    layer4_outputs(1572) <= a and b;
    layer4_outputs(1573) <= not (a or b);
    layer4_outputs(1574) <= not b;
    layer4_outputs(1575) <= not (a or b);
    layer4_outputs(1576) <= a and not b;
    layer4_outputs(1577) <= not (a and b);
    layer4_outputs(1578) <= b and not a;
    layer4_outputs(1579) <= a or b;
    layer4_outputs(1580) <= b;
    layer4_outputs(1581) <= not a or b;
    layer4_outputs(1582) <= 1'b0;
    layer4_outputs(1583) <= b;
    layer4_outputs(1584) <= not a or b;
    layer4_outputs(1585) <= not (a and b);
    layer4_outputs(1586) <= b and not a;
    layer4_outputs(1587) <= not b or a;
    layer4_outputs(1588) <= 1'b0;
    layer4_outputs(1589) <= 1'b1;
    layer4_outputs(1590) <= not b;
    layer4_outputs(1591) <= 1'b0;
    layer4_outputs(1592) <= a and b;
    layer4_outputs(1593) <= 1'b0;
    layer4_outputs(1594) <= not (a and b);
    layer4_outputs(1595) <= not a or b;
    layer4_outputs(1596) <= not b or a;
    layer4_outputs(1597) <= a or b;
    layer4_outputs(1598) <= a and not b;
    layer4_outputs(1599) <= not a or b;
    layer4_outputs(1600) <= b;
    layer4_outputs(1601) <= a or b;
    layer4_outputs(1602) <= not a or b;
    layer4_outputs(1603) <= not (a and b);
    layer4_outputs(1604) <= a and not b;
    layer4_outputs(1605) <= a or b;
    layer4_outputs(1606) <= a;
    layer4_outputs(1607) <= 1'b0;
    layer4_outputs(1608) <= 1'b0;
    layer4_outputs(1609) <= not b or a;
    layer4_outputs(1610) <= 1'b1;
    layer4_outputs(1611) <= a and not b;
    layer4_outputs(1612) <= a and b;
    layer4_outputs(1613) <= b and not a;
    layer4_outputs(1614) <= not b or a;
    layer4_outputs(1615) <= 1'b1;
    layer4_outputs(1616) <= 1'b0;
    layer4_outputs(1617) <= not a or b;
    layer4_outputs(1618) <= not b or a;
    layer4_outputs(1619) <= not a or b;
    layer4_outputs(1620) <= b;
    layer4_outputs(1621) <= a;
    layer4_outputs(1622) <= not b or a;
    layer4_outputs(1623) <= a and b;
    layer4_outputs(1624) <= a and not b;
    layer4_outputs(1625) <= not b;
    layer4_outputs(1626) <= not b or a;
    layer4_outputs(1627) <= a or b;
    layer4_outputs(1628) <= a;
    layer4_outputs(1629) <= a or b;
    layer4_outputs(1630) <= a or b;
    layer4_outputs(1631) <= 1'b1;
    layer4_outputs(1632) <= not a;
    layer4_outputs(1633) <= a and not b;
    layer4_outputs(1634) <= b and not a;
    layer4_outputs(1635) <= 1'b1;
    layer4_outputs(1636) <= not (a and b);
    layer4_outputs(1637) <= not a or b;
    layer4_outputs(1638) <= b;
    layer4_outputs(1639) <= a or b;
    layer4_outputs(1640) <= a or b;
    layer4_outputs(1641) <= not (a and b);
    layer4_outputs(1642) <= not (a and b);
    layer4_outputs(1643) <= a;
    layer4_outputs(1644) <= not a or b;
    layer4_outputs(1645) <= not (a or b);
    layer4_outputs(1646) <= not b or a;
    layer4_outputs(1647) <= not a or b;
    layer4_outputs(1648) <= 1'b1;
    layer4_outputs(1649) <= 1'b0;
    layer4_outputs(1650) <= 1'b0;
    layer4_outputs(1651) <= a and not b;
    layer4_outputs(1652) <= b;
    layer4_outputs(1653) <= 1'b1;
    layer4_outputs(1654) <= a and not b;
    layer4_outputs(1655) <= a or b;
    layer4_outputs(1656) <= not a or b;
    layer4_outputs(1657) <= not (a or b);
    layer4_outputs(1658) <= not a;
    layer4_outputs(1659) <= a and b;
    layer4_outputs(1660) <= not b or a;
    layer4_outputs(1661) <= not (a or b);
    layer4_outputs(1662) <= not (a and b);
    layer4_outputs(1663) <= not a or b;
    layer4_outputs(1664) <= not (a and b);
    layer4_outputs(1665) <= not a;
    layer4_outputs(1666) <= a and b;
    layer4_outputs(1667) <= 1'b0;
    layer4_outputs(1668) <= not b;
    layer4_outputs(1669) <= not a;
    layer4_outputs(1670) <= not (a xor b);
    layer4_outputs(1671) <= 1'b1;
    layer4_outputs(1672) <= b and not a;
    layer4_outputs(1673) <= b;
    layer4_outputs(1674) <= not (a and b);
    layer4_outputs(1675) <= not a;
    layer4_outputs(1676) <= b and not a;
    layer4_outputs(1677) <= not b;
    layer4_outputs(1678) <= b;
    layer4_outputs(1679) <= a and not b;
    layer4_outputs(1680) <= b;
    layer4_outputs(1681) <= 1'b0;
    layer4_outputs(1682) <= not a;
    layer4_outputs(1683) <= a;
    layer4_outputs(1684) <= not b or a;
    layer4_outputs(1685) <= a and not b;
    layer4_outputs(1686) <= not b or a;
    layer4_outputs(1687) <= not b;
    layer4_outputs(1688) <= not (a and b);
    layer4_outputs(1689) <= not b or a;
    layer4_outputs(1690) <= not (a or b);
    layer4_outputs(1691) <= a and b;
    layer4_outputs(1692) <= b;
    layer4_outputs(1693) <= b and not a;
    layer4_outputs(1694) <= a and b;
    layer4_outputs(1695) <= not (a or b);
    layer4_outputs(1696) <= not b or a;
    layer4_outputs(1697) <= not b;
    layer4_outputs(1698) <= b;
    layer4_outputs(1699) <= not (a xor b);
    layer4_outputs(1700) <= not a or b;
    layer4_outputs(1701) <= not (a and b);
    layer4_outputs(1702) <= b and not a;
    layer4_outputs(1703) <= b and not a;
    layer4_outputs(1704) <= not (a xor b);
    layer4_outputs(1705) <= not a;
    layer4_outputs(1706) <= 1'b0;
    layer4_outputs(1707) <= not a or b;
    layer4_outputs(1708) <= a;
    layer4_outputs(1709) <= not (a and b);
    layer4_outputs(1710) <= 1'b1;
    layer4_outputs(1711) <= a and b;
    layer4_outputs(1712) <= a and b;
    layer4_outputs(1713) <= 1'b1;
    layer4_outputs(1714) <= not a;
    layer4_outputs(1715) <= a and not b;
    layer4_outputs(1716) <= a;
    layer4_outputs(1717) <= not b or a;
    layer4_outputs(1718) <= b and not a;
    layer4_outputs(1719) <= b;
    layer4_outputs(1720) <= a;
    layer4_outputs(1721) <= b;
    layer4_outputs(1722) <= not (a xor b);
    layer4_outputs(1723) <= 1'b1;
    layer4_outputs(1724) <= a and b;
    layer4_outputs(1725) <= a;
    layer4_outputs(1726) <= not (a or b);
    layer4_outputs(1727) <= b;
    layer4_outputs(1728) <= 1'b0;
    layer4_outputs(1729) <= not (a and b);
    layer4_outputs(1730) <= not (a or b);
    layer4_outputs(1731) <= a xor b;
    layer4_outputs(1732) <= b and not a;
    layer4_outputs(1733) <= 1'b0;
    layer4_outputs(1734) <= not b;
    layer4_outputs(1735) <= 1'b0;
    layer4_outputs(1736) <= 1'b1;
    layer4_outputs(1737) <= not b or a;
    layer4_outputs(1738) <= a or b;
    layer4_outputs(1739) <= a xor b;
    layer4_outputs(1740) <= not (a or b);
    layer4_outputs(1741) <= a and b;
    layer4_outputs(1742) <= a and b;
    layer4_outputs(1743) <= a and not b;
    layer4_outputs(1744) <= b;
    layer4_outputs(1745) <= not a or b;
    layer4_outputs(1746) <= not a or b;
    layer4_outputs(1747) <= b;
    layer4_outputs(1748) <= not (a and b);
    layer4_outputs(1749) <= not b;
    layer4_outputs(1750) <= not (a and b);
    layer4_outputs(1751) <= b;
    layer4_outputs(1752) <= b;
    layer4_outputs(1753) <= not a or b;
    layer4_outputs(1754) <= 1'b1;
    layer4_outputs(1755) <= not b or a;
    layer4_outputs(1756) <= b;
    layer4_outputs(1757) <= a or b;
    layer4_outputs(1758) <= a and not b;
    layer4_outputs(1759) <= b;
    layer4_outputs(1760) <= a;
    layer4_outputs(1761) <= b;
    layer4_outputs(1762) <= a and not b;
    layer4_outputs(1763) <= 1'b0;
    layer4_outputs(1764) <= not (a or b);
    layer4_outputs(1765) <= 1'b1;
    layer4_outputs(1766) <= not (a or b);
    layer4_outputs(1767) <= not (a and b);
    layer4_outputs(1768) <= a and b;
    layer4_outputs(1769) <= b;
    layer4_outputs(1770) <= a;
    layer4_outputs(1771) <= 1'b0;
    layer4_outputs(1772) <= b;
    layer4_outputs(1773) <= not (a or b);
    layer4_outputs(1774) <= a and b;
    layer4_outputs(1775) <= not b;
    layer4_outputs(1776) <= not (a or b);
    layer4_outputs(1777) <= a and b;
    layer4_outputs(1778) <= not a or b;
    layer4_outputs(1779) <= b and not a;
    layer4_outputs(1780) <= not (a and b);
    layer4_outputs(1781) <= not b or a;
    layer4_outputs(1782) <= a or b;
    layer4_outputs(1783) <= a;
    layer4_outputs(1784) <= 1'b1;
    layer4_outputs(1785) <= a xor b;
    layer4_outputs(1786) <= b and not a;
    layer4_outputs(1787) <= b;
    layer4_outputs(1788) <= not b or a;
    layer4_outputs(1789) <= not (a or b);
    layer4_outputs(1790) <= not b;
    layer4_outputs(1791) <= a and not b;
    layer4_outputs(1792) <= b and not a;
    layer4_outputs(1793) <= 1'b1;
    layer4_outputs(1794) <= a or b;
    layer4_outputs(1795) <= 1'b0;
    layer4_outputs(1796) <= a;
    layer4_outputs(1797) <= a;
    layer4_outputs(1798) <= not a or b;
    layer4_outputs(1799) <= not a;
    layer4_outputs(1800) <= b and not a;
    layer4_outputs(1801) <= b;
    layer4_outputs(1802) <= a;
    layer4_outputs(1803) <= b and not a;
    layer4_outputs(1804) <= not b;
    layer4_outputs(1805) <= 1'b1;
    layer4_outputs(1806) <= a and b;
    layer4_outputs(1807) <= b;
    layer4_outputs(1808) <= 1'b1;
    layer4_outputs(1809) <= not (a or b);
    layer4_outputs(1810) <= a;
    layer4_outputs(1811) <= 1'b0;
    layer4_outputs(1812) <= not a or b;
    layer4_outputs(1813) <= a and b;
    layer4_outputs(1814) <= b and not a;
    layer4_outputs(1815) <= not a or b;
    layer4_outputs(1816) <= a;
    layer4_outputs(1817) <= b;
    layer4_outputs(1818) <= not a;
    layer4_outputs(1819) <= not b;
    layer4_outputs(1820) <= b;
    layer4_outputs(1821) <= b;
    layer4_outputs(1822) <= a or b;
    layer4_outputs(1823) <= b and not a;
    layer4_outputs(1824) <= a and not b;
    layer4_outputs(1825) <= not a;
    layer4_outputs(1826) <= a xor b;
    layer4_outputs(1827) <= a and not b;
    layer4_outputs(1828) <= not (a and b);
    layer4_outputs(1829) <= a and not b;
    layer4_outputs(1830) <= not a;
    layer4_outputs(1831) <= a and b;
    layer4_outputs(1832) <= a;
    layer4_outputs(1833) <= a;
    layer4_outputs(1834) <= not (a or b);
    layer4_outputs(1835) <= a or b;
    layer4_outputs(1836) <= not (a and b);
    layer4_outputs(1837) <= not a or b;
    layer4_outputs(1838) <= not (a and b);
    layer4_outputs(1839) <= b;
    layer4_outputs(1840) <= not b or a;
    layer4_outputs(1841) <= b;
    layer4_outputs(1842) <= a or b;
    layer4_outputs(1843) <= a xor b;
    layer4_outputs(1844) <= not (a xor b);
    layer4_outputs(1845) <= not (a xor b);
    layer4_outputs(1846) <= not a;
    layer4_outputs(1847) <= not (a xor b);
    layer4_outputs(1848) <= not (a or b);
    layer4_outputs(1849) <= not (a and b);
    layer4_outputs(1850) <= not a or b;
    layer4_outputs(1851) <= a and not b;
    layer4_outputs(1852) <= a and not b;
    layer4_outputs(1853) <= b;
    layer4_outputs(1854) <= 1'b0;
    layer4_outputs(1855) <= a and b;
    layer4_outputs(1856) <= 1'b0;
    layer4_outputs(1857) <= not b or a;
    layer4_outputs(1858) <= a xor b;
    layer4_outputs(1859) <= b;
    layer4_outputs(1860) <= a;
    layer4_outputs(1861) <= 1'b0;
    layer4_outputs(1862) <= a and b;
    layer4_outputs(1863) <= not b;
    layer4_outputs(1864) <= not b or a;
    layer4_outputs(1865) <= a;
    layer4_outputs(1866) <= a and b;
    layer4_outputs(1867) <= not b;
    layer4_outputs(1868) <= not b;
    layer4_outputs(1869) <= not (a and b);
    layer4_outputs(1870) <= b and not a;
    layer4_outputs(1871) <= not b;
    layer4_outputs(1872) <= a and not b;
    layer4_outputs(1873) <= not (a or b);
    layer4_outputs(1874) <= not b or a;
    layer4_outputs(1875) <= b;
    layer4_outputs(1876) <= not (a and b);
    layer4_outputs(1877) <= not (a or b);
    layer4_outputs(1878) <= not a or b;
    layer4_outputs(1879) <= a and not b;
    layer4_outputs(1880) <= not (a and b);
    layer4_outputs(1881) <= not (a or b);
    layer4_outputs(1882) <= a and b;
    layer4_outputs(1883) <= a or b;
    layer4_outputs(1884) <= a and not b;
    layer4_outputs(1885) <= b and not a;
    layer4_outputs(1886) <= a or b;
    layer4_outputs(1887) <= a or b;
    layer4_outputs(1888) <= a xor b;
    layer4_outputs(1889) <= b and not a;
    layer4_outputs(1890) <= not (a or b);
    layer4_outputs(1891) <= a or b;
    layer4_outputs(1892) <= a and b;
    layer4_outputs(1893) <= not (a and b);
    layer4_outputs(1894) <= b and not a;
    layer4_outputs(1895) <= not (a xor b);
    layer4_outputs(1896) <= not a or b;
    layer4_outputs(1897) <= b;
    layer4_outputs(1898) <= b and not a;
    layer4_outputs(1899) <= a and not b;
    layer4_outputs(1900) <= a or b;
    layer4_outputs(1901) <= not b;
    layer4_outputs(1902) <= b;
    layer4_outputs(1903) <= a or b;
    layer4_outputs(1904) <= 1'b1;
    layer4_outputs(1905) <= b and not a;
    layer4_outputs(1906) <= b and not a;
    layer4_outputs(1907) <= a;
    layer4_outputs(1908) <= 1'b1;
    layer4_outputs(1909) <= b and not a;
    layer4_outputs(1910) <= a and b;
    layer4_outputs(1911) <= b;
    layer4_outputs(1912) <= a and b;
    layer4_outputs(1913) <= b and not a;
    layer4_outputs(1914) <= a or b;
    layer4_outputs(1915) <= not a or b;
    layer4_outputs(1916) <= not (a xor b);
    layer4_outputs(1917) <= a and not b;
    layer4_outputs(1918) <= not a or b;
    layer4_outputs(1919) <= not a or b;
    layer4_outputs(1920) <= not b or a;
    layer4_outputs(1921) <= 1'b1;
    layer4_outputs(1922) <= not (a or b);
    layer4_outputs(1923) <= not b;
    layer4_outputs(1924) <= b;
    layer4_outputs(1925) <= b;
    layer4_outputs(1926) <= not (a and b);
    layer4_outputs(1927) <= a or b;
    layer4_outputs(1928) <= not a or b;
    layer4_outputs(1929) <= not (a or b);
    layer4_outputs(1930) <= a or b;
    layer4_outputs(1931) <= a;
    layer4_outputs(1932) <= not a or b;
    layer4_outputs(1933) <= not a or b;
    layer4_outputs(1934) <= not a;
    layer4_outputs(1935) <= not a;
    layer4_outputs(1936) <= a;
    layer4_outputs(1937) <= a;
    layer4_outputs(1938) <= a and b;
    layer4_outputs(1939) <= not b;
    layer4_outputs(1940) <= not b or a;
    layer4_outputs(1941) <= not (a and b);
    layer4_outputs(1942) <= a and b;
    layer4_outputs(1943) <= not (a and b);
    layer4_outputs(1944) <= b;
    layer4_outputs(1945) <= b;
    layer4_outputs(1946) <= a xor b;
    layer4_outputs(1947) <= b and not a;
    layer4_outputs(1948) <= a or b;
    layer4_outputs(1949) <= a and b;
    layer4_outputs(1950) <= b and not a;
    layer4_outputs(1951) <= not a;
    layer4_outputs(1952) <= 1'b1;
    layer4_outputs(1953) <= b and not a;
    layer4_outputs(1954) <= a and b;
    layer4_outputs(1955) <= a xor b;
    layer4_outputs(1956) <= not a or b;
    layer4_outputs(1957) <= a and not b;
    layer4_outputs(1958) <= a and not b;
    layer4_outputs(1959) <= not (a xor b);
    layer4_outputs(1960) <= a;
    layer4_outputs(1961) <= 1'b0;
    layer4_outputs(1962) <= 1'b1;
    layer4_outputs(1963) <= not b or a;
    layer4_outputs(1964) <= a and not b;
    layer4_outputs(1965) <= not a;
    layer4_outputs(1966) <= not (a or b);
    layer4_outputs(1967) <= not (a xor b);
    layer4_outputs(1968) <= b and not a;
    layer4_outputs(1969) <= not b;
    layer4_outputs(1970) <= not (a xor b);
    layer4_outputs(1971) <= a xor b;
    layer4_outputs(1972) <= not (a and b);
    layer4_outputs(1973) <= b and not a;
    layer4_outputs(1974) <= not a or b;
    layer4_outputs(1975) <= a and b;
    layer4_outputs(1976) <= not (a xor b);
    layer4_outputs(1977) <= a xor b;
    layer4_outputs(1978) <= not b or a;
    layer4_outputs(1979) <= not (a and b);
    layer4_outputs(1980) <= 1'b1;
    layer4_outputs(1981) <= not b;
    layer4_outputs(1982) <= 1'b1;
    layer4_outputs(1983) <= not (a or b);
    layer4_outputs(1984) <= b;
    layer4_outputs(1985) <= a;
    layer4_outputs(1986) <= not a;
    layer4_outputs(1987) <= not a;
    layer4_outputs(1988) <= a and b;
    layer4_outputs(1989) <= a xor b;
    layer4_outputs(1990) <= a;
    layer4_outputs(1991) <= 1'b0;
    layer4_outputs(1992) <= a;
    layer4_outputs(1993) <= not (a and b);
    layer4_outputs(1994) <= a xor b;
    layer4_outputs(1995) <= b;
    layer4_outputs(1996) <= not a;
    layer4_outputs(1997) <= b;
    layer4_outputs(1998) <= not (a xor b);
    layer4_outputs(1999) <= a;
    layer4_outputs(2000) <= not b;
    layer4_outputs(2001) <= not a or b;
    layer4_outputs(2002) <= 1'b1;
    layer4_outputs(2003) <= not (a xor b);
    layer4_outputs(2004) <= 1'b0;
    layer4_outputs(2005) <= not (a xor b);
    layer4_outputs(2006) <= not b;
    layer4_outputs(2007) <= not (a and b);
    layer4_outputs(2008) <= not (a or b);
    layer4_outputs(2009) <= a;
    layer4_outputs(2010) <= not a or b;
    layer4_outputs(2011) <= a and b;
    layer4_outputs(2012) <= a;
    layer4_outputs(2013) <= b;
    layer4_outputs(2014) <= b;
    layer4_outputs(2015) <= a;
    layer4_outputs(2016) <= b;
    layer4_outputs(2017) <= 1'b1;
    layer4_outputs(2018) <= a and not b;
    layer4_outputs(2019) <= not a;
    layer4_outputs(2020) <= 1'b1;
    layer4_outputs(2021) <= b;
    layer4_outputs(2022) <= a and b;
    layer4_outputs(2023) <= 1'b1;
    layer4_outputs(2024) <= b and not a;
    layer4_outputs(2025) <= a;
    layer4_outputs(2026) <= not (a or b);
    layer4_outputs(2027) <= a;
    layer4_outputs(2028) <= a and b;
    layer4_outputs(2029) <= a or b;
    layer4_outputs(2030) <= not b or a;
    layer4_outputs(2031) <= a xor b;
    layer4_outputs(2032) <= b;
    layer4_outputs(2033) <= not (a or b);
    layer4_outputs(2034) <= a or b;
    layer4_outputs(2035) <= a;
    layer4_outputs(2036) <= not b or a;
    layer4_outputs(2037) <= b;
    layer4_outputs(2038) <= a or b;
    layer4_outputs(2039) <= not (a and b);
    layer4_outputs(2040) <= not a or b;
    layer4_outputs(2041) <= 1'b1;
    layer4_outputs(2042) <= not a or b;
    layer4_outputs(2043) <= not (a and b);
    layer4_outputs(2044) <= not a or b;
    layer4_outputs(2045) <= a;
    layer4_outputs(2046) <= not b or a;
    layer4_outputs(2047) <= not b or a;
    layer4_outputs(2048) <= a and not b;
    layer4_outputs(2049) <= a;
    layer4_outputs(2050) <= a and not b;
    layer4_outputs(2051) <= not (a and b);
    layer4_outputs(2052) <= not b;
    layer4_outputs(2053) <= not a or b;
    layer4_outputs(2054) <= not b or a;
    layer4_outputs(2055) <= not a or b;
    layer4_outputs(2056) <= a and b;
    layer4_outputs(2057) <= 1'b0;
    layer4_outputs(2058) <= not (a or b);
    layer4_outputs(2059) <= a or b;
    layer4_outputs(2060) <= not b;
    layer4_outputs(2061) <= b and not a;
    layer4_outputs(2062) <= not b or a;
    layer4_outputs(2063) <= 1'b0;
    layer4_outputs(2064) <= a;
    layer4_outputs(2065) <= b;
    layer4_outputs(2066) <= a and not b;
    layer4_outputs(2067) <= not (a or b);
    layer4_outputs(2068) <= a;
    layer4_outputs(2069) <= not a;
    layer4_outputs(2070) <= not b or a;
    layer4_outputs(2071) <= not b;
    layer4_outputs(2072) <= not a or b;
    layer4_outputs(2073) <= not a or b;
    layer4_outputs(2074) <= a;
    layer4_outputs(2075) <= not (a or b);
    layer4_outputs(2076) <= not b;
    layer4_outputs(2077) <= not a;
    layer4_outputs(2078) <= a and b;
    layer4_outputs(2079) <= not b or a;
    layer4_outputs(2080) <= not b;
    layer4_outputs(2081) <= b;
    layer4_outputs(2082) <= not (a and b);
    layer4_outputs(2083) <= a or b;
    layer4_outputs(2084) <= a and not b;
    layer4_outputs(2085) <= not a;
    layer4_outputs(2086) <= not b;
    layer4_outputs(2087) <= not b or a;
    layer4_outputs(2088) <= 1'b1;
    layer4_outputs(2089) <= not b;
    layer4_outputs(2090) <= a or b;
    layer4_outputs(2091) <= a and not b;
    layer4_outputs(2092) <= a and b;
    layer4_outputs(2093) <= not (a and b);
    layer4_outputs(2094) <= b and not a;
    layer4_outputs(2095) <= not a;
    layer4_outputs(2096) <= a or b;
    layer4_outputs(2097) <= not a or b;
    layer4_outputs(2098) <= a and not b;
    layer4_outputs(2099) <= a and b;
    layer4_outputs(2100) <= a or b;
    layer4_outputs(2101) <= not (a and b);
    layer4_outputs(2102) <= not (a xor b);
    layer4_outputs(2103) <= not b;
    layer4_outputs(2104) <= b and not a;
    layer4_outputs(2105) <= a and not b;
    layer4_outputs(2106) <= 1'b0;
    layer4_outputs(2107) <= b;
    layer4_outputs(2108) <= 1'b1;
    layer4_outputs(2109) <= a and b;
    layer4_outputs(2110) <= a and b;
    layer4_outputs(2111) <= not (a and b);
    layer4_outputs(2112) <= a or b;
    layer4_outputs(2113) <= b and not a;
    layer4_outputs(2114) <= not b or a;
    layer4_outputs(2115) <= 1'b1;
    layer4_outputs(2116) <= a and b;
    layer4_outputs(2117) <= a;
    layer4_outputs(2118) <= not (a or b);
    layer4_outputs(2119) <= a and not b;
    layer4_outputs(2120) <= not (a and b);
    layer4_outputs(2121) <= 1'b0;
    layer4_outputs(2122) <= a;
    layer4_outputs(2123) <= 1'b1;
    layer4_outputs(2124) <= not a or b;
    layer4_outputs(2125) <= not b or a;
    layer4_outputs(2126) <= a or b;
    layer4_outputs(2127) <= a;
    layer4_outputs(2128) <= not b or a;
    layer4_outputs(2129) <= 1'b1;
    layer4_outputs(2130) <= b and not a;
    layer4_outputs(2131) <= not a;
    layer4_outputs(2132) <= a xor b;
    layer4_outputs(2133) <= not b or a;
    layer4_outputs(2134) <= a and b;
    layer4_outputs(2135) <= not (a and b);
    layer4_outputs(2136) <= not a or b;
    layer4_outputs(2137) <= not a;
    layer4_outputs(2138) <= not b or a;
    layer4_outputs(2139) <= b;
    layer4_outputs(2140) <= b and not a;
    layer4_outputs(2141) <= not a or b;
    layer4_outputs(2142) <= a and not b;
    layer4_outputs(2143) <= not b or a;
    layer4_outputs(2144) <= not (a and b);
    layer4_outputs(2145) <= not (a and b);
    layer4_outputs(2146) <= not b;
    layer4_outputs(2147) <= not b;
    layer4_outputs(2148) <= a or b;
    layer4_outputs(2149) <= not (a and b);
    layer4_outputs(2150) <= a or b;
    layer4_outputs(2151) <= b;
    layer4_outputs(2152) <= a;
    layer4_outputs(2153) <= 1'b0;
    layer4_outputs(2154) <= not (a xor b);
    layer4_outputs(2155) <= not (a xor b);
    layer4_outputs(2156) <= not b;
    layer4_outputs(2157) <= not (a xor b);
    layer4_outputs(2158) <= a and b;
    layer4_outputs(2159) <= not (a and b);
    layer4_outputs(2160) <= b;
    layer4_outputs(2161) <= a and b;
    layer4_outputs(2162) <= a xor b;
    layer4_outputs(2163) <= not b or a;
    layer4_outputs(2164) <= a and b;
    layer4_outputs(2165) <= a and not b;
    layer4_outputs(2166) <= a;
    layer4_outputs(2167) <= a;
    layer4_outputs(2168) <= 1'b0;
    layer4_outputs(2169) <= not (a or b);
    layer4_outputs(2170) <= not a;
    layer4_outputs(2171) <= not (a xor b);
    layer4_outputs(2172) <= 1'b1;
    layer4_outputs(2173) <= not a;
    layer4_outputs(2174) <= a;
    layer4_outputs(2175) <= not a or b;
    layer4_outputs(2176) <= not (a or b);
    layer4_outputs(2177) <= a;
    layer4_outputs(2178) <= b;
    layer4_outputs(2179) <= a xor b;
    layer4_outputs(2180) <= not (a and b);
    layer4_outputs(2181) <= 1'b1;
    layer4_outputs(2182) <= not (a or b);
    layer4_outputs(2183) <= not a;
    layer4_outputs(2184) <= a and b;
    layer4_outputs(2185) <= not a;
    layer4_outputs(2186) <= 1'b1;
    layer4_outputs(2187) <= not b;
    layer4_outputs(2188) <= a xor b;
    layer4_outputs(2189) <= b and not a;
    layer4_outputs(2190) <= not a;
    layer4_outputs(2191) <= a and not b;
    layer4_outputs(2192) <= a or b;
    layer4_outputs(2193) <= a;
    layer4_outputs(2194) <= a;
    layer4_outputs(2195) <= not a or b;
    layer4_outputs(2196) <= not (a and b);
    layer4_outputs(2197) <= a;
    layer4_outputs(2198) <= a or b;
    layer4_outputs(2199) <= a or b;
    layer4_outputs(2200) <= a and b;
    layer4_outputs(2201) <= not a or b;
    layer4_outputs(2202) <= b;
    layer4_outputs(2203) <= a or b;
    layer4_outputs(2204) <= b and not a;
    layer4_outputs(2205) <= not (a and b);
    layer4_outputs(2206) <= a;
    layer4_outputs(2207) <= a and b;
    layer4_outputs(2208) <= not a;
    layer4_outputs(2209) <= not a;
    layer4_outputs(2210) <= a xor b;
    layer4_outputs(2211) <= a or b;
    layer4_outputs(2212) <= not a;
    layer4_outputs(2213) <= not a;
    layer4_outputs(2214) <= not b or a;
    layer4_outputs(2215) <= not b or a;
    layer4_outputs(2216) <= not (a or b);
    layer4_outputs(2217) <= not (a or b);
    layer4_outputs(2218) <= not (a or b);
    layer4_outputs(2219) <= not a;
    layer4_outputs(2220) <= not a or b;
    layer4_outputs(2221) <= b;
    layer4_outputs(2222) <= b and not a;
    layer4_outputs(2223) <= a or b;
    layer4_outputs(2224) <= not a or b;
    layer4_outputs(2225) <= not a;
    layer4_outputs(2226) <= a xor b;
    layer4_outputs(2227) <= b and not a;
    layer4_outputs(2228) <= not a;
    layer4_outputs(2229) <= b and not a;
    layer4_outputs(2230) <= not (a and b);
    layer4_outputs(2231) <= not b or a;
    layer4_outputs(2232) <= 1'b0;
    layer4_outputs(2233) <= a and not b;
    layer4_outputs(2234) <= not b;
    layer4_outputs(2235) <= a and not b;
    layer4_outputs(2236) <= not a or b;
    layer4_outputs(2237) <= not b;
    layer4_outputs(2238) <= not a;
    layer4_outputs(2239) <= a;
    layer4_outputs(2240) <= b;
    layer4_outputs(2241) <= 1'b1;
    layer4_outputs(2242) <= not (a and b);
    layer4_outputs(2243) <= a or b;
    layer4_outputs(2244) <= 1'b0;
    layer4_outputs(2245) <= not a;
    layer4_outputs(2246) <= not a or b;
    layer4_outputs(2247) <= a and not b;
    layer4_outputs(2248) <= a and not b;
    layer4_outputs(2249) <= not b or a;
    layer4_outputs(2250) <= a or b;
    layer4_outputs(2251) <= not b or a;
    layer4_outputs(2252) <= 1'b0;
    layer4_outputs(2253) <= a and b;
    layer4_outputs(2254) <= not b;
    layer4_outputs(2255) <= not a or b;
    layer4_outputs(2256) <= a xor b;
    layer4_outputs(2257) <= b;
    layer4_outputs(2258) <= not a;
    layer4_outputs(2259) <= not b or a;
    layer4_outputs(2260) <= 1'b0;
    layer4_outputs(2261) <= 1'b0;
    layer4_outputs(2262) <= a or b;
    layer4_outputs(2263) <= b and not a;
    layer4_outputs(2264) <= not a;
    layer4_outputs(2265) <= a;
    layer4_outputs(2266) <= 1'b1;
    layer4_outputs(2267) <= b;
    layer4_outputs(2268) <= not b;
    layer4_outputs(2269) <= b and not a;
    layer4_outputs(2270) <= not (a xor b);
    layer4_outputs(2271) <= a and b;
    layer4_outputs(2272) <= not a;
    layer4_outputs(2273) <= not a;
    layer4_outputs(2274) <= a or b;
    layer4_outputs(2275) <= not a or b;
    layer4_outputs(2276) <= a and b;
    layer4_outputs(2277) <= a;
    layer4_outputs(2278) <= b;
    layer4_outputs(2279) <= a;
    layer4_outputs(2280) <= a;
    layer4_outputs(2281) <= not (a or b);
    layer4_outputs(2282) <= 1'b1;
    layer4_outputs(2283) <= not a or b;
    layer4_outputs(2284) <= a;
    layer4_outputs(2285) <= not b or a;
    layer4_outputs(2286) <= a;
    layer4_outputs(2287) <= b;
    layer4_outputs(2288) <= not (a and b);
    layer4_outputs(2289) <= not a;
    layer4_outputs(2290) <= a xor b;
    layer4_outputs(2291) <= not (a xor b);
    layer4_outputs(2292) <= b;
    layer4_outputs(2293) <= not a;
    layer4_outputs(2294) <= not a or b;
    layer4_outputs(2295) <= not a or b;
    layer4_outputs(2296) <= 1'b0;
    layer4_outputs(2297) <= not (a and b);
    layer4_outputs(2298) <= a;
    layer4_outputs(2299) <= a;
    layer4_outputs(2300) <= not (a and b);
    layer4_outputs(2301) <= 1'b1;
    layer4_outputs(2302) <= not (a xor b);
    layer4_outputs(2303) <= b;
    layer4_outputs(2304) <= a xor b;
    layer4_outputs(2305) <= not (a or b);
    layer4_outputs(2306) <= 1'b1;
    layer4_outputs(2307) <= not a or b;
    layer4_outputs(2308) <= not (a and b);
    layer4_outputs(2309) <= b and not a;
    layer4_outputs(2310) <= 1'b0;
    layer4_outputs(2311) <= not b;
    layer4_outputs(2312) <= not (a and b);
    layer4_outputs(2313) <= not b or a;
    layer4_outputs(2314) <= not a;
    layer4_outputs(2315) <= not (a or b);
    layer4_outputs(2316) <= b;
    layer4_outputs(2317) <= a;
    layer4_outputs(2318) <= a and b;
    layer4_outputs(2319) <= a or b;
    layer4_outputs(2320) <= a or b;
    layer4_outputs(2321) <= not b;
    layer4_outputs(2322) <= not a;
    layer4_outputs(2323) <= not a;
    layer4_outputs(2324) <= not b;
    layer4_outputs(2325) <= b and not a;
    layer4_outputs(2326) <= a or b;
    layer4_outputs(2327) <= b and not a;
    layer4_outputs(2328) <= a and not b;
    layer4_outputs(2329) <= not b or a;
    layer4_outputs(2330) <= not (a or b);
    layer4_outputs(2331) <= not a or b;
    layer4_outputs(2332) <= a and b;
    layer4_outputs(2333) <= not (a or b);
    layer4_outputs(2334) <= 1'b0;
    layer4_outputs(2335) <= b;
    layer4_outputs(2336) <= not b;
    layer4_outputs(2337) <= not (a and b);
    layer4_outputs(2338) <= not b or a;
    layer4_outputs(2339) <= a or b;
    layer4_outputs(2340) <= 1'b1;
    layer4_outputs(2341) <= not a;
    layer4_outputs(2342) <= not a or b;
    layer4_outputs(2343) <= not b;
    layer4_outputs(2344) <= a;
    layer4_outputs(2345) <= b;
    layer4_outputs(2346) <= b and not a;
    layer4_outputs(2347) <= a or b;
    layer4_outputs(2348) <= a and b;
    layer4_outputs(2349) <= not (a and b);
    layer4_outputs(2350) <= not (a or b);
    layer4_outputs(2351) <= not a;
    layer4_outputs(2352) <= 1'b1;
    layer4_outputs(2353) <= b;
    layer4_outputs(2354) <= b;
    layer4_outputs(2355) <= a and not b;
    layer4_outputs(2356) <= not a;
    layer4_outputs(2357) <= a;
    layer4_outputs(2358) <= a and b;
    layer4_outputs(2359) <= b;
    layer4_outputs(2360) <= not a or b;
    layer4_outputs(2361) <= not b;
    layer4_outputs(2362) <= a and b;
    layer4_outputs(2363) <= not a;
    layer4_outputs(2364) <= a;
    layer4_outputs(2365) <= a;
    layer4_outputs(2366) <= b;
    layer4_outputs(2367) <= 1'b0;
    layer4_outputs(2368) <= a and not b;
    layer4_outputs(2369) <= not b or a;
    layer4_outputs(2370) <= 1'b1;
    layer4_outputs(2371) <= not b or a;
    layer4_outputs(2372) <= b;
    layer4_outputs(2373) <= a xor b;
    layer4_outputs(2374) <= b;
    layer4_outputs(2375) <= b;
    layer4_outputs(2376) <= not (a and b);
    layer4_outputs(2377) <= 1'b1;
    layer4_outputs(2378) <= not (a xor b);
    layer4_outputs(2379) <= not a;
    layer4_outputs(2380) <= b;
    layer4_outputs(2381) <= not a;
    layer4_outputs(2382) <= a or b;
    layer4_outputs(2383) <= a and b;
    layer4_outputs(2384) <= 1'b1;
    layer4_outputs(2385) <= not a or b;
    layer4_outputs(2386) <= b and not a;
    layer4_outputs(2387) <= b and not a;
    layer4_outputs(2388) <= a and b;
    layer4_outputs(2389) <= a xor b;
    layer4_outputs(2390) <= 1'b0;
    layer4_outputs(2391) <= b and not a;
    layer4_outputs(2392) <= b;
    layer4_outputs(2393) <= not a or b;
    layer4_outputs(2394) <= not (a xor b);
    layer4_outputs(2395) <= not b or a;
    layer4_outputs(2396) <= a and b;
    layer4_outputs(2397) <= a or b;
    layer4_outputs(2398) <= not a or b;
    layer4_outputs(2399) <= not (a or b);
    layer4_outputs(2400) <= 1'b0;
    layer4_outputs(2401) <= not b;
    layer4_outputs(2402) <= not a or b;
    layer4_outputs(2403) <= not (a and b);
    layer4_outputs(2404) <= not a or b;
    layer4_outputs(2405) <= not a;
    layer4_outputs(2406) <= b and not a;
    layer4_outputs(2407) <= b;
    layer4_outputs(2408) <= not a or b;
    layer4_outputs(2409) <= b;
    layer4_outputs(2410) <= 1'b1;
    layer4_outputs(2411) <= 1'b1;
    layer4_outputs(2412) <= a xor b;
    layer4_outputs(2413) <= not b;
    layer4_outputs(2414) <= a xor b;
    layer4_outputs(2415) <= not a or b;
    layer4_outputs(2416) <= 1'b0;
    layer4_outputs(2417) <= not b;
    layer4_outputs(2418) <= a and not b;
    layer4_outputs(2419) <= 1'b0;
    layer4_outputs(2420) <= a;
    layer4_outputs(2421) <= not (a and b);
    layer4_outputs(2422) <= a or b;
    layer4_outputs(2423) <= a;
    layer4_outputs(2424) <= not a;
    layer4_outputs(2425) <= b;
    layer4_outputs(2426) <= not b or a;
    layer4_outputs(2427) <= 1'b1;
    layer4_outputs(2428) <= a and b;
    layer4_outputs(2429) <= a and not b;
    layer4_outputs(2430) <= a and b;
    layer4_outputs(2431) <= not a;
    layer4_outputs(2432) <= not a;
    layer4_outputs(2433) <= 1'b0;
    layer4_outputs(2434) <= a;
    layer4_outputs(2435) <= a;
    layer4_outputs(2436) <= 1'b0;
    layer4_outputs(2437) <= not a or b;
    layer4_outputs(2438) <= a and b;
    layer4_outputs(2439) <= b;
    layer4_outputs(2440) <= 1'b1;
    layer4_outputs(2441) <= a and not b;
    layer4_outputs(2442) <= not (a xor b);
    layer4_outputs(2443) <= a or b;
    layer4_outputs(2444) <= 1'b1;
    layer4_outputs(2445) <= not (a xor b);
    layer4_outputs(2446) <= a;
    layer4_outputs(2447) <= not b;
    layer4_outputs(2448) <= not (a and b);
    layer4_outputs(2449) <= 1'b1;
    layer4_outputs(2450) <= not a;
    layer4_outputs(2451) <= not a or b;
    layer4_outputs(2452) <= not b or a;
    layer4_outputs(2453) <= not b;
    layer4_outputs(2454) <= a and b;
    layer4_outputs(2455) <= 1'b0;
    layer4_outputs(2456) <= a and b;
    layer4_outputs(2457) <= b;
    layer4_outputs(2458) <= 1'b0;
    layer4_outputs(2459) <= not (a and b);
    layer4_outputs(2460) <= b and not a;
    layer4_outputs(2461) <= not b;
    layer4_outputs(2462) <= not (a or b);
    layer4_outputs(2463) <= a;
    layer4_outputs(2464) <= b and not a;
    layer4_outputs(2465) <= not b;
    layer4_outputs(2466) <= a or b;
    layer4_outputs(2467) <= not a or b;
    layer4_outputs(2468) <= b;
    layer4_outputs(2469) <= a and not b;
    layer4_outputs(2470) <= 1'b1;
    layer4_outputs(2471) <= 1'b0;
    layer4_outputs(2472) <= a and not b;
    layer4_outputs(2473) <= not a or b;
    layer4_outputs(2474) <= not b;
    layer4_outputs(2475) <= a and not b;
    layer4_outputs(2476) <= not a or b;
    layer4_outputs(2477) <= b;
    layer4_outputs(2478) <= not (a and b);
    layer4_outputs(2479) <= a and not b;
    layer4_outputs(2480) <= a and b;
    layer4_outputs(2481) <= not b or a;
    layer4_outputs(2482) <= a and b;
    layer4_outputs(2483) <= b and not a;
    layer4_outputs(2484) <= not a;
    layer4_outputs(2485) <= a and not b;
    layer4_outputs(2486) <= a and not b;
    layer4_outputs(2487) <= a;
    layer4_outputs(2488) <= 1'b0;
    layer4_outputs(2489) <= not a;
    layer4_outputs(2490) <= a and not b;
    layer4_outputs(2491) <= not (a and b);
    layer4_outputs(2492) <= a;
    layer4_outputs(2493) <= a and b;
    layer4_outputs(2494) <= 1'b0;
    layer4_outputs(2495) <= a and not b;
    layer4_outputs(2496) <= not b;
    layer4_outputs(2497) <= b;
    layer4_outputs(2498) <= b and not a;
    layer4_outputs(2499) <= not (a xor b);
    layer4_outputs(2500) <= not a;
    layer4_outputs(2501) <= not (a xor b);
    layer4_outputs(2502) <= b and not a;
    layer4_outputs(2503) <= 1'b1;
    layer4_outputs(2504) <= a or b;
    layer4_outputs(2505) <= not b or a;
    layer4_outputs(2506) <= b;
    layer4_outputs(2507) <= 1'b0;
    layer4_outputs(2508) <= a or b;
    layer4_outputs(2509) <= a and not b;
    layer4_outputs(2510) <= not a or b;
    layer4_outputs(2511) <= not (a or b);
    layer4_outputs(2512) <= a;
    layer4_outputs(2513) <= not a or b;
    layer4_outputs(2514) <= a;
    layer4_outputs(2515) <= b and not a;
    layer4_outputs(2516) <= a or b;
    layer4_outputs(2517) <= not a;
    layer4_outputs(2518) <= 1'b0;
    layer4_outputs(2519) <= a;
    layer4_outputs(2520) <= not a;
    layer4_outputs(2521) <= not (a or b);
    layer4_outputs(2522) <= a and b;
    layer4_outputs(2523) <= b;
    layer4_outputs(2524) <= not (a or b);
    layer4_outputs(2525) <= a;
    layer4_outputs(2526) <= 1'b1;
    layer4_outputs(2527) <= a;
    layer4_outputs(2528) <= not a;
    layer4_outputs(2529) <= 1'b1;
    layer4_outputs(2530) <= not b or a;
    layer4_outputs(2531) <= not a;
    layer4_outputs(2532) <= b;
    layer4_outputs(2533) <= 1'b0;
    layer4_outputs(2534) <= not a;
    layer4_outputs(2535) <= 1'b1;
    layer4_outputs(2536) <= not a or b;
    layer4_outputs(2537) <= a and not b;
    layer4_outputs(2538) <= 1'b1;
    layer4_outputs(2539) <= 1'b0;
    layer4_outputs(2540) <= not a or b;
    layer4_outputs(2541) <= not (a xor b);
    layer4_outputs(2542) <= a;
    layer4_outputs(2543) <= a or b;
    layer4_outputs(2544) <= not (a and b);
    layer4_outputs(2545) <= not (a or b);
    layer4_outputs(2546) <= 1'b0;
    layer4_outputs(2547) <= 1'b1;
    layer4_outputs(2548) <= a and b;
    layer4_outputs(2549) <= 1'b0;
    layer4_outputs(2550) <= a;
    layer4_outputs(2551) <= b and not a;
    layer4_outputs(2552) <= not (a and b);
    layer4_outputs(2553) <= b and not a;
    layer4_outputs(2554) <= a and b;
    layer4_outputs(2555) <= not a or b;
    layer4_outputs(2556) <= b;
    layer4_outputs(2557) <= a or b;
    layer4_outputs(2558) <= b and not a;
    layer4_outputs(2559) <= b and not a;
    layer4_outputs(2560) <= a and b;
    layer4_outputs(2561) <= not (a or b);
    layer4_outputs(2562) <= not b;
    layer4_outputs(2563) <= a and not b;
    layer4_outputs(2564) <= 1'b1;
    layer4_outputs(2565) <= not b;
    layer4_outputs(2566) <= not a;
    layer4_outputs(2567) <= not a or b;
    layer4_outputs(2568) <= not b;
    layer4_outputs(2569) <= not (a and b);
    layer4_outputs(2570) <= a and not b;
    layer4_outputs(2571) <= a and b;
    layer4_outputs(2572) <= not b;
    layer4_outputs(2573) <= b and not a;
    layer4_outputs(2574) <= a;
    layer4_outputs(2575) <= b;
    layer4_outputs(2576) <= not b;
    layer4_outputs(2577) <= not b;
    layer4_outputs(2578) <= not b or a;
    layer4_outputs(2579) <= not b or a;
    layer4_outputs(2580) <= b and not a;
    layer4_outputs(2581) <= 1'b1;
    layer4_outputs(2582) <= a;
    layer4_outputs(2583) <= not (a and b);
    layer4_outputs(2584) <= not b or a;
    layer4_outputs(2585) <= a and not b;
    layer4_outputs(2586) <= not a;
    layer4_outputs(2587) <= not (a and b);
    layer4_outputs(2588) <= b and not a;
    layer4_outputs(2589) <= not a;
    layer4_outputs(2590) <= not (a or b);
    layer4_outputs(2591) <= a and b;
    layer4_outputs(2592) <= not (a and b);
    layer4_outputs(2593) <= a;
    layer4_outputs(2594) <= not a;
    layer4_outputs(2595) <= a and b;
    layer4_outputs(2596) <= 1'b1;
    layer4_outputs(2597) <= not b;
    layer4_outputs(2598) <= not (a or b);
    layer4_outputs(2599) <= a or b;
    layer4_outputs(2600) <= not a or b;
    layer4_outputs(2601) <= b and not a;
    layer4_outputs(2602) <= a and b;
    layer4_outputs(2603) <= not (a and b);
    layer4_outputs(2604) <= b;
    layer4_outputs(2605) <= not (a and b);
    layer4_outputs(2606) <= not b or a;
    layer4_outputs(2607) <= not a;
    layer4_outputs(2608) <= not b or a;
    layer4_outputs(2609) <= a xor b;
    layer4_outputs(2610) <= a and not b;
    layer4_outputs(2611) <= not b;
    layer4_outputs(2612) <= not b or a;
    layer4_outputs(2613) <= not a or b;
    layer4_outputs(2614) <= a or b;
    layer4_outputs(2615) <= b and not a;
    layer4_outputs(2616) <= not (a and b);
    layer4_outputs(2617) <= b and not a;
    layer4_outputs(2618) <= not (a and b);
    layer4_outputs(2619) <= not a or b;
    layer4_outputs(2620) <= b;
    layer4_outputs(2621) <= not (a or b);
    layer4_outputs(2622) <= a;
    layer4_outputs(2623) <= a xor b;
    layer4_outputs(2624) <= not a;
    layer4_outputs(2625) <= 1'b1;
    layer4_outputs(2626) <= b;
    layer4_outputs(2627) <= a xor b;
    layer4_outputs(2628) <= b;
    layer4_outputs(2629) <= b and not a;
    layer4_outputs(2630) <= a and b;
    layer4_outputs(2631) <= a;
    layer4_outputs(2632) <= a and not b;
    layer4_outputs(2633) <= 1'b1;
    layer4_outputs(2634) <= not (a and b);
    layer4_outputs(2635) <= a or b;
    layer4_outputs(2636) <= b and not a;
    layer4_outputs(2637) <= not a;
    layer4_outputs(2638) <= not b;
    layer4_outputs(2639) <= a;
    layer4_outputs(2640) <= not b;
    layer4_outputs(2641) <= a and not b;
    layer4_outputs(2642) <= not a;
    layer4_outputs(2643) <= a and not b;
    layer4_outputs(2644) <= not (a or b);
    layer4_outputs(2645) <= 1'b0;
    layer4_outputs(2646) <= not b or a;
    layer4_outputs(2647) <= not (a and b);
    layer4_outputs(2648) <= not (a xor b);
    layer4_outputs(2649) <= not (a and b);
    layer4_outputs(2650) <= not a or b;
    layer4_outputs(2651) <= not a;
    layer4_outputs(2652) <= not a;
    layer4_outputs(2653) <= not (a and b);
    layer4_outputs(2654) <= a and b;
    layer4_outputs(2655) <= not (a or b);
    layer4_outputs(2656) <= a;
    layer4_outputs(2657) <= not b or a;
    layer4_outputs(2658) <= not (a or b);
    layer4_outputs(2659) <= not a;
    layer4_outputs(2660) <= a;
    layer4_outputs(2661) <= a xor b;
    layer4_outputs(2662) <= not a or b;
    layer4_outputs(2663) <= not a;
    layer4_outputs(2664) <= 1'b0;
    layer4_outputs(2665) <= a or b;
    layer4_outputs(2666) <= b and not a;
    layer4_outputs(2667) <= not (a xor b);
    layer4_outputs(2668) <= not (a and b);
    layer4_outputs(2669) <= a;
    layer4_outputs(2670) <= a and not b;
    layer4_outputs(2671) <= a and not b;
    layer4_outputs(2672) <= not (a and b);
    layer4_outputs(2673) <= b;
    layer4_outputs(2674) <= not b;
    layer4_outputs(2675) <= a or b;
    layer4_outputs(2676) <= a and not b;
    layer4_outputs(2677) <= not (a or b);
    layer4_outputs(2678) <= b;
    layer4_outputs(2679) <= not (a xor b);
    layer4_outputs(2680) <= not (a xor b);
    layer4_outputs(2681) <= a or b;
    layer4_outputs(2682) <= a or b;
    layer4_outputs(2683) <= a or b;
    layer4_outputs(2684) <= 1'b1;
    layer4_outputs(2685) <= 1'b0;
    layer4_outputs(2686) <= a or b;
    layer4_outputs(2687) <= a and b;
    layer4_outputs(2688) <= not a or b;
    layer4_outputs(2689) <= b;
    layer4_outputs(2690) <= not a;
    layer4_outputs(2691) <= a;
    layer4_outputs(2692) <= b and not a;
    layer4_outputs(2693) <= a xor b;
    layer4_outputs(2694) <= a or b;
    layer4_outputs(2695) <= a and b;
    layer4_outputs(2696) <= a and b;
    layer4_outputs(2697) <= not a;
    layer4_outputs(2698) <= not b or a;
    layer4_outputs(2699) <= not (a and b);
    layer4_outputs(2700) <= a or b;
    layer4_outputs(2701) <= a and not b;
    layer4_outputs(2702) <= b;
    layer4_outputs(2703) <= not (a or b);
    layer4_outputs(2704) <= b;
    layer4_outputs(2705) <= 1'b1;
    layer4_outputs(2706) <= not b or a;
    layer4_outputs(2707) <= a;
    layer4_outputs(2708) <= b and not a;
    layer4_outputs(2709) <= a xor b;
    layer4_outputs(2710) <= not a;
    layer4_outputs(2711) <= a and b;
    layer4_outputs(2712) <= not (a or b);
    layer4_outputs(2713) <= not a or b;
    layer4_outputs(2714) <= not a or b;
    layer4_outputs(2715) <= b;
    layer4_outputs(2716) <= a and not b;
    layer4_outputs(2717) <= not (a xor b);
    layer4_outputs(2718) <= 1'b0;
    layer4_outputs(2719) <= b;
    layer4_outputs(2720) <= 1'b0;
    layer4_outputs(2721) <= not (a or b);
    layer4_outputs(2722) <= not (a or b);
    layer4_outputs(2723) <= not a or b;
    layer4_outputs(2724) <= not a or b;
    layer4_outputs(2725) <= 1'b1;
    layer4_outputs(2726) <= not (a or b);
    layer4_outputs(2727) <= a and b;
    layer4_outputs(2728) <= b;
    layer4_outputs(2729) <= a and b;
    layer4_outputs(2730) <= a or b;
    layer4_outputs(2731) <= not a;
    layer4_outputs(2732) <= a or b;
    layer4_outputs(2733) <= a and not b;
    layer4_outputs(2734) <= 1'b0;
    layer4_outputs(2735) <= not (a or b);
    layer4_outputs(2736) <= a xor b;
    layer4_outputs(2737) <= not b;
    layer4_outputs(2738) <= not (a and b);
    layer4_outputs(2739) <= a and b;
    layer4_outputs(2740) <= not (a or b);
    layer4_outputs(2741) <= b and not a;
    layer4_outputs(2742) <= not (a xor b);
    layer4_outputs(2743) <= 1'b0;
    layer4_outputs(2744) <= a and not b;
    layer4_outputs(2745) <= b;
    layer4_outputs(2746) <= 1'b1;
    layer4_outputs(2747) <= a and not b;
    layer4_outputs(2748) <= not (a or b);
    layer4_outputs(2749) <= not a;
    layer4_outputs(2750) <= a or b;
    layer4_outputs(2751) <= not (a xor b);
    layer4_outputs(2752) <= not (a and b);
    layer4_outputs(2753) <= b and not a;
    layer4_outputs(2754) <= 1'b1;
    layer4_outputs(2755) <= b and not a;
    layer4_outputs(2756) <= a;
    layer4_outputs(2757) <= a or b;
    layer4_outputs(2758) <= a or b;
    layer4_outputs(2759) <= a and b;
    layer4_outputs(2760) <= not (a or b);
    layer4_outputs(2761) <= not b;
    layer4_outputs(2762) <= not (a and b);
    layer4_outputs(2763) <= b and not a;
    layer4_outputs(2764) <= a or b;
    layer4_outputs(2765) <= 1'b1;
    layer4_outputs(2766) <= not (a and b);
    layer4_outputs(2767) <= 1'b0;
    layer4_outputs(2768) <= b;
    layer4_outputs(2769) <= a;
    layer4_outputs(2770) <= not (a and b);
    layer4_outputs(2771) <= a xor b;
    layer4_outputs(2772) <= 1'b0;
    layer4_outputs(2773) <= not (a or b);
    layer4_outputs(2774) <= b;
    layer4_outputs(2775) <= 1'b0;
    layer4_outputs(2776) <= b and not a;
    layer4_outputs(2777) <= not (a or b);
    layer4_outputs(2778) <= a;
    layer4_outputs(2779) <= not (a xor b);
    layer4_outputs(2780) <= not (a and b);
    layer4_outputs(2781) <= a and b;
    layer4_outputs(2782) <= not a or b;
    layer4_outputs(2783) <= b and not a;
    layer4_outputs(2784) <= not b;
    layer4_outputs(2785) <= a and not b;
    layer4_outputs(2786) <= not (a or b);
    layer4_outputs(2787) <= b and not a;
    layer4_outputs(2788) <= a and not b;
    layer4_outputs(2789) <= not b;
    layer4_outputs(2790) <= 1'b1;
    layer4_outputs(2791) <= not (a and b);
    layer4_outputs(2792) <= not a or b;
    layer4_outputs(2793) <= not b or a;
    layer4_outputs(2794) <= 1'b0;
    layer4_outputs(2795) <= not (a or b);
    layer4_outputs(2796) <= 1'b1;
    layer4_outputs(2797) <= a;
    layer4_outputs(2798) <= b;
    layer4_outputs(2799) <= b;
    layer4_outputs(2800) <= a xor b;
    layer4_outputs(2801) <= not (a or b);
    layer4_outputs(2802) <= a;
    layer4_outputs(2803) <= a and b;
    layer4_outputs(2804) <= not (a and b);
    layer4_outputs(2805) <= b and not a;
    layer4_outputs(2806) <= not b or a;
    layer4_outputs(2807) <= b;
    layer4_outputs(2808) <= a and b;
    layer4_outputs(2809) <= not b;
    layer4_outputs(2810) <= not (a and b);
    layer4_outputs(2811) <= not b;
    layer4_outputs(2812) <= a;
    layer4_outputs(2813) <= a and not b;
    layer4_outputs(2814) <= not (a or b);
    layer4_outputs(2815) <= not (a and b);
    layer4_outputs(2816) <= a and b;
    layer4_outputs(2817) <= 1'b1;
    layer4_outputs(2818) <= not a;
    layer4_outputs(2819) <= a and not b;
    layer4_outputs(2820) <= a and not b;
    layer4_outputs(2821) <= b;
    layer4_outputs(2822) <= 1'b0;
    layer4_outputs(2823) <= not b or a;
    layer4_outputs(2824) <= not b;
    layer4_outputs(2825) <= a and b;
    layer4_outputs(2826) <= not (a and b);
    layer4_outputs(2827) <= not (a xor b);
    layer4_outputs(2828) <= 1'b0;
    layer4_outputs(2829) <= a and b;
    layer4_outputs(2830) <= not b;
    layer4_outputs(2831) <= b and not a;
    layer4_outputs(2832) <= 1'b0;
    layer4_outputs(2833) <= b and not a;
    layer4_outputs(2834) <= a or b;
    layer4_outputs(2835) <= a xor b;
    layer4_outputs(2836) <= 1'b0;
    layer4_outputs(2837) <= b and not a;
    layer4_outputs(2838) <= a and not b;
    layer4_outputs(2839) <= a and not b;
    layer4_outputs(2840) <= not (a or b);
    layer4_outputs(2841) <= not a;
    layer4_outputs(2842) <= 1'b1;
    layer4_outputs(2843) <= not (a or b);
    layer4_outputs(2844) <= a xor b;
    layer4_outputs(2845) <= b and not a;
    layer4_outputs(2846) <= not a or b;
    layer4_outputs(2847) <= not a or b;
    layer4_outputs(2848) <= not a;
    layer4_outputs(2849) <= not (a and b);
    layer4_outputs(2850) <= not (a and b);
    layer4_outputs(2851) <= not b;
    layer4_outputs(2852) <= a or b;
    layer4_outputs(2853) <= b;
    layer4_outputs(2854) <= not b;
    layer4_outputs(2855) <= 1'b1;
    layer4_outputs(2856) <= not b or a;
    layer4_outputs(2857) <= a and b;
    layer4_outputs(2858) <= 1'b0;
    layer4_outputs(2859) <= a and not b;
    layer4_outputs(2860) <= a and not b;
    layer4_outputs(2861) <= not a;
    layer4_outputs(2862) <= a;
    layer4_outputs(2863) <= b and not a;
    layer4_outputs(2864) <= a;
    layer4_outputs(2865) <= not (a or b);
    layer4_outputs(2866) <= a and not b;
    layer4_outputs(2867) <= not b or a;
    layer4_outputs(2868) <= not b or a;
    layer4_outputs(2869) <= a and not b;
    layer4_outputs(2870) <= not a;
    layer4_outputs(2871) <= not a;
    layer4_outputs(2872) <= not b or a;
    layer4_outputs(2873) <= not b;
    layer4_outputs(2874) <= b;
    layer4_outputs(2875) <= not b or a;
    layer4_outputs(2876) <= a and b;
    layer4_outputs(2877) <= 1'b0;
    layer4_outputs(2878) <= not a or b;
    layer4_outputs(2879) <= a;
    layer4_outputs(2880) <= not a;
    layer4_outputs(2881) <= b and not a;
    layer4_outputs(2882) <= not (a and b);
    layer4_outputs(2883) <= a and not b;
    layer4_outputs(2884) <= a;
    layer4_outputs(2885) <= not a or b;
    layer4_outputs(2886) <= not (a or b);
    layer4_outputs(2887) <= not b;
    layer4_outputs(2888) <= a and b;
    layer4_outputs(2889) <= b;
    layer4_outputs(2890) <= not a or b;
    layer4_outputs(2891) <= a xor b;
    layer4_outputs(2892) <= not a or b;
    layer4_outputs(2893) <= not b;
    layer4_outputs(2894) <= not a;
    layer4_outputs(2895) <= b;
    layer4_outputs(2896) <= b and not a;
    layer4_outputs(2897) <= not (a or b);
    layer4_outputs(2898) <= b;
    layer4_outputs(2899) <= not (a or b);
    layer4_outputs(2900) <= a and not b;
    layer4_outputs(2901) <= b;
    layer4_outputs(2902) <= not (a xor b);
    layer4_outputs(2903) <= not (a and b);
    layer4_outputs(2904) <= 1'b0;
    layer4_outputs(2905) <= not a;
    layer4_outputs(2906) <= not a;
    layer4_outputs(2907) <= 1'b1;
    layer4_outputs(2908) <= not (a or b);
    layer4_outputs(2909) <= 1'b1;
    layer4_outputs(2910) <= not (a or b);
    layer4_outputs(2911) <= b;
    layer4_outputs(2912) <= a and b;
    layer4_outputs(2913) <= 1'b1;
    layer4_outputs(2914) <= 1'b0;
    layer4_outputs(2915) <= b;
    layer4_outputs(2916) <= not a;
    layer4_outputs(2917) <= a;
    layer4_outputs(2918) <= b;
    layer4_outputs(2919) <= not (a and b);
    layer4_outputs(2920) <= a;
    layer4_outputs(2921) <= b and not a;
    layer4_outputs(2922) <= 1'b1;
    layer4_outputs(2923) <= a or b;
    layer4_outputs(2924) <= not a;
    layer4_outputs(2925) <= b and not a;
    layer4_outputs(2926) <= a or b;
    layer4_outputs(2927) <= b;
    layer4_outputs(2928) <= not a;
    layer4_outputs(2929) <= b;
    layer4_outputs(2930) <= not a or b;
    layer4_outputs(2931) <= a or b;
    layer4_outputs(2932) <= a and not b;
    layer4_outputs(2933) <= a or b;
    layer4_outputs(2934) <= a;
    layer4_outputs(2935) <= not a or b;
    layer4_outputs(2936) <= a or b;
    layer4_outputs(2937) <= 1'b1;
    layer4_outputs(2938) <= not a;
    layer4_outputs(2939) <= b;
    layer4_outputs(2940) <= a and b;
    layer4_outputs(2941) <= 1'b0;
    layer4_outputs(2942) <= not a or b;
    layer4_outputs(2943) <= 1'b0;
    layer4_outputs(2944) <= a and not b;
    layer4_outputs(2945) <= a and not b;
    layer4_outputs(2946) <= a and b;
    layer4_outputs(2947) <= not a;
    layer4_outputs(2948) <= not a;
    layer4_outputs(2949) <= 1'b0;
    layer4_outputs(2950) <= not (a and b);
    layer4_outputs(2951) <= not a or b;
    layer4_outputs(2952) <= not a;
    layer4_outputs(2953) <= not b;
    layer4_outputs(2954) <= not b or a;
    layer4_outputs(2955) <= not a;
    layer4_outputs(2956) <= a;
    layer4_outputs(2957) <= a;
    layer4_outputs(2958) <= a or b;
    layer4_outputs(2959) <= a or b;
    layer4_outputs(2960) <= not b or a;
    layer4_outputs(2961) <= not (a and b);
    layer4_outputs(2962) <= 1'b1;
    layer4_outputs(2963) <= not a or b;
    layer4_outputs(2964) <= b;
    layer4_outputs(2965) <= not b or a;
    layer4_outputs(2966) <= not b or a;
    layer4_outputs(2967) <= not a;
    layer4_outputs(2968) <= not a;
    layer4_outputs(2969) <= not a;
    layer4_outputs(2970) <= not a;
    layer4_outputs(2971) <= not (a or b);
    layer4_outputs(2972) <= a;
    layer4_outputs(2973) <= a or b;
    layer4_outputs(2974) <= b;
    layer4_outputs(2975) <= a or b;
    layer4_outputs(2976) <= a;
    layer4_outputs(2977) <= a;
    layer4_outputs(2978) <= 1'b0;
    layer4_outputs(2979) <= a or b;
    layer4_outputs(2980) <= a and b;
    layer4_outputs(2981) <= not (a and b);
    layer4_outputs(2982) <= not b or a;
    layer4_outputs(2983) <= b;
    layer4_outputs(2984) <= a xor b;
    layer4_outputs(2985) <= b;
    layer4_outputs(2986) <= a or b;
    layer4_outputs(2987) <= a and b;
    layer4_outputs(2988) <= not (a or b);
    layer4_outputs(2989) <= a;
    layer4_outputs(2990) <= a and b;
    layer4_outputs(2991) <= a;
    layer4_outputs(2992) <= b;
    layer4_outputs(2993) <= a or b;
    layer4_outputs(2994) <= not a;
    layer4_outputs(2995) <= 1'b0;
    layer4_outputs(2996) <= 1'b1;
    layer4_outputs(2997) <= not a;
    layer4_outputs(2998) <= not b or a;
    layer4_outputs(2999) <= not (a and b);
    layer4_outputs(3000) <= a and b;
    layer4_outputs(3001) <= a and b;
    layer4_outputs(3002) <= not (a or b);
    layer4_outputs(3003) <= a or b;
    layer4_outputs(3004) <= not b or a;
    layer4_outputs(3005) <= a or b;
    layer4_outputs(3006) <= b and not a;
    layer4_outputs(3007) <= not a;
    layer4_outputs(3008) <= a and b;
    layer4_outputs(3009) <= not (a and b);
    layer4_outputs(3010) <= b and not a;
    layer4_outputs(3011) <= 1'b1;
    layer4_outputs(3012) <= a and not b;
    layer4_outputs(3013) <= 1'b1;
    layer4_outputs(3014) <= a and b;
    layer4_outputs(3015) <= a;
    layer4_outputs(3016) <= a and b;
    layer4_outputs(3017) <= a xor b;
    layer4_outputs(3018) <= not (a or b);
    layer4_outputs(3019) <= not (a xor b);
    layer4_outputs(3020) <= 1'b1;
    layer4_outputs(3021) <= not b;
    layer4_outputs(3022) <= 1'b1;
    layer4_outputs(3023) <= a and b;
    layer4_outputs(3024) <= not b;
    layer4_outputs(3025) <= not (a or b);
    layer4_outputs(3026) <= a and not b;
    layer4_outputs(3027) <= not (a and b);
    layer4_outputs(3028) <= not (a or b);
    layer4_outputs(3029) <= a;
    layer4_outputs(3030) <= 1'b0;
    layer4_outputs(3031) <= not a;
    layer4_outputs(3032) <= a xor b;
    layer4_outputs(3033) <= not (a or b);
    layer4_outputs(3034) <= not a;
    layer4_outputs(3035) <= not a;
    layer4_outputs(3036) <= a and b;
    layer4_outputs(3037) <= b;
    layer4_outputs(3038) <= not b or a;
    layer4_outputs(3039) <= not a or b;
    layer4_outputs(3040) <= 1'b0;
    layer4_outputs(3041) <= a and b;
    layer4_outputs(3042) <= a or b;
    layer4_outputs(3043) <= 1'b1;
    layer4_outputs(3044) <= a;
    layer4_outputs(3045) <= not (a and b);
    layer4_outputs(3046) <= not (a and b);
    layer4_outputs(3047) <= not b;
    layer4_outputs(3048) <= not a or b;
    layer4_outputs(3049) <= not (a xor b);
    layer4_outputs(3050) <= not b or a;
    layer4_outputs(3051) <= not (a or b);
    layer4_outputs(3052) <= not (a or b);
    layer4_outputs(3053) <= a;
    layer4_outputs(3054) <= not a or b;
    layer4_outputs(3055) <= not b or a;
    layer4_outputs(3056) <= b;
    layer4_outputs(3057) <= a;
    layer4_outputs(3058) <= not b or a;
    layer4_outputs(3059) <= a and b;
    layer4_outputs(3060) <= not a or b;
    layer4_outputs(3061) <= 1'b1;
    layer4_outputs(3062) <= 1'b0;
    layer4_outputs(3063) <= not b;
    layer4_outputs(3064) <= b;
    layer4_outputs(3065) <= not a;
    layer4_outputs(3066) <= a;
    layer4_outputs(3067) <= b;
    layer4_outputs(3068) <= b and not a;
    layer4_outputs(3069) <= not b;
    layer4_outputs(3070) <= b and not a;
    layer4_outputs(3071) <= not b or a;
    layer4_outputs(3072) <= not b or a;
    layer4_outputs(3073) <= a and not b;
    layer4_outputs(3074) <= a xor b;
    layer4_outputs(3075) <= 1'b0;
    layer4_outputs(3076) <= a;
    layer4_outputs(3077) <= not a;
    layer4_outputs(3078) <= not b;
    layer4_outputs(3079) <= a and not b;
    layer4_outputs(3080) <= a;
    layer4_outputs(3081) <= a and b;
    layer4_outputs(3082) <= not (a or b);
    layer4_outputs(3083) <= 1'b0;
    layer4_outputs(3084) <= a and not b;
    layer4_outputs(3085) <= not (a and b);
    layer4_outputs(3086) <= not a or b;
    layer4_outputs(3087) <= not a or b;
    layer4_outputs(3088) <= not (a or b);
    layer4_outputs(3089) <= b;
    layer4_outputs(3090) <= not (a xor b);
    layer4_outputs(3091) <= a;
    layer4_outputs(3092) <= b and not a;
    layer4_outputs(3093) <= 1'b0;
    layer4_outputs(3094) <= not (a xor b);
    layer4_outputs(3095) <= a and not b;
    layer4_outputs(3096) <= not (a and b);
    layer4_outputs(3097) <= not b;
    layer4_outputs(3098) <= a;
    layer4_outputs(3099) <= a or b;
    layer4_outputs(3100) <= a and b;
    layer4_outputs(3101) <= not b;
    layer4_outputs(3102) <= not (a and b);
    layer4_outputs(3103) <= not b or a;
    layer4_outputs(3104) <= a and b;
    layer4_outputs(3105) <= b;
    layer4_outputs(3106) <= b and not a;
    layer4_outputs(3107) <= b;
    layer4_outputs(3108) <= not a;
    layer4_outputs(3109) <= not (a and b);
    layer4_outputs(3110) <= a xor b;
    layer4_outputs(3111) <= b;
    layer4_outputs(3112) <= b and not a;
    layer4_outputs(3113) <= not (a and b);
    layer4_outputs(3114) <= not (a or b);
    layer4_outputs(3115) <= not a;
    layer4_outputs(3116) <= b and not a;
    layer4_outputs(3117) <= a;
    layer4_outputs(3118) <= 1'b1;
    layer4_outputs(3119) <= not b;
    layer4_outputs(3120) <= not b;
    layer4_outputs(3121) <= 1'b1;
    layer4_outputs(3122) <= b and not a;
    layer4_outputs(3123) <= b;
    layer4_outputs(3124) <= b and not a;
    layer4_outputs(3125) <= b;
    layer4_outputs(3126) <= a or b;
    layer4_outputs(3127) <= b and not a;
    layer4_outputs(3128) <= a and not b;
    layer4_outputs(3129) <= a or b;
    layer4_outputs(3130) <= not a;
    layer4_outputs(3131) <= not a;
    layer4_outputs(3132) <= not a or b;
    layer4_outputs(3133) <= not b;
    layer4_outputs(3134) <= not a or b;
    layer4_outputs(3135) <= not (a xor b);
    layer4_outputs(3136) <= not a;
    layer4_outputs(3137) <= 1'b0;
    layer4_outputs(3138) <= 1'b1;
    layer4_outputs(3139) <= not a;
    layer4_outputs(3140) <= a xor b;
    layer4_outputs(3141) <= a and not b;
    layer4_outputs(3142) <= a or b;
    layer4_outputs(3143) <= not a;
    layer4_outputs(3144) <= not a or b;
    layer4_outputs(3145) <= b and not a;
    layer4_outputs(3146) <= b;
    layer4_outputs(3147) <= not b or a;
    layer4_outputs(3148) <= not (a or b);
    layer4_outputs(3149) <= a and b;
    layer4_outputs(3150) <= not b;
    layer4_outputs(3151) <= a and b;
    layer4_outputs(3152) <= 1'b0;
    layer4_outputs(3153) <= a and b;
    layer4_outputs(3154) <= not b;
    layer4_outputs(3155) <= a and b;
    layer4_outputs(3156) <= not b;
    layer4_outputs(3157) <= b and not a;
    layer4_outputs(3158) <= a and b;
    layer4_outputs(3159) <= a and not b;
    layer4_outputs(3160) <= a or b;
    layer4_outputs(3161) <= a or b;
    layer4_outputs(3162) <= 1'b0;
    layer4_outputs(3163) <= b and not a;
    layer4_outputs(3164) <= a;
    layer4_outputs(3165) <= not a or b;
    layer4_outputs(3166) <= not a or b;
    layer4_outputs(3167) <= a or b;
    layer4_outputs(3168) <= not b;
    layer4_outputs(3169) <= a and not b;
    layer4_outputs(3170) <= not (a or b);
    layer4_outputs(3171) <= not (a or b);
    layer4_outputs(3172) <= not (a or b);
    layer4_outputs(3173) <= 1'b0;
    layer4_outputs(3174) <= b;
    layer4_outputs(3175) <= b;
    layer4_outputs(3176) <= 1'b0;
    layer4_outputs(3177) <= not a;
    layer4_outputs(3178) <= not a or b;
    layer4_outputs(3179) <= a;
    layer4_outputs(3180) <= a and b;
    layer4_outputs(3181) <= a or b;
    layer4_outputs(3182) <= b;
    layer4_outputs(3183) <= not (a xor b);
    layer4_outputs(3184) <= not a or b;
    layer4_outputs(3185) <= a and b;
    layer4_outputs(3186) <= not (a or b);
    layer4_outputs(3187) <= a;
    layer4_outputs(3188) <= not b or a;
    layer4_outputs(3189) <= not a or b;
    layer4_outputs(3190) <= a xor b;
    layer4_outputs(3191) <= not (a and b);
    layer4_outputs(3192) <= a and b;
    layer4_outputs(3193) <= a;
    layer4_outputs(3194) <= 1'b0;
    layer4_outputs(3195) <= not b or a;
    layer4_outputs(3196) <= a or b;
    layer4_outputs(3197) <= 1'b0;
    layer4_outputs(3198) <= a;
    layer4_outputs(3199) <= b;
    layer4_outputs(3200) <= not (a and b);
    layer4_outputs(3201) <= not a;
    layer4_outputs(3202) <= a and b;
    layer4_outputs(3203) <= not (a and b);
    layer4_outputs(3204) <= a or b;
    layer4_outputs(3205) <= not b;
    layer4_outputs(3206) <= not (a or b);
    layer4_outputs(3207) <= not (a or b);
    layer4_outputs(3208) <= not b;
    layer4_outputs(3209) <= 1'b0;
    layer4_outputs(3210) <= not b or a;
    layer4_outputs(3211) <= a or b;
    layer4_outputs(3212) <= not (a xor b);
    layer4_outputs(3213) <= 1'b0;
    layer4_outputs(3214) <= 1'b0;
    layer4_outputs(3215) <= a or b;
    layer4_outputs(3216) <= a and b;
    layer4_outputs(3217) <= not b or a;
    layer4_outputs(3218) <= a and not b;
    layer4_outputs(3219) <= not b;
    layer4_outputs(3220) <= not (a and b);
    layer4_outputs(3221) <= not (a or b);
    layer4_outputs(3222) <= not a;
    layer4_outputs(3223) <= a and not b;
    layer4_outputs(3224) <= not a or b;
    layer4_outputs(3225) <= not (a xor b);
    layer4_outputs(3226) <= 1'b1;
    layer4_outputs(3227) <= 1'b1;
    layer4_outputs(3228) <= a xor b;
    layer4_outputs(3229) <= not (a xor b);
    layer4_outputs(3230) <= 1'b1;
    layer4_outputs(3231) <= not a;
    layer4_outputs(3232) <= not (a and b);
    layer4_outputs(3233) <= a;
    layer4_outputs(3234) <= a or b;
    layer4_outputs(3235) <= a and b;
    layer4_outputs(3236) <= a and not b;
    layer4_outputs(3237) <= b;
    layer4_outputs(3238) <= 1'b1;
    layer4_outputs(3239) <= b and not a;
    layer4_outputs(3240) <= a or b;
    layer4_outputs(3241) <= not (a xor b);
    layer4_outputs(3242) <= b;
    layer4_outputs(3243) <= a and b;
    layer4_outputs(3244) <= not a or b;
    layer4_outputs(3245) <= a and not b;
    layer4_outputs(3246) <= a and b;
    layer4_outputs(3247) <= not (a and b);
    layer4_outputs(3248) <= a;
    layer4_outputs(3249) <= b and not a;
    layer4_outputs(3250) <= 1'b0;
    layer4_outputs(3251) <= a;
    layer4_outputs(3252) <= a or b;
    layer4_outputs(3253) <= not (a and b);
    layer4_outputs(3254) <= not a or b;
    layer4_outputs(3255) <= not b or a;
    layer4_outputs(3256) <= not (a and b);
    layer4_outputs(3257) <= not a;
    layer4_outputs(3258) <= not b or a;
    layer4_outputs(3259) <= not b;
    layer4_outputs(3260) <= b;
    layer4_outputs(3261) <= not a;
    layer4_outputs(3262) <= not b or a;
    layer4_outputs(3263) <= 1'b0;
    layer4_outputs(3264) <= not b;
    layer4_outputs(3265) <= b;
    layer4_outputs(3266) <= not a;
    layer4_outputs(3267) <= not a or b;
    layer4_outputs(3268) <= b;
    layer4_outputs(3269) <= not a;
    layer4_outputs(3270) <= not b;
    layer4_outputs(3271) <= not b or a;
    layer4_outputs(3272) <= not a or b;
    layer4_outputs(3273) <= a or b;
    layer4_outputs(3274) <= not b;
    layer4_outputs(3275) <= a or b;
    layer4_outputs(3276) <= a and b;
    layer4_outputs(3277) <= b;
    layer4_outputs(3278) <= a;
    layer4_outputs(3279) <= b;
    layer4_outputs(3280) <= not b;
    layer4_outputs(3281) <= a and b;
    layer4_outputs(3282) <= not b;
    layer4_outputs(3283) <= 1'b0;
    layer4_outputs(3284) <= not a or b;
    layer4_outputs(3285) <= a and not b;
    layer4_outputs(3286) <= not (a or b);
    layer4_outputs(3287) <= not a;
    layer4_outputs(3288) <= a or b;
    layer4_outputs(3289) <= a xor b;
    layer4_outputs(3290) <= b;
    layer4_outputs(3291) <= a;
    layer4_outputs(3292) <= not (a or b);
    layer4_outputs(3293) <= 1'b1;
    layer4_outputs(3294) <= a;
    layer4_outputs(3295) <= 1'b0;
    layer4_outputs(3296) <= not (a or b);
    layer4_outputs(3297) <= a and not b;
    layer4_outputs(3298) <= not (a and b);
    layer4_outputs(3299) <= not a;
    layer4_outputs(3300) <= not a or b;
    layer4_outputs(3301) <= not (a and b);
    layer4_outputs(3302) <= a and b;
    layer4_outputs(3303) <= not b or a;
    layer4_outputs(3304) <= b and not a;
    layer4_outputs(3305) <= not b or a;
    layer4_outputs(3306) <= a and b;
    layer4_outputs(3307) <= a;
    layer4_outputs(3308) <= 1'b0;
    layer4_outputs(3309) <= 1'b1;
    layer4_outputs(3310) <= not a;
    layer4_outputs(3311) <= not b;
    layer4_outputs(3312) <= not (a and b);
    layer4_outputs(3313) <= a xor b;
    layer4_outputs(3314) <= not b;
    layer4_outputs(3315) <= not a or b;
    layer4_outputs(3316) <= not b or a;
    layer4_outputs(3317) <= a and b;
    layer4_outputs(3318) <= not (a or b);
    layer4_outputs(3319) <= b;
    layer4_outputs(3320) <= b and not a;
    layer4_outputs(3321) <= not a or b;
    layer4_outputs(3322) <= a and not b;
    layer4_outputs(3323) <= a and not b;
    layer4_outputs(3324) <= not (a or b);
    layer4_outputs(3325) <= not b;
    layer4_outputs(3326) <= not (a and b);
    layer4_outputs(3327) <= not b or a;
    layer4_outputs(3328) <= not b;
    layer4_outputs(3329) <= a or b;
    layer4_outputs(3330) <= a or b;
    layer4_outputs(3331) <= a or b;
    layer4_outputs(3332) <= b;
    layer4_outputs(3333) <= not b or a;
    layer4_outputs(3334) <= 1'b1;
    layer4_outputs(3335) <= a and b;
    layer4_outputs(3336) <= not b;
    layer4_outputs(3337) <= not a or b;
    layer4_outputs(3338) <= b;
    layer4_outputs(3339) <= b and not a;
    layer4_outputs(3340) <= b and not a;
    layer4_outputs(3341) <= not b;
    layer4_outputs(3342) <= 1'b0;
    layer4_outputs(3343) <= a or b;
    layer4_outputs(3344) <= not b or a;
    layer4_outputs(3345) <= not a;
    layer4_outputs(3346) <= a xor b;
    layer4_outputs(3347) <= a or b;
    layer4_outputs(3348) <= not b or a;
    layer4_outputs(3349) <= a;
    layer4_outputs(3350) <= 1'b1;
    layer4_outputs(3351) <= a xor b;
    layer4_outputs(3352) <= a;
    layer4_outputs(3353) <= 1'b1;
    layer4_outputs(3354) <= b;
    layer4_outputs(3355) <= not b;
    layer4_outputs(3356) <= not a or b;
    layer4_outputs(3357) <= a or b;
    layer4_outputs(3358) <= b;
    layer4_outputs(3359) <= b and not a;
    layer4_outputs(3360) <= a and b;
    layer4_outputs(3361) <= not (a xor b);
    layer4_outputs(3362) <= a or b;
    layer4_outputs(3363) <= a or b;
    layer4_outputs(3364) <= a and b;
    layer4_outputs(3365) <= b and not a;
    layer4_outputs(3366) <= not (a or b);
    layer4_outputs(3367) <= a and not b;
    layer4_outputs(3368) <= not a or b;
    layer4_outputs(3369) <= b;
    layer4_outputs(3370) <= 1'b1;
    layer4_outputs(3371) <= b;
    layer4_outputs(3372) <= a and not b;
    layer4_outputs(3373) <= 1'b0;
    layer4_outputs(3374) <= not a;
    layer4_outputs(3375) <= a and not b;
    layer4_outputs(3376) <= a and b;
    layer4_outputs(3377) <= a;
    layer4_outputs(3378) <= not b;
    layer4_outputs(3379) <= a and b;
    layer4_outputs(3380) <= b;
    layer4_outputs(3381) <= 1'b1;
    layer4_outputs(3382) <= 1'b1;
    layer4_outputs(3383) <= 1'b1;
    layer4_outputs(3384) <= b;
    layer4_outputs(3385) <= not (a and b);
    layer4_outputs(3386) <= b and not a;
    layer4_outputs(3387) <= a or b;
    layer4_outputs(3388) <= a or b;
    layer4_outputs(3389) <= 1'b1;
    layer4_outputs(3390) <= 1'b1;
    layer4_outputs(3391) <= b and not a;
    layer4_outputs(3392) <= a;
    layer4_outputs(3393) <= not a or b;
    layer4_outputs(3394) <= a xor b;
    layer4_outputs(3395) <= a and not b;
    layer4_outputs(3396) <= b;
    layer4_outputs(3397) <= 1'b0;
    layer4_outputs(3398) <= a xor b;
    layer4_outputs(3399) <= b;
    layer4_outputs(3400) <= 1'b0;
    layer4_outputs(3401) <= a and not b;
    layer4_outputs(3402) <= b;
    layer4_outputs(3403) <= a or b;
    layer4_outputs(3404) <= not a;
    layer4_outputs(3405) <= a;
    layer4_outputs(3406) <= a xor b;
    layer4_outputs(3407) <= b;
    layer4_outputs(3408) <= a or b;
    layer4_outputs(3409) <= a or b;
    layer4_outputs(3410) <= not (a or b);
    layer4_outputs(3411) <= not b or a;
    layer4_outputs(3412) <= not (a and b);
    layer4_outputs(3413) <= b;
    layer4_outputs(3414) <= a and b;
    layer4_outputs(3415) <= a and b;
    layer4_outputs(3416) <= not b or a;
    layer4_outputs(3417) <= not a or b;
    layer4_outputs(3418) <= a and not b;
    layer4_outputs(3419) <= a and not b;
    layer4_outputs(3420) <= not (a or b);
    layer4_outputs(3421) <= a;
    layer4_outputs(3422) <= not (a and b);
    layer4_outputs(3423) <= not a;
    layer4_outputs(3424) <= a or b;
    layer4_outputs(3425) <= b;
    layer4_outputs(3426) <= not a;
    layer4_outputs(3427) <= not a;
    layer4_outputs(3428) <= a xor b;
    layer4_outputs(3429) <= not (a or b);
    layer4_outputs(3430) <= a and not b;
    layer4_outputs(3431) <= b;
    layer4_outputs(3432) <= not b or a;
    layer4_outputs(3433) <= b;
    layer4_outputs(3434) <= not b;
    layer4_outputs(3435) <= not a;
    layer4_outputs(3436) <= not b;
    layer4_outputs(3437) <= a or b;
    layer4_outputs(3438) <= not (a and b);
    layer4_outputs(3439) <= not a;
    layer4_outputs(3440) <= not a;
    layer4_outputs(3441) <= 1'b0;
    layer4_outputs(3442) <= 1'b0;
    layer4_outputs(3443) <= a or b;
    layer4_outputs(3444) <= a or b;
    layer4_outputs(3445) <= not a or b;
    layer4_outputs(3446) <= a;
    layer4_outputs(3447) <= not b or a;
    layer4_outputs(3448) <= b and not a;
    layer4_outputs(3449) <= 1'b1;
    layer4_outputs(3450) <= not a or b;
    layer4_outputs(3451) <= not a;
    layer4_outputs(3452) <= 1'b0;
    layer4_outputs(3453) <= not b;
    layer4_outputs(3454) <= not (a xor b);
    layer4_outputs(3455) <= not a or b;
    layer4_outputs(3456) <= not (a and b);
    layer4_outputs(3457) <= a;
    layer4_outputs(3458) <= 1'b1;
    layer4_outputs(3459) <= a xor b;
    layer4_outputs(3460) <= b;
    layer4_outputs(3461) <= a;
    layer4_outputs(3462) <= b and not a;
    layer4_outputs(3463) <= 1'b1;
    layer4_outputs(3464) <= 1'b0;
    layer4_outputs(3465) <= not (a and b);
    layer4_outputs(3466) <= a;
    layer4_outputs(3467) <= not a or b;
    layer4_outputs(3468) <= a and b;
    layer4_outputs(3469) <= not (a xor b);
    layer4_outputs(3470) <= not a;
    layer4_outputs(3471) <= not b;
    layer4_outputs(3472) <= not b or a;
    layer4_outputs(3473) <= b;
    layer4_outputs(3474) <= a xor b;
    layer4_outputs(3475) <= not a or b;
    layer4_outputs(3476) <= not a or b;
    layer4_outputs(3477) <= not (a and b);
    layer4_outputs(3478) <= a or b;
    layer4_outputs(3479) <= a and not b;
    layer4_outputs(3480) <= not b;
    layer4_outputs(3481) <= not a or b;
    layer4_outputs(3482) <= a;
    layer4_outputs(3483) <= a and not b;
    layer4_outputs(3484) <= a and not b;
    layer4_outputs(3485) <= not (a xor b);
    layer4_outputs(3486) <= a and b;
    layer4_outputs(3487) <= not a or b;
    layer4_outputs(3488) <= not (a and b);
    layer4_outputs(3489) <= a and not b;
    layer4_outputs(3490) <= not b;
    layer4_outputs(3491) <= not (a or b);
    layer4_outputs(3492) <= a and not b;
    layer4_outputs(3493) <= not a;
    layer4_outputs(3494) <= a and b;
    layer4_outputs(3495) <= b;
    layer4_outputs(3496) <= not b or a;
    layer4_outputs(3497) <= not b or a;
    layer4_outputs(3498) <= b and not a;
    layer4_outputs(3499) <= not (a or b);
    layer4_outputs(3500) <= not a or b;
    layer4_outputs(3501) <= not (a xor b);
    layer4_outputs(3502) <= a or b;
    layer4_outputs(3503) <= not b or a;
    layer4_outputs(3504) <= a and not b;
    layer4_outputs(3505) <= not a or b;
    layer4_outputs(3506) <= a and b;
    layer4_outputs(3507) <= not b or a;
    layer4_outputs(3508) <= 1'b1;
    layer4_outputs(3509) <= not a or b;
    layer4_outputs(3510) <= not (a xor b);
    layer4_outputs(3511) <= not a or b;
    layer4_outputs(3512) <= not a or b;
    layer4_outputs(3513) <= not b;
    layer4_outputs(3514) <= not a or b;
    layer4_outputs(3515) <= a or b;
    layer4_outputs(3516) <= b;
    layer4_outputs(3517) <= a and not b;
    layer4_outputs(3518) <= not (a or b);
    layer4_outputs(3519) <= not (a or b);
    layer4_outputs(3520) <= not a;
    layer4_outputs(3521) <= a;
    layer4_outputs(3522) <= a;
    layer4_outputs(3523) <= not a;
    layer4_outputs(3524) <= 1'b1;
    layer4_outputs(3525) <= a or b;
    layer4_outputs(3526) <= a xor b;
    layer4_outputs(3527) <= a and b;
    layer4_outputs(3528) <= a and not b;
    layer4_outputs(3529) <= a and not b;
    layer4_outputs(3530) <= not b;
    layer4_outputs(3531) <= not a or b;
    layer4_outputs(3532) <= b and not a;
    layer4_outputs(3533) <= b and not a;
    layer4_outputs(3534) <= not b or a;
    layer4_outputs(3535) <= not (a and b);
    layer4_outputs(3536) <= not b or a;
    layer4_outputs(3537) <= a and b;
    layer4_outputs(3538) <= not (a and b);
    layer4_outputs(3539) <= b and not a;
    layer4_outputs(3540) <= b;
    layer4_outputs(3541) <= b;
    layer4_outputs(3542) <= not b or a;
    layer4_outputs(3543) <= not b;
    layer4_outputs(3544) <= a;
    layer4_outputs(3545) <= not a;
    layer4_outputs(3546) <= not (a and b);
    layer4_outputs(3547) <= not b;
    layer4_outputs(3548) <= not b or a;
    layer4_outputs(3549) <= not (a or b);
    layer4_outputs(3550) <= 1'b0;
    layer4_outputs(3551) <= a and not b;
    layer4_outputs(3552) <= 1'b1;
    layer4_outputs(3553) <= a;
    layer4_outputs(3554) <= not (a and b);
    layer4_outputs(3555) <= not a or b;
    layer4_outputs(3556) <= 1'b0;
    layer4_outputs(3557) <= not a;
    layer4_outputs(3558) <= not b or a;
    layer4_outputs(3559) <= a and b;
    layer4_outputs(3560) <= not a;
    layer4_outputs(3561) <= 1'b1;
    layer4_outputs(3562) <= a and b;
    layer4_outputs(3563) <= a;
    layer4_outputs(3564) <= not (a and b);
    layer4_outputs(3565) <= 1'b0;
    layer4_outputs(3566) <= not b;
    layer4_outputs(3567) <= not a;
    layer4_outputs(3568) <= not a;
    layer4_outputs(3569) <= a and b;
    layer4_outputs(3570) <= a;
    layer4_outputs(3571) <= a or b;
    layer4_outputs(3572) <= not (a or b);
    layer4_outputs(3573) <= 1'b1;
    layer4_outputs(3574) <= a;
    layer4_outputs(3575) <= not (a or b);
    layer4_outputs(3576) <= a and not b;
    layer4_outputs(3577) <= not a;
    layer4_outputs(3578) <= a and b;
    layer4_outputs(3579) <= a;
    layer4_outputs(3580) <= a or b;
    layer4_outputs(3581) <= not a;
    layer4_outputs(3582) <= b;
    layer4_outputs(3583) <= not (a xor b);
    layer4_outputs(3584) <= not a or b;
    layer4_outputs(3585) <= not b;
    layer4_outputs(3586) <= a and b;
    layer4_outputs(3587) <= 1'b1;
    layer4_outputs(3588) <= not a;
    layer4_outputs(3589) <= not b or a;
    layer4_outputs(3590) <= not b;
    layer4_outputs(3591) <= 1'b1;
    layer4_outputs(3592) <= a or b;
    layer4_outputs(3593) <= a and b;
    layer4_outputs(3594) <= not b;
    layer4_outputs(3595) <= not a or b;
    layer4_outputs(3596) <= a and b;
    layer4_outputs(3597) <= not b;
    layer4_outputs(3598) <= not (a or b);
    layer4_outputs(3599) <= b and not a;
    layer4_outputs(3600) <= not a or b;
    layer4_outputs(3601) <= a and not b;
    layer4_outputs(3602) <= not a;
    layer4_outputs(3603) <= not a;
    layer4_outputs(3604) <= b and not a;
    layer4_outputs(3605) <= not (a or b);
    layer4_outputs(3606) <= a or b;
    layer4_outputs(3607) <= not (a and b);
    layer4_outputs(3608) <= a;
    layer4_outputs(3609) <= not (a and b);
    layer4_outputs(3610) <= b and not a;
    layer4_outputs(3611) <= a;
    layer4_outputs(3612) <= not b or a;
    layer4_outputs(3613) <= not a or b;
    layer4_outputs(3614) <= a and b;
    layer4_outputs(3615) <= not b;
    layer4_outputs(3616) <= not b or a;
    layer4_outputs(3617) <= not (a or b);
    layer4_outputs(3618) <= a;
    layer4_outputs(3619) <= b and not a;
    layer4_outputs(3620) <= not b;
    layer4_outputs(3621) <= not b;
    layer4_outputs(3622) <= a;
    layer4_outputs(3623) <= not a;
    layer4_outputs(3624) <= 1'b0;
    layer4_outputs(3625) <= not (a or b);
    layer4_outputs(3626) <= not b;
    layer4_outputs(3627) <= b;
    layer4_outputs(3628) <= a or b;
    layer4_outputs(3629) <= not b;
    layer4_outputs(3630) <= not (a xor b);
    layer4_outputs(3631) <= not (a or b);
    layer4_outputs(3632) <= not a or b;
    layer4_outputs(3633) <= a and not b;
    layer4_outputs(3634) <= b;
    layer4_outputs(3635) <= b;
    layer4_outputs(3636) <= a and not b;
    layer4_outputs(3637) <= a and b;
    layer4_outputs(3638) <= a or b;
    layer4_outputs(3639) <= not (a or b);
    layer4_outputs(3640) <= not a;
    layer4_outputs(3641) <= not b;
    layer4_outputs(3642) <= a;
    layer4_outputs(3643) <= b and not a;
    layer4_outputs(3644) <= not (a and b);
    layer4_outputs(3645) <= not b or a;
    layer4_outputs(3646) <= not (a and b);
    layer4_outputs(3647) <= not (a or b);
    layer4_outputs(3648) <= not (a or b);
    layer4_outputs(3649) <= a and b;
    layer4_outputs(3650) <= 1'b0;
    layer4_outputs(3651) <= not b or a;
    layer4_outputs(3652) <= not a or b;
    layer4_outputs(3653) <= not b or a;
    layer4_outputs(3654) <= not b or a;
    layer4_outputs(3655) <= not a;
    layer4_outputs(3656) <= not (a or b);
    layer4_outputs(3657) <= b and not a;
    layer4_outputs(3658) <= 1'b1;
    layer4_outputs(3659) <= not b;
    layer4_outputs(3660) <= a and b;
    layer4_outputs(3661) <= 1'b1;
    layer4_outputs(3662) <= a;
    layer4_outputs(3663) <= not b;
    layer4_outputs(3664) <= a and b;
    layer4_outputs(3665) <= not b or a;
    layer4_outputs(3666) <= a or b;
    layer4_outputs(3667) <= a and b;
    layer4_outputs(3668) <= not b;
    layer4_outputs(3669) <= a and b;
    layer4_outputs(3670) <= not b;
    layer4_outputs(3671) <= not (a or b);
    layer4_outputs(3672) <= not b;
    layer4_outputs(3673) <= not a;
    layer4_outputs(3674) <= a and b;
    layer4_outputs(3675) <= not (a xor b);
    layer4_outputs(3676) <= not (a and b);
    layer4_outputs(3677) <= 1'b0;
    layer4_outputs(3678) <= not b;
    layer4_outputs(3679) <= a or b;
    layer4_outputs(3680) <= 1'b1;
    layer4_outputs(3681) <= 1'b1;
    layer4_outputs(3682) <= 1'b1;
    layer4_outputs(3683) <= a xor b;
    layer4_outputs(3684) <= a xor b;
    layer4_outputs(3685) <= not b;
    layer4_outputs(3686) <= not (a and b);
    layer4_outputs(3687) <= a and not b;
    layer4_outputs(3688) <= not a;
    layer4_outputs(3689) <= not b;
    layer4_outputs(3690) <= not (a or b);
    layer4_outputs(3691) <= not b;
    layer4_outputs(3692) <= a and not b;
    layer4_outputs(3693) <= not a or b;
    layer4_outputs(3694) <= not b or a;
    layer4_outputs(3695) <= not (a and b);
    layer4_outputs(3696) <= not b or a;
    layer4_outputs(3697) <= a and not b;
    layer4_outputs(3698) <= not a or b;
    layer4_outputs(3699) <= a and b;
    layer4_outputs(3700) <= not a or b;
    layer4_outputs(3701) <= not a or b;
    layer4_outputs(3702) <= not a or b;
    layer4_outputs(3703) <= not (a or b);
    layer4_outputs(3704) <= 1'b0;
    layer4_outputs(3705) <= not a;
    layer4_outputs(3706) <= a xor b;
    layer4_outputs(3707) <= not b or a;
    layer4_outputs(3708) <= a and not b;
    layer4_outputs(3709) <= b and not a;
    layer4_outputs(3710) <= b;
    layer4_outputs(3711) <= 1'b0;
    layer4_outputs(3712) <= a;
    layer4_outputs(3713) <= b and not a;
    layer4_outputs(3714) <= not a;
    layer4_outputs(3715) <= not (a xor b);
    layer4_outputs(3716) <= 1'b1;
    layer4_outputs(3717) <= not (a and b);
    layer4_outputs(3718) <= not (a or b);
    layer4_outputs(3719) <= a and b;
    layer4_outputs(3720) <= 1'b1;
    layer4_outputs(3721) <= 1'b1;
    layer4_outputs(3722) <= 1'b0;
    layer4_outputs(3723) <= b;
    layer4_outputs(3724) <= a;
    layer4_outputs(3725) <= 1'b0;
    layer4_outputs(3726) <= b and not a;
    layer4_outputs(3727) <= not (a and b);
    layer4_outputs(3728) <= a and not b;
    layer4_outputs(3729) <= 1'b1;
    layer4_outputs(3730) <= a;
    layer4_outputs(3731) <= not b or a;
    layer4_outputs(3732) <= not b;
    layer4_outputs(3733) <= b and not a;
    layer4_outputs(3734) <= not a or b;
    layer4_outputs(3735) <= a or b;
    layer4_outputs(3736) <= not b;
    layer4_outputs(3737) <= a xor b;
    layer4_outputs(3738) <= a;
    layer4_outputs(3739) <= a and b;
    layer4_outputs(3740) <= not b;
    layer4_outputs(3741) <= not (a and b);
    layer4_outputs(3742) <= not b or a;
    layer4_outputs(3743) <= a and not b;
    layer4_outputs(3744) <= not b;
    layer4_outputs(3745) <= not (a and b);
    layer4_outputs(3746) <= not (a or b);
    layer4_outputs(3747) <= not a;
    layer4_outputs(3748) <= not (a and b);
    layer4_outputs(3749) <= b and not a;
    layer4_outputs(3750) <= not b or a;
    layer4_outputs(3751) <= a and b;
    layer4_outputs(3752) <= not (a or b);
    layer4_outputs(3753) <= a and b;
    layer4_outputs(3754) <= not (a or b);
    layer4_outputs(3755) <= a;
    layer4_outputs(3756) <= not b;
    layer4_outputs(3757) <= a and b;
    layer4_outputs(3758) <= a;
    layer4_outputs(3759) <= a;
    layer4_outputs(3760) <= a and not b;
    layer4_outputs(3761) <= a and not b;
    layer4_outputs(3762) <= b and not a;
    layer4_outputs(3763) <= a and not b;
    layer4_outputs(3764) <= 1'b1;
    layer4_outputs(3765) <= b;
    layer4_outputs(3766) <= a and b;
    layer4_outputs(3767) <= 1'b1;
    layer4_outputs(3768) <= a and b;
    layer4_outputs(3769) <= a;
    layer4_outputs(3770) <= a;
    layer4_outputs(3771) <= not a or b;
    layer4_outputs(3772) <= not a or b;
    layer4_outputs(3773) <= 1'b0;
    layer4_outputs(3774) <= 1'b0;
    layer4_outputs(3775) <= b and not a;
    layer4_outputs(3776) <= a or b;
    layer4_outputs(3777) <= b;
    layer4_outputs(3778) <= a xor b;
    layer4_outputs(3779) <= a and b;
    layer4_outputs(3780) <= 1'b0;
    layer4_outputs(3781) <= b;
    layer4_outputs(3782) <= b;
    layer4_outputs(3783) <= not a or b;
    layer4_outputs(3784) <= not b;
    layer4_outputs(3785) <= not a;
    layer4_outputs(3786) <= a;
    layer4_outputs(3787) <= not a or b;
    layer4_outputs(3788) <= not (a or b);
    layer4_outputs(3789) <= a and not b;
    layer4_outputs(3790) <= a and b;
    layer4_outputs(3791) <= a;
    layer4_outputs(3792) <= not b;
    layer4_outputs(3793) <= a and b;
    layer4_outputs(3794) <= not a;
    layer4_outputs(3795) <= b and not a;
    layer4_outputs(3796) <= a and b;
    layer4_outputs(3797) <= a and b;
    layer4_outputs(3798) <= not (a or b);
    layer4_outputs(3799) <= a and not b;
    layer4_outputs(3800) <= not (a xor b);
    layer4_outputs(3801) <= a and b;
    layer4_outputs(3802) <= 1'b0;
    layer4_outputs(3803) <= a;
    layer4_outputs(3804) <= a xor b;
    layer4_outputs(3805) <= a and not b;
    layer4_outputs(3806) <= not a;
    layer4_outputs(3807) <= not a;
    layer4_outputs(3808) <= not b;
    layer4_outputs(3809) <= not b or a;
    layer4_outputs(3810) <= 1'b0;
    layer4_outputs(3811) <= not b;
    layer4_outputs(3812) <= not (a or b);
    layer4_outputs(3813) <= a or b;
    layer4_outputs(3814) <= a;
    layer4_outputs(3815) <= not (a xor b);
    layer4_outputs(3816) <= a and b;
    layer4_outputs(3817) <= not b;
    layer4_outputs(3818) <= a;
    layer4_outputs(3819) <= b and not a;
    layer4_outputs(3820) <= a or b;
    layer4_outputs(3821) <= not b;
    layer4_outputs(3822) <= not (a and b);
    layer4_outputs(3823) <= not (a and b);
    layer4_outputs(3824) <= a or b;
    layer4_outputs(3825) <= not a;
    layer4_outputs(3826) <= b and not a;
    layer4_outputs(3827) <= not (a and b);
    layer4_outputs(3828) <= not b or a;
    layer4_outputs(3829) <= b and not a;
    layer4_outputs(3830) <= not a or b;
    layer4_outputs(3831) <= b and not a;
    layer4_outputs(3832) <= not (a xor b);
    layer4_outputs(3833) <= not a;
    layer4_outputs(3834) <= not a or b;
    layer4_outputs(3835) <= not (a and b);
    layer4_outputs(3836) <= not a or b;
    layer4_outputs(3837) <= not (a and b);
    layer4_outputs(3838) <= b and not a;
    layer4_outputs(3839) <= not (a or b);
    layer4_outputs(3840) <= b;
    layer4_outputs(3841) <= 1'b0;
    layer4_outputs(3842) <= not (a or b);
    layer4_outputs(3843) <= not b;
    layer4_outputs(3844) <= b and not a;
    layer4_outputs(3845) <= not b;
    layer4_outputs(3846) <= not a;
    layer4_outputs(3847) <= a and not b;
    layer4_outputs(3848) <= not b;
    layer4_outputs(3849) <= 1'b0;
    layer4_outputs(3850) <= a and b;
    layer4_outputs(3851) <= not b or a;
    layer4_outputs(3852) <= 1'b0;
    layer4_outputs(3853) <= a;
    layer4_outputs(3854) <= b and not a;
    layer4_outputs(3855) <= a and b;
    layer4_outputs(3856) <= not a or b;
    layer4_outputs(3857) <= a and not b;
    layer4_outputs(3858) <= a or b;
    layer4_outputs(3859) <= b and not a;
    layer4_outputs(3860) <= not (a and b);
    layer4_outputs(3861) <= a or b;
    layer4_outputs(3862) <= not b or a;
    layer4_outputs(3863) <= not (a or b);
    layer4_outputs(3864) <= a and not b;
    layer4_outputs(3865) <= b;
    layer4_outputs(3866) <= 1'b1;
    layer4_outputs(3867) <= not (a or b);
    layer4_outputs(3868) <= not (a xor b);
    layer4_outputs(3869) <= a;
    layer4_outputs(3870) <= b and not a;
    layer4_outputs(3871) <= 1'b0;
    layer4_outputs(3872) <= b;
    layer4_outputs(3873) <= 1'b0;
    layer4_outputs(3874) <= not a;
    layer4_outputs(3875) <= not (a or b);
    layer4_outputs(3876) <= not b;
    layer4_outputs(3877) <= a and not b;
    layer4_outputs(3878) <= not (a or b);
    layer4_outputs(3879) <= a and b;
    layer4_outputs(3880) <= 1'b1;
    layer4_outputs(3881) <= a xor b;
    layer4_outputs(3882) <= b and not a;
    layer4_outputs(3883) <= not (a xor b);
    layer4_outputs(3884) <= b and not a;
    layer4_outputs(3885) <= not (a or b);
    layer4_outputs(3886) <= a;
    layer4_outputs(3887) <= not a or b;
    layer4_outputs(3888) <= a;
    layer4_outputs(3889) <= not a;
    layer4_outputs(3890) <= not b or a;
    layer4_outputs(3891) <= a and not b;
    layer4_outputs(3892) <= b and not a;
    layer4_outputs(3893) <= 1'b1;
    layer4_outputs(3894) <= b;
    layer4_outputs(3895) <= not b or a;
    layer4_outputs(3896) <= a;
    layer4_outputs(3897) <= b;
    layer4_outputs(3898) <= not b;
    layer4_outputs(3899) <= b and not a;
    layer4_outputs(3900) <= a;
    layer4_outputs(3901) <= not b;
    layer4_outputs(3902) <= 1'b1;
    layer4_outputs(3903) <= not (a or b);
    layer4_outputs(3904) <= 1'b0;
    layer4_outputs(3905) <= 1'b1;
    layer4_outputs(3906) <= not a or b;
    layer4_outputs(3907) <= 1'b1;
    layer4_outputs(3908) <= b and not a;
    layer4_outputs(3909) <= b;
    layer4_outputs(3910) <= not a;
    layer4_outputs(3911) <= not b;
    layer4_outputs(3912) <= 1'b0;
    layer4_outputs(3913) <= a and not b;
    layer4_outputs(3914) <= a xor b;
    layer4_outputs(3915) <= a;
    layer4_outputs(3916) <= b and not a;
    layer4_outputs(3917) <= not (a and b);
    layer4_outputs(3918) <= not (a or b);
    layer4_outputs(3919) <= b and not a;
    layer4_outputs(3920) <= not b or a;
    layer4_outputs(3921) <= 1'b1;
    layer4_outputs(3922) <= b and not a;
    layer4_outputs(3923) <= a or b;
    layer4_outputs(3924) <= not b or a;
    layer4_outputs(3925) <= 1'b1;
    layer4_outputs(3926) <= a and b;
    layer4_outputs(3927) <= a;
    layer4_outputs(3928) <= a or b;
    layer4_outputs(3929) <= a;
    layer4_outputs(3930) <= 1'b0;
    layer4_outputs(3931) <= not b;
    layer4_outputs(3932) <= b;
    layer4_outputs(3933) <= b;
    layer4_outputs(3934) <= not (a xor b);
    layer4_outputs(3935) <= not (a and b);
    layer4_outputs(3936) <= not b or a;
    layer4_outputs(3937) <= not (a and b);
    layer4_outputs(3938) <= 1'b0;
    layer4_outputs(3939) <= a xor b;
    layer4_outputs(3940) <= not a or b;
    layer4_outputs(3941) <= not (a xor b);
    layer4_outputs(3942) <= not (a and b);
    layer4_outputs(3943) <= 1'b1;
    layer4_outputs(3944) <= not (a or b);
    layer4_outputs(3945) <= 1'b0;
    layer4_outputs(3946) <= not (a or b);
    layer4_outputs(3947) <= 1'b0;
    layer4_outputs(3948) <= a or b;
    layer4_outputs(3949) <= not b;
    layer4_outputs(3950) <= b;
    layer4_outputs(3951) <= a or b;
    layer4_outputs(3952) <= b and not a;
    layer4_outputs(3953) <= a and not b;
    layer4_outputs(3954) <= not a or b;
    layer4_outputs(3955) <= not a;
    layer4_outputs(3956) <= b and not a;
    layer4_outputs(3957) <= a;
    layer4_outputs(3958) <= not (a or b);
    layer4_outputs(3959) <= a;
    layer4_outputs(3960) <= b and not a;
    layer4_outputs(3961) <= a or b;
    layer4_outputs(3962) <= b and not a;
    layer4_outputs(3963) <= not b or a;
    layer4_outputs(3964) <= not (a and b);
    layer4_outputs(3965) <= a or b;
    layer4_outputs(3966) <= a or b;
    layer4_outputs(3967) <= a and not b;
    layer4_outputs(3968) <= 1'b0;
    layer4_outputs(3969) <= a and not b;
    layer4_outputs(3970) <= not (a or b);
    layer4_outputs(3971) <= not (a and b);
    layer4_outputs(3972) <= a or b;
    layer4_outputs(3973) <= b and not a;
    layer4_outputs(3974) <= a and not b;
    layer4_outputs(3975) <= not b;
    layer4_outputs(3976) <= not b;
    layer4_outputs(3977) <= not b;
    layer4_outputs(3978) <= b;
    layer4_outputs(3979) <= a and not b;
    layer4_outputs(3980) <= b;
    layer4_outputs(3981) <= b;
    layer4_outputs(3982) <= not a or b;
    layer4_outputs(3983) <= a;
    layer4_outputs(3984) <= b and not a;
    layer4_outputs(3985) <= a or b;
    layer4_outputs(3986) <= not a;
    layer4_outputs(3987) <= not (a and b);
    layer4_outputs(3988) <= not (a and b);
    layer4_outputs(3989) <= b and not a;
    layer4_outputs(3990) <= not b or a;
    layer4_outputs(3991) <= a or b;
    layer4_outputs(3992) <= a;
    layer4_outputs(3993) <= not a;
    layer4_outputs(3994) <= a;
    layer4_outputs(3995) <= b;
    layer4_outputs(3996) <= a and not b;
    layer4_outputs(3997) <= 1'b1;
    layer4_outputs(3998) <= b and not a;
    layer4_outputs(3999) <= b and not a;
    layer4_outputs(4000) <= not (a or b);
    layer4_outputs(4001) <= a;
    layer4_outputs(4002) <= a and not b;
    layer4_outputs(4003) <= a;
    layer4_outputs(4004) <= not b or a;
    layer4_outputs(4005) <= a or b;
    layer4_outputs(4006) <= not b or a;
    layer4_outputs(4007) <= not a;
    layer4_outputs(4008) <= not a;
    layer4_outputs(4009) <= b and not a;
    layer4_outputs(4010) <= 1'b1;
    layer4_outputs(4011) <= 1'b1;
    layer4_outputs(4012) <= a;
    layer4_outputs(4013) <= not a;
    layer4_outputs(4014) <= a or b;
    layer4_outputs(4015) <= not b;
    layer4_outputs(4016) <= 1'b0;
    layer4_outputs(4017) <= a;
    layer4_outputs(4018) <= a;
    layer4_outputs(4019) <= a;
    layer4_outputs(4020) <= a and b;
    layer4_outputs(4021) <= not a;
    layer4_outputs(4022) <= not (a and b);
    layer4_outputs(4023) <= 1'b1;
    layer4_outputs(4024) <= a;
    layer4_outputs(4025) <= a xor b;
    layer4_outputs(4026) <= b;
    layer4_outputs(4027) <= b;
    layer4_outputs(4028) <= a and not b;
    layer4_outputs(4029) <= 1'b0;
    layer4_outputs(4030) <= b;
    layer4_outputs(4031) <= not a;
    layer4_outputs(4032) <= a or b;
    layer4_outputs(4033) <= 1'b1;
    layer4_outputs(4034) <= b;
    layer4_outputs(4035) <= 1'b1;
    layer4_outputs(4036) <= not a or b;
    layer4_outputs(4037) <= not (a or b);
    layer4_outputs(4038) <= 1'b0;
    layer4_outputs(4039) <= a and not b;
    layer4_outputs(4040) <= 1'b0;
    layer4_outputs(4041) <= not b;
    layer4_outputs(4042) <= a;
    layer4_outputs(4043) <= 1'b1;
    layer4_outputs(4044) <= not b;
    layer4_outputs(4045) <= not b;
    layer4_outputs(4046) <= not a;
    layer4_outputs(4047) <= not (a or b);
    layer4_outputs(4048) <= not (a or b);
    layer4_outputs(4049) <= a or b;
    layer4_outputs(4050) <= a xor b;
    layer4_outputs(4051) <= a;
    layer4_outputs(4052) <= a and b;
    layer4_outputs(4053) <= not (a or b);
    layer4_outputs(4054) <= not a or b;
    layer4_outputs(4055) <= not b or a;
    layer4_outputs(4056) <= b and not a;
    layer4_outputs(4057) <= not b or a;
    layer4_outputs(4058) <= a;
    layer4_outputs(4059) <= b and not a;
    layer4_outputs(4060) <= a and not b;
    layer4_outputs(4061) <= not (a or b);
    layer4_outputs(4062) <= a or b;
    layer4_outputs(4063) <= not b or a;
    layer4_outputs(4064) <= b;
    layer4_outputs(4065) <= b;
    layer4_outputs(4066) <= a or b;
    layer4_outputs(4067) <= b;
    layer4_outputs(4068) <= a;
    layer4_outputs(4069) <= not (a and b);
    layer4_outputs(4070) <= not b or a;
    layer4_outputs(4071) <= not (a and b);
    layer4_outputs(4072) <= not b or a;
    layer4_outputs(4073) <= a and b;
    layer4_outputs(4074) <= a or b;
    layer4_outputs(4075) <= not (a or b);
    layer4_outputs(4076) <= 1'b0;
    layer4_outputs(4077) <= not (a or b);
    layer4_outputs(4078) <= not a;
    layer4_outputs(4079) <= a or b;
    layer4_outputs(4080) <= b and not a;
    layer4_outputs(4081) <= b;
    layer4_outputs(4082) <= b;
    layer4_outputs(4083) <= not a;
    layer4_outputs(4084) <= a;
    layer4_outputs(4085) <= a and not b;
    layer4_outputs(4086) <= not b or a;
    layer4_outputs(4087) <= a and not b;
    layer4_outputs(4088) <= not b;
    layer4_outputs(4089) <= not b or a;
    layer4_outputs(4090) <= 1'b1;
    layer4_outputs(4091) <= 1'b0;
    layer4_outputs(4092) <= not b;
    layer4_outputs(4093) <= not a or b;
    layer4_outputs(4094) <= b;
    layer4_outputs(4095) <= b and not a;
    layer4_outputs(4096) <= not (a or b);
    layer4_outputs(4097) <= not (a and b);
    layer4_outputs(4098) <= 1'b1;
    layer4_outputs(4099) <= a or b;
    layer4_outputs(4100) <= not b or a;
    layer4_outputs(4101) <= 1'b1;
    layer4_outputs(4102) <= 1'b0;
    layer4_outputs(4103) <= b and not a;
    layer4_outputs(4104) <= not b;
    layer4_outputs(4105) <= a;
    layer4_outputs(4106) <= not a;
    layer4_outputs(4107) <= not b;
    layer4_outputs(4108) <= b and not a;
    layer4_outputs(4109) <= not (a or b);
    layer4_outputs(4110) <= not (a or b);
    layer4_outputs(4111) <= b;
    layer4_outputs(4112) <= not b;
    layer4_outputs(4113) <= b and not a;
    layer4_outputs(4114) <= 1'b1;
    layer4_outputs(4115) <= not b or a;
    layer4_outputs(4116) <= not b;
    layer4_outputs(4117) <= not b or a;
    layer4_outputs(4118) <= a;
    layer4_outputs(4119) <= a;
    layer4_outputs(4120) <= not b;
    layer4_outputs(4121) <= a and not b;
    layer4_outputs(4122) <= not a or b;
    layer4_outputs(4123) <= not (a or b);
    layer4_outputs(4124) <= not b or a;
    layer4_outputs(4125) <= 1'b1;
    layer4_outputs(4126) <= 1'b1;
    layer4_outputs(4127) <= a and not b;
    layer4_outputs(4128) <= not a or b;
    layer4_outputs(4129) <= b and not a;
    layer4_outputs(4130) <= 1'b1;
    layer4_outputs(4131) <= a;
    layer4_outputs(4132) <= 1'b1;
    layer4_outputs(4133) <= 1'b1;
    layer4_outputs(4134) <= b;
    layer4_outputs(4135) <= b;
    layer4_outputs(4136) <= not (a xor b);
    layer4_outputs(4137) <= b;
    layer4_outputs(4138) <= 1'b1;
    layer4_outputs(4139) <= a xor b;
    layer4_outputs(4140) <= not a or b;
    layer4_outputs(4141) <= a;
    layer4_outputs(4142) <= not a;
    layer4_outputs(4143) <= a and not b;
    layer4_outputs(4144) <= a;
    layer4_outputs(4145) <= not (a or b);
    layer4_outputs(4146) <= not a or b;
    layer4_outputs(4147) <= not b or a;
    layer4_outputs(4148) <= a xor b;
    layer4_outputs(4149) <= not (a and b);
    layer4_outputs(4150) <= not b or a;
    layer4_outputs(4151) <= a or b;
    layer4_outputs(4152) <= not a;
    layer4_outputs(4153) <= not (a and b);
    layer4_outputs(4154) <= not (a and b);
    layer4_outputs(4155) <= a;
    layer4_outputs(4156) <= 1'b0;
    layer4_outputs(4157) <= 1'b1;
    layer4_outputs(4158) <= a and b;
    layer4_outputs(4159) <= a and b;
    layer4_outputs(4160) <= a and not b;
    layer4_outputs(4161) <= 1'b0;
    layer4_outputs(4162) <= a or b;
    layer4_outputs(4163) <= a and b;
    layer4_outputs(4164) <= not (a and b);
    layer4_outputs(4165) <= a and not b;
    layer4_outputs(4166) <= not (a and b);
    layer4_outputs(4167) <= not a or b;
    layer4_outputs(4168) <= a xor b;
    layer4_outputs(4169) <= 1'b0;
    layer4_outputs(4170) <= not a or b;
    layer4_outputs(4171) <= not a or b;
    layer4_outputs(4172) <= b and not a;
    layer4_outputs(4173) <= b;
    layer4_outputs(4174) <= not (a or b);
    layer4_outputs(4175) <= b;
    layer4_outputs(4176) <= not (a and b);
    layer4_outputs(4177) <= a and not b;
    layer4_outputs(4178) <= not (a or b);
    layer4_outputs(4179) <= 1'b1;
    layer4_outputs(4180) <= not a;
    layer4_outputs(4181) <= not (a or b);
    layer4_outputs(4182) <= a and b;
    layer4_outputs(4183) <= not b;
    layer4_outputs(4184) <= not b;
    layer4_outputs(4185) <= b;
    layer4_outputs(4186) <= b;
    layer4_outputs(4187) <= not b;
    layer4_outputs(4188) <= not (a xor b);
    layer4_outputs(4189) <= not b or a;
    layer4_outputs(4190) <= b;
    layer4_outputs(4191) <= not (a xor b);
    layer4_outputs(4192) <= not a;
    layer4_outputs(4193) <= not a;
    layer4_outputs(4194) <= not (a or b);
    layer4_outputs(4195) <= not b or a;
    layer4_outputs(4196) <= not a;
    layer4_outputs(4197) <= b and not a;
    layer4_outputs(4198) <= b and not a;
    layer4_outputs(4199) <= a and not b;
    layer4_outputs(4200) <= 1'b1;
    layer4_outputs(4201) <= not b;
    layer4_outputs(4202) <= 1'b1;
    layer4_outputs(4203) <= not b or a;
    layer4_outputs(4204) <= a and b;
    layer4_outputs(4205) <= 1'b1;
    layer4_outputs(4206) <= b;
    layer4_outputs(4207) <= a;
    layer4_outputs(4208) <= not a or b;
    layer4_outputs(4209) <= a and b;
    layer4_outputs(4210) <= b;
    layer4_outputs(4211) <= a and not b;
    layer4_outputs(4212) <= a and b;
    layer4_outputs(4213) <= a xor b;
    layer4_outputs(4214) <= a;
    layer4_outputs(4215) <= not (a and b);
    layer4_outputs(4216) <= a;
    layer4_outputs(4217) <= not a or b;
    layer4_outputs(4218) <= not b;
    layer4_outputs(4219) <= not (a or b);
    layer4_outputs(4220) <= not (a and b);
    layer4_outputs(4221) <= not a;
    layer4_outputs(4222) <= not a or b;
    layer4_outputs(4223) <= not b or a;
    layer4_outputs(4224) <= not (a or b);
    layer4_outputs(4225) <= a and b;
    layer4_outputs(4226) <= a and not b;
    layer4_outputs(4227) <= 1'b0;
    layer4_outputs(4228) <= b and not a;
    layer4_outputs(4229) <= not b or a;
    layer4_outputs(4230) <= a xor b;
    layer4_outputs(4231) <= 1'b0;
    layer4_outputs(4232) <= not a or b;
    layer4_outputs(4233) <= not b;
    layer4_outputs(4234) <= not b;
    layer4_outputs(4235) <= b;
    layer4_outputs(4236) <= a and b;
    layer4_outputs(4237) <= not a or b;
    layer4_outputs(4238) <= b and not a;
    layer4_outputs(4239) <= not b;
    layer4_outputs(4240) <= 1'b0;
    layer4_outputs(4241) <= not (a or b);
    layer4_outputs(4242) <= a;
    layer4_outputs(4243) <= 1'b0;
    layer4_outputs(4244) <= b;
    layer4_outputs(4245) <= 1'b1;
    layer4_outputs(4246) <= 1'b1;
    layer4_outputs(4247) <= not a or b;
    layer4_outputs(4248) <= a xor b;
    layer4_outputs(4249) <= not a or b;
    layer4_outputs(4250) <= 1'b1;
    layer4_outputs(4251) <= a;
    layer4_outputs(4252) <= a and b;
    layer4_outputs(4253) <= not a or b;
    layer4_outputs(4254) <= a and b;
    layer4_outputs(4255) <= not a;
    layer4_outputs(4256) <= a;
    layer4_outputs(4257) <= a;
    layer4_outputs(4258) <= a;
    layer4_outputs(4259) <= a or b;
    layer4_outputs(4260) <= a and b;
    layer4_outputs(4261) <= b;
    layer4_outputs(4262) <= a and b;
    layer4_outputs(4263) <= b;
    layer4_outputs(4264) <= not a;
    layer4_outputs(4265) <= 1'b1;
    layer4_outputs(4266) <= a xor b;
    layer4_outputs(4267) <= a and not b;
    layer4_outputs(4268) <= not b or a;
    layer4_outputs(4269) <= a xor b;
    layer4_outputs(4270) <= b;
    layer4_outputs(4271) <= not (a or b);
    layer4_outputs(4272) <= not a;
    layer4_outputs(4273) <= not a or b;
    layer4_outputs(4274) <= b;
    layer4_outputs(4275) <= not (a and b);
    layer4_outputs(4276) <= not b;
    layer4_outputs(4277) <= a;
    layer4_outputs(4278) <= not b or a;
    layer4_outputs(4279) <= b;
    layer4_outputs(4280) <= not (a or b);
    layer4_outputs(4281) <= not b or a;
    layer4_outputs(4282) <= a and b;
    layer4_outputs(4283) <= not a;
    layer4_outputs(4284) <= not (a or b);
    layer4_outputs(4285) <= not (a or b);
    layer4_outputs(4286) <= not a or b;
    layer4_outputs(4287) <= not a;
    layer4_outputs(4288) <= not a or b;
    layer4_outputs(4289) <= b;
    layer4_outputs(4290) <= 1'b1;
    layer4_outputs(4291) <= a xor b;
    layer4_outputs(4292) <= 1'b1;
    layer4_outputs(4293) <= not a;
    layer4_outputs(4294) <= b and not a;
    layer4_outputs(4295) <= not (a and b);
    layer4_outputs(4296) <= a and b;
    layer4_outputs(4297) <= not (a xor b);
    layer4_outputs(4298) <= not a;
    layer4_outputs(4299) <= a or b;
    layer4_outputs(4300) <= a or b;
    layer4_outputs(4301) <= a and not b;
    layer4_outputs(4302) <= 1'b1;
    layer4_outputs(4303) <= not (a or b);
    layer4_outputs(4304) <= a or b;
    layer4_outputs(4305) <= not (a or b);
    layer4_outputs(4306) <= 1'b0;
    layer4_outputs(4307) <= not (a and b);
    layer4_outputs(4308) <= b;
    layer4_outputs(4309) <= not b or a;
    layer4_outputs(4310) <= 1'b0;
    layer4_outputs(4311) <= b and not a;
    layer4_outputs(4312) <= b and not a;
    layer4_outputs(4313) <= a and b;
    layer4_outputs(4314) <= not (a xor b);
    layer4_outputs(4315) <= b;
    layer4_outputs(4316) <= 1'b0;
    layer4_outputs(4317) <= b and not a;
    layer4_outputs(4318) <= not a;
    layer4_outputs(4319) <= not (a or b);
    layer4_outputs(4320) <= a or b;
    layer4_outputs(4321) <= b;
    layer4_outputs(4322) <= a;
    layer4_outputs(4323) <= not b;
    layer4_outputs(4324) <= b and not a;
    layer4_outputs(4325) <= a and not b;
    layer4_outputs(4326) <= not a;
    layer4_outputs(4327) <= a or b;
    layer4_outputs(4328) <= 1'b0;
    layer4_outputs(4329) <= not a or b;
    layer4_outputs(4330) <= not b;
    layer4_outputs(4331) <= b;
    layer4_outputs(4332) <= a and not b;
    layer4_outputs(4333) <= b and not a;
    layer4_outputs(4334) <= not b or a;
    layer4_outputs(4335) <= not (a or b);
    layer4_outputs(4336) <= not (a or b);
    layer4_outputs(4337) <= not b;
    layer4_outputs(4338) <= a and b;
    layer4_outputs(4339) <= not (a or b);
    layer4_outputs(4340) <= b and not a;
    layer4_outputs(4341) <= not (a and b);
    layer4_outputs(4342) <= not b;
    layer4_outputs(4343) <= not (a or b);
    layer4_outputs(4344) <= a;
    layer4_outputs(4345) <= not (a and b);
    layer4_outputs(4346) <= not a or b;
    layer4_outputs(4347) <= a and b;
    layer4_outputs(4348) <= not b;
    layer4_outputs(4349) <= a xor b;
    layer4_outputs(4350) <= 1'b0;
    layer4_outputs(4351) <= not a;
    layer4_outputs(4352) <= not a or b;
    layer4_outputs(4353) <= a or b;
    layer4_outputs(4354) <= not b;
    layer4_outputs(4355) <= not (a and b);
    layer4_outputs(4356) <= not (a and b);
    layer4_outputs(4357) <= not (a xor b);
    layer4_outputs(4358) <= b;
    layer4_outputs(4359) <= a and b;
    layer4_outputs(4360) <= b and not a;
    layer4_outputs(4361) <= not a;
    layer4_outputs(4362) <= a and b;
    layer4_outputs(4363) <= a and b;
    layer4_outputs(4364) <= not a or b;
    layer4_outputs(4365) <= 1'b1;
    layer4_outputs(4366) <= 1'b1;
    layer4_outputs(4367) <= a or b;
    layer4_outputs(4368) <= not b;
    layer4_outputs(4369) <= a and not b;
    layer4_outputs(4370) <= not a;
    layer4_outputs(4371) <= not a;
    layer4_outputs(4372) <= a and not b;
    layer4_outputs(4373) <= not b;
    layer4_outputs(4374) <= not (a or b);
    layer4_outputs(4375) <= b;
    layer4_outputs(4376) <= a or b;
    layer4_outputs(4377) <= not b;
    layer4_outputs(4378) <= a and b;
    layer4_outputs(4379) <= not b or a;
    layer4_outputs(4380) <= a;
    layer4_outputs(4381) <= a or b;
    layer4_outputs(4382) <= a and b;
    layer4_outputs(4383) <= not (a and b);
    layer4_outputs(4384) <= not (a and b);
    layer4_outputs(4385) <= b and not a;
    layer4_outputs(4386) <= not (a and b);
    layer4_outputs(4387) <= not (a or b);
    layer4_outputs(4388) <= not a or b;
    layer4_outputs(4389) <= a and b;
    layer4_outputs(4390) <= not a;
    layer4_outputs(4391) <= a and b;
    layer4_outputs(4392) <= not (a xor b);
    layer4_outputs(4393) <= a or b;
    layer4_outputs(4394) <= not (a and b);
    layer4_outputs(4395) <= not (a and b);
    layer4_outputs(4396) <= b and not a;
    layer4_outputs(4397) <= 1'b1;
    layer4_outputs(4398) <= not b or a;
    layer4_outputs(4399) <= not a;
    layer4_outputs(4400) <= not (a and b);
    layer4_outputs(4401) <= a;
    layer4_outputs(4402) <= not b or a;
    layer4_outputs(4403) <= b;
    layer4_outputs(4404) <= b;
    layer4_outputs(4405) <= a xor b;
    layer4_outputs(4406) <= a and b;
    layer4_outputs(4407) <= 1'b0;
    layer4_outputs(4408) <= 1'b1;
    layer4_outputs(4409) <= not a;
    layer4_outputs(4410) <= not a;
    layer4_outputs(4411) <= not a;
    layer4_outputs(4412) <= a;
    layer4_outputs(4413) <= not (a or b);
    layer4_outputs(4414) <= b;
    layer4_outputs(4415) <= b;
    layer4_outputs(4416) <= not b;
    layer4_outputs(4417) <= not (a or b);
    layer4_outputs(4418) <= a;
    layer4_outputs(4419) <= not b or a;
    layer4_outputs(4420) <= 1'b0;
    layer4_outputs(4421) <= not a;
    layer4_outputs(4422) <= not a or b;
    layer4_outputs(4423) <= b;
    layer4_outputs(4424) <= b and not a;
    layer4_outputs(4425) <= not b;
    layer4_outputs(4426) <= a and b;
    layer4_outputs(4427) <= not b or a;
    layer4_outputs(4428) <= not (a and b);
    layer4_outputs(4429) <= 1'b1;
    layer4_outputs(4430) <= a and b;
    layer4_outputs(4431) <= a xor b;
    layer4_outputs(4432) <= a and not b;
    layer4_outputs(4433) <= not (a and b);
    layer4_outputs(4434) <= b;
    layer4_outputs(4435) <= not a or b;
    layer4_outputs(4436) <= a;
    layer4_outputs(4437) <= 1'b0;
    layer4_outputs(4438) <= not a;
    layer4_outputs(4439) <= b and not a;
    layer4_outputs(4440) <= b;
    layer4_outputs(4441) <= not a;
    layer4_outputs(4442) <= not b;
    layer4_outputs(4443) <= not (a and b);
    layer4_outputs(4444) <= not b;
    layer4_outputs(4445) <= a;
    layer4_outputs(4446) <= not (a or b);
    layer4_outputs(4447) <= not (a xor b);
    layer4_outputs(4448) <= not b;
    layer4_outputs(4449) <= not b or a;
    layer4_outputs(4450) <= 1'b1;
    layer4_outputs(4451) <= a xor b;
    layer4_outputs(4452) <= b and not a;
    layer4_outputs(4453) <= 1'b1;
    layer4_outputs(4454) <= a xor b;
    layer4_outputs(4455) <= not (a or b);
    layer4_outputs(4456) <= a and not b;
    layer4_outputs(4457) <= b and not a;
    layer4_outputs(4458) <= a;
    layer4_outputs(4459) <= a or b;
    layer4_outputs(4460) <= a or b;
    layer4_outputs(4461) <= a or b;
    layer4_outputs(4462) <= not a;
    layer4_outputs(4463) <= not b;
    layer4_outputs(4464) <= not (a or b);
    layer4_outputs(4465) <= not a;
    layer4_outputs(4466) <= not a;
    layer4_outputs(4467) <= 1'b0;
    layer4_outputs(4468) <= not a or b;
    layer4_outputs(4469) <= a or b;
    layer4_outputs(4470) <= a;
    layer4_outputs(4471) <= a xor b;
    layer4_outputs(4472) <= not b or a;
    layer4_outputs(4473) <= 1'b0;
    layer4_outputs(4474) <= not a or b;
    layer4_outputs(4475) <= not b or a;
    layer4_outputs(4476) <= not (a and b);
    layer4_outputs(4477) <= not a;
    layer4_outputs(4478) <= a or b;
    layer4_outputs(4479) <= a;
    layer4_outputs(4480) <= a and not b;
    layer4_outputs(4481) <= a;
    layer4_outputs(4482) <= not (a and b);
    layer4_outputs(4483) <= a;
    layer4_outputs(4484) <= a and b;
    layer4_outputs(4485) <= not (a xor b);
    layer4_outputs(4486) <= a xor b;
    layer4_outputs(4487) <= not b;
    layer4_outputs(4488) <= not (a and b);
    layer4_outputs(4489) <= a or b;
    layer4_outputs(4490) <= a or b;
    layer4_outputs(4491) <= a;
    layer4_outputs(4492) <= a and b;
    layer4_outputs(4493) <= not (a or b);
    layer4_outputs(4494) <= not b;
    layer4_outputs(4495) <= not (a xor b);
    layer4_outputs(4496) <= a and b;
    layer4_outputs(4497) <= not a or b;
    layer4_outputs(4498) <= not b or a;
    layer4_outputs(4499) <= not a;
    layer4_outputs(4500) <= not a;
    layer4_outputs(4501) <= 1'b1;
    layer4_outputs(4502) <= not b;
    layer4_outputs(4503) <= not (a and b);
    layer4_outputs(4504) <= not b;
    layer4_outputs(4505) <= not (a or b);
    layer4_outputs(4506) <= b;
    layer4_outputs(4507) <= not a;
    layer4_outputs(4508) <= not b;
    layer4_outputs(4509) <= not (a xor b);
    layer4_outputs(4510) <= b;
    layer4_outputs(4511) <= not b;
    layer4_outputs(4512) <= not (a or b);
    layer4_outputs(4513) <= not (a and b);
    layer4_outputs(4514) <= not b or a;
    layer4_outputs(4515) <= not (a or b);
    layer4_outputs(4516) <= b and not a;
    layer4_outputs(4517) <= b;
    layer4_outputs(4518) <= a xor b;
    layer4_outputs(4519) <= a and b;
    layer4_outputs(4520) <= a and b;
    layer4_outputs(4521) <= b and not a;
    layer4_outputs(4522) <= not b or a;
    layer4_outputs(4523) <= not (a or b);
    layer4_outputs(4524) <= not (a xor b);
    layer4_outputs(4525) <= a and b;
    layer4_outputs(4526) <= not (a and b);
    layer4_outputs(4527) <= 1'b0;
    layer4_outputs(4528) <= not b or a;
    layer4_outputs(4529) <= b;
    layer4_outputs(4530) <= not (a or b);
    layer4_outputs(4531) <= a and b;
    layer4_outputs(4532) <= b;
    layer4_outputs(4533) <= 1'b0;
    layer4_outputs(4534) <= a xor b;
    layer4_outputs(4535) <= not b or a;
    layer4_outputs(4536) <= a or b;
    layer4_outputs(4537) <= not (a and b);
    layer4_outputs(4538) <= not b;
    layer4_outputs(4539) <= not a;
    layer4_outputs(4540) <= 1'b1;
    layer4_outputs(4541) <= a or b;
    layer4_outputs(4542) <= not b;
    layer4_outputs(4543) <= not a or b;
    layer4_outputs(4544) <= not b;
    layer4_outputs(4545) <= 1'b1;
    layer4_outputs(4546) <= not (a and b);
    layer4_outputs(4547) <= a or b;
    layer4_outputs(4548) <= b;
    layer4_outputs(4549) <= not b or a;
    layer4_outputs(4550) <= a;
    layer4_outputs(4551) <= a or b;
    layer4_outputs(4552) <= not a;
    layer4_outputs(4553) <= b and not a;
    layer4_outputs(4554) <= a and not b;
    layer4_outputs(4555) <= b and not a;
    layer4_outputs(4556) <= not a or b;
    layer4_outputs(4557) <= 1'b1;
    layer4_outputs(4558) <= not (a or b);
    layer4_outputs(4559) <= 1'b1;
    layer4_outputs(4560) <= b;
    layer4_outputs(4561) <= b and not a;
    layer4_outputs(4562) <= a and b;
    layer4_outputs(4563) <= not b;
    layer4_outputs(4564) <= b;
    layer4_outputs(4565) <= not (a xor b);
    layer4_outputs(4566) <= not b or a;
    layer4_outputs(4567) <= not (a and b);
    layer4_outputs(4568) <= not a or b;
    layer4_outputs(4569) <= 1'b0;
    layer4_outputs(4570) <= not (a or b);
    layer4_outputs(4571) <= 1'b0;
    layer4_outputs(4572) <= a;
    layer4_outputs(4573) <= not a or b;
    layer4_outputs(4574) <= b;
    layer4_outputs(4575) <= 1'b1;
    layer4_outputs(4576) <= not b;
    layer4_outputs(4577) <= not b or a;
    layer4_outputs(4578) <= b;
    layer4_outputs(4579) <= not a;
    layer4_outputs(4580) <= a and b;
    layer4_outputs(4581) <= a or b;
    layer4_outputs(4582) <= not (a or b);
    layer4_outputs(4583) <= not a;
    layer4_outputs(4584) <= not (a xor b);
    layer4_outputs(4585) <= a and not b;
    layer4_outputs(4586) <= a;
    layer4_outputs(4587) <= a and not b;
    layer4_outputs(4588) <= not (a or b);
    layer4_outputs(4589) <= a;
    layer4_outputs(4590) <= 1'b0;
    layer4_outputs(4591) <= not (a or b);
    layer4_outputs(4592) <= not a;
    layer4_outputs(4593) <= b and not a;
    layer4_outputs(4594) <= not (a and b);
    layer4_outputs(4595) <= 1'b1;
    layer4_outputs(4596) <= 1'b1;
    layer4_outputs(4597) <= a or b;
    layer4_outputs(4598) <= 1'b0;
    layer4_outputs(4599) <= not (a or b);
    layer4_outputs(4600) <= 1'b0;
    layer4_outputs(4601) <= not b;
    layer4_outputs(4602) <= not a;
    layer4_outputs(4603) <= not a;
    layer4_outputs(4604) <= a and not b;
    layer4_outputs(4605) <= b;
    layer4_outputs(4606) <= a or b;
    layer4_outputs(4607) <= 1'b1;
    layer4_outputs(4608) <= b;
    layer4_outputs(4609) <= not b;
    layer4_outputs(4610) <= not b or a;
    layer4_outputs(4611) <= b and not a;
    layer4_outputs(4612) <= not b;
    layer4_outputs(4613) <= a;
    layer4_outputs(4614) <= not a or b;
    layer4_outputs(4615) <= a or b;
    layer4_outputs(4616) <= not a or b;
    layer4_outputs(4617) <= b;
    layer4_outputs(4618) <= a and b;
    layer4_outputs(4619) <= not b or a;
    layer4_outputs(4620) <= not b or a;
    layer4_outputs(4621) <= a xor b;
    layer4_outputs(4622) <= not b or a;
    layer4_outputs(4623) <= not b;
    layer4_outputs(4624) <= not b or a;
    layer4_outputs(4625) <= not a;
    layer4_outputs(4626) <= a and not b;
    layer4_outputs(4627) <= b and not a;
    layer4_outputs(4628) <= 1'b1;
    layer4_outputs(4629) <= a or b;
    layer4_outputs(4630) <= not (a or b);
    layer4_outputs(4631) <= a;
    layer4_outputs(4632) <= b;
    layer4_outputs(4633) <= 1'b0;
    layer4_outputs(4634) <= not (a and b);
    layer4_outputs(4635) <= 1'b0;
    layer4_outputs(4636) <= a or b;
    layer4_outputs(4637) <= 1'b0;
    layer4_outputs(4638) <= b and not a;
    layer4_outputs(4639) <= a;
    layer4_outputs(4640) <= a xor b;
    layer4_outputs(4641) <= not a or b;
    layer4_outputs(4642) <= not a;
    layer4_outputs(4643) <= not b or a;
    layer4_outputs(4644) <= not (a and b);
    layer4_outputs(4645) <= b and not a;
    layer4_outputs(4646) <= a and not b;
    layer4_outputs(4647) <= a and b;
    layer4_outputs(4648) <= b and not a;
    layer4_outputs(4649) <= not b;
    layer4_outputs(4650) <= not a;
    layer4_outputs(4651) <= b;
    layer4_outputs(4652) <= not (a and b);
    layer4_outputs(4653) <= a and not b;
    layer4_outputs(4654) <= a;
    layer4_outputs(4655) <= not (a or b);
    layer4_outputs(4656) <= not a;
    layer4_outputs(4657) <= not (a and b);
    layer4_outputs(4658) <= a;
    layer4_outputs(4659) <= b;
    layer4_outputs(4660) <= b and not a;
    layer4_outputs(4661) <= not b;
    layer4_outputs(4662) <= not a or b;
    layer4_outputs(4663) <= a xor b;
    layer4_outputs(4664) <= a and not b;
    layer4_outputs(4665) <= a and not b;
    layer4_outputs(4666) <= not a or b;
    layer4_outputs(4667) <= 1'b0;
    layer4_outputs(4668) <= a and b;
    layer4_outputs(4669) <= a;
    layer4_outputs(4670) <= a and b;
    layer4_outputs(4671) <= not (a and b);
    layer4_outputs(4672) <= not a;
    layer4_outputs(4673) <= not a;
    layer4_outputs(4674) <= not (a and b);
    layer4_outputs(4675) <= not b;
    layer4_outputs(4676) <= 1'b0;
    layer4_outputs(4677) <= b;
    layer4_outputs(4678) <= not a or b;
    layer4_outputs(4679) <= not b or a;
    layer4_outputs(4680) <= b;
    layer4_outputs(4681) <= 1'b0;
    layer4_outputs(4682) <= b;
    layer4_outputs(4683) <= not a or b;
    layer4_outputs(4684) <= not a;
    layer4_outputs(4685) <= a and b;
    layer4_outputs(4686) <= not a or b;
    layer4_outputs(4687) <= not a;
    layer4_outputs(4688) <= not a or b;
    layer4_outputs(4689) <= a and b;
    layer4_outputs(4690) <= not a or b;
    layer4_outputs(4691) <= 1'b1;
    layer4_outputs(4692) <= a and not b;
    layer4_outputs(4693) <= a and b;
    layer4_outputs(4694) <= not a;
    layer4_outputs(4695) <= a and b;
    layer4_outputs(4696) <= not (a and b);
    layer4_outputs(4697) <= a or b;
    layer4_outputs(4698) <= not b;
    layer4_outputs(4699) <= 1'b1;
    layer4_outputs(4700) <= not (a or b);
    layer4_outputs(4701) <= not a or b;
    layer4_outputs(4702) <= b;
    layer4_outputs(4703) <= not a;
    layer4_outputs(4704) <= not (a and b);
    layer4_outputs(4705) <= a xor b;
    layer4_outputs(4706) <= not (a and b);
    layer4_outputs(4707) <= a or b;
    layer4_outputs(4708) <= not a;
    layer4_outputs(4709) <= not b or a;
    layer4_outputs(4710) <= a or b;
    layer4_outputs(4711) <= a xor b;
    layer4_outputs(4712) <= not a;
    layer4_outputs(4713) <= not b or a;
    layer4_outputs(4714) <= a;
    layer4_outputs(4715) <= 1'b0;
    layer4_outputs(4716) <= 1'b0;
    layer4_outputs(4717) <= not b;
    layer4_outputs(4718) <= a;
    layer4_outputs(4719) <= a xor b;
    layer4_outputs(4720) <= not a or b;
    layer4_outputs(4721) <= b and not a;
    layer4_outputs(4722) <= 1'b1;
    layer4_outputs(4723) <= a and not b;
    layer4_outputs(4724) <= not (a xor b);
    layer4_outputs(4725) <= not (a xor b);
    layer4_outputs(4726) <= not b;
    layer4_outputs(4727) <= not a;
    layer4_outputs(4728) <= 1'b1;
    layer4_outputs(4729) <= not b;
    layer4_outputs(4730) <= a;
    layer4_outputs(4731) <= not b or a;
    layer4_outputs(4732) <= a;
    layer4_outputs(4733) <= a and not b;
    layer4_outputs(4734) <= a and not b;
    layer4_outputs(4735) <= not b;
    layer4_outputs(4736) <= a;
    layer4_outputs(4737) <= not (a or b);
    layer4_outputs(4738) <= not (a xor b);
    layer4_outputs(4739) <= not b;
    layer4_outputs(4740) <= not b or a;
    layer4_outputs(4741) <= 1'b0;
    layer4_outputs(4742) <= a and b;
    layer4_outputs(4743) <= 1'b1;
    layer4_outputs(4744) <= not (a and b);
    layer4_outputs(4745) <= a and b;
    layer4_outputs(4746) <= not b;
    layer4_outputs(4747) <= a;
    layer4_outputs(4748) <= not b or a;
    layer4_outputs(4749) <= a and b;
    layer4_outputs(4750) <= b;
    layer4_outputs(4751) <= not (a xor b);
    layer4_outputs(4752) <= a and not b;
    layer4_outputs(4753) <= a and b;
    layer4_outputs(4754) <= a and b;
    layer4_outputs(4755) <= not (a xor b);
    layer4_outputs(4756) <= a and b;
    layer4_outputs(4757) <= b;
    layer4_outputs(4758) <= not (a and b);
    layer4_outputs(4759) <= not (a and b);
    layer4_outputs(4760) <= b and not a;
    layer4_outputs(4761) <= not b;
    layer4_outputs(4762) <= a or b;
    layer4_outputs(4763) <= a xor b;
    layer4_outputs(4764) <= b and not a;
    layer4_outputs(4765) <= b;
    layer4_outputs(4766) <= a and not b;
    layer4_outputs(4767) <= not (a or b);
    layer4_outputs(4768) <= a xor b;
    layer4_outputs(4769) <= 1'b1;
    layer4_outputs(4770) <= not a or b;
    layer4_outputs(4771) <= not b or a;
    layer4_outputs(4772) <= a or b;
    layer4_outputs(4773) <= a;
    layer4_outputs(4774) <= a and not b;
    layer4_outputs(4775) <= 1'b1;
    layer4_outputs(4776) <= b and not a;
    layer4_outputs(4777) <= a xor b;
    layer4_outputs(4778) <= a or b;
    layer4_outputs(4779) <= a or b;
    layer4_outputs(4780) <= not (a or b);
    layer4_outputs(4781) <= 1'b0;
    layer4_outputs(4782) <= not a or b;
    layer4_outputs(4783) <= not (a or b);
    layer4_outputs(4784) <= not b or a;
    layer4_outputs(4785) <= b;
    layer4_outputs(4786) <= not a;
    layer4_outputs(4787) <= not (a and b);
    layer4_outputs(4788) <= not b or a;
    layer4_outputs(4789) <= 1'b0;
    layer4_outputs(4790) <= a and not b;
    layer4_outputs(4791) <= a and not b;
    layer4_outputs(4792) <= not (a or b);
    layer4_outputs(4793) <= not (a xor b);
    layer4_outputs(4794) <= a and not b;
    layer4_outputs(4795) <= not a;
    layer4_outputs(4796) <= b;
    layer4_outputs(4797) <= not b or a;
    layer4_outputs(4798) <= 1'b0;
    layer4_outputs(4799) <= a or b;
    layer4_outputs(4800) <= not a;
    layer4_outputs(4801) <= b and not a;
    layer4_outputs(4802) <= not b or a;
    layer4_outputs(4803) <= a or b;
    layer4_outputs(4804) <= a and b;
    layer4_outputs(4805) <= not b or a;
    layer4_outputs(4806) <= a and not b;
    layer4_outputs(4807) <= 1'b1;
    layer4_outputs(4808) <= not b;
    layer4_outputs(4809) <= a and b;
    layer4_outputs(4810) <= 1'b1;
    layer4_outputs(4811) <= 1'b1;
    layer4_outputs(4812) <= not (a or b);
    layer4_outputs(4813) <= a or b;
    layer4_outputs(4814) <= b;
    layer4_outputs(4815) <= 1'b1;
    layer4_outputs(4816) <= not (a and b);
    layer4_outputs(4817) <= not (a or b);
    layer4_outputs(4818) <= a and not b;
    layer4_outputs(4819) <= a or b;
    layer4_outputs(4820) <= not b or a;
    layer4_outputs(4821) <= not a or b;
    layer4_outputs(4822) <= a;
    layer4_outputs(4823) <= not b or a;
    layer4_outputs(4824) <= a;
    layer4_outputs(4825) <= not a or b;
    layer4_outputs(4826) <= a;
    layer4_outputs(4827) <= not (a or b);
    layer4_outputs(4828) <= not a;
    layer4_outputs(4829) <= b;
    layer4_outputs(4830) <= not b;
    layer4_outputs(4831) <= b and not a;
    layer4_outputs(4832) <= not (a and b);
    layer4_outputs(4833) <= a xor b;
    layer4_outputs(4834) <= b and not a;
    layer4_outputs(4835) <= 1'b0;
    layer4_outputs(4836) <= a;
    layer4_outputs(4837) <= not (a or b);
    layer4_outputs(4838) <= b;
    layer4_outputs(4839) <= a or b;
    layer4_outputs(4840) <= a;
    layer4_outputs(4841) <= 1'b0;
    layer4_outputs(4842) <= a or b;
    layer4_outputs(4843) <= not a or b;
    layer4_outputs(4844) <= b and not a;
    layer4_outputs(4845) <= not b;
    layer4_outputs(4846) <= not b or a;
    layer4_outputs(4847) <= b and not a;
    layer4_outputs(4848) <= a;
    layer4_outputs(4849) <= a;
    layer4_outputs(4850) <= not b;
    layer4_outputs(4851) <= not (a xor b);
    layer4_outputs(4852) <= not b;
    layer4_outputs(4853) <= a xor b;
    layer4_outputs(4854) <= not (a or b);
    layer4_outputs(4855) <= not b;
    layer4_outputs(4856) <= a;
    layer4_outputs(4857) <= a;
    layer4_outputs(4858) <= a and b;
    layer4_outputs(4859) <= a;
    layer4_outputs(4860) <= b;
    layer4_outputs(4861) <= 1'b1;
    layer4_outputs(4862) <= not a;
    layer4_outputs(4863) <= b and not a;
    layer4_outputs(4864) <= not a;
    layer4_outputs(4865) <= b;
    layer4_outputs(4866) <= not (a or b);
    layer4_outputs(4867) <= not b;
    layer4_outputs(4868) <= not (a and b);
    layer4_outputs(4869) <= a and not b;
    layer4_outputs(4870) <= not b;
    layer4_outputs(4871) <= a xor b;
    layer4_outputs(4872) <= not b or a;
    layer4_outputs(4873) <= a and b;
    layer4_outputs(4874) <= a and b;
    layer4_outputs(4875) <= a or b;
    layer4_outputs(4876) <= b and not a;
    layer4_outputs(4877) <= b;
    layer4_outputs(4878) <= a;
    layer4_outputs(4879) <= not b;
    layer4_outputs(4880) <= not b;
    layer4_outputs(4881) <= not (a or b);
    layer4_outputs(4882) <= a;
    layer4_outputs(4883) <= a and b;
    layer4_outputs(4884) <= not b or a;
    layer4_outputs(4885) <= not a or b;
    layer4_outputs(4886) <= not a;
    layer4_outputs(4887) <= b and not a;
    layer4_outputs(4888) <= a and not b;
    layer4_outputs(4889) <= b and not a;
    layer4_outputs(4890) <= not a or b;
    layer4_outputs(4891) <= a and b;
    layer4_outputs(4892) <= not a;
    layer4_outputs(4893) <= not (a or b);
    layer4_outputs(4894) <= a and b;
    layer4_outputs(4895) <= not b or a;
    layer4_outputs(4896) <= a or b;
    layer4_outputs(4897) <= not a;
    layer4_outputs(4898) <= 1'b0;
    layer4_outputs(4899) <= not a;
    layer4_outputs(4900) <= b and not a;
    layer4_outputs(4901) <= not a or b;
    layer4_outputs(4902) <= not b;
    layer4_outputs(4903) <= a or b;
    layer4_outputs(4904) <= b and not a;
    layer4_outputs(4905) <= 1'b0;
    layer4_outputs(4906) <= b;
    layer4_outputs(4907) <= a;
    layer4_outputs(4908) <= not b or a;
    layer4_outputs(4909) <= 1'b0;
    layer4_outputs(4910) <= a or b;
    layer4_outputs(4911) <= not b;
    layer4_outputs(4912) <= a or b;
    layer4_outputs(4913) <= a and b;
    layer4_outputs(4914) <= not b or a;
    layer4_outputs(4915) <= not a or b;
    layer4_outputs(4916) <= not a or b;
    layer4_outputs(4917) <= a or b;
    layer4_outputs(4918) <= not b;
    layer4_outputs(4919) <= not a;
    layer4_outputs(4920) <= a and b;
    layer4_outputs(4921) <= not a;
    layer4_outputs(4922) <= not (a or b);
    layer4_outputs(4923) <= not b;
    layer4_outputs(4924) <= a xor b;
    layer4_outputs(4925) <= a and not b;
    layer4_outputs(4926) <= 1'b0;
    layer4_outputs(4927) <= not b;
    layer4_outputs(4928) <= b and not a;
    layer4_outputs(4929) <= a or b;
    layer4_outputs(4930) <= a xor b;
    layer4_outputs(4931) <= not a;
    layer4_outputs(4932) <= b and not a;
    layer4_outputs(4933) <= 1'b1;
    layer4_outputs(4934) <= a;
    layer4_outputs(4935) <= a;
    layer4_outputs(4936) <= b;
    layer4_outputs(4937) <= not (a or b);
    layer4_outputs(4938) <= not (a or b);
    layer4_outputs(4939) <= not b;
    layer4_outputs(4940) <= not (a and b);
    layer4_outputs(4941) <= 1'b0;
    layer4_outputs(4942) <= a;
    layer4_outputs(4943) <= not a or b;
    layer4_outputs(4944) <= not (a xor b);
    layer4_outputs(4945) <= a and not b;
    layer4_outputs(4946) <= a and not b;
    layer4_outputs(4947) <= not (a and b);
    layer4_outputs(4948) <= a xor b;
    layer4_outputs(4949) <= a and not b;
    layer4_outputs(4950) <= a;
    layer4_outputs(4951) <= 1'b0;
    layer4_outputs(4952) <= b;
    layer4_outputs(4953) <= 1'b1;
    layer4_outputs(4954) <= b and not a;
    layer4_outputs(4955) <= b;
    layer4_outputs(4956) <= a;
    layer4_outputs(4957) <= not b or a;
    layer4_outputs(4958) <= not a;
    layer4_outputs(4959) <= 1'b1;
    layer4_outputs(4960) <= b;
    layer4_outputs(4961) <= not a or b;
    layer4_outputs(4962) <= not a or b;
    layer4_outputs(4963) <= a or b;
    layer4_outputs(4964) <= a or b;
    layer4_outputs(4965) <= not a or b;
    layer4_outputs(4966) <= b and not a;
    layer4_outputs(4967) <= not (a or b);
    layer4_outputs(4968) <= not (a and b);
    layer4_outputs(4969) <= not b;
    layer4_outputs(4970) <= b and not a;
    layer4_outputs(4971) <= not (a or b);
    layer4_outputs(4972) <= not a;
    layer4_outputs(4973) <= 1'b1;
    layer4_outputs(4974) <= not b or a;
    layer4_outputs(4975) <= a xor b;
    layer4_outputs(4976) <= not (a or b);
    layer4_outputs(4977) <= not (a xor b);
    layer4_outputs(4978) <= not a;
    layer4_outputs(4979) <= not b;
    layer4_outputs(4980) <= a;
    layer4_outputs(4981) <= not a;
    layer4_outputs(4982) <= not (a and b);
    layer4_outputs(4983) <= a and b;
    layer4_outputs(4984) <= b;
    layer4_outputs(4985) <= 1'b0;
    layer4_outputs(4986) <= b and not a;
    layer4_outputs(4987) <= not (a and b);
    layer4_outputs(4988) <= not b;
    layer4_outputs(4989) <= 1'b0;
    layer4_outputs(4990) <= b;
    layer4_outputs(4991) <= not b;
    layer4_outputs(4992) <= not (a and b);
    layer4_outputs(4993) <= not (a and b);
    layer4_outputs(4994) <= b and not a;
    layer4_outputs(4995) <= a xor b;
    layer4_outputs(4996) <= a;
    layer4_outputs(4997) <= a and b;
    layer4_outputs(4998) <= not b;
    layer4_outputs(4999) <= not b;
    layer4_outputs(5000) <= b and not a;
    layer4_outputs(5001) <= not b;
    layer4_outputs(5002) <= not a or b;
    layer4_outputs(5003) <= a xor b;
    layer4_outputs(5004) <= not (a and b);
    layer4_outputs(5005) <= 1'b1;
    layer4_outputs(5006) <= a;
    layer4_outputs(5007) <= a or b;
    layer4_outputs(5008) <= b;
    layer4_outputs(5009) <= a;
    layer4_outputs(5010) <= not b or a;
    layer4_outputs(5011) <= a;
    layer4_outputs(5012) <= b;
    layer4_outputs(5013) <= not a or b;
    layer4_outputs(5014) <= not b or a;
    layer4_outputs(5015) <= 1'b0;
    layer4_outputs(5016) <= b;
    layer4_outputs(5017) <= not b;
    layer4_outputs(5018) <= b and not a;
    layer4_outputs(5019) <= a and not b;
    layer4_outputs(5020) <= not b;
    layer4_outputs(5021) <= a or b;
    layer4_outputs(5022) <= a and not b;
    layer4_outputs(5023) <= 1'b0;
    layer4_outputs(5024) <= not b;
    layer4_outputs(5025) <= 1'b1;
    layer4_outputs(5026) <= a or b;
    layer4_outputs(5027) <= 1'b0;
    layer4_outputs(5028) <= a and not b;
    layer4_outputs(5029) <= not b or a;
    layer4_outputs(5030) <= not (a or b);
    layer4_outputs(5031) <= not b or a;
    layer4_outputs(5032) <= 1'b0;
    layer4_outputs(5033) <= not (a xor b);
    layer4_outputs(5034) <= a or b;
    layer4_outputs(5035) <= a xor b;
    layer4_outputs(5036) <= a and b;
    layer4_outputs(5037) <= b and not a;
    layer4_outputs(5038) <= not (a or b);
    layer4_outputs(5039) <= a;
    layer4_outputs(5040) <= not a or b;
    layer4_outputs(5041) <= not (a or b);
    layer4_outputs(5042) <= not (a or b);
    layer4_outputs(5043) <= 1'b1;
    layer4_outputs(5044) <= not (a and b);
    layer4_outputs(5045) <= not b;
    layer4_outputs(5046) <= not b;
    layer4_outputs(5047) <= b and not a;
    layer4_outputs(5048) <= a and not b;
    layer4_outputs(5049) <= b;
    layer4_outputs(5050) <= b and not a;
    layer4_outputs(5051) <= a;
    layer4_outputs(5052) <= not a;
    layer4_outputs(5053) <= 1'b0;
    layer4_outputs(5054) <= 1'b1;
    layer4_outputs(5055) <= a xor b;
    layer4_outputs(5056) <= not a;
    layer4_outputs(5057) <= not (a or b);
    layer4_outputs(5058) <= a or b;
    layer4_outputs(5059) <= not b;
    layer4_outputs(5060) <= not a;
    layer4_outputs(5061) <= a or b;
    layer4_outputs(5062) <= not a or b;
    layer4_outputs(5063) <= 1'b0;
    layer4_outputs(5064) <= not (a and b);
    layer4_outputs(5065) <= b;
    layer4_outputs(5066) <= a and not b;
    layer4_outputs(5067) <= a;
    layer4_outputs(5068) <= b;
    layer4_outputs(5069) <= 1'b1;
    layer4_outputs(5070) <= not (a xor b);
    layer4_outputs(5071) <= a and not b;
    layer4_outputs(5072) <= not a;
    layer4_outputs(5073) <= a and not b;
    layer4_outputs(5074) <= b;
    layer4_outputs(5075) <= a and not b;
    layer4_outputs(5076) <= a and b;
    layer4_outputs(5077) <= a xor b;
    layer4_outputs(5078) <= not b;
    layer4_outputs(5079) <= not a;
    layer4_outputs(5080) <= a and not b;
    layer4_outputs(5081) <= not (a or b);
    layer4_outputs(5082) <= a or b;
    layer4_outputs(5083) <= not b;
    layer4_outputs(5084) <= a xor b;
    layer4_outputs(5085) <= b and not a;
    layer4_outputs(5086) <= not b;
    layer4_outputs(5087) <= a;
    layer4_outputs(5088) <= b;
    layer4_outputs(5089) <= 1'b0;
    layer4_outputs(5090) <= not b or a;
    layer4_outputs(5091) <= a and not b;
    layer4_outputs(5092) <= not (a xor b);
    layer4_outputs(5093) <= a or b;
    layer4_outputs(5094) <= b and not a;
    layer4_outputs(5095) <= 1'b0;
    layer4_outputs(5096) <= b and not a;
    layer4_outputs(5097) <= a and not b;
    layer4_outputs(5098) <= not a or b;
    layer4_outputs(5099) <= not a;
    layer4_outputs(5100) <= a and not b;
    layer4_outputs(5101) <= not b or a;
    layer4_outputs(5102) <= b and not a;
    layer4_outputs(5103) <= a and b;
    layer4_outputs(5104) <= not (a and b);
    layer4_outputs(5105) <= a;
    layer4_outputs(5106) <= not a or b;
    layer4_outputs(5107) <= not a or b;
    layer4_outputs(5108) <= not b or a;
    layer4_outputs(5109) <= b;
    layer4_outputs(5110) <= 1'b1;
    layer4_outputs(5111) <= not a;
    layer4_outputs(5112) <= a and b;
    layer4_outputs(5113) <= a xor b;
    layer4_outputs(5114) <= a and not b;
    layer4_outputs(5115) <= not b or a;
    layer4_outputs(5116) <= a or b;
    layer4_outputs(5117) <= b;
    layer4_outputs(5118) <= not (a xor b);
    layer4_outputs(5119) <= not a or b;
    layer4_outputs(5120) <= not (a and b);
    layer4_outputs(5121) <= not b;
    layer4_outputs(5122) <= not b;
    layer4_outputs(5123) <= not b or a;
    layer4_outputs(5124) <= not (a and b);
    layer4_outputs(5125) <= not b;
    layer4_outputs(5126) <= not (a or b);
    layer4_outputs(5127) <= a;
    layer4_outputs(5128) <= a;
    layer4_outputs(5129) <= a;
    layer4_outputs(5130) <= 1'b1;
    layer4_outputs(5131) <= not b;
    layer4_outputs(5132) <= b;
    layer4_outputs(5133) <= a and b;
    layer4_outputs(5134) <= not (a and b);
    layer4_outputs(5135) <= not (a and b);
    layer4_outputs(5136) <= a and b;
    layer4_outputs(5137) <= not a or b;
    layer4_outputs(5138) <= 1'b0;
    layer4_outputs(5139) <= not (a xor b);
    layer4_outputs(5140) <= a or b;
    layer4_outputs(5141) <= not a;
    layer4_outputs(5142) <= b and not a;
    layer4_outputs(5143) <= a;
    layer4_outputs(5144) <= not a;
    layer4_outputs(5145) <= not (a or b);
    layer4_outputs(5146) <= a and not b;
    layer4_outputs(5147) <= not b;
    layer4_outputs(5148) <= not b or a;
    layer4_outputs(5149) <= not b;
    layer4_outputs(5150) <= a or b;
    layer4_outputs(5151) <= 1'b1;
    layer4_outputs(5152) <= not (a and b);
    layer4_outputs(5153) <= not a or b;
    layer4_outputs(5154) <= 1'b1;
    layer4_outputs(5155) <= not a;
    layer4_outputs(5156) <= not a or b;
    layer4_outputs(5157) <= a;
    layer4_outputs(5158) <= a;
    layer4_outputs(5159) <= a and b;
    layer4_outputs(5160) <= a and not b;
    layer4_outputs(5161) <= a;
    layer4_outputs(5162) <= a and not b;
    layer4_outputs(5163) <= a and not b;
    layer4_outputs(5164) <= not b;
    layer4_outputs(5165) <= not (a and b);
    layer4_outputs(5166) <= not (a and b);
    layer4_outputs(5167) <= 1'b1;
    layer4_outputs(5168) <= not (a and b);
    layer4_outputs(5169) <= not a;
    layer4_outputs(5170) <= a;
    layer4_outputs(5171) <= b and not a;
    layer4_outputs(5172) <= not a;
    layer4_outputs(5173) <= a and b;
    layer4_outputs(5174) <= a;
    layer4_outputs(5175) <= a and b;
    layer4_outputs(5176) <= b and not a;
    layer4_outputs(5177) <= not b;
    layer4_outputs(5178) <= 1'b0;
    layer4_outputs(5179) <= a or b;
    layer4_outputs(5180) <= b;
    layer4_outputs(5181) <= b;
    layer4_outputs(5182) <= a and b;
    layer4_outputs(5183) <= not a or b;
    layer4_outputs(5184) <= not (a xor b);
    layer4_outputs(5185) <= a and b;
    layer4_outputs(5186) <= not a;
    layer4_outputs(5187) <= 1'b0;
    layer4_outputs(5188) <= not (a xor b);
    layer4_outputs(5189) <= a;
    layer4_outputs(5190) <= b;
    layer4_outputs(5191) <= b and not a;
    layer4_outputs(5192) <= b;
    layer4_outputs(5193) <= a xor b;
    layer4_outputs(5194) <= not (a and b);
    layer4_outputs(5195) <= b;
    layer4_outputs(5196) <= a and b;
    layer4_outputs(5197) <= 1'b1;
    layer4_outputs(5198) <= not b or a;
    layer4_outputs(5199) <= not (a xor b);
    layer4_outputs(5200) <= a;
    layer4_outputs(5201) <= not (a or b);
    layer4_outputs(5202) <= b;
    layer4_outputs(5203) <= b;
    layer4_outputs(5204) <= not b;
    layer4_outputs(5205) <= not b or a;
    layer4_outputs(5206) <= a and not b;
    layer4_outputs(5207) <= a or b;
    layer4_outputs(5208) <= a xor b;
    layer4_outputs(5209) <= not (a xor b);
    layer4_outputs(5210) <= 1'b1;
    layer4_outputs(5211) <= a and not b;
    layer4_outputs(5212) <= a and not b;
    layer4_outputs(5213) <= not b or a;
    layer4_outputs(5214) <= b and not a;
    layer4_outputs(5215) <= b;
    layer4_outputs(5216) <= b and not a;
    layer4_outputs(5217) <= a and b;
    layer4_outputs(5218) <= 1'b1;
    layer4_outputs(5219) <= b;
    layer4_outputs(5220) <= not b;
    layer4_outputs(5221) <= not b or a;
    layer4_outputs(5222) <= not (a or b);
    layer4_outputs(5223) <= a;
    layer4_outputs(5224) <= a or b;
    layer4_outputs(5225) <= a and b;
    layer4_outputs(5226) <= b;
    layer4_outputs(5227) <= not (a and b);
    layer4_outputs(5228) <= not b;
    layer4_outputs(5229) <= a;
    layer4_outputs(5230) <= not a or b;
    layer4_outputs(5231) <= a xor b;
    layer4_outputs(5232) <= not (a or b);
    layer4_outputs(5233) <= not (a or b);
    layer4_outputs(5234) <= not (a or b);
    layer4_outputs(5235) <= not a or b;
    layer4_outputs(5236) <= a;
    layer4_outputs(5237) <= not a;
    layer4_outputs(5238) <= not (a and b);
    layer4_outputs(5239) <= not (a or b);
    layer4_outputs(5240) <= not b;
    layer4_outputs(5241) <= not (a xor b);
    layer4_outputs(5242) <= not a or b;
    layer4_outputs(5243) <= a;
    layer4_outputs(5244) <= 1'b0;
    layer4_outputs(5245) <= not b;
    layer4_outputs(5246) <= not a or b;
    layer4_outputs(5247) <= not b;
    layer4_outputs(5248) <= not a;
    layer4_outputs(5249) <= b;
    layer4_outputs(5250) <= 1'b0;
    layer4_outputs(5251) <= 1'b0;
    layer4_outputs(5252) <= 1'b0;
    layer4_outputs(5253) <= not a;
    layer4_outputs(5254) <= not (a or b);
    layer4_outputs(5255) <= 1'b1;
    layer4_outputs(5256) <= not b or a;
    layer4_outputs(5257) <= a xor b;
    layer4_outputs(5258) <= not (a and b);
    layer4_outputs(5259) <= not a or b;
    layer4_outputs(5260) <= not a;
    layer4_outputs(5261) <= not b or a;
    layer4_outputs(5262) <= a;
    layer4_outputs(5263) <= b;
    layer4_outputs(5264) <= 1'b0;
    layer4_outputs(5265) <= not a;
    layer4_outputs(5266) <= a;
    layer4_outputs(5267) <= not b;
    layer4_outputs(5268) <= not a or b;
    layer4_outputs(5269) <= 1'b1;
    layer4_outputs(5270) <= not a or b;
    layer4_outputs(5271) <= a xor b;
    layer4_outputs(5272) <= a xor b;
    layer4_outputs(5273) <= not b or a;
    layer4_outputs(5274) <= a or b;
    layer4_outputs(5275) <= a or b;
    layer4_outputs(5276) <= not (a xor b);
    layer4_outputs(5277) <= a and b;
    layer4_outputs(5278) <= not (a or b);
    layer4_outputs(5279) <= b and not a;
    layer4_outputs(5280) <= a or b;
    layer4_outputs(5281) <= not b;
    layer4_outputs(5282) <= b and not a;
    layer4_outputs(5283) <= not b;
    layer4_outputs(5284) <= not a;
    layer4_outputs(5285) <= not (a and b);
    layer4_outputs(5286) <= not b;
    layer4_outputs(5287) <= not b or a;
    layer4_outputs(5288) <= not (a or b);
    layer4_outputs(5289) <= not a or b;
    layer4_outputs(5290) <= 1'b0;
    layer4_outputs(5291) <= not (a and b);
    layer4_outputs(5292) <= 1'b0;
    layer4_outputs(5293) <= not (a and b);
    layer4_outputs(5294) <= b;
    layer4_outputs(5295) <= a or b;
    layer4_outputs(5296) <= not (a or b);
    layer4_outputs(5297) <= a or b;
    layer4_outputs(5298) <= not a;
    layer4_outputs(5299) <= not b or a;
    layer4_outputs(5300) <= 1'b0;
    layer4_outputs(5301) <= not b;
    layer4_outputs(5302) <= not a;
    layer4_outputs(5303) <= not b;
    layer4_outputs(5304) <= a;
    layer4_outputs(5305) <= a and not b;
    layer4_outputs(5306) <= not b;
    layer4_outputs(5307) <= a and b;
    layer4_outputs(5308) <= not a or b;
    layer4_outputs(5309) <= 1'b0;
    layer4_outputs(5310) <= not (a xor b);
    layer4_outputs(5311) <= b and not a;
    layer4_outputs(5312) <= a and b;
    layer4_outputs(5313) <= not (a or b);
    layer4_outputs(5314) <= a and b;
    layer4_outputs(5315) <= not (a and b);
    layer4_outputs(5316) <= not b or a;
    layer4_outputs(5317) <= a;
    layer4_outputs(5318) <= not a;
    layer4_outputs(5319) <= not a;
    layer4_outputs(5320) <= 1'b1;
    layer4_outputs(5321) <= 1'b0;
    layer4_outputs(5322) <= a and b;
    layer4_outputs(5323) <= b;
    layer4_outputs(5324) <= 1'b0;
    layer4_outputs(5325) <= b and not a;
    layer4_outputs(5326) <= a and b;
    layer4_outputs(5327) <= not a or b;
    layer4_outputs(5328) <= not b;
    layer4_outputs(5329) <= b;
    layer4_outputs(5330) <= b and not a;
    layer4_outputs(5331) <= b and not a;
    layer4_outputs(5332) <= not (a xor b);
    layer4_outputs(5333) <= b and not a;
    layer4_outputs(5334) <= 1'b1;
    layer4_outputs(5335) <= a or b;
    layer4_outputs(5336) <= not a;
    layer4_outputs(5337) <= a and not b;
    layer4_outputs(5338) <= not a;
    layer4_outputs(5339) <= a;
    layer4_outputs(5340) <= not a;
    layer4_outputs(5341) <= not a;
    layer4_outputs(5342) <= a and not b;
    layer4_outputs(5343) <= a and b;
    layer4_outputs(5344) <= a or b;
    layer4_outputs(5345) <= not b or a;
    layer4_outputs(5346) <= not (a and b);
    layer4_outputs(5347) <= a and b;
    layer4_outputs(5348) <= a or b;
    layer4_outputs(5349) <= not b or a;
    layer4_outputs(5350) <= a xor b;
    layer4_outputs(5351) <= b and not a;
    layer4_outputs(5352) <= a;
    layer4_outputs(5353) <= 1'b0;
    layer4_outputs(5354) <= a and not b;
    layer4_outputs(5355) <= a and b;
    layer4_outputs(5356) <= a or b;
    layer4_outputs(5357) <= 1'b0;
    layer4_outputs(5358) <= a xor b;
    layer4_outputs(5359) <= a or b;
    layer4_outputs(5360) <= 1'b1;
    layer4_outputs(5361) <= b;
    layer4_outputs(5362) <= not b;
    layer4_outputs(5363) <= a;
    layer4_outputs(5364) <= a and not b;
    layer4_outputs(5365) <= not b;
    layer4_outputs(5366) <= not a or b;
    layer4_outputs(5367) <= a;
    layer4_outputs(5368) <= not b;
    layer4_outputs(5369) <= not b;
    layer4_outputs(5370) <= a xor b;
    layer4_outputs(5371) <= not (a and b);
    layer4_outputs(5372) <= a xor b;
    layer4_outputs(5373) <= not a or b;
    layer4_outputs(5374) <= not a or b;
    layer4_outputs(5375) <= b;
    layer4_outputs(5376) <= b and not a;
    layer4_outputs(5377) <= not a;
    layer4_outputs(5378) <= not b;
    layer4_outputs(5379) <= a or b;
    layer4_outputs(5380) <= a;
    layer4_outputs(5381) <= 1'b0;
    layer4_outputs(5382) <= 1'b1;
    layer4_outputs(5383) <= not (a or b);
    layer4_outputs(5384) <= a or b;
    layer4_outputs(5385) <= a and b;
    layer4_outputs(5386) <= a and b;
    layer4_outputs(5387) <= not (a xor b);
    layer4_outputs(5388) <= not b;
    layer4_outputs(5389) <= b;
    layer4_outputs(5390) <= a and b;
    layer4_outputs(5391) <= b;
    layer4_outputs(5392) <= 1'b0;
    layer4_outputs(5393) <= 1'b0;
    layer4_outputs(5394) <= b and not a;
    layer4_outputs(5395) <= not b or a;
    layer4_outputs(5396) <= not a;
    layer4_outputs(5397) <= not a or b;
    layer4_outputs(5398) <= a;
    layer4_outputs(5399) <= not a or b;
    layer4_outputs(5400) <= 1'b0;
    layer4_outputs(5401) <= not a;
    layer4_outputs(5402) <= not (a and b);
    layer4_outputs(5403) <= not b or a;
    layer4_outputs(5404) <= 1'b0;
    layer4_outputs(5405) <= not a or b;
    layer4_outputs(5406) <= b and not a;
    layer4_outputs(5407) <= not a;
    layer4_outputs(5408) <= 1'b0;
    layer4_outputs(5409) <= not b or a;
    layer4_outputs(5410) <= a or b;
    layer4_outputs(5411) <= not (a or b);
    layer4_outputs(5412) <= a;
    layer4_outputs(5413) <= b;
    layer4_outputs(5414) <= a or b;
    layer4_outputs(5415) <= 1'b0;
    layer4_outputs(5416) <= not (a and b);
    layer4_outputs(5417) <= a or b;
    layer4_outputs(5418) <= not (a xor b);
    layer4_outputs(5419) <= a;
    layer4_outputs(5420) <= not b or a;
    layer4_outputs(5421) <= b;
    layer4_outputs(5422) <= not (a or b);
    layer4_outputs(5423) <= b;
    layer4_outputs(5424) <= a and b;
    layer4_outputs(5425) <= not (a or b);
    layer4_outputs(5426) <= b and not a;
    layer4_outputs(5427) <= b and not a;
    layer4_outputs(5428) <= 1'b1;
    layer4_outputs(5429) <= a or b;
    layer4_outputs(5430) <= b and not a;
    layer4_outputs(5431) <= a;
    layer4_outputs(5432) <= a;
    layer4_outputs(5433) <= b and not a;
    layer4_outputs(5434) <= not b or a;
    layer4_outputs(5435) <= not a or b;
    layer4_outputs(5436) <= 1'b0;
    layer4_outputs(5437) <= not (a xor b);
    layer4_outputs(5438) <= not b or a;
    layer4_outputs(5439) <= b;
    layer4_outputs(5440) <= not (a xor b);
    layer4_outputs(5441) <= 1'b1;
    layer4_outputs(5442) <= a and not b;
    layer4_outputs(5443) <= a and not b;
    layer4_outputs(5444) <= not (a xor b);
    layer4_outputs(5445) <= a and not b;
    layer4_outputs(5446) <= a or b;
    layer4_outputs(5447) <= not a;
    layer4_outputs(5448) <= b and not a;
    layer4_outputs(5449) <= not (a and b);
    layer4_outputs(5450) <= a and not b;
    layer4_outputs(5451) <= a and b;
    layer4_outputs(5452) <= 1'b1;
    layer4_outputs(5453) <= b;
    layer4_outputs(5454) <= a or b;
    layer4_outputs(5455) <= not (a and b);
    layer4_outputs(5456) <= b;
    layer4_outputs(5457) <= b;
    layer4_outputs(5458) <= not (a and b);
    layer4_outputs(5459) <= not (a or b);
    layer4_outputs(5460) <= not a;
    layer4_outputs(5461) <= not (a or b);
    layer4_outputs(5462) <= a;
    layer4_outputs(5463) <= not b;
    layer4_outputs(5464) <= not a;
    layer4_outputs(5465) <= not a;
    layer4_outputs(5466) <= not b or a;
    layer4_outputs(5467) <= a and b;
    layer4_outputs(5468) <= b;
    layer4_outputs(5469) <= a and b;
    layer4_outputs(5470) <= a or b;
    layer4_outputs(5471) <= a;
    layer4_outputs(5472) <= a and not b;
    layer4_outputs(5473) <= not (a or b);
    layer4_outputs(5474) <= not a;
    layer4_outputs(5475) <= not (a and b);
    layer4_outputs(5476) <= not (a or b);
    layer4_outputs(5477) <= a and not b;
    layer4_outputs(5478) <= a or b;
    layer4_outputs(5479) <= a xor b;
    layer4_outputs(5480) <= not (a or b);
    layer4_outputs(5481) <= not a;
    layer4_outputs(5482) <= a and not b;
    layer4_outputs(5483) <= not b or a;
    layer4_outputs(5484) <= a and b;
    layer4_outputs(5485) <= not a;
    layer4_outputs(5486) <= not b;
    layer4_outputs(5487) <= not a;
    layer4_outputs(5488) <= not a;
    layer4_outputs(5489) <= not a;
    layer4_outputs(5490) <= not (a and b);
    layer4_outputs(5491) <= a and not b;
    layer4_outputs(5492) <= not a or b;
    layer4_outputs(5493) <= a;
    layer4_outputs(5494) <= not (a or b);
    layer4_outputs(5495) <= not b or a;
    layer4_outputs(5496) <= a and b;
    layer4_outputs(5497) <= not a;
    layer4_outputs(5498) <= not b or a;
    layer4_outputs(5499) <= a and not b;
    layer4_outputs(5500) <= b;
    layer4_outputs(5501) <= a or b;
    layer4_outputs(5502) <= 1'b0;
    layer4_outputs(5503) <= b;
    layer4_outputs(5504) <= a and b;
    layer4_outputs(5505) <= b and not a;
    layer4_outputs(5506) <= not a or b;
    layer4_outputs(5507) <= 1'b0;
    layer4_outputs(5508) <= b and not a;
    layer4_outputs(5509) <= not b;
    layer4_outputs(5510) <= not a or b;
    layer4_outputs(5511) <= not a or b;
    layer4_outputs(5512) <= a xor b;
    layer4_outputs(5513) <= not (a and b);
    layer4_outputs(5514) <= a xor b;
    layer4_outputs(5515) <= b and not a;
    layer4_outputs(5516) <= 1'b1;
    layer4_outputs(5517) <= a and b;
    layer4_outputs(5518) <= a and b;
    layer4_outputs(5519) <= a or b;
    layer4_outputs(5520) <= a;
    layer4_outputs(5521) <= not a or b;
    layer4_outputs(5522) <= a and not b;
    layer4_outputs(5523) <= b and not a;
    layer4_outputs(5524) <= a;
    layer4_outputs(5525) <= not (a xor b);
    layer4_outputs(5526) <= b;
    layer4_outputs(5527) <= not a;
    layer4_outputs(5528) <= a xor b;
    layer4_outputs(5529) <= a;
    layer4_outputs(5530) <= not (a or b);
    layer4_outputs(5531) <= 1'b0;
    layer4_outputs(5532) <= a and not b;
    layer4_outputs(5533) <= 1'b1;
    layer4_outputs(5534) <= a or b;
    layer4_outputs(5535) <= a or b;
    layer4_outputs(5536) <= not a;
    layer4_outputs(5537) <= not b or a;
    layer4_outputs(5538) <= a or b;
    layer4_outputs(5539) <= a;
    layer4_outputs(5540) <= b and not a;
    layer4_outputs(5541) <= not b or a;
    layer4_outputs(5542) <= not b or a;
    layer4_outputs(5543) <= not b or a;
    layer4_outputs(5544) <= a or b;
    layer4_outputs(5545) <= 1'b0;
    layer4_outputs(5546) <= b;
    layer4_outputs(5547) <= b and not a;
    layer4_outputs(5548) <= a and not b;
    layer4_outputs(5549) <= b and not a;
    layer4_outputs(5550) <= not b;
    layer4_outputs(5551) <= a or b;
    layer4_outputs(5552) <= not a;
    layer4_outputs(5553) <= not b;
    layer4_outputs(5554) <= not a or b;
    layer4_outputs(5555) <= a xor b;
    layer4_outputs(5556) <= not b;
    layer4_outputs(5557) <= not a or b;
    layer4_outputs(5558) <= a and b;
    layer4_outputs(5559) <= not a or b;
    layer4_outputs(5560) <= 1'b1;
    layer4_outputs(5561) <= a and b;
    layer4_outputs(5562) <= not (a or b);
    layer4_outputs(5563) <= a and b;
    layer4_outputs(5564) <= a and not b;
    layer4_outputs(5565) <= not a;
    layer4_outputs(5566) <= not (a and b);
    layer4_outputs(5567) <= a and not b;
    layer4_outputs(5568) <= a and b;
    layer4_outputs(5569) <= 1'b1;
    layer4_outputs(5570) <= a and not b;
    layer4_outputs(5571) <= a and not b;
    layer4_outputs(5572) <= a and b;
    layer4_outputs(5573) <= not b or a;
    layer4_outputs(5574) <= not a;
    layer4_outputs(5575) <= not (a xor b);
    layer4_outputs(5576) <= a or b;
    layer4_outputs(5577) <= a or b;
    layer4_outputs(5578) <= 1'b0;
    layer4_outputs(5579) <= a;
    layer4_outputs(5580) <= not (a and b);
    layer4_outputs(5581) <= not a;
    layer4_outputs(5582) <= 1'b0;
    layer4_outputs(5583) <= b;
    layer4_outputs(5584) <= not (a and b);
    layer4_outputs(5585) <= not a or b;
    layer4_outputs(5586) <= a and not b;
    layer4_outputs(5587) <= not b;
    layer4_outputs(5588) <= a and b;
    layer4_outputs(5589) <= not b or a;
    layer4_outputs(5590) <= a;
    layer4_outputs(5591) <= not (a and b);
    layer4_outputs(5592) <= not (a and b);
    layer4_outputs(5593) <= a;
    layer4_outputs(5594) <= not (a xor b);
    layer4_outputs(5595) <= not b;
    layer4_outputs(5596) <= not a or b;
    layer4_outputs(5597) <= not b;
    layer4_outputs(5598) <= a and b;
    layer4_outputs(5599) <= not (a or b);
    layer4_outputs(5600) <= a;
    layer4_outputs(5601) <= a and not b;
    layer4_outputs(5602) <= a and b;
    layer4_outputs(5603) <= 1'b1;
    layer4_outputs(5604) <= not (a or b);
    layer4_outputs(5605) <= b;
    layer4_outputs(5606) <= not (a or b);
    layer4_outputs(5607) <= 1'b1;
    layer4_outputs(5608) <= a and b;
    layer4_outputs(5609) <= a and not b;
    layer4_outputs(5610) <= a and b;
    layer4_outputs(5611) <= not a;
    layer4_outputs(5612) <= a and b;
    layer4_outputs(5613) <= a;
    layer4_outputs(5614) <= a and b;
    layer4_outputs(5615) <= a or b;
    layer4_outputs(5616) <= b and not a;
    layer4_outputs(5617) <= 1'b0;
    layer4_outputs(5618) <= a;
    layer4_outputs(5619) <= 1'b1;
    layer4_outputs(5620) <= not b;
    layer4_outputs(5621) <= 1'b0;
    layer4_outputs(5622) <= a xor b;
    layer4_outputs(5623) <= a and b;
    layer4_outputs(5624) <= not (a and b);
    layer4_outputs(5625) <= 1'b0;
    layer4_outputs(5626) <= not (a xor b);
    layer4_outputs(5627) <= b and not a;
    layer4_outputs(5628) <= b and not a;
    layer4_outputs(5629) <= not a;
    layer4_outputs(5630) <= 1'b1;
    layer4_outputs(5631) <= not (a or b);
    layer4_outputs(5632) <= not (a xor b);
    layer4_outputs(5633) <= 1'b0;
    layer4_outputs(5634) <= a or b;
    layer4_outputs(5635) <= a and not b;
    layer4_outputs(5636) <= not a;
    layer4_outputs(5637) <= a and b;
    layer4_outputs(5638) <= b;
    layer4_outputs(5639) <= not (a or b);
    layer4_outputs(5640) <= 1'b0;
    layer4_outputs(5641) <= 1'b1;
    layer4_outputs(5642) <= a and not b;
    layer4_outputs(5643) <= not b or a;
    layer4_outputs(5644) <= a xor b;
    layer4_outputs(5645) <= not (a or b);
    layer4_outputs(5646) <= not b or a;
    layer4_outputs(5647) <= 1'b1;
    layer4_outputs(5648) <= 1'b1;
    layer4_outputs(5649) <= a and not b;
    layer4_outputs(5650) <= not (a or b);
    layer4_outputs(5651) <= not (a and b);
    layer4_outputs(5652) <= a and not b;
    layer4_outputs(5653) <= a;
    layer4_outputs(5654) <= not (a or b);
    layer4_outputs(5655) <= not a or b;
    layer4_outputs(5656) <= not a or b;
    layer4_outputs(5657) <= a;
    layer4_outputs(5658) <= not (a or b);
    layer4_outputs(5659) <= not b;
    layer4_outputs(5660) <= not b or a;
    layer4_outputs(5661) <= not b;
    layer4_outputs(5662) <= a or b;
    layer4_outputs(5663) <= not (a and b);
    layer4_outputs(5664) <= not b;
    layer4_outputs(5665) <= a;
    layer4_outputs(5666) <= a;
    layer4_outputs(5667) <= b and not a;
    layer4_outputs(5668) <= not b or a;
    layer4_outputs(5669) <= b;
    layer4_outputs(5670) <= not a;
    layer4_outputs(5671) <= b;
    layer4_outputs(5672) <= not (a or b);
    layer4_outputs(5673) <= 1'b1;
    layer4_outputs(5674) <= a;
    layer4_outputs(5675) <= b and not a;
    layer4_outputs(5676) <= not a or b;
    layer4_outputs(5677) <= a and b;
    layer4_outputs(5678) <= 1'b1;
    layer4_outputs(5679) <= not (a or b);
    layer4_outputs(5680) <= not (a and b);
    layer4_outputs(5681) <= 1'b1;
    layer4_outputs(5682) <= not b;
    layer4_outputs(5683) <= not a;
    layer4_outputs(5684) <= not a or b;
    layer4_outputs(5685) <= b and not a;
    layer4_outputs(5686) <= 1'b0;
    layer4_outputs(5687) <= not a;
    layer4_outputs(5688) <= a xor b;
    layer4_outputs(5689) <= 1'b1;
    layer4_outputs(5690) <= a;
    layer4_outputs(5691) <= not (a and b);
    layer4_outputs(5692) <= 1'b0;
    layer4_outputs(5693) <= a and not b;
    layer4_outputs(5694) <= not b or a;
    layer4_outputs(5695) <= not a;
    layer4_outputs(5696) <= not (a or b);
    layer4_outputs(5697) <= 1'b1;
    layer4_outputs(5698) <= b;
    layer4_outputs(5699) <= not a;
    layer4_outputs(5700) <= b and not a;
    layer4_outputs(5701) <= a;
    layer4_outputs(5702) <= not (a or b);
    layer4_outputs(5703) <= a and b;
    layer4_outputs(5704) <= not a or b;
    layer4_outputs(5705) <= not a;
    layer4_outputs(5706) <= 1'b1;
    layer4_outputs(5707) <= not b;
    layer4_outputs(5708) <= a and not b;
    layer4_outputs(5709) <= not a or b;
    layer4_outputs(5710) <= not a or b;
    layer4_outputs(5711) <= not (a or b);
    layer4_outputs(5712) <= not b or a;
    layer4_outputs(5713) <= not b;
    layer4_outputs(5714) <= not (a xor b);
    layer4_outputs(5715) <= a xor b;
    layer4_outputs(5716) <= a and b;
    layer4_outputs(5717) <= a and not b;
    layer4_outputs(5718) <= a or b;
    layer4_outputs(5719) <= not a or b;
    layer4_outputs(5720) <= 1'b0;
    layer4_outputs(5721) <= not b;
    layer4_outputs(5722) <= not b or a;
    layer4_outputs(5723) <= not a;
    layer4_outputs(5724) <= not b;
    layer4_outputs(5725) <= b;
    layer4_outputs(5726) <= not (a or b);
    layer4_outputs(5727) <= a;
    layer4_outputs(5728) <= b;
    layer4_outputs(5729) <= not b or a;
    layer4_outputs(5730) <= not (a or b);
    layer4_outputs(5731) <= a and b;
    layer4_outputs(5732) <= not (a and b);
    layer4_outputs(5733) <= b and not a;
    layer4_outputs(5734) <= not a or b;
    layer4_outputs(5735) <= not b or a;
    layer4_outputs(5736) <= not a;
    layer4_outputs(5737) <= not (a and b);
    layer4_outputs(5738) <= a and b;
    layer4_outputs(5739) <= a;
    layer4_outputs(5740) <= a;
    layer4_outputs(5741) <= not a or b;
    layer4_outputs(5742) <= b;
    layer4_outputs(5743) <= not (a and b);
    layer4_outputs(5744) <= a;
    layer4_outputs(5745) <= not b;
    layer4_outputs(5746) <= 1'b0;
    layer4_outputs(5747) <= not a or b;
    layer4_outputs(5748) <= b and not a;
    layer4_outputs(5749) <= not (a or b);
    layer4_outputs(5750) <= a;
    layer4_outputs(5751) <= not a;
    layer4_outputs(5752) <= not a or b;
    layer4_outputs(5753) <= a;
    layer4_outputs(5754) <= a and b;
    layer4_outputs(5755) <= 1'b0;
    layer4_outputs(5756) <= b and not a;
    layer4_outputs(5757) <= b and not a;
    layer4_outputs(5758) <= b and not a;
    layer4_outputs(5759) <= not a;
    layer4_outputs(5760) <= not (a and b);
    layer4_outputs(5761) <= not (a or b);
    layer4_outputs(5762) <= not a or b;
    layer4_outputs(5763) <= not (a and b);
    layer4_outputs(5764) <= not a or b;
    layer4_outputs(5765) <= 1'b1;
    layer4_outputs(5766) <= 1'b0;
    layer4_outputs(5767) <= a and not b;
    layer4_outputs(5768) <= 1'b0;
    layer4_outputs(5769) <= b and not a;
    layer4_outputs(5770) <= a and b;
    layer4_outputs(5771) <= a and b;
    layer4_outputs(5772) <= not (a and b);
    layer4_outputs(5773) <= not (a xor b);
    layer4_outputs(5774) <= not (a and b);
    layer4_outputs(5775) <= not (a or b);
    layer4_outputs(5776) <= 1'b0;
    layer4_outputs(5777) <= not b or a;
    layer4_outputs(5778) <= 1'b0;
    layer4_outputs(5779) <= not a;
    layer4_outputs(5780) <= not b or a;
    layer4_outputs(5781) <= a or b;
    layer4_outputs(5782) <= not (a and b);
    layer4_outputs(5783) <= not b;
    layer4_outputs(5784) <= a or b;
    layer4_outputs(5785) <= not a;
    layer4_outputs(5786) <= not (a or b);
    layer4_outputs(5787) <= not (a and b);
    layer4_outputs(5788) <= a and b;
    layer4_outputs(5789) <= 1'b0;
    layer4_outputs(5790) <= not b or a;
    layer4_outputs(5791) <= not b;
    layer4_outputs(5792) <= not (a and b);
    layer4_outputs(5793) <= a xor b;
    layer4_outputs(5794) <= a;
    layer4_outputs(5795) <= 1'b1;
    layer4_outputs(5796) <= 1'b0;
    layer4_outputs(5797) <= 1'b1;
    layer4_outputs(5798) <= a and not b;
    layer4_outputs(5799) <= b;
    layer4_outputs(5800) <= not a or b;
    layer4_outputs(5801) <= a or b;
    layer4_outputs(5802) <= not (a or b);
    layer4_outputs(5803) <= 1'b1;
    layer4_outputs(5804) <= 1'b0;
    layer4_outputs(5805) <= 1'b1;
    layer4_outputs(5806) <= not (a xor b);
    layer4_outputs(5807) <= a xor b;
    layer4_outputs(5808) <= 1'b1;
    layer4_outputs(5809) <= 1'b0;
    layer4_outputs(5810) <= a or b;
    layer4_outputs(5811) <= not b or a;
    layer4_outputs(5812) <= not a;
    layer4_outputs(5813) <= not b or a;
    layer4_outputs(5814) <= b;
    layer4_outputs(5815) <= b;
    layer4_outputs(5816) <= not a;
    layer4_outputs(5817) <= b and not a;
    layer4_outputs(5818) <= not a;
    layer4_outputs(5819) <= not a;
    layer4_outputs(5820) <= a or b;
    layer4_outputs(5821) <= not a or b;
    layer4_outputs(5822) <= a;
    layer4_outputs(5823) <= a or b;
    layer4_outputs(5824) <= a;
    layer4_outputs(5825) <= 1'b0;
    layer4_outputs(5826) <= b and not a;
    layer4_outputs(5827) <= a xor b;
    layer4_outputs(5828) <= b;
    layer4_outputs(5829) <= a and b;
    layer4_outputs(5830) <= not b;
    layer4_outputs(5831) <= a and not b;
    layer4_outputs(5832) <= 1'b0;
    layer4_outputs(5833) <= a and not b;
    layer4_outputs(5834) <= a xor b;
    layer4_outputs(5835) <= a;
    layer4_outputs(5836) <= not (a and b);
    layer4_outputs(5837) <= a;
    layer4_outputs(5838) <= not a;
    layer4_outputs(5839) <= not (a or b);
    layer4_outputs(5840) <= not b or a;
    layer4_outputs(5841) <= 1'b1;
    layer4_outputs(5842) <= not b;
    layer4_outputs(5843) <= a and not b;
    layer4_outputs(5844) <= a and b;
    layer4_outputs(5845) <= a and not b;
    layer4_outputs(5846) <= 1'b1;
    layer4_outputs(5847) <= not b or a;
    layer4_outputs(5848) <= not (a or b);
    layer4_outputs(5849) <= a or b;
    layer4_outputs(5850) <= not b or a;
    layer4_outputs(5851) <= 1'b0;
    layer4_outputs(5852) <= not b;
    layer4_outputs(5853) <= not a;
    layer4_outputs(5854) <= not b;
    layer4_outputs(5855) <= b and not a;
    layer4_outputs(5856) <= 1'b0;
    layer4_outputs(5857) <= b;
    layer4_outputs(5858) <= not a;
    layer4_outputs(5859) <= not (a and b);
    layer4_outputs(5860) <= 1'b1;
    layer4_outputs(5861) <= not a or b;
    layer4_outputs(5862) <= not (a or b);
    layer4_outputs(5863) <= b and not a;
    layer4_outputs(5864) <= b;
    layer4_outputs(5865) <= not a or b;
    layer4_outputs(5866) <= b and not a;
    layer4_outputs(5867) <= 1'b0;
    layer4_outputs(5868) <= 1'b0;
    layer4_outputs(5869) <= b;
    layer4_outputs(5870) <= not (a or b);
    layer4_outputs(5871) <= 1'b0;
    layer4_outputs(5872) <= a or b;
    layer4_outputs(5873) <= not b;
    layer4_outputs(5874) <= not b;
    layer4_outputs(5875) <= not (a and b);
    layer4_outputs(5876) <= not a;
    layer4_outputs(5877) <= a;
    layer4_outputs(5878) <= b;
    layer4_outputs(5879) <= 1'b0;
    layer4_outputs(5880) <= not (a and b);
    layer4_outputs(5881) <= not (a and b);
    layer4_outputs(5882) <= b and not a;
    layer4_outputs(5883) <= not b;
    layer4_outputs(5884) <= not a;
    layer4_outputs(5885) <= a and not b;
    layer4_outputs(5886) <= a xor b;
    layer4_outputs(5887) <= a or b;
    layer4_outputs(5888) <= 1'b0;
    layer4_outputs(5889) <= a or b;
    layer4_outputs(5890) <= not a or b;
    layer4_outputs(5891) <= not a or b;
    layer4_outputs(5892) <= 1'b0;
    layer4_outputs(5893) <= not b;
    layer4_outputs(5894) <= not (a and b);
    layer4_outputs(5895) <= not (a or b);
    layer4_outputs(5896) <= 1'b1;
    layer4_outputs(5897) <= a;
    layer4_outputs(5898) <= a xor b;
    layer4_outputs(5899) <= not a;
    layer4_outputs(5900) <= 1'b0;
    layer4_outputs(5901) <= not a;
    layer4_outputs(5902) <= not a;
    layer4_outputs(5903) <= not (a and b);
    layer4_outputs(5904) <= not a or b;
    layer4_outputs(5905) <= a and b;
    layer4_outputs(5906) <= b;
    layer4_outputs(5907) <= not b;
    layer4_outputs(5908) <= a;
    layer4_outputs(5909) <= not b;
    layer4_outputs(5910) <= b and not a;
    layer4_outputs(5911) <= not b or a;
    layer4_outputs(5912) <= b and not a;
    layer4_outputs(5913) <= not b;
    layer4_outputs(5914) <= not (a and b);
    layer4_outputs(5915) <= 1'b0;
    layer4_outputs(5916) <= not (a xor b);
    layer4_outputs(5917) <= not (a or b);
    layer4_outputs(5918) <= not b or a;
    layer4_outputs(5919) <= a;
    layer4_outputs(5920) <= b;
    layer4_outputs(5921) <= 1'b0;
    layer4_outputs(5922) <= a;
    layer4_outputs(5923) <= not (a xor b);
    layer4_outputs(5924) <= a and not b;
    layer4_outputs(5925) <= not a;
    layer4_outputs(5926) <= b;
    layer4_outputs(5927) <= a;
    layer4_outputs(5928) <= a and b;
    layer4_outputs(5929) <= not b or a;
    layer4_outputs(5930) <= b;
    layer4_outputs(5931) <= a;
    layer4_outputs(5932) <= a;
    layer4_outputs(5933) <= not (a and b);
    layer4_outputs(5934) <= not b or a;
    layer4_outputs(5935) <= 1'b0;
    layer4_outputs(5936) <= not a;
    layer4_outputs(5937) <= a;
    layer4_outputs(5938) <= 1'b1;
    layer4_outputs(5939) <= not (a or b);
    layer4_outputs(5940) <= b and not a;
    layer4_outputs(5941) <= a or b;
    layer4_outputs(5942) <= not b;
    layer4_outputs(5943) <= b;
    layer4_outputs(5944) <= a;
    layer4_outputs(5945) <= not (a and b);
    layer4_outputs(5946) <= 1'b1;
    layer4_outputs(5947) <= b;
    layer4_outputs(5948) <= not a or b;
    layer4_outputs(5949) <= 1'b0;
    layer4_outputs(5950) <= a or b;
    layer4_outputs(5951) <= b and not a;
    layer4_outputs(5952) <= b;
    layer4_outputs(5953) <= not b or a;
    layer4_outputs(5954) <= not (a and b);
    layer4_outputs(5955) <= a xor b;
    layer4_outputs(5956) <= not a;
    layer4_outputs(5957) <= 1'b1;
    layer4_outputs(5958) <= not a or b;
    layer4_outputs(5959) <= a or b;
    layer4_outputs(5960) <= not b or a;
    layer4_outputs(5961) <= a and b;
    layer4_outputs(5962) <= a and not b;
    layer4_outputs(5963) <= not b;
    layer4_outputs(5964) <= not b;
    layer4_outputs(5965) <= not (a and b);
    layer4_outputs(5966) <= not (a or b);
    layer4_outputs(5967) <= a;
    layer4_outputs(5968) <= not b or a;
    layer4_outputs(5969) <= not (a or b);
    layer4_outputs(5970) <= not a;
    layer4_outputs(5971) <= not a or b;
    layer4_outputs(5972) <= not a or b;
    layer4_outputs(5973) <= a and b;
    layer4_outputs(5974) <= a and b;
    layer4_outputs(5975) <= 1'b0;
    layer4_outputs(5976) <= not b;
    layer4_outputs(5977) <= not a or b;
    layer4_outputs(5978) <= not a or b;
    layer4_outputs(5979) <= not a;
    layer4_outputs(5980) <= not a or b;
    layer4_outputs(5981) <= 1'b1;
    layer4_outputs(5982) <= not a;
    layer4_outputs(5983) <= a and b;
    layer4_outputs(5984) <= not (a and b);
    layer4_outputs(5985) <= b;
    layer4_outputs(5986) <= a;
    layer4_outputs(5987) <= not (a or b);
    layer4_outputs(5988) <= not (a and b);
    layer4_outputs(5989) <= 1'b0;
    layer4_outputs(5990) <= not b or a;
    layer4_outputs(5991) <= not a;
    layer4_outputs(5992) <= not b;
    layer4_outputs(5993) <= b and not a;
    layer4_outputs(5994) <= not a or b;
    layer4_outputs(5995) <= a and not b;
    layer4_outputs(5996) <= a;
    layer4_outputs(5997) <= b and not a;
    layer4_outputs(5998) <= 1'b0;
    layer4_outputs(5999) <= not a;
    layer4_outputs(6000) <= not a;
    layer4_outputs(6001) <= a or b;
    layer4_outputs(6002) <= not a or b;
    layer4_outputs(6003) <= b and not a;
    layer4_outputs(6004) <= b;
    layer4_outputs(6005) <= not b;
    layer4_outputs(6006) <= b;
    layer4_outputs(6007) <= not a or b;
    layer4_outputs(6008) <= a and not b;
    layer4_outputs(6009) <= a and b;
    layer4_outputs(6010) <= a;
    layer4_outputs(6011) <= b and not a;
    layer4_outputs(6012) <= not a or b;
    layer4_outputs(6013) <= not (a and b);
    layer4_outputs(6014) <= a and not b;
    layer4_outputs(6015) <= not a;
    layer4_outputs(6016) <= not b;
    layer4_outputs(6017) <= not a or b;
    layer4_outputs(6018) <= b;
    layer4_outputs(6019) <= not b or a;
    layer4_outputs(6020) <= a xor b;
    layer4_outputs(6021) <= 1'b1;
    layer4_outputs(6022) <= a and b;
    layer4_outputs(6023) <= not (a xor b);
    layer4_outputs(6024) <= b;
    layer4_outputs(6025) <= not (a and b);
    layer4_outputs(6026) <= b;
    layer4_outputs(6027) <= not b or a;
    layer4_outputs(6028) <= not a;
    layer4_outputs(6029) <= not b;
    layer4_outputs(6030) <= not a;
    layer4_outputs(6031) <= not b;
    layer4_outputs(6032) <= not b;
    layer4_outputs(6033) <= not a or b;
    layer4_outputs(6034) <= not (a and b);
    layer4_outputs(6035) <= not a or b;
    layer4_outputs(6036) <= 1'b0;
    layer4_outputs(6037) <= not (a xor b);
    layer4_outputs(6038) <= a or b;
    layer4_outputs(6039) <= a and not b;
    layer4_outputs(6040) <= a and not b;
    layer4_outputs(6041) <= 1'b0;
    layer4_outputs(6042) <= b and not a;
    layer4_outputs(6043) <= a;
    layer4_outputs(6044) <= not (a and b);
    layer4_outputs(6045) <= b;
    layer4_outputs(6046) <= not a or b;
    layer4_outputs(6047) <= not b or a;
    layer4_outputs(6048) <= a;
    layer4_outputs(6049) <= not (a xor b);
    layer4_outputs(6050) <= not (a or b);
    layer4_outputs(6051) <= a and b;
    layer4_outputs(6052) <= not b;
    layer4_outputs(6053) <= not b or a;
    layer4_outputs(6054) <= not (a or b);
    layer4_outputs(6055) <= b and not a;
    layer4_outputs(6056) <= a or b;
    layer4_outputs(6057) <= b;
    layer4_outputs(6058) <= not b;
    layer4_outputs(6059) <= not b or a;
    layer4_outputs(6060) <= a;
    layer4_outputs(6061) <= a and not b;
    layer4_outputs(6062) <= a or b;
    layer4_outputs(6063) <= a and b;
    layer4_outputs(6064) <= not b or a;
    layer4_outputs(6065) <= not (a xor b);
    layer4_outputs(6066) <= not (a xor b);
    layer4_outputs(6067) <= not b;
    layer4_outputs(6068) <= not a or b;
    layer4_outputs(6069) <= a and not b;
    layer4_outputs(6070) <= a;
    layer4_outputs(6071) <= b;
    layer4_outputs(6072) <= 1'b1;
    layer4_outputs(6073) <= not b;
    layer4_outputs(6074) <= a;
    layer4_outputs(6075) <= a or b;
    layer4_outputs(6076) <= not b;
    layer4_outputs(6077) <= not (a or b);
    layer4_outputs(6078) <= not (a and b);
    layer4_outputs(6079) <= not a or b;
    layer4_outputs(6080) <= not b or a;
    layer4_outputs(6081) <= a xor b;
    layer4_outputs(6082) <= a and not b;
    layer4_outputs(6083) <= 1'b0;
    layer4_outputs(6084) <= 1'b1;
    layer4_outputs(6085) <= a and b;
    layer4_outputs(6086) <= 1'b0;
    layer4_outputs(6087) <= not (a or b);
    layer4_outputs(6088) <= a and b;
    layer4_outputs(6089) <= a and not b;
    layer4_outputs(6090) <= not (a or b);
    layer4_outputs(6091) <= not a or b;
    layer4_outputs(6092) <= not a;
    layer4_outputs(6093) <= a;
    layer4_outputs(6094) <= 1'b1;
    layer4_outputs(6095) <= a;
    layer4_outputs(6096) <= b;
    layer4_outputs(6097) <= a;
    layer4_outputs(6098) <= b and not a;
    layer4_outputs(6099) <= 1'b0;
    layer4_outputs(6100) <= a xor b;
    layer4_outputs(6101) <= b;
    layer4_outputs(6102) <= not (a xor b);
    layer4_outputs(6103) <= b;
    layer4_outputs(6104) <= not b or a;
    layer4_outputs(6105) <= a and not b;
    layer4_outputs(6106) <= not a;
    layer4_outputs(6107) <= not (a xor b);
    layer4_outputs(6108) <= a;
    layer4_outputs(6109) <= a or b;
    layer4_outputs(6110) <= a;
    layer4_outputs(6111) <= 1'b0;
    layer4_outputs(6112) <= not (a xor b);
    layer4_outputs(6113) <= a or b;
    layer4_outputs(6114) <= 1'b1;
    layer4_outputs(6115) <= not (a and b);
    layer4_outputs(6116) <= not b or a;
    layer4_outputs(6117) <= a;
    layer4_outputs(6118) <= not b or a;
    layer4_outputs(6119) <= not (a xor b);
    layer4_outputs(6120) <= 1'b0;
    layer4_outputs(6121) <= a xor b;
    layer4_outputs(6122) <= not (a or b);
    layer4_outputs(6123) <= 1'b1;
    layer4_outputs(6124) <= not a;
    layer4_outputs(6125) <= not (a or b);
    layer4_outputs(6126) <= b;
    layer4_outputs(6127) <= a;
    layer4_outputs(6128) <= not a;
    layer4_outputs(6129) <= 1'b0;
    layer4_outputs(6130) <= not a;
    layer4_outputs(6131) <= a and not b;
    layer4_outputs(6132) <= a or b;
    layer4_outputs(6133) <= a and b;
    layer4_outputs(6134) <= 1'b0;
    layer4_outputs(6135) <= not a or b;
    layer4_outputs(6136) <= not a or b;
    layer4_outputs(6137) <= not (a and b);
    layer4_outputs(6138) <= not b;
    layer4_outputs(6139) <= b;
    layer4_outputs(6140) <= a and b;
    layer4_outputs(6141) <= not b;
    layer4_outputs(6142) <= not (a and b);
    layer4_outputs(6143) <= not (a xor b);
    layer4_outputs(6144) <= 1'b0;
    layer4_outputs(6145) <= b and not a;
    layer4_outputs(6146) <= a;
    layer4_outputs(6147) <= a and b;
    layer4_outputs(6148) <= a or b;
    layer4_outputs(6149) <= a or b;
    layer4_outputs(6150) <= b;
    layer4_outputs(6151) <= b and not a;
    layer4_outputs(6152) <= a or b;
    layer4_outputs(6153) <= a and b;
    layer4_outputs(6154) <= not (a or b);
    layer4_outputs(6155) <= not (a xor b);
    layer4_outputs(6156) <= not (a or b);
    layer4_outputs(6157) <= a and not b;
    layer4_outputs(6158) <= a;
    layer4_outputs(6159) <= a or b;
    layer4_outputs(6160) <= b and not a;
    layer4_outputs(6161) <= 1'b1;
    layer4_outputs(6162) <= not a or b;
    layer4_outputs(6163) <= a;
    layer4_outputs(6164) <= not a;
    layer4_outputs(6165) <= not b or a;
    layer4_outputs(6166) <= a;
    layer4_outputs(6167) <= not b;
    layer4_outputs(6168) <= 1'b1;
    layer4_outputs(6169) <= not (a or b);
    layer4_outputs(6170) <= 1'b0;
    layer4_outputs(6171) <= not b;
    layer4_outputs(6172) <= b;
    layer4_outputs(6173) <= b and not a;
    layer4_outputs(6174) <= a;
    layer4_outputs(6175) <= b;
    layer4_outputs(6176) <= not a or b;
    layer4_outputs(6177) <= not a or b;
    layer4_outputs(6178) <= a and b;
    layer4_outputs(6179) <= not b or a;
    layer4_outputs(6180) <= a;
    layer4_outputs(6181) <= not (a or b);
    layer4_outputs(6182) <= a and not b;
    layer4_outputs(6183) <= not b;
    layer4_outputs(6184) <= not (a or b);
    layer4_outputs(6185) <= b and not a;
    layer4_outputs(6186) <= not a or b;
    layer4_outputs(6187) <= a and b;
    layer4_outputs(6188) <= not b or a;
    layer4_outputs(6189) <= a and b;
    layer4_outputs(6190) <= b;
    layer4_outputs(6191) <= 1'b0;
    layer4_outputs(6192) <= not b;
    layer4_outputs(6193) <= not (a or b);
    layer4_outputs(6194) <= a xor b;
    layer4_outputs(6195) <= not b or a;
    layer4_outputs(6196) <= not a;
    layer4_outputs(6197) <= not a or b;
    layer4_outputs(6198) <= b;
    layer4_outputs(6199) <= a or b;
    layer4_outputs(6200) <= a;
    layer4_outputs(6201) <= not (a or b);
    layer4_outputs(6202) <= 1'b1;
    layer4_outputs(6203) <= b and not a;
    layer4_outputs(6204) <= a;
    layer4_outputs(6205) <= 1'b1;
    layer4_outputs(6206) <= a or b;
    layer4_outputs(6207) <= b and not a;
    layer4_outputs(6208) <= 1'b0;
    layer4_outputs(6209) <= not b;
    layer4_outputs(6210) <= a and not b;
    layer4_outputs(6211) <= b;
    layer4_outputs(6212) <= a;
    layer4_outputs(6213) <= a;
    layer4_outputs(6214) <= not b;
    layer4_outputs(6215) <= b and not a;
    layer4_outputs(6216) <= a and not b;
    layer4_outputs(6217) <= a and not b;
    layer4_outputs(6218) <= not (a xor b);
    layer4_outputs(6219) <= a or b;
    layer4_outputs(6220) <= not b;
    layer4_outputs(6221) <= 1'b0;
    layer4_outputs(6222) <= not (a or b);
    layer4_outputs(6223) <= a or b;
    layer4_outputs(6224) <= not a or b;
    layer4_outputs(6225) <= b and not a;
    layer4_outputs(6226) <= not (a or b);
    layer4_outputs(6227) <= not (a and b);
    layer4_outputs(6228) <= not (a and b);
    layer4_outputs(6229) <= b and not a;
    layer4_outputs(6230) <= a and not b;
    layer4_outputs(6231) <= not a or b;
    layer4_outputs(6232) <= a;
    layer4_outputs(6233) <= a and not b;
    layer4_outputs(6234) <= not (a and b);
    layer4_outputs(6235) <= not b;
    layer4_outputs(6236) <= a;
    layer4_outputs(6237) <= not a;
    layer4_outputs(6238) <= b;
    layer4_outputs(6239) <= b;
    layer4_outputs(6240) <= not b or a;
    layer4_outputs(6241) <= not a;
    layer4_outputs(6242) <= not b or a;
    layer4_outputs(6243) <= not a;
    layer4_outputs(6244) <= not b;
    layer4_outputs(6245) <= not (a or b);
    layer4_outputs(6246) <= not (a and b);
    layer4_outputs(6247) <= b;
    layer4_outputs(6248) <= not a;
    layer4_outputs(6249) <= a and not b;
    layer4_outputs(6250) <= not b or a;
    layer4_outputs(6251) <= b and not a;
    layer4_outputs(6252) <= a;
    layer4_outputs(6253) <= 1'b1;
    layer4_outputs(6254) <= 1'b1;
    layer4_outputs(6255) <= not a or b;
    layer4_outputs(6256) <= not a or b;
    layer4_outputs(6257) <= a or b;
    layer4_outputs(6258) <= not a or b;
    layer4_outputs(6259) <= not b;
    layer4_outputs(6260) <= a and b;
    layer4_outputs(6261) <= not (a or b);
    layer4_outputs(6262) <= not a;
    layer4_outputs(6263) <= not (a or b);
    layer4_outputs(6264) <= not (a or b);
    layer4_outputs(6265) <= b;
    layer4_outputs(6266) <= a xor b;
    layer4_outputs(6267) <= a and b;
    layer4_outputs(6268) <= not a or b;
    layer4_outputs(6269) <= 1'b1;
    layer4_outputs(6270) <= b and not a;
    layer4_outputs(6271) <= not (a and b);
    layer4_outputs(6272) <= not b or a;
    layer4_outputs(6273) <= b;
    layer4_outputs(6274) <= a and b;
    layer4_outputs(6275) <= a xor b;
    layer4_outputs(6276) <= a or b;
    layer4_outputs(6277) <= a or b;
    layer4_outputs(6278) <= a xor b;
    layer4_outputs(6279) <= not a or b;
    layer4_outputs(6280) <= not b or a;
    layer4_outputs(6281) <= a and not b;
    layer4_outputs(6282) <= 1'b0;
    layer4_outputs(6283) <= a;
    layer4_outputs(6284) <= not b or a;
    layer4_outputs(6285) <= not b;
    layer4_outputs(6286) <= not (a or b);
    layer4_outputs(6287) <= a and not b;
    layer4_outputs(6288) <= not b;
    layer4_outputs(6289) <= a or b;
    layer4_outputs(6290) <= a and b;
    layer4_outputs(6291) <= b and not a;
    layer4_outputs(6292) <= not (a or b);
    layer4_outputs(6293) <= 1'b1;
    layer4_outputs(6294) <= b;
    layer4_outputs(6295) <= not b;
    layer4_outputs(6296) <= a or b;
    layer4_outputs(6297) <= not b;
    layer4_outputs(6298) <= not (a and b);
    layer4_outputs(6299) <= not a or b;
    layer4_outputs(6300) <= a;
    layer4_outputs(6301) <= not (a and b);
    layer4_outputs(6302) <= b;
    layer4_outputs(6303) <= not (a or b);
    layer4_outputs(6304) <= not (a xor b);
    layer4_outputs(6305) <= not a or b;
    layer4_outputs(6306) <= a;
    layer4_outputs(6307) <= a;
    layer4_outputs(6308) <= not a or b;
    layer4_outputs(6309) <= not (a or b);
    layer4_outputs(6310) <= not a or b;
    layer4_outputs(6311) <= not b;
    layer4_outputs(6312) <= not (a and b);
    layer4_outputs(6313) <= a and b;
    layer4_outputs(6314) <= b and not a;
    layer4_outputs(6315) <= 1'b0;
    layer4_outputs(6316) <= b and not a;
    layer4_outputs(6317) <= b;
    layer4_outputs(6318) <= not a;
    layer4_outputs(6319) <= a and not b;
    layer4_outputs(6320) <= 1'b1;
    layer4_outputs(6321) <= a and b;
    layer4_outputs(6322) <= not b;
    layer4_outputs(6323) <= a and not b;
    layer4_outputs(6324) <= not b or a;
    layer4_outputs(6325) <= not a or b;
    layer4_outputs(6326) <= a and not b;
    layer4_outputs(6327) <= a or b;
    layer4_outputs(6328) <= not a;
    layer4_outputs(6329) <= b;
    layer4_outputs(6330) <= 1'b1;
    layer4_outputs(6331) <= a and not b;
    layer4_outputs(6332) <= 1'b0;
    layer4_outputs(6333) <= not a or b;
    layer4_outputs(6334) <= b;
    layer4_outputs(6335) <= b;
    layer4_outputs(6336) <= not a or b;
    layer4_outputs(6337) <= not b or a;
    layer4_outputs(6338) <= a or b;
    layer4_outputs(6339) <= not (a or b);
    layer4_outputs(6340) <= not a or b;
    layer4_outputs(6341) <= a and not b;
    layer4_outputs(6342) <= not b or a;
    layer4_outputs(6343) <= not b or a;
    layer4_outputs(6344) <= not (a and b);
    layer4_outputs(6345) <= not b;
    layer4_outputs(6346) <= not (a or b);
    layer4_outputs(6347) <= not b;
    layer4_outputs(6348) <= not b or a;
    layer4_outputs(6349) <= not b;
    layer4_outputs(6350) <= not (a or b);
    layer4_outputs(6351) <= a and not b;
    layer4_outputs(6352) <= a and b;
    layer4_outputs(6353) <= not b;
    layer4_outputs(6354) <= not a or b;
    layer4_outputs(6355) <= not (a and b);
    layer4_outputs(6356) <= b;
    layer4_outputs(6357) <= not b;
    layer4_outputs(6358) <= a;
    layer4_outputs(6359) <= not (a or b);
    layer4_outputs(6360) <= not b or a;
    layer4_outputs(6361) <= a or b;
    layer4_outputs(6362) <= not (a or b);
    layer4_outputs(6363) <= not a or b;
    layer4_outputs(6364) <= b and not a;
    layer4_outputs(6365) <= a and b;
    layer4_outputs(6366) <= not b;
    layer4_outputs(6367) <= not b;
    layer4_outputs(6368) <= not (a xor b);
    layer4_outputs(6369) <= a;
    layer4_outputs(6370) <= 1'b1;
    layer4_outputs(6371) <= not a;
    layer4_outputs(6372) <= a or b;
    layer4_outputs(6373) <= not a;
    layer4_outputs(6374) <= a;
    layer4_outputs(6375) <= a or b;
    layer4_outputs(6376) <= a;
    layer4_outputs(6377) <= a;
    layer4_outputs(6378) <= not a or b;
    layer4_outputs(6379) <= not (a or b);
    layer4_outputs(6380) <= not b;
    layer4_outputs(6381) <= not a;
    layer4_outputs(6382) <= not b;
    layer4_outputs(6383) <= not a or b;
    layer4_outputs(6384) <= a and not b;
    layer4_outputs(6385) <= not b;
    layer4_outputs(6386) <= not b or a;
    layer4_outputs(6387) <= a or b;
    layer4_outputs(6388) <= a and not b;
    layer4_outputs(6389) <= a or b;
    layer4_outputs(6390) <= b and not a;
    layer4_outputs(6391) <= a and b;
    layer4_outputs(6392) <= b;
    layer4_outputs(6393) <= a xor b;
    layer4_outputs(6394) <= not (a and b);
    layer4_outputs(6395) <= not a or b;
    layer4_outputs(6396) <= b;
    layer4_outputs(6397) <= not (a and b);
    layer4_outputs(6398) <= not (a and b);
    layer4_outputs(6399) <= not a or b;
    layer4_outputs(6400) <= a and b;
    layer4_outputs(6401) <= not a or b;
    layer4_outputs(6402) <= a or b;
    layer4_outputs(6403) <= not a;
    layer4_outputs(6404) <= b;
    layer4_outputs(6405) <= a or b;
    layer4_outputs(6406) <= not a or b;
    layer4_outputs(6407) <= a and b;
    layer4_outputs(6408) <= b and not a;
    layer4_outputs(6409) <= not a or b;
    layer4_outputs(6410) <= a xor b;
    layer4_outputs(6411) <= not a or b;
    layer4_outputs(6412) <= not a or b;
    layer4_outputs(6413) <= not a;
    layer4_outputs(6414) <= not (a or b);
    layer4_outputs(6415) <= b;
    layer4_outputs(6416) <= not (a or b);
    layer4_outputs(6417) <= not (a xor b);
    layer4_outputs(6418) <= a and not b;
    layer4_outputs(6419) <= a and not b;
    layer4_outputs(6420) <= 1'b0;
    layer4_outputs(6421) <= not a or b;
    layer4_outputs(6422) <= 1'b1;
    layer4_outputs(6423) <= 1'b1;
    layer4_outputs(6424) <= a or b;
    layer4_outputs(6425) <= not a;
    layer4_outputs(6426) <= b and not a;
    layer4_outputs(6427) <= not b or a;
    layer4_outputs(6428) <= a and b;
    layer4_outputs(6429) <= b;
    layer4_outputs(6430) <= a;
    layer4_outputs(6431) <= b;
    layer4_outputs(6432) <= b;
    layer4_outputs(6433) <= b;
    layer4_outputs(6434) <= b and not a;
    layer4_outputs(6435) <= a and not b;
    layer4_outputs(6436) <= a or b;
    layer4_outputs(6437) <= a or b;
    layer4_outputs(6438) <= b;
    layer4_outputs(6439) <= not (a or b);
    layer4_outputs(6440) <= a or b;
    layer4_outputs(6441) <= a and b;
    layer4_outputs(6442) <= a or b;
    layer4_outputs(6443) <= a or b;
    layer4_outputs(6444) <= not (a xor b);
    layer4_outputs(6445) <= 1'b1;
    layer4_outputs(6446) <= a;
    layer4_outputs(6447) <= a;
    layer4_outputs(6448) <= 1'b0;
    layer4_outputs(6449) <= a and not b;
    layer4_outputs(6450) <= b and not a;
    layer4_outputs(6451) <= not a;
    layer4_outputs(6452) <= a and not b;
    layer4_outputs(6453) <= a and not b;
    layer4_outputs(6454) <= not (a xor b);
    layer4_outputs(6455) <= b and not a;
    layer4_outputs(6456) <= not b;
    layer4_outputs(6457) <= 1'b1;
    layer4_outputs(6458) <= not b or a;
    layer4_outputs(6459) <= a and b;
    layer4_outputs(6460) <= not b;
    layer4_outputs(6461) <= a and b;
    layer4_outputs(6462) <= not a or b;
    layer4_outputs(6463) <= a;
    layer4_outputs(6464) <= not a or b;
    layer4_outputs(6465) <= b;
    layer4_outputs(6466) <= 1'b0;
    layer4_outputs(6467) <= not (a xor b);
    layer4_outputs(6468) <= a and b;
    layer4_outputs(6469) <= b;
    layer4_outputs(6470) <= not a or b;
    layer4_outputs(6471) <= not (a or b);
    layer4_outputs(6472) <= not a;
    layer4_outputs(6473) <= not a or b;
    layer4_outputs(6474) <= a and b;
    layer4_outputs(6475) <= a and b;
    layer4_outputs(6476) <= a;
    layer4_outputs(6477) <= b and not a;
    layer4_outputs(6478) <= not b or a;
    layer4_outputs(6479) <= not b;
    layer4_outputs(6480) <= a and b;
    layer4_outputs(6481) <= not b or a;
    layer4_outputs(6482) <= not b;
    layer4_outputs(6483) <= not (a and b);
    layer4_outputs(6484) <= 1'b1;
    layer4_outputs(6485) <= b and not a;
    layer4_outputs(6486) <= a or b;
    layer4_outputs(6487) <= not b;
    layer4_outputs(6488) <= 1'b1;
    layer4_outputs(6489) <= 1'b1;
    layer4_outputs(6490) <= 1'b0;
    layer4_outputs(6491) <= not a or b;
    layer4_outputs(6492) <= not b or a;
    layer4_outputs(6493) <= b and not a;
    layer4_outputs(6494) <= a or b;
    layer4_outputs(6495) <= not b;
    layer4_outputs(6496) <= b;
    layer4_outputs(6497) <= a;
    layer4_outputs(6498) <= not (a or b);
    layer4_outputs(6499) <= a;
    layer4_outputs(6500) <= not a;
    layer4_outputs(6501) <= a;
    layer4_outputs(6502) <= a xor b;
    layer4_outputs(6503) <= not b or a;
    layer4_outputs(6504) <= a;
    layer4_outputs(6505) <= b and not a;
    layer4_outputs(6506) <= a and b;
    layer4_outputs(6507) <= a;
    layer4_outputs(6508) <= not (a and b);
    layer4_outputs(6509) <= a xor b;
    layer4_outputs(6510) <= 1'b1;
    layer4_outputs(6511) <= a or b;
    layer4_outputs(6512) <= 1'b0;
    layer4_outputs(6513) <= a or b;
    layer4_outputs(6514) <= not a or b;
    layer4_outputs(6515) <= b;
    layer4_outputs(6516) <= not (a xor b);
    layer4_outputs(6517) <= not (a xor b);
    layer4_outputs(6518) <= a and b;
    layer4_outputs(6519) <= a;
    layer4_outputs(6520) <= 1'b0;
    layer4_outputs(6521) <= not a or b;
    layer4_outputs(6522) <= not a;
    layer4_outputs(6523) <= a and not b;
    layer4_outputs(6524) <= not (a or b);
    layer4_outputs(6525) <= not a or b;
    layer4_outputs(6526) <= not b or a;
    layer4_outputs(6527) <= 1'b0;
    layer4_outputs(6528) <= b;
    layer4_outputs(6529) <= a;
    layer4_outputs(6530) <= a and not b;
    layer4_outputs(6531) <= not a;
    layer4_outputs(6532) <= b and not a;
    layer4_outputs(6533) <= b;
    layer4_outputs(6534) <= not a or b;
    layer4_outputs(6535) <= 1'b1;
    layer4_outputs(6536) <= a xor b;
    layer4_outputs(6537) <= a and not b;
    layer4_outputs(6538) <= 1'b1;
    layer4_outputs(6539) <= 1'b1;
    layer4_outputs(6540) <= not a;
    layer4_outputs(6541) <= not (a or b);
    layer4_outputs(6542) <= b;
    layer4_outputs(6543) <= not (a and b);
    layer4_outputs(6544) <= a and not b;
    layer4_outputs(6545) <= a or b;
    layer4_outputs(6546) <= 1'b1;
    layer4_outputs(6547) <= not a;
    layer4_outputs(6548) <= 1'b1;
    layer4_outputs(6549) <= not a or b;
    layer4_outputs(6550) <= 1'b1;
    layer4_outputs(6551) <= b;
    layer4_outputs(6552) <= a and b;
    layer4_outputs(6553) <= not (a or b);
    layer4_outputs(6554) <= not (a or b);
    layer4_outputs(6555) <= a xor b;
    layer4_outputs(6556) <= not a or b;
    layer4_outputs(6557) <= not b;
    layer4_outputs(6558) <= a and not b;
    layer4_outputs(6559) <= 1'b1;
    layer4_outputs(6560) <= not b;
    layer4_outputs(6561) <= a or b;
    layer4_outputs(6562) <= b and not a;
    layer4_outputs(6563) <= a and not b;
    layer4_outputs(6564) <= not a or b;
    layer4_outputs(6565) <= not (a and b);
    layer4_outputs(6566) <= not a or b;
    layer4_outputs(6567) <= a and not b;
    layer4_outputs(6568) <= not (a and b);
    layer4_outputs(6569) <= not (a and b);
    layer4_outputs(6570) <= a;
    layer4_outputs(6571) <= a and b;
    layer4_outputs(6572) <= not a or b;
    layer4_outputs(6573) <= not a or b;
    layer4_outputs(6574) <= not a;
    layer4_outputs(6575) <= not (a or b);
    layer4_outputs(6576) <= 1'b0;
    layer4_outputs(6577) <= not a;
    layer4_outputs(6578) <= a;
    layer4_outputs(6579) <= 1'b0;
    layer4_outputs(6580) <= b and not a;
    layer4_outputs(6581) <= not b;
    layer4_outputs(6582) <= not (a or b);
    layer4_outputs(6583) <= b;
    layer4_outputs(6584) <= 1'b0;
    layer4_outputs(6585) <= a and not b;
    layer4_outputs(6586) <= not a;
    layer4_outputs(6587) <= 1'b0;
    layer4_outputs(6588) <= not a or b;
    layer4_outputs(6589) <= not a;
    layer4_outputs(6590) <= not (a and b);
    layer4_outputs(6591) <= a and b;
    layer4_outputs(6592) <= a or b;
    layer4_outputs(6593) <= b and not a;
    layer4_outputs(6594) <= a xor b;
    layer4_outputs(6595) <= not a or b;
    layer4_outputs(6596) <= b and not a;
    layer4_outputs(6597) <= a or b;
    layer4_outputs(6598) <= 1'b1;
    layer4_outputs(6599) <= not (a and b);
    layer4_outputs(6600) <= a and b;
    layer4_outputs(6601) <= not (a and b);
    layer4_outputs(6602) <= not (a xor b);
    layer4_outputs(6603) <= a and b;
    layer4_outputs(6604) <= not a or b;
    layer4_outputs(6605) <= b and not a;
    layer4_outputs(6606) <= a or b;
    layer4_outputs(6607) <= not a;
    layer4_outputs(6608) <= not (a or b);
    layer4_outputs(6609) <= not (a xor b);
    layer4_outputs(6610) <= a or b;
    layer4_outputs(6611) <= b and not a;
    layer4_outputs(6612) <= b;
    layer4_outputs(6613) <= a and b;
    layer4_outputs(6614) <= a and not b;
    layer4_outputs(6615) <= b;
    layer4_outputs(6616) <= not a or b;
    layer4_outputs(6617) <= not a;
    layer4_outputs(6618) <= 1'b0;
    layer4_outputs(6619) <= b;
    layer4_outputs(6620) <= b and not a;
    layer4_outputs(6621) <= b;
    layer4_outputs(6622) <= b and not a;
    layer4_outputs(6623) <= a;
    layer4_outputs(6624) <= a and b;
    layer4_outputs(6625) <= not (a or b);
    layer4_outputs(6626) <= not (a xor b);
    layer4_outputs(6627) <= not a;
    layer4_outputs(6628) <= not a;
    layer4_outputs(6629) <= not a;
    layer4_outputs(6630) <= 1'b0;
    layer4_outputs(6631) <= not b;
    layer4_outputs(6632) <= 1'b1;
    layer4_outputs(6633) <= a or b;
    layer4_outputs(6634) <= a or b;
    layer4_outputs(6635) <= a and not b;
    layer4_outputs(6636) <= not b or a;
    layer4_outputs(6637) <= a;
    layer4_outputs(6638) <= not (a or b);
    layer4_outputs(6639) <= not a;
    layer4_outputs(6640) <= b and not a;
    layer4_outputs(6641) <= not (a and b);
    layer4_outputs(6642) <= a or b;
    layer4_outputs(6643) <= 1'b0;
    layer4_outputs(6644) <= not (a or b);
    layer4_outputs(6645) <= not a;
    layer4_outputs(6646) <= a and not b;
    layer4_outputs(6647) <= 1'b1;
    layer4_outputs(6648) <= b;
    layer4_outputs(6649) <= b;
    layer4_outputs(6650) <= not (a and b);
    layer4_outputs(6651) <= not (a and b);
    layer4_outputs(6652) <= a and b;
    layer4_outputs(6653) <= a;
    layer4_outputs(6654) <= b and not a;
    layer4_outputs(6655) <= not b or a;
    layer4_outputs(6656) <= not (a or b);
    layer4_outputs(6657) <= not a or b;
    layer4_outputs(6658) <= 1'b0;
    layer4_outputs(6659) <= b and not a;
    layer4_outputs(6660) <= not a;
    layer4_outputs(6661) <= b and not a;
    layer4_outputs(6662) <= 1'b1;
    layer4_outputs(6663) <= a or b;
    layer4_outputs(6664) <= 1'b1;
    layer4_outputs(6665) <= a;
    layer4_outputs(6666) <= a and b;
    layer4_outputs(6667) <= a or b;
    layer4_outputs(6668) <= a or b;
    layer4_outputs(6669) <= not (a or b);
    layer4_outputs(6670) <= a or b;
    layer4_outputs(6671) <= a or b;
    layer4_outputs(6672) <= not a;
    layer4_outputs(6673) <= not a or b;
    layer4_outputs(6674) <= not b;
    layer4_outputs(6675) <= b and not a;
    layer4_outputs(6676) <= a xor b;
    layer4_outputs(6677) <= not (a xor b);
    layer4_outputs(6678) <= not b or a;
    layer4_outputs(6679) <= a and b;
    layer4_outputs(6680) <= b and not a;
    layer4_outputs(6681) <= a;
    layer4_outputs(6682) <= a;
    layer4_outputs(6683) <= b;
    layer4_outputs(6684) <= b and not a;
    layer4_outputs(6685) <= not a;
    layer4_outputs(6686) <= 1'b0;
    layer4_outputs(6687) <= not (a or b);
    layer4_outputs(6688) <= not b;
    layer4_outputs(6689) <= b and not a;
    layer4_outputs(6690) <= a and b;
    layer4_outputs(6691) <= not (a xor b);
    layer4_outputs(6692) <= 1'b1;
    layer4_outputs(6693) <= a;
    layer4_outputs(6694) <= a and not b;
    layer4_outputs(6695) <= not (a or b);
    layer4_outputs(6696) <= not (a and b);
    layer4_outputs(6697) <= a;
    layer4_outputs(6698) <= a xor b;
    layer4_outputs(6699) <= a and b;
    layer4_outputs(6700) <= b;
    layer4_outputs(6701) <= a and not b;
    layer4_outputs(6702) <= 1'b0;
    layer4_outputs(6703) <= a;
    layer4_outputs(6704) <= a or b;
    layer4_outputs(6705) <= not a;
    layer4_outputs(6706) <= not a or b;
    layer4_outputs(6707) <= not b or a;
    layer4_outputs(6708) <= a;
    layer4_outputs(6709) <= a;
    layer4_outputs(6710) <= not (a and b);
    layer4_outputs(6711) <= b;
    layer4_outputs(6712) <= b and not a;
    layer4_outputs(6713) <= not (a or b);
    layer4_outputs(6714) <= not (a or b);
    layer4_outputs(6715) <= b;
    layer4_outputs(6716) <= b and not a;
    layer4_outputs(6717) <= 1'b1;
    layer4_outputs(6718) <= not b or a;
    layer4_outputs(6719) <= not (a xor b);
    layer4_outputs(6720) <= not (a and b);
    layer4_outputs(6721) <= a;
    layer4_outputs(6722) <= not a;
    layer4_outputs(6723) <= not b;
    layer4_outputs(6724) <= 1'b0;
    layer4_outputs(6725) <= b;
    layer4_outputs(6726) <= b;
    layer4_outputs(6727) <= not b;
    layer4_outputs(6728) <= not a;
    layer4_outputs(6729) <= not (a and b);
    layer4_outputs(6730) <= not a or b;
    layer4_outputs(6731) <= not b;
    layer4_outputs(6732) <= not (a or b);
    layer4_outputs(6733) <= 1'b1;
    layer4_outputs(6734) <= not b;
    layer4_outputs(6735) <= 1'b0;
    layer4_outputs(6736) <= b and not a;
    layer4_outputs(6737) <= a or b;
    layer4_outputs(6738) <= not (a or b);
    layer4_outputs(6739) <= not a;
    layer4_outputs(6740) <= b;
    layer4_outputs(6741) <= not b;
    layer4_outputs(6742) <= a and not b;
    layer4_outputs(6743) <= 1'b1;
    layer4_outputs(6744) <= a;
    layer4_outputs(6745) <= not a;
    layer4_outputs(6746) <= not (a and b);
    layer4_outputs(6747) <= b and not a;
    layer4_outputs(6748) <= a and not b;
    layer4_outputs(6749) <= not b or a;
    layer4_outputs(6750) <= a;
    layer4_outputs(6751) <= not (a and b);
    layer4_outputs(6752) <= b and not a;
    layer4_outputs(6753) <= not (a and b);
    layer4_outputs(6754) <= a;
    layer4_outputs(6755) <= a and not b;
    layer4_outputs(6756) <= 1'b0;
    layer4_outputs(6757) <= a and b;
    layer4_outputs(6758) <= a;
    layer4_outputs(6759) <= not b;
    layer4_outputs(6760) <= not a;
    layer4_outputs(6761) <= not (a xor b);
    layer4_outputs(6762) <= a;
    layer4_outputs(6763) <= a;
    layer4_outputs(6764) <= a and b;
    layer4_outputs(6765) <= 1'b1;
    layer4_outputs(6766) <= b and not a;
    layer4_outputs(6767) <= b;
    layer4_outputs(6768) <= 1'b0;
    layer4_outputs(6769) <= a and b;
    layer4_outputs(6770) <= not a;
    layer4_outputs(6771) <= not b or a;
    layer4_outputs(6772) <= not b;
    layer4_outputs(6773) <= a;
    layer4_outputs(6774) <= a and not b;
    layer4_outputs(6775) <= not (a and b);
    layer4_outputs(6776) <= not (a or b);
    layer4_outputs(6777) <= not a or b;
    layer4_outputs(6778) <= 1'b1;
    layer4_outputs(6779) <= a and b;
    layer4_outputs(6780) <= not (a or b);
    layer4_outputs(6781) <= a;
    layer4_outputs(6782) <= a and b;
    layer4_outputs(6783) <= a;
    layer4_outputs(6784) <= b;
    layer4_outputs(6785) <= b and not a;
    layer4_outputs(6786) <= 1'b1;
    layer4_outputs(6787) <= not (a and b);
    layer4_outputs(6788) <= a;
    layer4_outputs(6789) <= 1'b0;
    layer4_outputs(6790) <= not (a or b);
    layer4_outputs(6791) <= b;
    layer4_outputs(6792) <= not b;
    layer4_outputs(6793) <= not (a or b);
    layer4_outputs(6794) <= not b or a;
    layer4_outputs(6795) <= b;
    layer4_outputs(6796) <= a;
    layer4_outputs(6797) <= not a or b;
    layer4_outputs(6798) <= not (a or b);
    layer4_outputs(6799) <= not a or b;
    layer4_outputs(6800) <= 1'b1;
    layer4_outputs(6801) <= not a;
    layer4_outputs(6802) <= not (a and b);
    layer4_outputs(6803) <= b;
    layer4_outputs(6804) <= not b;
    layer4_outputs(6805) <= not b;
    layer4_outputs(6806) <= not (a xor b);
    layer4_outputs(6807) <= a or b;
    layer4_outputs(6808) <= not b;
    layer4_outputs(6809) <= a;
    layer4_outputs(6810) <= not a or b;
    layer4_outputs(6811) <= a and not b;
    layer4_outputs(6812) <= not a;
    layer4_outputs(6813) <= 1'b1;
    layer4_outputs(6814) <= 1'b0;
    layer4_outputs(6815) <= not a;
    layer4_outputs(6816) <= 1'b1;
    layer4_outputs(6817) <= not a;
    layer4_outputs(6818) <= a and not b;
    layer4_outputs(6819) <= b and not a;
    layer4_outputs(6820) <= a;
    layer4_outputs(6821) <= b and not a;
    layer4_outputs(6822) <= a;
    layer4_outputs(6823) <= 1'b0;
    layer4_outputs(6824) <= not (a and b);
    layer4_outputs(6825) <= a or b;
    layer4_outputs(6826) <= not (a and b);
    layer4_outputs(6827) <= not (a xor b);
    layer4_outputs(6828) <= a and not b;
    layer4_outputs(6829) <= a or b;
    layer4_outputs(6830) <= not a;
    layer4_outputs(6831) <= 1'b0;
    layer4_outputs(6832) <= a and not b;
    layer4_outputs(6833) <= 1'b0;
    layer4_outputs(6834) <= 1'b0;
    layer4_outputs(6835) <= b and not a;
    layer4_outputs(6836) <= not b or a;
    layer4_outputs(6837) <= 1'b1;
    layer4_outputs(6838) <= not (a and b);
    layer4_outputs(6839) <= b and not a;
    layer4_outputs(6840) <= not b;
    layer4_outputs(6841) <= 1'b0;
    layer4_outputs(6842) <= a;
    layer4_outputs(6843) <= not (a and b);
    layer4_outputs(6844) <= not (a xor b);
    layer4_outputs(6845) <= not (a and b);
    layer4_outputs(6846) <= a xor b;
    layer4_outputs(6847) <= a and b;
    layer4_outputs(6848) <= not b or a;
    layer4_outputs(6849) <= not (a or b);
    layer4_outputs(6850) <= b and not a;
    layer4_outputs(6851) <= 1'b0;
    layer4_outputs(6852) <= b;
    layer4_outputs(6853) <= b and not a;
    layer4_outputs(6854) <= b;
    layer4_outputs(6855) <= not b or a;
    layer4_outputs(6856) <= not (a and b);
    layer4_outputs(6857) <= a and not b;
    layer4_outputs(6858) <= a or b;
    layer4_outputs(6859) <= not a or b;
    layer4_outputs(6860) <= b;
    layer4_outputs(6861) <= not (a and b);
    layer4_outputs(6862) <= b;
    layer4_outputs(6863) <= not b;
    layer4_outputs(6864) <= b;
    layer4_outputs(6865) <= b;
    layer4_outputs(6866) <= not b or a;
    layer4_outputs(6867) <= not b;
    layer4_outputs(6868) <= not b or a;
    layer4_outputs(6869) <= a;
    layer4_outputs(6870) <= a or b;
    layer4_outputs(6871) <= 1'b1;
    layer4_outputs(6872) <= not b;
    layer4_outputs(6873) <= not (a or b);
    layer4_outputs(6874) <= not a;
    layer4_outputs(6875) <= b;
    layer4_outputs(6876) <= b;
    layer4_outputs(6877) <= not a or b;
    layer4_outputs(6878) <= not (a and b);
    layer4_outputs(6879) <= not a;
    layer4_outputs(6880) <= a;
    layer4_outputs(6881) <= a or b;
    layer4_outputs(6882) <= not (a or b);
    layer4_outputs(6883) <= not b;
    layer4_outputs(6884) <= a and not b;
    layer4_outputs(6885) <= 1'b0;
    layer4_outputs(6886) <= 1'b0;
    layer4_outputs(6887) <= 1'b0;
    layer4_outputs(6888) <= a;
    layer4_outputs(6889) <= 1'b1;
    layer4_outputs(6890) <= b and not a;
    layer4_outputs(6891) <= not b;
    layer4_outputs(6892) <= 1'b1;
    layer4_outputs(6893) <= a;
    layer4_outputs(6894) <= not a or b;
    layer4_outputs(6895) <= a or b;
    layer4_outputs(6896) <= not (a xor b);
    layer4_outputs(6897) <= a and b;
    layer4_outputs(6898) <= b and not a;
    layer4_outputs(6899) <= b;
    layer4_outputs(6900) <= 1'b1;
    layer4_outputs(6901) <= 1'b0;
    layer4_outputs(6902) <= a;
    layer4_outputs(6903) <= 1'b0;
    layer4_outputs(6904) <= not (a xor b);
    layer4_outputs(6905) <= not b;
    layer4_outputs(6906) <= a and not b;
    layer4_outputs(6907) <= not (a and b);
    layer4_outputs(6908) <= not b or a;
    layer4_outputs(6909) <= not a;
    layer4_outputs(6910) <= not b;
    layer4_outputs(6911) <= b;
    layer4_outputs(6912) <= b and not a;
    layer4_outputs(6913) <= b and not a;
    layer4_outputs(6914) <= a and not b;
    layer4_outputs(6915) <= a;
    layer4_outputs(6916) <= a xor b;
    layer4_outputs(6917) <= b;
    layer4_outputs(6918) <= a and not b;
    layer4_outputs(6919) <= b;
    layer4_outputs(6920) <= not (a or b);
    layer4_outputs(6921) <= not (a and b);
    layer4_outputs(6922) <= a and b;
    layer4_outputs(6923) <= a xor b;
    layer4_outputs(6924) <= a and not b;
    layer4_outputs(6925) <= not a or b;
    layer4_outputs(6926) <= b and not a;
    layer4_outputs(6927) <= a;
    layer4_outputs(6928) <= not b;
    layer4_outputs(6929) <= b and not a;
    layer4_outputs(6930) <= not (a and b);
    layer4_outputs(6931) <= b;
    layer4_outputs(6932) <= a and b;
    layer4_outputs(6933) <= 1'b1;
    layer4_outputs(6934) <= not a;
    layer4_outputs(6935) <= not a;
    layer4_outputs(6936) <= not a;
    layer4_outputs(6937) <= not b;
    layer4_outputs(6938) <= not b;
    layer4_outputs(6939) <= b and not a;
    layer4_outputs(6940) <= not (a and b);
    layer4_outputs(6941) <= not (a and b);
    layer4_outputs(6942) <= 1'b1;
    layer4_outputs(6943) <= a;
    layer4_outputs(6944) <= b;
    layer4_outputs(6945) <= not a;
    layer4_outputs(6946) <= 1'b1;
    layer4_outputs(6947) <= 1'b1;
    layer4_outputs(6948) <= not a;
    layer4_outputs(6949) <= not (a xor b);
    layer4_outputs(6950) <= 1'b0;
    layer4_outputs(6951) <= not a or b;
    layer4_outputs(6952) <= 1'b1;
    layer4_outputs(6953) <= not a;
    layer4_outputs(6954) <= a or b;
    layer4_outputs(6955) <= not (a or b);
    layer4_outputs(6956) <= not a;
    layer4_outputs(6957) <= not a;
    layer4_outputs(6958) <= not (a or b);
    layer4_outputs(6959) <= b and not a;
    layer4_outputs(6960) <= not a or b;
    layer4_outputs(6961) <= not a;
    layer4_outputs(6962) <= not b;
    layer4_outputs(6963) <= 1'b1;
    layer4_outputs(6964) <= not (a and b);
    layer4_outputs(6965) <= not a or b;
    layer4_outputs(6966) <= b and not a;
    layer4_outputs(6967) <= not b or a;
    layer4_outputs(6968) <= b;
    layer4_outputs(6969) <= not (a or b);
    layer4_outputs(6970) <= not a or b;
    layer4_outputs(6971) <= not b or a;
    layer4_outputs(6972) <= not (a or b);
    layer4_outputs(6973) <= not a;
    layer4_outputs(6974) <= a xor b;
    layer4_outputs(6975) <= a and not b;
    layer4_outputs(6976) <= not b;
    layer4_outputs(6977) <= not b;
    layer4_outputs(6978) <= not (a and b);
    layer4_outputs(6979) <= not b or a;
    layer4_outputs(6980) <= not (a and b);
    layer4_outputs(6981) <= not a;
    layer4_outputs(6982) <= b and not a;
    layer4_outputs(6983) <= b;
    layer4_outputs(6984) <= not b or a;
    layer4_outputs(6985) <= not a;
    layer4_outputs(6986) <= a or b;
    layer4_outputs(6987) <= not (a xor b);
    layer4_outputs(6988) <= a and not b;
    layer4_outputs(6989) <= not b;
    layer4_outputs(6990) <= a;
    layer4_outputs(6991) <= not b;
    layer4_outputs(6992) <= not (a or b);
    layer4_outputs(6993) <= a and not b;
    layer4_outputs(6994) <= a or b;
    layer4_outputs(6995) <= not b or a;
    layer4_outputs(6996) <= not b;
    layer4_outputs(6997) <= not (a or b);
    layer4_outputs(6998) <= not (a and b);
    layer4_outputs(6999) <= 1'b1;
    layer4_outputs(7000) <= not b;
    layer4_outputs(7001) <= 1'b1;
    layer4_outputs(7002) <= not (a xor b);
    layer4_outputs(7003) <= not (a xor b);
    layer4_outputs(7004) <= not a;
    layer4_outputs(7005) <= 1'b1;
    layer4_outputs(7006) <= 1'b1;
    layer4_outputs(7007) <= 1'b1;
    layer4_outputs(7008) <= a and b;
    layer4_outputs(7009) <= a or b;
    layer4_outputs(7010) <= a xor b;
    layer4_outputs(7011) <= not (a and b);
    layer4_outputs(7012) <= not a or b;
    layer4_outputs(7013) <= not b;
    layer4_outputs(7014) <= b and not a;
    layer4_outputs(7015) <= not a or b;
    layer4_outputs(7016) <= not a;
    layer4_outputs(7017) <= a and not b;
    layer4_outputs(7018) <= not b or a;
    layer4_outputs(7019) <= a;
    layer4_outputs(7020) <= not b;
    layer4_outputs(7021) <= a or b;
    layer4_outputs(7022) <= not b or a;
    layer4_outputs(7023) <= not a;
    layer4_outputs(7024) <= not b;
    layer4_outputs(7025) <= not (a or b);
    layer4_outputs(7026) <= not a or b;
    layer4_outputs(7027) <= not b;
    layer4_outputs(7028) <= a or b;
    layer4_outputs(7029) <= a;
    layer4_outputs(7030) <= b and not a;
    layer4_outputs(7031) <= a;
    layer4_outputs(7032) <= not b;
    layer4_outputs(7033) <= not a;
    layer4_outputs(7034) <= b;
    layer4_outputs(7035) <= not (a or b);
    layer4_outputs(7036) <= b and not a;
    layer4_outputs(7037) <= 1'b0;
    layer4_outputs(7038) <= not a;
    layer4_outputs(7039) <= 1'b1;
    layer4_outputs(7040) <= not b;
    layer4_outputs(7041) <= not a;
    layer4_outputs(7042) <= 1'b1;
    layer4_outputs(7043) <= not b;
    layer4_outputs(7044) <= not a or b;
    layer4_outputs(7045) <= a or b;
    layer4_outputs(7046) <= not b;
    layer4_outputs(7047) <= not a or b;
    layer4_outputs(7048) <= not b or a;
    layer4_outputs(7049) <= 1'b1;
    layer4_outputs(7050) <= a and not b;
    layer4_outputs(7051) <= not a or b;
    layer4_outputs(7052) <= a and not b;
    layer4_outputs(7053) <= not a;
    layer4_outputs(7054) <= not b or a;
    layer4_outputs(7055) <= not b;
    layer4_outputs(7056) <= b;
    layer4_outputs(7057) <= a;
    layer4_outputs(7058) <= a;
    layer4_outputs(7059) <= not a;
    layer4_outputs(7060) <= not a or b;
    layer4_outputs(7061) <= a;
    layer4_outputs(7062) <= not a or b;
    layer4_outputs(7063) <= b and not a;
    layer4_outputs(7064) <= b;
    layer4_outputs(7065) <= a or b;
    layer4_outputs(7066) <= not a;
    layer4_outputs(7067) <= not (a or b);
    layer4_outputs(7068) <= a and b;
    layer4_outputs(7069) <= a and not b;
    layer4_outputs(7070) <= not a;
    layer4_outputs(7071) <= not (a and b);
    layer4_outputs(7072) <= 1'b0;
    layer4_outputs(7073) <= a and not b;
    layer4_outputs(7074) <= not (a and b);
    layer4_outputs(7075) <= b and not a;
    layer4_outputs(7076) <= 1'b0;
    layer4_outputs(7077) <= a;
    layer4_outputs(7078) <= b;
    layer4_outputs(7079) <= b and not a;
    layer4_outputs(7080) <= a or b;
    layer4_outputs(7081) <= not a or b;
    layer4_outputs(7082) <= 1'b1;
    layer4_outputs(7083) <= 1'b0;
    layer4_outputs(7084) <= not b;
    layer4_outputs(7085) <= a xor b;
    layer4_outputs(7086) <= b and not a;
    layer4_outputs(7087) <= not (a and b);
    layer4_outputs(7088) <= not a or b;
    layer4_outputs(7089) <= 1'b1;
    layer4_outputs(7090) <= a and b;
    layer4_outputs(7091) <= not a or b;
    layer4_outputs(7092) <= a xor b;
    layer4_outputs(7093) <= not a;
    layer4_outputs(7094) <= not a or b;
    layer4_outputs(7095) <= a or b;
    layer4_outputs(7096) <= 1'b1;
    layer4_outputs(7097) <= not b or a;
    layer4_outputs(7098) <= 1'b1;
    layer4_outputs(7099) <= a and b;
    layer4_outputs(7100) <= not b or a;
    layer4_outputs(7101) <= not b or a;
    layer4_outputs(7102) <= a;
    layer4_outputs(7103) <= 1'b0;
    layer4_outputs(7104) <= b and not a;
    layer4_outputs(7105) <= 1'b1;
    layer4_outputs(7106) <= not a;
    layer4_outputs(7107) <= not b or a;
    layer4_outputs(7108) <= a xor b;
    layer4_outputs(7109) <= not (a or b);
    layer4_outputs(7110) <= b and not a;
    layer4_outputs(7111) <= b;
    layer4_outputs(7112) <= a and b;
    layer4_outputs(7113) <= not b;
    layer4_outputs(7114) <= not b;
    layer4_outputs(7115) <= not a;
    layer4_outputs(7116) <= a and b;
    layer4_outputs(7117) <= b;
    layer4_outputs(7118) <= not (a and b);
    layer4_outputs(7119) <= b;
    layer4_outputs(7120) <= a and b;
    layer4_outputs(7121) <= a and b;
    layer4_outputs(7122) <= a;
    layer4_outputs(7123) <= a or b;
    layer4_outputs(7124) <= not b;
    layer4_outputs(7125) <= b and not a;
    layer4_outputs(7126) <= a and b;
    layer4_outputs(7127) <= a;
    layer4_outputs(7128) <= not b;
    layer4_outputs(7129) <= 1'b1;
    layer4_outputs(7130) <= a;
    layer4_outputs(7131) <= 1'b0;
    layer4_outputs(7132) <= a and not b;
    layer4_outputs(7133) <= not b;
    layer4_outputs(7134) <= not a or b;
    layer4_outputs(7135) <= a and not b;
    layer4_outputs(7136) <= not (a and b);
    layer4_outputs(7137) <= a and b;
    layer4_outputs(7138) <= a and b;
    layer4_outputs(7139) <= 1'b0;
    layer4_outputs(7140) <= a or b;
    layer4_outputs(7141) <= b;
    layer4_outputs(7142) <= not (a or b);
    layer4_outputs(7143) <= not a;
    layer4_outputs(7144) <= not a or b;
    layer4_outputs(7145) <= not b or a;
    layer4_outputs(7146) <= a or b;
    layer4_outputs(7147) <= not b or a;
    layer4_outputs(7148) <= a and not b;
    layer4_outputs(7149) <= 1'b0;
    layer4_outputs(7150) <= not b or a;
    layer4_outputs(7151) <= not a;
    layer4_outputs(7152) <= 1'b0;
    layer4_outputs(7153) <= a and not b;
    layer4_outputs(7154) <= a and not b;
    layer4_outputs(7155) <= b;
    layer4_outputs(7156) <= not a or b;
    layer4_outputs(7157) <= not a;
    layer4_outputs(7158) <= a and b;
    layer4_outputs(7159) <= b;
    layer4_outputs(7160) <= a and not b;
    layer4_outputs(7161) <= not (a and b);
    layer4_outputs(7162) <= a or b;
    layer4_outputs(7163) <= not b;
    layer4_outputs(7164) <= not b;
    layer4_outputs(7165) <= not (a and b);
    layer4_outputs(7166) <= not b;
    layer4_outputs(7167) <= 1'b0;
    layer4_outputs(7168) <= a and b;
    layer4_outputs(7169) <= a and b;
    layer4_outputs(7170) <= 1'b1;
    layer4_outputs(7171) <= 1'b0;
    layer4_outputs(7172) <= not b;
    layer4_outputs(7173) <= a;
    layer4_outputs(7174) <= 1'b1;
    layer4_outputs(7175) <= not (a or b);
    layer4_outputs(7176) <= not (a xor b);
    layer4_outputs(7177) <= not (a xor b);
    layer4_outputs(7178) <= a and not b;
    layer4_outputs(7179) <= 1'b1;
    layer4_outputs(7180) <= not a;
    layer4_outputs(7181) <= a;
    layer4_outputs(7182) <= a or b;
    layer4_outputs(7183) <= 1'b1;
    layer4_outputs(7184) <= 1'b1;
    layer4_outputs(7185) <= a or b;
    layer4_outputs(7186) <= a;
    layer4_outputs(7187) <= not (a or b);
    layer4_outputs(7188) <= 1'b1;
    layer4_outputs(7189) <= not (a or b);
    layer4_outputs(7190) <= a;
    layer4_outputs(7191) <= a or b;
    layer4_outputs(7192) <= not (a and b);
    layer4_outputs(7193) <= 1'b0;
    layer4_outputs(7194) <= not b or a;
    layer4_outputs(7195) <= b;
    layer4_outputs(7196) <= 1'b0;
    layer4_outputs(7197) <= not (a or b);
    layer4_outputs(7198) <= not (a and b);
    layer4_outputs(7199) <= b;
    layer4_outputs(7200) <= b and not a;
    layer4_outputs(7201) <= 1'b0;
    layer4_outputs(7202) <= a;
    layer4_outputs(7203) <= 1'b1;
    layer4_outputs(7204) <= not a;
    layer4_outputs(7205) <= not (a or b);
    layer4_outputs(7206) <= b;
    layer4_outputs(7207) <= not (a or b);
    layer4_outputs(7208) <= b and not a;
    layer4_outputs(7209) <= b and not a;
    layer4_outputs(7210) <= not (a and b);
    layer4_outputs(7211) <= a or b;
    layer4_outputs(7212) <= not a or b;
    layer4_outputs(7213) <= b and not a;
    layer4_outputs(7214) <= a;
    layer4_outputs(7215) <= a and b;
    layer4_outputs(7216) <= not a or b;
    layer4_outputs(7217) <= not (a and b);
    layer4_outputs(7218) <= not a or b;
    layer4_outputs(7219) <= b;
    layer4_outputs(7220) <= 1'b0;
    layer4_outputs(7221) <= a xor b;
    layer4_outputs(7222) <= not (a and b);
    layer4_outputs(7223) <= not b or a;
    layer4_outputs(7224) <= a and b;
    layer4_outputs(7225) <= b;
    layer4_outputs(7226) <= not (a or b);
    layer4_outputs(7227) <= not (a and b);
    layer4_outputs(7228) <= a or b;
    layer4_outputs(7229) <= a and not b;
    layer4_outputs(7230) <= not a;
    layer4_outputs(7231) <= not b;
    layer4_outputs(7232) <= b;
    layer4_outputs(7233) <= a and b;
    layer4_outputs(7234) <= a and not b;
    layer4_outputs(7235) <= not a;
    layer4_outputs(7236) <= a and b;
    layer4_outputs(7237) <= not (a or b);
    layer4_outputs(7238) <= not b;
    layer4_outputs(7239) <= not (a or b);
    layer4_outputs(7240) <= not (a or b);
    layer4_outputs(7241) <= not (a and b);
    layer4_outputs(7242) <= a;
    layer4_outputs(7243) <= not b;
    layer4_outputs(7244) <= a and b;
    layer4_outputs(7245) <= b;
    layer4_outputs(7246) <= a;
    layer4_outputs(7247) <= not b;
    layer4_outputs(7248) <= b;
    layer4_outputs(7249) <= a;
    layer4_outputs(7250) <= 1'b0;
    layer4_outputs(7251) <= b and not a;
    layer4_outputs(7252) <= not (a and b);
    layer4_outputs(7253) <= a and b;
    layer4_outputs(7254) <= not a;
    layer4_outputs(7255) <= not a;
    layer4_outputs(7256) <= not b or a;
    layer4_outputs(7257) <= not a or b;
    layer4_outputs(7258) <= a and not b;
    layer4_outputs(7259) <= b;
    layer4_outputs(7260) <= a xor b;
    layer4_outputs(7261) <= b;
    layer4_outputs(7262) <= a and b;
    layer4_outputs(7263) <= a;
    layer4_outputs(7264) <= a;
    layer4_outputs(7265) <= a or b;
    layer4_outputs(7266) <= a and not b;
    layer4_outputs(7267) <= a and not b;
    layer4_outputs(7268) <= not b or a;
    layer4_outputs(7269) <= 1'b1;
    layer4_outputs(7270) <= not (a or b);
    layer4_outputs(7271) <= a or b;
    layer4_outputs(7272) <= not (a xor b);
    layer4_outputs(7273) <= 1'b0;
    layer4_outputs(7274) <= not a;
    layer4_outputs(7275) <= not a or b;
    layer4_outputs(7276) <= not a;
    layer4_outputs(7277) <= a;
    layer4_outputs(7278) <= 1'b0;
    layer4_outputs(7279) <= b and not a;
    layer4_outputs(7280) <= a or b;
    layer4_outputs(7281) <= not (a and b);
    layer4_outputs(7282) <= 1'b0;
    layer4_outputs(7283) <= not b;
    layer4_outputs(7284) <= b and not a;
    layer4_outputs(7285) <= not a or b;
    layer4_outputs(7286) <= a;
    layer4_outputs(7287) <= b;
    layer4_outputs(7288) <= 1'b0;
    layer4_outputs(7289) <= not (a and b);
    layer4_outputs(7290) <= not a;
    layer4_outputs(7291) <= a and b;
    layer4_outputs(7292) <= not (a and b);
    layer4_outputs(7293) <= a xor b;
    layer4_outputs(7294) <= b and not a;
    layer4_outputs(7295) <= a and b;
    layer4_outputs(7296) <= a xor b;
    layer4_outputs(7297) <= not b or a;
    layer4_outputs(7298) <= b;
    layer4_outputs(7299) <= not (a or b);
    layer4_outputs(7300) <= 1'b1;
    layer4_outputs(7301) <= not b;
    layer4_outputs(7302) <= b;
    layer4_outputs(7303) <= b;
    layer4_outputs(7304) <= a;
    layer4_outputs(7305) <= a and b;
    layer4_outputs(7306) <= 1'b0;
    layer4_outputs(7307) <= b;
    layer4_outputs(7308) <= not a or b;
    layer4_outputs(7309) <= b;
    layer4_outputs(7310) <= not b or a;
    layer4_outputs(7311) <= not a;
    layer4_outputs(7312) <= a;
    layer4_outputs(7313) <= not a;
    layer4_outputs(7314) <= a xor b;
    layer4_outputs(7315) <= not (a xor b);
    layer4_outputs(7316) <= a and b;
    layer4_outputs(7317) <= a and b;
    layer4_outputs(7318) <= not b or a;
    layer4_outputs(7319) <= not b or a;
    layer4_outputs(7320) <= a and not b;
    layer4_outputs(7321) <= not a;
    layer4_outputs(7322) <= not a or b;
    layer4_outputs(7323) <= a or b;
    layer4_outputs(7324) <= not (a and b);
    layer4_outputs(7325) <= not a;
    layer4_outputs(7326) <= not (a xor b);
    layer4_outputs(7327) <= a or b;
    layer4_outputs(7328) <= not (a and b);
    layer4_outputs(7329) <= a and not b;
    layer4_outputs(7330) <= not (a and b);
    layer4_outputs(7331) <= not (a and b);
    layer4_outputs(7332) <= 1'b0;
    layer4_outputs(7333) <= not b;
    layer4_outputs(7334) <= a or b;
    layer4_outputs(7335) <= a xor b;
    layer4_outputs(7336) <= 1'b1;
    layer4_outputs(7337) <= not b or a;
    layer4_outputs(7338) <= a and b;
    layer4_outputs(7339) <= 1'b1;
    layer4_outputs(7340) <= not a;
    layer4_outputs(7341) <= 1'b0;
    layer4_outputs(7342) <= not a;
    layer4_outputs(7343) <= a;
    layer4_outputs(7344) <= a;
    layer4_outputs(7345) <= not a;
    layer4_outputs(7346) <= not b;
    layer4_outputs(7347) <= not a;
    layer4_outputs(7348) <= a or b;
    layer4_outputs(7349) <= not b;
    layer4_outputs(7350) <= not b;
    layer4_outputs(7351) <= not a or b;
    layer4_outputs(7352) <= b;
    layer4_outputs(7353) <= 1'b0;
    layer4_outputs(7354) <= not a;
    layer4_outputs(7355) <= 1'b1;
    layer4_outputs(7356) <= a;
    layer4_outputs(7357) <= a and b;
    layer4_outputs(7358) <= not (a xor b);
    layer4_outputs(7359) <= not (a or b);
    layer4_outputs(7360) <= not (a and b);
    layer4_outputs(7361) <= a and not b;
    layer4_outputs(7362) <= not b or a;
    layer4_outputs(7363) <= not (a and b);
    layer4_outputs(7364) <= b and not a;
    layer4_outputs(7365) <= not a or b;
    layer4_outputs(7366) <= a;
    layer4_outputs(7367) <= a xor b;
    layer4_outputs(7368) <= not (a and b);
    layer4_outputs(7369) <= a;
    layer4_outputs(7370) <= b;
    layer4_outputs(7371) <= 1'b1;
    layer4_outputs(7372) <= b;
    layer4_outputs(7373) <= b;
    layer4_outputs(7374) <= a xor b;
    layer4_outputs(7375) <= 1'b0;
    layer4_outputs(7376) <= b and not a;
    layer4_outputs(7377) <= a or b;
    layer4_outputs(7378) <= 1'b0;
    layer4_outputs(7379) <= a and not b;
    layer4_outputs(7380) <= not (a and b);
    layer4_outputs(7381) <= a xor b;
    layer4_outputs(7382) <= a xor b;
    layer4_outputs(7383) <= not a or b;
    layer4_outputs(7384) <= a and b;
    layer4_outputs(7385) <= not (a or b);
    layer4_outputs(7386) <= b;
    layer4_outputs(7387) <= a and b;
    layer4_outputs(7388) <= not b;
    layer4_outputs(7389) <= not a or b;
    layer4_outputs(7390) <= b;
    layer4_outputs(7391) <= not (a xor b);
    layer4_outputs(7392) <= a or b;
    layer4_outputs(7393) <= a;
    layer4_outputs(7394) <= not b or a;
    layer4_outputs(7395) <= a and not b;
    layer4_outputs(7396) <= not a or b;
    layer4_outputs(7397) <= not a;
    layer4_outputs(7398) <= a or b;
    layer4_outputs(7399) <= a and not b;
    layer4_outputs(7400) <= a xor b;
    layer4_outputs(7401) <= b and not a;
    layer4_outputs(7402) <= not b or a;
    layer4_outputs(7403) <= a;
    layer4_outputs(7404) <= a;
    layer4_outputs(7405) <= 1'b1;
    layer4_outputs(7406) <= not b or a;
    layer4_outputs(7407) <= a or b;
    layer4_outputs(7408) <= a and b;
    layer4_outputs(7409) <= a;
    layer4_outputs(7410) <= a and not b;
    layer4_outputs(7411) <= not a or b;
    layer4_outputs(7412) <= 1'b0;
    layer4_outputs(7413) <= 1'b0;
    layer4_outputs(7414) <= not a or b;
    layer4_outputs(7415) <= not a or b;
    layer4_outputs(7416) <= a;
    layer4_outputs(7417) <= a or b;
    layer4_outputs(7418) <= not a or b;
    layer4_outputs(7419) <= a and not b;
    layer4_outputs(7420) <= b and not a;
    layer4_outputs(7421) <= not a;
    layer4_outputs(7422) <= not b;
    layer4_outputs(7423) <= not b or a;
    layer4_outputs(7424) <= a xor b;
    layer4_outputs(7425) <= not b;
    layer4_outputs(7426) <= not a;
    layer4_outputs(7427) <= b;
    layer4_outputs(7428) <= 1'b0;
    layer4_outputs(7429) <= a or b;
    layer4_outputs(7430) <= 1'b1;
    layer4_outputs(7431) <= a or b;
    layer4_outputs(7432) <= not (a and b);
    layer4_outputs(7433) <= a;
    layer4_outputs(7434) <= 1'b0;
    layer4_outputs(7435) <= 1'b0;
    layer4_outputs(7436) <= not a or b;
    layer4_outputs(7437) <= not (a and b);
    layer4_outputs(7438) <= b and not a;
    layer4_outputs(7439) <= not b;
    layer4_outputs(7440) <= a or b;
    layer4_outputs(7441) <= a or b;
    layer4_outputs(7442) <= not b or a;
    layer4_outputs(7443) <= not (a and b);
    layer4_outputs(7444) <= b and not a;
    layer4_outputs(7445) <= a xor b;
    layer4_outputs(7446) <= a and not b;
    layer4_outputs(7447) <= not (a and b);
    layer4_outputs(7448) <= not a;
    layer4_outputs(7449) <= not a;
    layer4_outputs(7450) <= a xor b;
    layer4_outputs(7451) <= 1'b0;
    layer4_outputs(7452) <= not a;
    layer4_outputs(7453) <= not (a and b);
    layer4_outputs(7454) <= 1'b1;
    layer4_outputs(7455) <= not (a and b);
    layer4_outputs(7456) <= not a or b;
    layer4_outputs(7457) <= not (a and b);
    layer4_outputs(7458) <= 1'b1;
    layer4_outputs(7459) <= not b or a;
    layer4_outputs(7460) <= a or b;
    layer4_outputs(7461) <= not a or b;
    layer4_outputs(7462) <= a and b;
    layer4_outputs(7463) <= not a or b;
    layer4_outputs(7464) <= not b;
    layer4_outputs(7465) <= 1'b0;
    layer4_outputs(7466) <= not b;
    layer4_outputs(7467) <= not a;
    layer4_outputs(7468) <= a xor b;
    layer4_outputs(7469) <= not a;
    layer4_outputs(7470) <= not a;
    layer4_outputs(7471) <= not b;
    layer4_outputs(7472) <= 1'b1;
    layer4_outputs(7473) <= 1'b0;
    layer4_outputs(7474) <= not a or b;
    layer4_outputs(7475) <= a and not b;
    layer4_outputs(7476) <= 1'b1;
    layer4_outputs(7477) <= not (a or b);
    layer4_outputs(7478) <= not (a and b);
    layer4_outputs(7479) <= 1'b0;
    layer4_outputs(7480) <= not a or b;
    layer4_outputs(7481) <= a and not b;
    layer4_outputs(7482) <= not b;
    layer4_outputs(7483) <= 1'b1;
    layer4_outputs(7484) <= not a;
    layer4_outputs(7485) <= a and not b;
    layer4_outputs(7486) <= not a or b;
    layer4_outputs(7487) <= not b;
    layer4_outputs(7488) <= not b or a;
    layer4_outputs(7489) <= a and not b;
    layer4_outputs(7490) <= 1'b1;
    layer4_outputs(7491) <= not (a and b);
    layer4_outputs(7492) <= b;
    layer4_outputs(7493) <= b;
    layer4_outputs(7494) <= not (a or b);
    layer4_outputs(7495) <= a or b;
    layer4_outputs(7496) <= not b;
    layer4_outputs(7497) <= a;
    layer4_outputs(7498) <= not b or a;
    layer4_outputs(7499) <= a;
    layer4_outputs(7500) <= not b;
    layer4_outputs(7501) <= not b or a;
    layer4_outputs(7502) <= not (a or b);
    layer4_outputs(7503) <= a or b;
    layer4_outputs(7504) <= b and not a;
    layer4_outputs(7505) <= 1'b0;
    layer4_outputs(7506) <= a and b;
    layer4_outputs(7507) <= a and b;
    layer4_outputs(7508) <= b;
    layer4_outputs(7509) <= a xor b;
    layer4_outputs(7510) <= not b;
    layer4_outputs(7511) <= a or b;
    layer4_outputs(7512) <= not (a and b);
    layer4_outputs(7513) <= 1'b0;
    layer4_outputs(7514) <= not (a and b);
    layer4_outputs(7515) <= 1'b0;
    layer4_outputs(7516) <= a or b;
    layer4_outputs(7517) <= a or b;
    layer4_outputs(7518) <= not (a and b);
    layer4_outputs(7519) <= a;
    layer4_outputs(7520) <= not (a and b);
    layer4_outputs(7521) <= a;
    layer4_outputs(7522) <= b;
    layer4_outputs(7523) <= a and b;
    layer4_outputs(7524) <= 1'b1;
    layer4_outputs(7525) <= b and not a;
    layer4_outputs(7526) <= not (a xor b);
    layer4_outputs(7527) <= a and b;
    layer4_outputs(7528) <= not b;
    layer4_outputs(7529) <= not b or a;
    layer4_outputs(7530) <= not b or a;
    layer4_outputs(7531) <= not a;
    layer4_outputs(7532) <= not a;
    layer4_outputs(7533) <= not (a and b);
    layer4_outputs(7534) <= a xor b;
    layer4_outputs(7535) <= 1'b1;
    layer4_outputs(7536) <= not a;
    layer4_outputs(7537) <= b and not a;
    layer4_outputs(7538) <= a;
    layer4_outputs(7539) <= not a or b;
    layer4_outputs(7540) <= a and b;
    layer4_outputs(7541) <= a or b;
    layer4_outputs(7542) <= a;
    layer4_outputs(7543) <= a or b;
    layer4_outputs(7544) <= a;
    layer4_outputs(7545) <= a;
    layer4_outputs(7546) <= not (a and b);
    layer4_outputs(7547) <= a and not b;
    layer4_outputs(7548) <= a and b;
    layer4_outputs(7549) <= not b or a;
    layer4_outputs(7550) <= not a;
    layer4_outputs(7551) <= b;
    layer4_outputs(7552) <= not a or b;
    layer4_outputs(7553) <= not (a and b);
    layer4_outputs(7554) <= not (a xor b);
    layer4_outputs(7555) <= 1'b0;
    layer4_outputs(7556) <= not a;
    layer4_outputs(7557) <= a and b;
    layer4_outputs(7558) <= 1'b1;
    layer4_outputs(7559) <= not (a or b);
    layer4_outputs(7560) <= not a or b;
    layer4_outputs(7561) <= a or b;
    layer4_outputs(7562) <= a and not b;
    layer4_outputs(7563) <= b;
    layer4_outputs(7564) <= b;
    layer4_outputs(7565) <= not (a and b);
    layer4_outputs(7566) <= a and b;
    layer4_outputs(7567) <= 1'b1;
    layer4_outputs(7568) <= not b or a;
    layer4_outputs(7569) <= b and not a;
    layer4_outputs(7570) <= a;
    layer4_outputs(7571) <= not a;
    layer4_outputs(7572) <= not (a and b);
    layer4_outputs(7573) <= b and not a;
    layer4_outputs(7574) <= 1'b0;
    layer4_outputs(7575) <= not a;
    layer4_outputs(7576) <= a and not b;
    layer4_outputs(7577) <= a;
    layer4_outputs(7578) <= b and not a;
    layer4_outputs(7579) <= a;
    layer4_outputs(7580) <= not a;
    layer4_outputs(7581) <= not (a and b);
    layer4_outputs(7582) <= not b or a;
    layer4_outputs(7583) <= a and not b;
    layer4_outputs(7584) <= not a or b;
    layer4_outputs(7585) <= not a;
    layer4_outputs(7586) <= not a or b;
    layer4_outputs(7587) <= a xor b;
    layer4_outputs(7588) <= a and not b;
    layer4_outputs(7589) <= not a;
    layer4_outputs(7590) <= a or b;
    layer4_outputs(7591) <= 1'b0;
    layer4_outputs(7592) <= not a or b;
    layer4_outputs(7593) <= a and not b;
    layer4_outputs(7594) <= not a or b;
    layer4_outputs(7595) <= a or b;
    layer4_outputs(7596) <= not b;
    layer4_outputs(7597) <= a and b;
    layer4_outputs(7598) <= not (a and b);
    layer4_outputs(7599) <= a or b;
    layer4_outputs(7600) <= a;
    layer4_outputs(7601) <= not (a or b);
    layer4_outputs(7602) <= a and not b;
    layer4_outputs(7603) <= a;
    layer4_outputs(7604) <= b and not a;
    layer4_outputs(7605) <= not (a or b);
    layer4_outputs(7606) <= a;
    layer4_outputs(7607) <= not (a or b);
    layer4_outputs(7608) <= 1'b1;
    layer4_outputs(7609) <= b;
    layer4_outputs(7610) <= not a or b;
    layer4_outputs(7611) <= not a or b;
    layer4_outputs(7612) <= a and not b;
    layer4_outputs(7613) <= a;
    layer4_outputs(7614) <= not b;
    layer4_outputs(7615) <= not a;
    layer4_outputs(7616) <= a;
    layer4_outputs(7617) <= not a;
    layer4_outputs(7618) <= not a or b;
    layer4_outputs(7619) <= not (a or b);
    layer4_outputs(7620) <= not a;
    layer4_outputs(7621) <= not (a xor b);
    layer4_outputs(7622) <= b;
    layer4_outputs(7623) <= not a;
    layer4_outputs(7624) <= not b;
    layer4_outputs(7625) <= a and not b;
    layer4_outputs(7626) <= 1'b0;
    layer4_outputs(7627) <= not b;
    layer4_outputs(7628) <= not a;
    layer4_outputs(7629) <= 1'b0;
    layer4_outputs(7630) <= 1'b1;
    layer4_outputs(7631) <= not (a or b);
    layer4_outputs(7632) <= not b or a;
    layer4_outputs(7633) <= a;
    layer4_outputs(7634) <= 1'b1;
    layer4_outputs(7635) <= a or b;
    layer4_outputs(7636) <= a and b;
    layer4_outputs(7637) <= b;
    layer4_outputs(7638) <= 1'b1;
    layer4_outputs(7639) <= not a;
    layer4_outputs(7640) <= b;
    layer4_outputs(7641) <= not a or b;
    layer4_outputs(7642) <= not b or a;
    layer4_outputs(7643) <= 1'b1;
    layer4_outputs(7644) <= a or b;
    layer4_outputs(7645) <= not a or b;
    layer4_outputs(7646) <= not a or b;
    layer4_outputs(7647) <= a and not b;
    layer4_outputs(7648) <= not a;
    layer4_outputs(7649) <= a and b;
    layer4_outputs(7650) <= not (a xor b);
    layer4_outputs(7651) <= not a or b;
    layer4_outputs(7652) <= not b or a;
    layer4_outputs(7653) <= a and b;
    layer4_outputs(7654) <= not (a or b);
    layer4_outputs(7655) <= not (a and b);
    layer4_outputs(7656) <= 1'b0;
    layer4_outputs(7657) <= b;
    layer4_outputs(7658) <= a;
    layer4_outputs(7659) <= not (a or b);
    layer4_outputs(7660) <= not b or a;
    layer4_outputs(7661) <= not a or b;
    layer4_outputs(7662) <= not b;
    layer4_outputs(7663) <= not (a or b);
    layer4_outputs(7664) <= a;
    layer4_outputs(7665) <= 1'b1;
    layer4_outputs(7666) <= 1'b0;
    layer4_outputs(7667) <= b and not a;
    layer4_outputs(7668) <= b;
    layer4_outputs(7669) <= a and b;
    layer4_outputs(7670) <= a;
    layer4_outputs(7671) <= not b;
    layer4_outputs(7672) <= 1'b1;
    layer4_outputs(7673) <= not b;
    layer4_outputs(7674) <= a or b;
    layer4_outputs(7675) <= b;
    layer4_outputs(7676) <= not (a or b);
    layer4_outputs(7677) <= b;
    layer4_outputs(7678) <= not (a or b);
    layer4_outputs(7679) <= not a;
    layer4_outputs(7680) <= a xor b;
    layer4_outputs(7681) <= not (a or b);
    layer4_outputs(7682) <= 1'b1;
    layer4_outputs(7683) <= a or b;
    layer4_outputs(7684) <= a and not b;
    layer4_outputs(7685) <= b and not a;
    layer4_outputs(7686) <= a and b;
    layer4_outputs(7687) <= b;
    layer4_outputs(7688) <= not (a and b);
    layer4_outputs(7689) <= not (a and b);
    layer4_outputs(7690) <= b and not a;
    layer4_outputs(7691) <= a;
    layer4_outputs(7692) <= 1'b1;
    layer4_outputs(7693) <= a and b;
    layer4_outputs(7694) <= 1'b0;
    layer4_outputs(7695) <= a and b;
    layer4_outputs(7696) <= a;
    layer4_outputs(7697) <= not (a xor b);
    layer4_outputs(7698) <= not b or a;
    layer4_outputs(7699) <= not a or b;
    layer4_outputs(7700) <= a;
    layer4_outputs(7701) <= 1'b1;
    layer4_outputs(7702) <= not a;
    layer4_outputs(7703) <= not a or b;
    layer4_outputs(7704) <= a xor b;
    layer4_outputs(7705) <= a and not b;
    layer4_outputs(7706) <= a and b;
    layer4_outputs(7707) <= a and not b;
    layer4_outputs(7708) <= not a or b;
    layer4_outputs(7709) <= not a or b;
    layer4_outputs(7710) <= not a;
    layer4_outputs(7711) <= not (a and b);
    layer4_outputs(7712) <= a xor b;
    layer4_outputs(7713) <= b and not a;
    layer4_outputs(7714) <= 1'b0;
    layer4_outputs(7715) <= b and not a;
    layer4_outputs(7716) <= 1'b0;
    layer4_outputs(7717) <= a and b;
    layer4_outputs(7718) <= not (a and b);
    layer4_outputs(7719) <= b;
    layer4_outputs(7720) <= not (a and b);
    layer4_outputs(7721) <= b;
    layer4_outputs(7722) <= not b;
    layer4_outputs(7723) <= a;
    layer4_outputs(7724) <= not a or b;
    layer4_outputs(7725) <= not b;
    layer4_outputs(7726) <= not (a and b);
    layer4_outputs(7727) <= not b;
    layer4_outputs(7728) <= 1'b0;
    layer4_outputs(7729) <= not (a and b);
    layer4_outputs(7730) <= a;
    layer4_outputs(7731) <= a xor b;
    layer4_outputs(7732) <= a or b;
    layer4_outputs(7733) <= not b or a;
    layer4_outputs(7734) <= not (a and b);
    layer4_outputs(7735) <= not a;
    layer4_outputs(7736) <= b and not a;
    layer4_outputs(7737) <= not a;
    layer4_outputs(7738) <= not a or b;
    layer4_outputs(7739) <= 1'b1;
    layer4_outputs(7740) <= 1'b0;
    layer4_outputs(7741) <= a or b;
    layer4_outputs(7742) <= not a or b;
    layer4_outputs(7743) <= a and b;
    layer4_outputs(7744) <= not a;
    layer4_outputs(7745) <= 1'b0;
    layer4_outputs(7746) <= a and b;
    layer4_outputs(7747) <= 1'b1;
    layer4_outputs(7748) <= a or b;
    layer4_outputs(7749) <= a;
    layer4_outputs(7750) <= not b;
    layer4_outputs(7751) <= b;
    layer4_outputs(7752) <= not (a or b);
    layer4_outputs(7753) <= a;
    layer4_outputs(7754) <= not b;
    layer4_outputs(7755) <= not (a xor b);
    layer4_outputs(7756) <= 1'b1;
    layer4_outputs(7757) <= b and not a;
    layer4_outputs(7758) <= b and not a;
    layer4_outputs(7759) <= not a;
    layer4_outputs(7760) <= not (a xor b);
    layer4_outputs(7761) <= 1'b1;
    layer4_outputs(7762) <= b;
    layer4_outputs(7763) <= a and b;
    layer4_outputs(7764) <= 1'b0;
    layer4_outputs(7765) <= b and not a;
    layer4_outputs(7766) <= a and b;
    layer4_outputs(7767) <= not b or a;
    layer4_outputs(7768) <= a and not b;
    layer4_outputs(7769) <= a or b;
    layer4_outputs(7770) <= not (a or b);
    layer4_outputs(7771) <= not a or b;
    layer4_outputs(7772) <= not b;
    layer4_outputs(7773) <= b and not a;
    layer4_outputs(7774) <= not (a and b);
    layer4_outputs(7775) <= a or b;
    layer4_outputs(7776) <= b;
    layer4_outputs(7777) <= a xor b;
    layer4_outputs(7778) <= 1'b1;
    layer4_outputs(7779) <= b and not a;
    layer4_outputs(7780) <= 1'b1;
    layer4_outputs(7781) <= a;
    layer4_outputs(7782) <= a;
    layer4_outputs(7783) <= b;
    layer4_outputs(7784) <= 1'b1;
    layer4_outputs(7785) <= a or b;
    layer4_outputs(7786) <= not b or a;
    layer4_outputs(7787) <= not (a or b);
    layer4_outputs(7788) <= not a or b;
    layer4_outputs(7789) <= not (a or b);
    layer4_outputs(7790) <= a and b;
    layer4_outputs(7791) <= 1'b0;
    layer4_outputs(7792) <= a;
    layer4_outputs(7793) <= b and not a;
    layer4_outputs(7794) <= 1'b1;
    layer4_outputs(7795) <= not b;
    layer4_outputs(7796) <= a or b;
    layer4_outputs(7797) <= not (a or b);
    layer4_outputs(7798) <= a;
    layer4_outputs(7799) <= a or b;
    layer4_outputs(7800) <= a;
    layer4_outputs(7801) <= a;
    layer4_outputs(7802) <= not (a and b);
    layer4_outputs(7803) <= a and b;
    layer4_outputs(7804) <= b and not a;
    layer4_outputs(7805) <= not (a or b);
    layer4_outputs(7806) <= a xor b;
    layer4_outputs(7807) <= b and not a;
    layer4_outputs(7808) <= a or b;
    layer4_outputs(7809) <= b and not a;
    layer4_outputs(7810) <= not a or b;
    layer4_outputs(7811) <= 1'b0;
    layer4_outputs(7812) <= 1'b1;
    layer4_outputs(7813) <= not (a and b);
    layer4_outputs(7814) <= a or b;
    layer4_outputs(7815) <= a and not b;
    layer4_outputs(7816) <= not (a or b);
    layer4_outputs(7817) <= a or b;
    layer4_outputs(7818) <= 1'b0;
    layer4_outputs(7819) <= a and not b;
    layer4_outputs(7820) <= a xor b;
    layer4_outputs(7821) <= a xor b;
    layer4_outputs(7822) <= 1'b1;
    layer4_outputs(7823) <= a;
    layer4_outputs(7824) <= a;
    layer4_outputs(7825) <= a or b;
    layer4_outputs(7826) <= not (a or b);
    layer4_outputs(7827) <= a and not b;
    layer4_outputs(7828) <= not b;
    layer4_outputs(7829) <= 1'b0;
    layer4_outputs(7830) <= not (a or b);
    layer4_outputs(7831) <= 1'b0;
    layer4_outputs(7832) <= 1'b1;
    layer4_outputs(7833) <= 1'b1;
    layer4_outputs(7834) <= not b;
    layer4_outputs(7835) <= a xor b;
    layer4_outputs(7836) <= a;
    layer4_outputs(7837) <= 1'b0;
    layer4_outputs(7838) <= a and b;
    layer4_outputs(7839) <= not b or a;
    layer4_outputs(7840) <= a;
    layer4_outputs(7841) <= not (a and b);
    layer4_outputs(7842) <= not a;
    layer4_outputs(7843) <= not b or a;
    layer4_outputs(7844) <= a or b;
    layer4_outputs(7845) <= a and b;
    layer4_outputs(7846) <= 1'b1;
    layer4_outputs(7847) <= 1'b0;
    layer4_outputs(7848) <= b and not a;
    layer4_outputs(7849) <= 1'b1;
    layer4_outputs(7850) <= not b;
    layer4_outputs(7851) <= not (a or b);
    layer4_outputs(7852) <= a;
    layer4_outputs(7853) <= a;
    layer4_outputs(7854) <= 1'b1;
    layer4_outputs(7855) <= b;
    layer4_outputs(7856) <= 1'b0;
    layer4_outputs(7857) <= 1'b0;
    layer4_outputs(7858) <= not a;
    layer4_outputs(7859) <= a and b;
    layer4_outputs(7860) <= b;
    layer4_outputs(7861) <= not b or a;
    layer4_outputs(7862) <= not b or a;
    layer4_outputs(7863) <= a and not b;
    layer4_outputs(7864) <= not a;
    layer4_outputs(7865) <= not b or a;
    layer4_outputs(7866) <= 1'b1;
    layer4_outputs(7867) <= not a or b;
    layer4_outputs(7868) <= b;
    layer4_outputs(7869) <= not b;
    layer4_outputs(7870) <= a and not b;
    layer4_outputs(7871) <= not a;
    layer4_outputs(7872) <= not (a or b);
    layer4_outputs(7873) <= not b;
    layer4_outputs(7874) <= not (a or b);
    layer4_outputs(7875) <= not a;
    layer4_outputs(7876) <= not b;
    layer4_outputs(7877) <= a;
    layer4_outputs(7878) <= 1'b0;
    layer4_outputs(7879) <= not (a and b);
    layer4_outputs(7880) <= not a;
    layer4_outputs(7881) <= not b or a;
    layer4_outputs(7882) <= b;
    layer4_outputs(7883) <= not a;
    layer4_outputs(7884) <= not b;
    layer4_outputs(7885) <= not b;
    layer4_outputs(7886) <= a or b;
    layer4_outputs(7887) <= not (a or b);
    layer4_outputs(7888) <= not a or b;
    layer4_outputs(7889) <= not a or b;
    layer4_outputs(7890) <= not a or b;
    layer4_outputs(7891) <= not (a or b);
    layer4_outputs(7892) <= not b or a;
    layer4_outputs(7893) <= a and b;
    layer4_outputs(7894) <= a or b;
    layer4_outputs(7895) <= a and b;
    layer4_outputs(7896) <= a xor b;
    layer4_outputs(7897) <= b;
    layer4_outputs(7898) <= a;
    layer4_outputs(7899) <= not (a or b);
    layer4_outputs(7900) <= a and b;
    layer4_outputs(7901) <= not (a and b);
    layer4_outputs(7902) <= b and not a;
    layer4_outputs(7903) <= b;
    layer4_outputs(7904) <= a and b;
    layer4_outputs(7905) <= a and b;
    layer4_outputs(7906) <= a;
    layer4_outputs(7907) <= a and not b;
    layer4_outputs(7908) <= b;
    layer4_outputs(7909) <= 1'b1;
    layer4_outputs(7910) <= a and not b;
    layer4_outputs(7911) <= 1'b1;
    layer4_outputs(7912) <= b and not a;
    layer4_outputs(7913) <= not (a and b);
    layer4_outputs(7914) <= 1'b1;
    layer4_outputs(7915) <= not b;
    layer4_outputs(7916) <= 1'b0;
    layer4_outputs(7917) <= a;
    layer4_outputs(7918) <= a xor b;
    layer4_outputs(7919) <= a;
    layer4_outputs(7920) <= a xor b;
    layer4_outputs(7921) <= 1'b0;
    layer4_outputs(7922) <= a;
    layer4_outputs(7923) <= b;
    layer4_outputs(7924) <= a or b;
    layer4_outputs(7925) <= 1'b1;
    layer4_outputs(7926) <= not a or b;
    layer4_outputs(7927) <= a and b;
    layer4_outputs(7928) <= b;
    layer4_outputs(7929) <= not a or b;
    layer4_outputs(7930) <= not a;
    layer4_outputs(7931) <= not (a or b);
    layer4_outputs(7932) <= b;
    layer4_outputs(7933) <= not b;
    layer4_outputs(7934) <= not (a or b);
    layer4_outputs(7935) <= not (a or b);
    layer4_outputs(7936) <= b and not a;
    layer4_outputs(7937) <= 1'b0;
    layer4_outputs(7938) <= not b or a;
    layer4_outputs(7939) <= not (a or b);
    layer4_outputs(7940) <= 1'b1;
    layer4_outputs(7941) <= 1'b0;
    layer4_outputs(7942) <= 1'b1;
    layer4_outputs(7943) <= b;
    layer4_outputs(7944) <= a and b;
    layer4_outputs(7945) <= a and b;
    layer4_outputs(7946) <= not b or a;
    layer4_outputs(7947) <= a and not b;
    layer4_outputs(7948) <= b and not a;
    layer4_outputs(7949) <= not a;
    layer4_outputs(7950) <= a;
    layer4_outputs(7951) <= not (a xor b);
    layer4_outputs(7952) <= not a;
    layer4_outputs(7953) <= a;
    layer4_outputs(7954) <= b and not a;
    layer4_outputs(7955) <= 1'b0;
    layer4_outputs(7956) <= a xor b;
    layer4_outputs(7957) <= a and b;
    layer4_outputs(7958) <= not a;
    layer4_outputs(7959) <= 1'b0;
    layer4_outputs(7960) <= not (a or b);
    layer4_outputs(7961) <= not (a or b);
    layer4_outputs(7962) <= not b;
    layer4_outputs(7963) <= not a;
    layer4_outputs(7964) <= not (a and b);
    layer4_outputs(7965) <= not (a or b);
    layer4_outputs(7966) <= not b or a;
    layer4_outputs(7967) <= 1'b0;
    layer4_outputs(7968) <= not (a and b);
    layer4_outputs(7969) <= 1'b0;
    layer4_outputs(7970) <= not a;
    layer4_outputs(7971) <= not (a or b);
    layer4_outputs(7972) <= not a or b;
    layer4_outputs(7973) <= not b;
    layer4_outputs(7974) <= not a or b;
    layer4_outputs(7975) <= not a or b;
    layer4_outputs(7976) <= not b;
    layer4_outputs(7977) <= not a;
    layer4_outputs(7978) <= a xor b;
    layer4_outputs(7979) <= b;
    layer4_outputs(7980) <= not b;
    layer4_outputs(7981) <= not (a and b);
    layer4_outputs(7982) <= not b;
    layer4_outputs(7983) <= not a or b;
    layer4_outputs(7984) <= not (a and b);
    layer4_outputs(7985) <= a or b;
    layer4_outputs(7986) <= b;
    layer4_outputs(7987) <= not (a and b);
    layer4_outputs(7988) <= a and not b;
    layer4_outputs(7989) <= b and not a;
    layer4_outputs(7990) <= not a;
    layer4_outputs(7991) <= 1'b1;
    layer4_outputs(7992) <= a and not b;
    layer4_outputs(7993) <= a and not b;
    layer4_outputs(7994) <= a and b;
    layer4_outputs(7995) <= a;
    layer4_outputs(7996) <= not (a xor b);
    layer4_outputs(7997) <= not (a or b);
    layer4_outputs(7998) <= a and b;
    layer4_outputs(7999) <= 1'b0;
    layer4_outputs(8000) <= a and b;
    layer4_outputs(8001) <= a or b;
    layer4_outputs(8002) <= 1'b0;
    layer4_outputs(8003) <= a or b;
    layer4_outputs(8004) <= not b;
    layer4_outputs(8005) <= not a;
    layer4_outputs(8006) <= a or b;
    layer4_outputs(8007) <= a and not b;
    layer4_outputs(8008) <= not (a xor b);
    layer4_outputs(8009) <= b and not a;
    layer4_outputs(8010) <= a xor b;
    layer4_outputs(8011) <= 1'b1;
    layer4_outputs(8012) <= a;
    layer4_outputs(8013) <= not b or a;
    layer4_outputs(8014) <= not b or a;
    layer4_outputs(8015) <= not a;
    layer4_outputs(8016) <= not (a and b);
    layer4_outputs(8017) <= a and not b;
    layer4_outputs(8018) <= b and not a;
    layer4_outputs(8019) <= not b;
    layer4_outputs(8020) <= 1'b1;
    layer4_outputs(8021) <= not (a or b);
    layer4_outputs(8022) <= not (a or b);
    layer4_outputs(8023) <= not a;
    layer4_outputs(8024) <= a and b;
    layer4_outputs(8025) <= a xor b;
    layer4_outputs(8026) <= a and not b;
    layer4_outputs(8027) <= a and not b;
    layer4_outputs(8028) <= 1'b0;
    layer4_outputs(8029) <= not (a or b);
    layer4_outputs(8030) <= a or b;
    layer4_outputs(8031) <= not b or a;
    layer4_outputs(8032) <= a or b;
    layer4_outputs(8033) <= not a;
    layer4_outputs(8034) <= b and not a;
    layer4_outputs(8035) <= 1'b0;
    layer4_outputs(8036) <= not b or a;
    layer4_outputs(8037) <= a xor b;
    layer4_outputs(8038) <= not b;
    layer4_outputs(8039) <= a and b;
    layer4_outputs(8040) <= a;
    layer4_outputs(8041) <= 1'b0;
    layer4_outputs(8042) <= not a or b;
    layer4_outputs(8043) <= a;
    layer4_outputs(8044) <= a and b;
    layer4_outputs(8045) <= a and b;
    layer4_outputs(8046) <= a or b;
    layer4_outputs(8047) <= a or b;
    layer4_outputs(8048) <= not a;
    layer4_outputs(8049) <= 1'b0;
    layer4_outputs(8050) <= b and not a;
    layer4_outputs(8051) <= a;
    layer4_outputs(8052) <= 1'b0;
    layer4_outputs(8053) <= a;
    layer4_outputs(8054) <= not (a xor b);
    layer4_outputs(8055) <= not b or a;
    layer4_outputs(8056) <= b;
    layer4_outputs(8057) <= not b;
    layer4_outputs(8058) <= not a;
    layer4_outputs(8059) <= a or b;
    layer4_outputs(8060) <= 1'b1;
    layer4_outputs(8061) <= a;
    layer4_outputs(8062) <= a and not b;
    layer4_outputs(8063) <= not (a and b);
    layer4_outputs(8064) <= not b;
    layer4_outputs(8065) <= not a or b;
    layer4_outputs(8066) <= not (a and b);
    layer4_outputs(8067) <= a and b;
    layer4_outputs(8068) <= a;
    layer4_outputs(8069) <= not (a and b);
    layer4_outputs(8070) <= not b;
    layer4_outputs(8071) <= a and b;
    layer4_outputs(8072) <= b and not a;
    layer4_outputs(8073) <= a and not b;
    layer4_outputs(8074) <= not a;
    layer4_outputs(8075) <= b;
    layer4_outputs(8076) <= 1'b1;
    layer4_outputs(8077) <= not (a and b);
    layer4_outputs(8078) <= not (a and b);
    layer4_outputs(8079) <= b;
    layer4_outputs(8080) <= not (a and b);
    layer4_outputs(8081) <= a or b;
    layer4_outputs(8082) <= not a;
    layer4_outputs(8083) <= not b;
    layer4_outputs(8084) <= b;
    layer4_outputs(8085) <= b;
    layer4_outputs(8086) <= not a or b;
    layer4_outputs(8087) <= a;
    layer4_outputs(8088) <= b;
    layer4_outputs(8089) <= not a or b;
    layer4_outputs(8090) <= a xor b;
    layer4_outputs(8091) <= b and not a;
    layer4_outputs(8092) <= not a or b;
    layer4_outputs(8093) <= b;
    layer4_outputs(8094) <= a xor b;
    layer4_outputs(8095) <= a and b;
    layer4_outputs(8096) <= not (a and b);
    layer4_outputs(8097) <= b;
    layer4_outputs(8098) <= not a or b;
    layer4_outputs(8099) <= not b;
    layer4_outputs(8100) <= a;
    layer4_outputs(8101) <= a xor b;
    layer4_outputs(8102) <= not (a or b);
    layer4_outputs(8103) <= a and b;
    layer4_outputs(8104) <= not b or a;
    layer4_outputs(8105) <= a xor b;
    layer4_outputs(8106) <= not (a or b);
    layer4_outputs(8107) <= b and not a;
    layer4_outputs(8108) <= not (a or b);
    layer4_outputs(8109) <= not b or a;
    layer4_outputs(8110) <= not a;
    layer4_outputs(8111) <= not b or a;
    layer4_outputs(8112) <= a and b;
    layer4_outputs(8113) <= 1'b1;
    layer4_outputs(8114) <= not (a and b);
    layer4_outputs(8115) <= b;
    layer4_outputs(8116) <= a;
    layer4_outputs(8117) <= a and b;
    layer4_outputs(8118) <= a xor b;
    layer4_outputs(8119) <= a or b;
    layer4_outputs(8120) <= a and not b;
    layer4_outputs(8121) <= not b or a;
    layer4_outputs(8122) <= not (a or b);
    layer4_outputs(8123) <= a;
    layer4_outputs(8124) <= 1'b0;
    layer4_outputs(8125) <= a and b;
    layer4_outputs(8126) <= b and not a;
    layer4_outputs(8127) <= not b;
    layer4_outputs(8128) <= not b;
    layer4_outputs(8129) <= not b or a;
    layer4_outputs(8130) <= a and b;
    layer4_outputs(8131) <= not b;
    layer4_outputs(8132) <= 1'b1;
    layer4_outputs(8133) <= not b or a;
    layer4_outputs(8134) <= not (a xor b);
    layer4_outputs(8135) <= a;
    layer4_outputs(8136) <= not a;
    layer4_outputs(8137) <= not (a xor b);
    layer4_outputs(8138) <= a and b;
    layer4_outputs(8139) <= not a;
    layer4_outputs(8140) <= not a or b;
    layer4_outputs(8141) <= not (a and b);
    layer4_outputs(8142) <= 1'b1;
    layer4_outputs(8143) <= not (a and b);
    layer4_outputs(8144) <= b and not a;
    layer4_outputs(8145) <= a and not b;
    layer4_outputs(8146) <= b;
    layer4_outputs(8147) <= not a;
    layer4_outputs(8148) <= 1'b0;
    layer4_outputs(8149) <= a and not b;
    layer4_outputs(8150) <= a or b;
    layer4_outputs(8151) <= a and b;
    layer4_outputs(8152) <= a xor b;
    layer4_outputs(8153) <= not b;
    layer4_outputs(8154) <= not a;
    layer4_outputs(8155) <= b;
    layer4_outputs(8156) <= not a or b;
    layer4_outputs(8157) <= a and not b;
    layer4_outputs(8158) <= not (a or b);
    layer4_outputs(8159) <= 1'b1;
    layer4_outputs(8160) <= 1'b0;
    layer4_outputs(8161) <= a and not b;
    layer4_outputs(8162) <= not a or b;
    layer4_outputs(8163) <= not (a and b);
    layer4_outputs(8164) <= not a or b;
    layer4_outputs(8165) <= a or b;
    layer4_outputs(8166) <= a;
    layer4_outputs(8167) <= not (a xor b);
    layer4_outputs(8168) <= b;
    layer4_outputs(8169) <= not b;
    layer4_outputs(8170) <= a and not b;
    layer4_outputs(8171) <= not a;
    layer4_outputs(8172) <= 1'b1;
    layer4_outputs(8173) <= a and b;
    layer4_outputs(8174) <= not a or b;
    layer4_outputs(8175) <= 1'b1;
    layer4_outputs(8176) <= not a;
    layer4_outputs(8177) <= not (a and b);
    layer4_outputs(8178) <= b and not a;
    layer4_outputs(8179) <= a or b;
    layer4_outputs(8180) <= not a;
    layer4_outputs(8181) <= not a or b;
    layer4_outputs(8182) <= not (a xor b);
    layer4_outputs(8183) <= b and not a;
    layer4_outputs(8184) <= b;
    layer4_outputs(8185) <= not a or b;
    layer4_outputs(8186) <= not b;
    layer4_outputs(8187) <= 1'b1;
    layer4_outputs(8188) <= not a or b;
    layer4_outputs(8189) <= 1'b1;
    layer4_outputs(8190) <= not b;
    layer4_outputs(8191) <= not (a and b);
    layer4_outputs(8192) <= not a;
    layer4_outputs(8193) <= a;
    layer4_outputs(8194) <= a or b;
    layer4_outputs(8195) <= a and b;
    layer4_outputs(8196) <= a or b;
    layer4_outputs(8197) <= a and not b;
    layer4_outputs(8198) <= 1'b1;
    layer4_outputs(8199) <= b and not a;
    layer4_outputs(8200) <= not b or a;
    layer4_outputs(8201) <= 1'b1;
    layer4_outputs(8202) <= not b;
    layer4_outputs(8203) <= a xor b;
    layer4_outputs(8204) <= a or b;
    layer4_outputs(8205) <= not (a and b);
    layer4_outputs(8206) <= a and b;
    layer4_outputs(8207) <= not a;
    layer4_outputs(8208) <= not b or a;
    layer4_outputs(8209) <= not b;
    layer4_outputs(8210) <= 1'b1;
    layer4_outputs(8211) <= a and b;
    layer4_outputs(8212) <= a or b;
    layer4_outputs(8213) <= b and not a;
    layer4_outputs(8214) <= not b;
    layer4_outputs(8215) <= 1'b1;
    layer4_outputs(8216) <= b;
    layer4_outputs(8217) <= not (a and b);
    layer4_outputs(8218) <= a or b;
    layer4_outputs(8219) <= not (a xor b);
    layer4_outputs(8220) <= not (a xor b);
    layer4_outputs(8221) <= a and not b;
    layer4_outputs(8222) <= a or b;
    layer4_outputs(8223) <= not (a or b);
    layer4_outputs(8224) <= 1'b1;
    layer4_outputs(8225) <= b and not a;
    layer4_outputs(8226) <= 1'b0;
    layer4_outputs(8227) <= not b;
    layer4_outputs(8228) <= a and b;
    layer4_outputs(8229) <= a or b;
    layer4_outputs(8230) <= not a or b;
    layer4_outputs(8231) <= b;
    layer4_outputs(8232) <= a;
    layer4_outputs(8233) <= not (a or b);
    layer4_outputs(8234) <= b;
    layer4_outputs(8235) <= a and not b;
    layer4_outputs(8236) <= not a or b;
    layer4_outputs(8237) <= not (a and b);
    layer4_outputs(8238) <= a;
    layer4_outputs(8239) <= a;
    layer4_outputs(8240) <= b and not a;
    layer4_outputs(8241) <= not (a xor b);
    layer4_outputs(8242) <= b;
    layer4_outputs(8243) <= b;
    layer4_outputs(8244) <= not a;
    layer4_outputs(8245) <= not a;
    layer4_outputs(8246) <= not a or b;
    layer4_outputs(8247) <= a;
    layer4_outputs(8248) <= a and b;
    layer4_outputs(8249) <= not a or b;
    layer4_outputs(8250) <= b and not a;
    layer4_outputs(8251) <= a and not b;
    layer4_outputs(8252) <= not b;
    layer4_outputs(8253) <= not (a or b);
    layer4_outputs(8254) <= not a;
    layer4_outputs(8255) <= not (a or b);
    layer4_outputs(8256) <= a xor b;
    layer4_outputs(8257) <= 1'b0;
    layer4_outputs(8258) <= a xor b;
    layer4_outputs(8259) <= not (a or b);
    layer4_outputs(8260) <= not (a or b);
    layer4_outputs(8261) <= a or b;
    layer4_outputs(8262) <= not b;
    layer4_outputs(8263) <= a and not b;
    layer4_outputs(8264) <= not a or b;
    layer4_outputs(8265) <= a and b;
    layer4_outputs(8266) <= 1'b0;
    layer4_outputs(8267) <= b;
    layer4_outputs(8268) <= a;
    layer4_outputs(8269) <= b;
    layer4_outputs(8270) <= 1'b0;
    layer4_outputs(8271) <= a;
    layer4_outputs(8272) <= not (a xor b);
    layer4_outputs(8273) <= not a or b;
    layer4_outputs(8274) <= a or b;
    layer4_outputs(8275) <= not a or b;
    layer4_outputs(8276) <= b and not a;
    layer4_outputs(8277) <= a and b;
    layer4_outputs(8278) <= not b;
    layer4_outputs(8279) <= a or b;
    layer4_outputs(8280) <= not b;
    layer4_outputs(8281) <= not (a or b);
    layer4_outputs(8282) <= b;
    layer4_outputs(8283) <= not (a xor b);
    layer4_outputs(8284) <= not (a and b);
    layer4_outputs(8285) <= a xor b;
    layer4_outputs(8286) <= 1'b0;
    layer4_outputs(8287) <= not a;
    layer4_outputs(8288) <= 1'b1;
    layer4_outputs(8289) <= not a;
    layer4_outputs(8290) <= not b;
    layer4_outputs(8291) <= b and not a;
    layer4_outputs(8292) <= not a;
    layer4_outputs(8293) <= b and not a;
    layer4_outputs(8294) <= a xor b;
    layer4_outputs(8295) <= not (a and b);
    layer4_outputs(8296) <= a and not b;
    layer4_outputs(8297) <= b;
    layer4_outputs(8298) <= a and b;
    layer4_outputs(8299) <= not (a and b);
    layer4_outputs(8300) <= b;
    layer4_outputs(8301) <= not a or b;
    layer4_outputs(8302) <= a or b;
    layer4_outputs(8303) <= b and not a;
    layer4_outputs(8304) <= not (a or b);
    layer4_outputs(8305) <= not (a or b);
    layer4_outputs(8306) <= not a or b;
    layer4_outputs(8307) <= 1'b0;
    layer4_outputs(8308) <= a;
    layer4_outputs(8309) <= b;
    layer4_outputs(8310) <= a and b;
    layer4_outputs(8311) <= 1'b1;
    layer4_outputs(8312) <= 1'b0;
    layer4_outputs(8313) <= not a or b;
    layer4_outputs(8314) <= not a;
    layer4_outputs(8315) <= not b;
    layer4_outputs(8316) <= not a;
    layer4_outputs(8317) <= a and not b;
    layer4_outputs(8318) <= not b;
    layer4_outputs(8319) <= a or b;
    layer4_outputs(8320) <= b and not a;
    layer4_outputs(8321) <= a;
    layer4_outputs(8322) <= b and not a;
    layer4_outputs(8323) <= not (a and b);
    layer4_outputs(8324) <= 1'b0;
    layer4_outputs(8325) <= 1'b1;
    layer4_outputs(8326) <= b;
    layer4_outputs(8327) <= 1'b1;
    layer4_outputs(8328) <= b;
    layer4_outputs(8329) <= b;
    layer4_outputs(8330) <= 1'b1;
    layer4_outputs(8331) <= not b or a;
    layer4_outputs(8332) <= not b;
    layer4_outputs(8333) <= a and not b;
    layer4_outputs(8334) <= not b or a;
    layer4_outputs(8335) <= not (a or b);
    layer4_outputs(8336) <= b;
    layer4_outputs(8337) <= not b;
    layer4_outputs(8338) <= a or b;
    layer4_outputs(8339) <= not a;
    layer4_outputs(8340) <= b;
    layer4_outputs(8341) <= not a;
    layer4_outputs(8342) <= a;
    layer4_outputs(8343) <= 1'b0;
    layer4_outputs(8344) <= b;
    layer4_outputs(8345) <= not (a and b);
    layer4_outputs(8346) <= 1'b1;
    layer4_outputs(8347) <= a;
    layer4_outputs(8348) <= 1'b1;
    layer4_outputs(8349) <= 1'b0;
    layer4_outputs(8350) <= 1'b0;
    layer4_outputs(8351) <= b and not a;
    layer4_outputs(8352) <= not b;
    layer4_outputs(8353) <= a or b;
    layer4_outputs(8354) <= a;
    layer4_outputs(8355) <= b;
    layer4_outputs(8356) <= not (a xor b);
    layer4_outputs(8357) <= a and not b;
    layer4_outputs(8358) <= b and not a;
    layer4_outputs(8359) <= b and not a;
    layer4_outputs(8360) <= not (a or b);
    layer4_outputs(8361) <= not b or a;
    layer4_outputs(8362) <= 1'b1;
    layer4_outputs(8363) <= 1'b1;
    layer4_outputs(8364) <= not (a or b);
    layer4_outputs(8365) <= a and not b;
    layer4_outputs(8366) <= not a;
    layer4_outputs(8367) <= not b;
    layer4_outputs(8368) <= not (a and b);
    layer4_outputs(8369) <= not b;
    layer4_outputs(8370) <= a xor b;
    layer4_outputs(8371) <= 1'b1;
    layer4_outputs(8372) <= not (a or b);
    layer4_outputs(8373) <= not a;
    layer4_outputs(8374) <= not b or a;
    layer4_outputs(8375) <= not b;
    layer4_outputs(8376) <= a and b;
    layer4_outputs(8377) <= not (a xor b);
    layer4_outputs(8378) <= not (a or b);
    layer4_outputs(8379) <= not b or a;
    layer4_outputs(8380) <= not (a xor b);
    layer4_outputs(8381) <= a and not b;
    layer4_outputs(8382) <= b and not a;
    layer4_outputs(8383) <= not a or b;
    layer4_outputs(8384) <= b;
    layer4_outputs(8385) <= b;
    layer4_outputs(8386) <= not a;
    layer4_outputs(8387) <= not a;
    layer4_outputs(8388) <= b and not a;
    layer4_outputs(8389) <= a and b;
    layer4_outputs(8390) <= not a or b;
    layer4_outputs(8391) <= not (a or b);
    layer4_outputs(8392) <= 1'b0;
    layer4_outputs(8393) <= a or b;
    layer4_outputs(8394) <= 1'b0;
    layer4_outputs(8395) <= a;
    layer4_outputs(8396) <= not (a and b);
    layer4_outputs(8397) <= not a;
    layer4_outputs(8398) <= b and not a;
    layer4_outputs(8399) <= b;
    layer4_outputs(8400) <= not a;
    layer4_outputs(8401) <= 1'b0;
    layer4_outputs(8402) <= b and not a;
    layer4_outputs(8403) <= not a;
    layer4_outputs(8404) <= a and b;
    layer4_outputs(8405) <= not b;
    layer4_outputs(8406) <= not a or b;
    layer4_outputs(8407) <= not a;
    layer4_outputs(8408) <= not (a xor b);
    layer4_outputs(8409) <= not a or b;
    layer4_outputs(8410) <= a;
    layer4_outputs(8411) <= a;
    layer4_outputs(8412) <= b and not a;
    layer4_outputs(8413) <= not a;
    layer4_outputs(8414) <= b;
    layer4_outputs(8415) <= not b;
    layer4_outputs(8416) <= a and not b;
    layer4_outputs(8417) <= a and b;
    layer4_outputs(8418) <= not b;
    layer4_outputs(8419) <= not a;
    layer4_outputs(8420) <= not a;
    layer4_outputs(8421) <= not (a or b);
    layer4_outputs(8422) <= not a;
    layer4_outputs(8423) <= a and b;
    layer4_outputs(8424) <= b;
    layer4_outputs(8425) <= a;
    layer4_outputs(8426) <= not (a and b);
    layer4_outputs(8427) <= a xor b;
    layer4_outputs(8428) <= 1'b0;
    layer4_outputs(8429) <= not b;
    layer4_outputs(8430) <= not a or b;
    layer4_outputs(8431) <= not (a or b);
    layer4_outputs(8432) <= not (a or b);
    layer4_outputs(8433) <= not b;
    layer4_outputs(8434) <= b;
    layer4_outputs(8435) <= not b;
    layer4_outputs(8436) <= not b or a;
    layer4_outputs(8437) <= not a or b;
    layer4_outputs(8438) <= 1'b0;
    layer4_outputs(8439) <= a and b;
    layer4_outputs(8440) <= a or b;
    layer4_outputs(8441) <= not b;
    layer4_outputs(8442) <= a and not b;
    layer4_outputs(8443) <= not a or b;
    layer4_outputs(8444) <= not b or a;
    layer4_outputs(8445) <= a and not b;
    layer4_outputs(8446) <= a and not b;
    layer4_outputs(8447) <= not b or a;
    layer4_outputs(8448) <= a xor b;
    layer4_outputs(8449) <= b;
    layer4_outputs(8450) <= not b;
    layer4_outputs(8451) <= a;
    layer4_outputs(8452) <= not a or b;
    layer4_outputs(8453) <= not b;
    layer4_outputs(8454) <= a;
    layer4_outputs(8455) <= 1'b0;
    layer4_outputs(8456) <= not a or b;
    layer4_outputs(8457) <= 1'b0;
    layer4_outputs(8458) <= not a;
    layer4_outputs(8459) <= a and b;
    layer4_outputs(8460) <= 1'b0;
    layer4_outputs(8461) <= a and not b;
    layer4_outputs(8462) <= not b or a;
    layer4_outputs(8463) <= a and b;
    layer4_outputs(8464) <= a and b;
    layer4_outputs(8465) <= not a or b;
    layer4_outputs(8466) <= not a or b;
    layer4_outputs(8467) <= a or b;
    layer4_outputs(8468) <= 1'b1;
    layer4_outputs(8469) <= a;
    layer4_outputs(8470) <= not a or b;
    layer4_outputs(8471) <= 1'b0;
    layer4_outputs(8472) <= not a;
    layer4_outputs(8473) <= a and b;
    layer4_outputs(8474) <= a;
    layer4_outputs(8475) <= b and not a;
    layer4_outputs(8476) <= b;
    layer4_outputs(8477) <= 1'b0;
    layer4_outputs(8478) <= a and b;
    layer4_outputs(8479) <= b;
    layer4_outputs(8480) <= b;
    layer4_outputs(8481) <= not a;
    layer4_outputs(8482) <= 1'b0;
    layer4_outputs(8483) <= not (a and b);
    layer4_outputs(8484) <= a and b;
    layer4_outputs(8485) <= b and not a;
    layer4_outputs(8486) <= not b;
    layer4_outputs(8487) <= a;
    layer4_outputs(8488) <= 1'b0;
    layer4_outputs(8489) <= 1'b1;
    layer4_outputs(8490) <= a or b;
    layer4_outputs(8491) <= not a or b;
    layer4_outputs(8492) <= not (a or b);
    layer4_outputs(8493) <= 1'b1;
    layer4_outputs(8494) <= not (a xor b);
    layer4_outputs(8495) <= not a or b;
    layer4_outputs(8496) <= a and b;
    layer4_outputs(8497) <= b and not a;
    layer4_outputs(8498) <= not (a or b);
    layer4_outputs(8499) <= b and not a;
    layer4_outputs(8500) <= not (a or b);
    layer4_outputs(8501) <= a or b;
    layer4_outputs(8502) <= not b;
    layer4_outputs(8503) <= not a or b;
    layer4_outputs(8504) <= a or b;
    layer4_outputs(8505) <= a and b;
    layer4_outputs(8506) <= b and not a;
    layer4_outputs(8507) <= b;
    layer4_outputs(8508) <= not (a or b);
    layer4_outputs(8509) <= not b;
    layer4_outputs(8510) <= b and not a;
    layer4_outputs(8511) <= a and not b;
    layer4_outputs(8512) <= not a or b;
    layer4_outputs(8513) <= b and not a;
    layer4_outputs(8514) <= 1'b0;
    layer4_outputs(8515) <= not (a or b);
    layer4_outputs(8516) <= 1'b1;
    layer4_outputs(8517) <= not b;
    layer4_outputs(8518) <= b and not a;
    layer4_outputs(8519) <= a;
    layer4_outputs(8520) <= 1'b1;
    layer4_outputs(8521) <= not b;
    layer4_outputs(8522) <= a xor b;
    layer4_outputs(8523) <= not (a or b);
    layer4_outputs(8524) <= a or b;
    layer4_outputs(8525) <= not a or b;
    layer4_outputs(8526) <= not (a or b);
    layer4_outputs(8527) <= b;
    layer4_outputs(8528) <= a xor b;
    layer4_outputs(8529) <= b and not a;
    layer4_outputs(8530) <= a and not b;
    layer4_outputs(8531) <= 1'b1;
    layer4_outputs(8532) <= a and not b;
    layer4_outputs(8533) <= a;
    layer4_outputs(8534) <= not a or b;
    layer4_outputs(8535) <= b;
    layer4_outputs(8536) <= a;
    layer4_outputs(8537) <= a and not b;
    layer4_outputs(8538) <= not (a or b);
    layer4_outputs(8539) <= b;
    layer4_outputs(8540) <= b;
    layer4_outputs(8541) <= b and not a;
    layer4_outputs(8542) <= b;
    layer4_outputs(8543) <= b;
    layer4_outputs(8544) <= not b;
    layer4_outputs(8545) <= not (a and b);
    layer4_outputs(8546) <= a;
    layer4_outputs(8547) <= a and not b;
    layer4_outputs(8548) <= a and not b;
    layer4_outputs(8549) <= 1'b0;
    layer4_outputs(8550) <= b;
    layer4_outputs(8551) <= not b or a;
    layer4_outputs(8552) <= a;
    layer4_outputs(8553) <= b and not a;
    layer4_outputs(8554) <= not (a or b);
    layer4_outputs(8555) <= 1'b0;
    layer4_outputs(8556) <= a and not b;
    layer4_outputs(8557) <= not a;
    layer4_outputs(8558) <= a;
    layer4_outputs(8559) <= not a or b;
    layer4_outputs(8560) <= a and b;
    layer4_outputs(8561) <= not b;
    layer4_outputs(8562) <= 1'b0;
    layer4_outputs(8563) <= 1'b1;
    layer4_outputs(8564) <= not (a or b);
    layer4_outputs(8565) <= a and b;
    layer4_outputs(8566) <= b;
    layer4_outputs(8567) <= not b;
    layer4_outputs(8568) <= b;
    layer4_outputs(8569) <= not a or b;
    layer4_outputs(8570) <= not b;
    layer4_outputs(8571) <= 1'b0;
    layer4_outputs(8572) <= 1'b1;
    layer4_outputs(8573) <= a;
    layer4_outputs(8574) <= b and not a;
    layer4_outputs(8575) <= not a;
    layer4_outputs(8576) <= b;
    layer4_outputs(8577) <= b;
    layer4_outputs(8578) <= not (a and b);
    layer4_outputs(8579) <= not b or a;
    layer4_outputs(8580) <= not a or b;
    layer4_outputs(8581) <= 1'b1;
    layer4_outputs(8582) <= not a or b;
    layer4_outputs(8583) <= not (a and b);
    layer4_outputs(8584) <= not (a and b);
    layer4_outputs(8585) <= a xor b;
    layer4_outputs(8586) <= a or b;
    layer4_outputs(8587) <= a or b;
    layer4_outputs(8588) <= not b or a;
    layer4_outputs(8589) <= 1'b0;
    layer4_outputs(8590) <= a and not b;
    layer4_outputs(8591) <= not b;
    layer4_outputs(8592) <= a xor b;
    layer4_outputs(8593) <= 1'b1;
    layer4_outputs(8594) <= 1'b0;
    layer4_outputs(8595) <= a or b;
    layer4_outputs(8596) <= not (a or b);
    layer4_outputs(8597) <= a and b;
    layer4_outputs(8598) <= not (a and b);
    layer4_outputs(8599) <= not (a xor b);
    layer4_outputs(8600) <= b and not a;
    layer4_outputs(8601) <= not (a or b);
    layer4_outputs(8602) <= not b or a;
    layer4_outputs(8603) <= a or b;
    layer4_outputs(8604) <= 1'b1;
    layer4_outputs(8605) <= a;
    layer4_outputs(8606) <= not b or a;
    layer4_outputs(8607) <= a or b;
    layer4_outputs(8608) <= b and not a;
    layer4_outputs(8609) <= a;
    layer4_outputs(8610) <= not (a or b);
    layer4_outputs(8611) <= not b;
    layer4_outputs(8612) <= 1'b0;
    layer4_outputs(8613) <= not a;
    layer4_outputs(8614) <= b and not a;
    layer4_outputs(8615) <= not b;
    layer4_outputs(8616) <= b;
    layer4_outputs(8617) <= 1'b1;
    layer4_outputs(8618) <= a;
    layer4_outputs(8619) <= a and not b;
    layer4_outputs(8620) <= not b or a;
    layer4_outputs(8621) <= not (a and b);
    layer4_outputs(8622) <= not b;
    layer4_outputs(8623) <= not a;
    layer4_outputs(8624) <= a and not b;
    layer4_outputs(8625) <= a and not b;
    layer4_outputs(8626) <= a;
    layer4_outputs(8627) <= not b;
    layer4_outputs(8628) <= not a or b;
    layer4_outputs(8629) <= not b or a;
    layer4_outputs(8630) <= not (a or b);
    layer4_outputs(8631) <= not b;
    layer4_outputs(8632) <= b and not a;
    layer4_outputs(8633) <= not b;
    layer4_outputs(8634) <= not (a xor b);
    layer4_outputs(8635) <= a;
    layer4_outputs(8636) <= a or b;
    layer4_outputs(8637) <= a;
    layer4_outputs(8638) <= not b or a;
    layer4_outputs(8639) <= not a;
    layer4_outputs(8640) <= a and not b;
    layer4_outputs(8641) <= a;
    layer4_outputs(8642) <= not b;
    layer4_outputs(8643) <= not (a or b);
    layer4_outputs(8644) <= a and b;
    layer4_outputs(8645) <= not b;
    layer4_outputs(8646) <= a or b;
    layer4_outputs(8647) <= b and not a;
    layer4_outputs(8648) <= not (a or b);
    layer4_outputs(8649) <= a and not b;
    layer4_outputs(8650) <= not a;
    layer4_outputs(8651) <= b and not a;
    layer4_outputs(8652) <= b;
    layer4_outputs(8653) <= b and not a;
    layer4_outputs(8654) <= a;
    layer4_outputs(8655) <= a;
    layer4_outputs(8656) <= a or b;
    layer4_outputs(8657) <= not a;
    layer4_outputs(8658) <= a or b;
    layer4_outputs(8659) <= a and not b;
    layer4_outputs(8660) <= a and b;
    layer4_outputs(8661) <= not (a and b);
    layer4_outputs(8662) <= b;
    layer4_outputs(8663) <= a or b;
    layer4_outputs(8664) <= b;
    layer4_outputs(8665) <= not b or a;
    layer4_outputs(8666) <= not b;
    layer4_outputs(8667) <= a or b;
    layer4_outputs(8668) <= not (a and b);
    layer4_outputs(8669) <= not (a and b);
    layer4_outputs(8670) <= not a;
    layer4_outputs(8671) <= b and not a;
    layer4_outputs(8672) <= not a or b;
    layer4_outputs(8673) <= not a;
    layer4_outputs(8674) <= a or b;
    layer4_outputs(8675) <= a and not b;
    layer4_outputs(8676) <= not b;
    layer4_outputs(8677) <= a or b;
    layer4_outputs(8678) <= not (a and b);
    layer4_outputs(8679) <= not b;
    layer4_outputs(8680) <= not b;
    layer4_outputs(8681) <= 1'b0;
    layer4_outputs(8682) <= b;
    layer4_outputs(8683) <= a and not b;
    layer4_outputs(8684) <= not b;
    layer4_outputs(8685) <= a and not b;
    layer4_outputs(8686) <= a and b;
    layer4_outputs(8687) <= a;
    layer4_outputs(8688) <= not b or a;
    layer4_outputs(8689) <= not a or b;
    layer4_outputs(8690) <= a and not b;
    layer4_outputs(8691) <= not a;
    layer4_outputs(8692) <= b and not a;
    layer4_outputs(8693) <= 1'b0;
    layer4_outputs(8694) <= a;
    layer4_outputs(8695) <= not (a and b);
    layer4_outputs(8696) <= 1'b0;
    layer4_outputs(8697) <= not b;
    layer4_outputs(8698) <= b;
    layer4_outputs(8699) <= not b or a;
    layer4_outputs(8700) <= not (a or b);
    layer4_outputs(8701) <= a and not b;
    layer4_outputs(8702) <= a and not b;
    layer4_outputs(8703) <= not b or a;
    layer4_outputs(8704) <= a and b;
    layer4_outputs(8705) <= not a;
    layer4_outputs(8706) <= a;
    layer4_outputs(8707) <= not a;
    layer4_outputs(8708) <= not (a or b);
    layer4_outputs(8709) <= a;
    layer4_outputs(8710) <= a or b;
    layer4_outputs(8711) <= not b or a;
    layer4_outputs(8712) <= a and not b;
    layer4_outputs(8713) <= a and b;
    layer4_outputs(8714) <= a and not b;
    layer4_outputs(8715) <= a or b;
    layer4_outputs(8716) <= 1'b1;
    layer4_outputs(8717) <= not a or b;
    layer4_outputs(8718) <= not b;
    layer4_outputs(8719) <= not b or a;
    layer4_outputs(8720) <= a and not b;
    layer4_outputs(8721) <= a or b;
    layer4_outputs(8722) <= not a;
    layer4_outputs(8723) <= not a;
    layer4_outputs(8724) <= b;
    layer4_outputs(8725) <= 1'b0;
    layer4_outputs(8726) <= a xor b;
    layer4_outputs(8727) <= 1'b1;
    layer4_outputs(8728) <= a or b;
    layer4_outputs(8729) <= a and not b;
    layer4_outputs(8730) <= not (a and b);
    layer4_outputs(8731) <= b;
    layer4_outputs(8732) <= not b or a;
    layer4_outputs(8733) <= not a or b;
    layer4_outputs(8734) <= b;
    layer4_outputs(8735) <= a and b;
    layer4_outputs(8736) <= 1'b0;
    layer4_outputs(8737) <= b and not a;
    layer4_outputs(8738) <= a or b;
    layer4_outputs(8739) <= a and not b;
    layer4_outputs(8740) <= b and not a;
    layer4_outputs(8741) <= 1'b0;
    layer4_outputs(8742) <= b and not a;
    layer4_outputs(8743) <= b;
    layer4_outputs(8744) <= a;
    layer4_outputs(8745) <= a and b;
    layer4_outputs(8746) <= b and not a;
    layer4_outputs(8747) <= 1'b1;
    layer4_outputs(8748) <= not (a and b);
    layer4_outputs(8749) <= not (a or b);
    layer4_outputs(8750) <= not (a and b);
    layer4_outputs(8751) <= not a;
    layer4_outputs(8752) <= not a or b;
    layer4_outputs(8753) <= not (a and b);
    layer4_outputs(8754) <= not b;
    layer4_outputs(8755) <= not b;
    layer4_outputs(8756) <= not (a or b);
    layer4_outputs(8757) <= not b or a;
    layer4_outputs(8758) <= b;
    layer4_outputs(8759) <= not (a or b);
    layer4_outputs(8760) <= not b or a;
    layer4_outputs(8761) <= a or b;
    layer4_outputs(8762) <= not a or b;
    layer4_outputs(8763) <= 1'b0;
    layer4_outputs(8764) <= a and not b;
    layer4_outputs(8765) <= not b;
    layer4_outputs(8766) <= not a;
    layer4_outputs(8767) <= a and b;
    layer4_outputs(8768) <= a and b;
    layer4_outputs(8769) <= not b;
    layer4_outputs(8770) <= not (a or b);
    layer4_outputs(8771) <= not a or b;
    layer4_outputs(8772) <= not (a xor b);
    layer4_outputs(8773) <= 1'b1;
    layer4_outputs(8774) <= a;
    layer4_outputs(8775) <= b and not a;
    layer4_outputs(8776) <= not a;
    layer4_outputs(8777) <= b and not a;
    layer4_outputs(8778) <= not (a and b);
    layer4_outputs(8779) <= not (a and b);
    layer4_outputs(8780) <= a or b;
    layer4_outputs(8781) <= not (a and b);
    layer4_outputs(8782) <= a and b;
    layer4_outputs(8783) <= not (a or b);
    layer4_outputs(8784) <= 1'b0;
    layer4_outputs(8785) <= a and b;
    layer4_outputs(8786) <= b and not a;
    layer4_outputs(8787) <= b and not a;
    layer4_outputs(8788) <= not (a xor b);
    layer4_outputs(8789) <= a;
    layer4_outputs(8790) <= a and not b;
    layer4_outputs(8791) <= a;
    layer4_outputs(8792) <= 1'b1;
    layer4_outputs(8793) <= 1'b1;
    layer4_outputs(8794) <= 1'b0;
    layer4_outputs(8795) <= not (a or b);
    layer4_outputs(8796) <= 1'b1;
    layer4_outputs(8797) <= not (a and b);
    layer4_outputs(8798) <= 1'b0;
    layer4_outputs(8799) <= b;
    layer4_outputs(8800) <= a or b;
    layer4_outputs(8801) <= 1'b1;
    layer4_outputs(8802) <= a or b;
    layer4_outputs(8803) <= not a or b;
    layer4_outputs(8804) <= not (a or b);
    layer4_outputs(8805) <= 1'b1;
    layer4_outputs(8806) <= not a or b;
    layer4_outputs(8807) <= a and b;
    layer4_outputs(8808) <= not a or b;
    layer4_outputs(8809) <= not b or a;
    layer4_outputs(8810) <= a;
    layer4_outputs(8811) <= b;
    layer4_outputs(8812) <= not a or b;
    layer4_outputs(8813) <= a and not b;
    layer4_outputs(8814) <= a or b;
    layer4_outputs(8815) <= a;
    layer4_outputs(8816) <= a;
    layer4_outputs(8817) <= a;
    layer4_outputs(8818) <= not a or b;
    layer4_outputs(8819) <= b and not a;
    layer4_outputs(8820) <= not b;
    layer4_outputs(8821) <= not a or b;
    layer4_outputs(8822) <= a or b;
    layer4_outputs(8823) <= a and not b;
    layer4_outputs(8824) <= not a;
    layer4_outputs(8825) <= b;
    layer4_outputs(8826) <= b;
    layer4_outputs(8827) <= 1'b1;
    layer4_outputs(8828) <= 1'b1;
    layer4_outputs(8829) <= a xor b;
    layer4_outputs(8830) <= a xor b;
    layer4_outputs(8831) <= not b or a;
    layer4_outputs(8832) <= not (a and b);
    layer4_outputs(8833) <= not (a and b);
    layer4_outputs(8834) <= a and b;
    layer4_outputs(8835) <= a and not b;
    layer4_outputs(8836) <= 1'b1;
    layer4_outputs(8837) <= not (a xor b);
    layer4_outputs(8838) <= b;
    layer4_outputs(8839) <= b;
    layer4_outputs(8840) <= not b or a;
    layer4_outputs(8841) <= not a or b;
    layer4_outputs(8842) <= 1'b1;
    layer4_outputs(8843) <= not a;
    layer4_outputs(8844) <= b and not a;
    layer4_outputs(8845) <= b and not a;
    layer4_outputs(8846) <= not a or b;
    layer4_outputs(8847) <= b and not a;
    layer4_outputs(8848) <= not (a or b);
    layer4_outputs(8849) <= not b;
    layer4_outputs(8850) <= not b;
    layer4_outputs(8851) <= not b or a;
    layer4_outputs(8852) <= not (a and b);
    layer4_outputs(8853) <= not b;
    layer4_outputs(8854) <= a and b;
    layer4_outputs(8855) <= a and not b;
    layer4_outputs(8856) <= 1'b0;
    layer4_outputs(8857) <= not (a and b);
    layer4_outputs(8858) <= a and b;
    layer4_outputs(8859) <= not (a or b);
    layer4_outputs(8860) <= a xor b;
    layer4_outputs(8861) <= not b or a;
    layer4_outputs(8862) <= a and b;
    layer4_outputs(8863) <= 1'b1;
    layer4_outputs(8864) <= a;
    layer4_outputs(8865) <= a xor b;
    layer4_outputs(8866) <= b and not a;
    layer4_outputs(8867) <= a and not b;
    layer4_outputs(8868) <= not b or a;
    layer4_outputs(8869) <= not a or b;
    layer4_outputs(8870) <= not a or b;
    layer4_outputs(8871) <= not a;
    layer4_outputs(8872) <= not (a and b);
    layer4_outputs(8873) <= not b or a;
    layer4_outputs(8874) <= not (a and b);
    layer4_outputs(8875) <= b and not a;
    layer4_outputs(8876) <= not a;
    layer4_outputs(8877) <= not a;
    layer4_outputs(8878) <= not a;
    layer4_outputs(8879) <= a and not b;
    layer4_outputs(8880) <= b;
    layer4_outputs(8881) <= 1'b1;
    layer4_outputs(8882) <= not b;
    layer4_outputs(8883) <= not (a or b);
    layer4_outputs(8884) <= not b or a;
    layer4_outputs(8885) <= not b or a;
    layer4_outputs(8886) <= a;
    layer4_outputs(8887) <= not (a and b);
    layer4_outputs(8888) <= 1'b1;
    layer4_outputs(8889) <= a xor b;
    layer4_outputs(8890) <= a and b;
    layer4_outputs(8891) <= not (a and b);
    layer4_outputs(8892) <= a;
    layer4_outputs(8893) <= not b;
    layer4_outputs(8894) <= a;
    layer4_outputs(8895) <= a;
    layer4_outputs(8896) <= a or b;
    layer4_outputs(8897) <= not (a or b);
    layer4_outputs(8898) <= not (a and b);
    layer4_outputs(8899) <= a or b;
    layer4_outputs(8900) <= a or b;
    layer4_outputs(8901) <= b;
    layer4_outputs(8902) <= b;
    layer4_outputs(8903) <= not (a or b);
    layer4_outputs(8904) <= not b;
    layer4_outputs(8905) <= a;
    layer4_outputs(8906) <= a;
    layer4_outputs(8907) <= b and not a;
    layer4_outputs(8908) <= b;
    layer4_outputs(8909) <= not (a xor b);
    layer4_outputs(8910) <= a and not b;
    layer4_outputs(8911) <= 1'b1;
    layer4_outputs(8912) <= 1'b0;
    layer4_outputs(8913) <= not a;
    layer4_outputs(8914) <= b;
    layer4_outputs(8915) <= not a or b;
    layer4_outputs(8916) <= 1'b0;
    layer4_outputs(8917) <= a and b;
    layer4_outputs(8918) <= a xor b;
    layer4_outputs(8919) <= not (a and b);
    layer4_outputs(8920) <= not b or a;
    layer4_outputs(8921) <= not a or b;
    layer4_outputs(8922) <= a and not b;
    layer4_outputs(8923) <= not b or a;
    layer4_outputs(8924) <= not a;
    layer4_outputs(8925) <= a xor b;
    layer4_outputs(8926) <= a and b;
    layer4_outputs(8927) <= a or b;
    layer4_outputs(8928) <= not (a or b);
    layer4_outputs(8929) <= a and not b;
    layer4_outputs(8930) <= a or b;
    layer4_outputs(8931) <= b;
    layer4_outputs(8932) <= b and not a;
    layer4_outputs(8933) <= not a;
    layer4_outputs(8934) <= b and not a;
    layer4_outputs(8935) <= not b;
    layer4_outputs(8936) <= a xor b;
    layer4_outputs(8937) <= not (a and b);
    layer4_outputs(8938) <= not (a xor b);
    layer4_outputs(8939) <= a;
    layer4_outputs(8940) <= a and b;
    layer4_outputs(8941) <= b;
    layer4_outputs(8942) <= not a or b;
    layer4_outputs(8943) <= b;
    layer4_outputs(8944) <= 1'b1;
    layer4_outputs(8945) <= b and not a;
    layer4_outputs(8946) <= a and not b;
    layer4_outputs(8947) <= a and not b;
    layer4_outputs(8948) <= not b;
    layer4_outputs(8949) <= 1'b1;
    layer4_outputs(8950) <= a or b;
    layer4_outputs(8951) <= a and b;
    layer4_outputs(8952) <= not b;
    layer4_outputs(8953) <= not a or b;
    layer4_outputs(8954) <= not a;
    layer4_outputs(8955) <= 1'b0;
    layer4_outputs(8956) <= not a or b;
    layer4_outputs(8957) <= not a;
    layer4_outputs(8958) <= not (a and b);
    layer4_outputs(8959) <= a xor b;
    layer4_outputs(8960) <= a and not b;
    layer4_outputs(8961) <= a and not b;
    layer4_outputs(8962) <= b;
    layer4_outputs(8963) <= a;
    layer4_outputs(8964) <= not b;
    layer4_outputs(8965) <= not a;
    layer4_outputs(8966) <= not (a and b);
    layer4_outputs(8967) <= a;
    layer4_outputs(8968) <= 1'b0;
    layer4_outputs(8969) <= not b;
    layer4_outputs(8970) <= a or b;
    layer4_outputs(8971) <= a and b;
    layer4_outputs(8972) <= not a;
    layer4_outputs(8973) <= not a or b;
    layer4_outputs(8974) <= a and not b;
    layer4_outputs(8975) <= not (a and b);
    layer4_outputs(8976) <= not (a and b);
    layer4_outputs(8977) <= b;
    layer4_outputs(8978) <= a and not b;
    layer4_outputs(8979) <= 1'b1;
    layer4_outputs(8980) <= b and not a;
    layer4_outputs(8981) <= a and not b;
    layer4_outputs(8982) <= b;
    layer4_outputs(8983) <= not (a and b);
    layer4_outputs(8984) <= a and b;
    layer4_outputs(8985) <= a or b;
    layer4_outputs(8986) <= a and b;
    layer4_outputs(8987) <= not (a and b);
    layer4_outputs(8988) <= not a;
    layer4_outputs(8989) <= b and not a;
    layer4_outputs(8990) <= a xor b;
    layer4_outputs(8991) <= not (a and b);
    layer4_outputs(8992) <= b;
    layer4_outputs(8993) <= b;
    layer4_outputs(8994) <= not (a xor b);
    layer4_outputs(8995) <= not (a or b);
    layer4_outputs(8996) <= not a or b;
    layer4_outputs(8997) <= not a;
    layer4_outputs(8998) <= b and not a;
    layer4_outputs(8999) <= 1'b1;
    layer4_outputs(9000) <= a;
    layer4_outputs(9001) <= a or b;
    layer4_outputs(9002) <= a and not b;
    layer4_outputs(9003) <= a and not b;
    layer4_outputs(9004) <= not (a and b);
    layer4_outputs(9005) <= not (a or b);
    layer4_outputs(9006) <= not a or b;
    layer4_outputs(9007) <= 1'b0;
    layer4_outputs(9008) <= a;
    layer4_outputs(9009) <= a;
    layer4_outputs(9010) <= not b;
    layer4_outputs(9011) <= not a;
    layer4_outputs(9012) <= not a;
    layer4_outputs(9013) <= a and not b;
    layer4_outputs(9014) <= not b or a;
    layer4_outputs(9015) <= not b or a;
    layer4_outputs(9016) <= 1'b1;
    layer4_outputs(9017) <= not b or a;
    layer4_outputs(9018) <= a;
    layer4_outputs(9019) <= not b or a;
    layer4_outputs(9020) <= 1'b0;
    layer4_outputs(9021) <= a or b;
    layer4_outputs(9022) <= not a or b;
    layer4_outputs(9023) <= 1'b0;
    layer4_outputs(9024) <= not (a and b);
    layer4_outputs(9025) <= not b;
    layer4_outputs(9026) <= 1'b1;
    layer4_outputs(9027) <= not a or b;
    layer4_outputs(9028) <= 1'b1;
    layer4_outputs(9029) <= 1'b0;
    layer4_outputs(9030) <= 1'b1;
    layer4_outputs(9031) <= not b or a;
    layer4_outputs(9032) <= not (a and b);
    layer4_outputs(9033) <= not a or b;
    layer4_outputs(9034) <= not (a xor b);
    layer4_outputs(9035) <= not a;
    layer4_outputs(9036) <= not a or b;
    layer4_outputs(9037) <= not b;
    layer4_outputs(9038) <= a;
    layer4_outputs(9039) <= not a;
    layer4_outputs(9040) <= a;
    layer4_outputs(9041) <= a;
    layer4_outputs(9042) <= not (a or b);
    layer4_outputs(9043) <= a xor b;
    layer4_outputs(9044) <= not a;
    layer4_outputs(9045) <= b;
    layer4_outputs(9046) <= b;
    layer4_outputs(9047) <= a and b;
    layer4_outputs(9048) <= not (a xor b);
    layer4_outputs(9049) <= 1'b1;
    layer4_outputs(9050) <= not a or b;
    layer4_outputs(9051) <= b;
    layer4_outputs(9052) <= b;
    layer4_outputs(9053) <= not b or a;
    layer4_outputs(9054) <= a;
    layer4_outputs(9055) <= b;
    layer4_outputs(9056) <= not (a and b);
    layer4_outputs(9057) <= b;
    layer4_outputs(9058) <= b;
    layer4_outputs(9059) <= a and b;
    layer4_outputs(9060) <= not a or b;
    layer4_outputs(9061) <= b and not a;
    layer4_outputs(9062) <= not (a or b);
    layer4_outputs(9063) <= not b or a;
    layer4_outputs(9064) <= b and not a;
    layer4_outputs(9065) <= b;
    layer4_outputs(9066) <= 1'b0;
    layer4_outputs(9067) <= a;
    layer4_outputs(9068) <= not b or a;
    layer4_outputs(9069) <= a or b;
    layer4_outputs(9070) <= a and not b;
    layer4_outputs(9071) <= a xor b;
    layer4_outputs(9072) <= a;
    layer4_outputs(9073) <= not (a or b);
    layer4_outputs(9074) <= a or b;
    layer4_outputs(9075) <= not (a or b);
    layer4_outputs(9076) <= b and not a;
    layer4_outputs(9077) <= a or b;
    layer4_outputs(9078) <= not (a xor b);
    layer4_outputs(9079) <= b;
    layer4_outputs(9080) <= not a or b;
    layer4_outputs(9081) <= b;
    layer4_outputs(9082) <= not b or a;
    layer4_outputs(9083) <= 1'b1;
    layer4_outputs(9084) <= a;
    layer4_outputs(9085) <= not b;
    layer4_outputs(9086) <= 1'b0;
    layer4_outputs(9087) <= b and not a;
    layer4_outputs(9088) <= a or b;
    layer4_outputs(9089) <= not (a xor b);
    layer4_outputs(9090) <= a and b;
    layer4_outputs(9091) <= a and not b;
    layer4_outputs(9092) <= b;
    layer4_outputs(9093) <= b and not a;
    layer4_outputs(9094) <= not a;
    layer4_outputs(9095) <= not a;
    layer4_outputs(9096) <= not (a or b);
    layer4_outputs(9097) <= a or b;
    layer4_outputs(9098) <= not b or a;
    layer4_outputs(9099) <= 1'b1;
    layer4_outputs(9100) <= a xor b;
    layer4_outputs(9101) <= not (a or b);
    layer4_outputs(9102) <= not (a xor b);
    layer4_outputs(9103) <= a;
    layer4_outputs(9104) <= not (a or b);
    layer4_outputs(9105) <= 1'b0;
    layer4_outputs(9106) <= a;
    layer4_outputs(9107) <= not a;
    layer4_outputs(9108) <= not b;
    layer4_outputs(9109) <= not a;
    layer4_outputs(9110) <= not b;
    layer4_outputs(9111) <= 1'b0;
    layer4_outputs(9112) <= not b or a;
    layer4_outputs(9113) <= a and not b;
    layer4_outputs(9114) <= not a or b;
    layer4_outputs(9115) <= not (a and b);
    layer4_outputs(9116) <= a or b;
    layer4_outputs(9117) <= 1'b0;
    layer4_outputs(9118) <= a and b;
    layer4_outputs(9119) <= not b;
    layer4_outputs(9120) <= not (a and b);
    layer4_outputs(9121) <= a or b;
    layer4_outputs(9122) <= b;
    layer4_outputs(9123) <= not a;
    layer4_outputs(9124) <= b;
    layer4_outputs(9125) <= not a or b;
    layer4_outputs(9126) <= not b or a;
    layer4_outputs(9127) <= not (a and b);
    layer4_outputs(9128) <= not a;
    layer4_outputs(9129) <= not (a or b);
    layer4_outputs(9130) <= a;
    layer4_outputs(9131) <= a;
    layer4_outputs(9132) <= a or b;
    layer4_outputs(9133) <= not b or a;
    layer4_outputs(9134) <= not b or a;
    layer4_outputs(9135) <= not a or b;
    layer4_outputs(9136) <= a and not b;
    layer4_outputs(9137) <= not b;
    layer4_outputs(9138) <= not (a or b);
    layer4_outputs(9139) <= not a or b;
    layer4_outputs(9140) <= not a;
    layer4_outputs(9141) <= 1'b1;
    layer4_outputs(9142) <= not a or b;
    layer4_outputs(9143) <= 1'b0;
    layer4_outputs(9144) <= not a;
    layer4_outputs(9145) <= a and not b;
    layer4_outputs(9146) <= a xor b;
    layer4_outputs(9147) <= b and not a;
    layer4_outputs(9148) <= b;
    layer4_outputs(9149) <= b;
    layer4_outputs(9150) <= a;
    layer4_outputs(9151) <= a xor b;
    layer4_outputs(9152) <= not a or b;
    layer4_outputs(9153) <= b;
    layer4_outputs(9154) <= not a or b;
    layer4_outputs(9155) <= b;
    layer4_outputs(9156) <= 1'b1;
    layer4_outputs(9157) <= 1'b0;
    layer4_outputs(9158) <= a and not b;
    layer4_outputs(9159) <= not a;
    layer4_outputs(9160) <= b;
    layer4_outputs(9161) <= a or b;
    layer4_outputs(9162) <= not a;
    layer4_outputs(9163) <= a and not b;
    layer4_outputs(9164) <= 1'b1;
    layer4_outputs(9165) <= not (a and b);
    layer4_outputs(9166) <= not (a and b);
    layer4_outputs(9167) <= not (a or b);
    layer4_outputs(9168) <= a or b;
    layer4_outputs(9169) <= b;
    layer4_outputs(9170) <= not b or a;
    layer4_outputs(9171) <= b and not a;
    layer4_outputs(9172) <= a xor b;
    layer4_outputs(9173) <= not b or a;
    layer4_outputs(9174) <= a or b;
    layer4_outputs(9175) <= 1'b0;
    layer4_outputs(9176) <= not b;
    layer4_outputs(9177) <= b;
    layer4_outputs(9178) <= a xor b;
    layer4_outputs(9179) <= b;
    layer4_outputs(9180) <= not a;
    layer4_outputs(9181) <= a and b;
    layer4_outputs(9182) <= not (a or b);
    layer4_outputs(9183) <= not (a and b);
    layer4_outputs(9184) <= not (a and b);
    layer4_outputs(9185) <= not b or a;
    layer4_outputs(9186) <= a and not b;
    layer4_outputs(9187) <= not a or b;
    layer4_outputs(9188) <= not (a xor b);
    layer4_outputs(9189) <= not (a or b);
    layer4_outputs(9190) <= not (a or b);
    layer4_outputs(9191) <= not a or b;
    layer4_outputs(9192) <= not a or b;
    layer4_outputs(9193) <= not a or b;
    layer4_outputs(9194) <= 1'b0;
    layer4_outputs(9195) <= 1'b1;
    layer4_outputs(9196) <= not (a and b);
    layer4_outputs(9197) <= a and b;
    layer4_outputs(9198) <= b;
    layer4_outputs(9199) <= not a or b;
    layer4_outputs(9200) <= a or b;
    layer4_outputs(9201) <= not a;
    layer4_outputs(9202) <= b;
    layer4_outputs(9203) <= not a or b;
    layer4_outputs(9204) <= not b or a;
    layer4_outputs(9205) <= not b;
    layer4_outputs(9206) <= a;
    layer4_outputs(9207) <= not (a or b);
    layer4_outputs(9208) <= b and not a;
    layer4_outputs(9209) <= not b or a;
    layer4_outputs(9210) <= b and not a;
    layer4_outputs(9211) <= a xor b;
    layer4_outputs(9212) <= a and b;
    layer4_outputs(9213) <= a or b;
    layer4_outputs(9214) <= a or b;
    layer4_outputs(9215) <= not b or a;
    layer4_outputs(9216) <= a xor b;
    layer4_outputs(9217) <= not b or a;
    layer4_outputs(9218) <= not a;
    layer4_outputs(9219) <= not b;
    layer4_outputs(9220) <= a or b;
    layer4_outputs(9221) <= a;
    layer4_outputs(9222) <= not b;
    layer4_outputs(9223) <= a or b;
    layer4_outputs(9224) <= a;
    layer4_outputs(9225) <= not a;
    layer4_outputs(9226) <= 1'b0;
    layer4_outputs(9227) <= not a or b;
    layer4_outputs(9228) <= b and not a;
    layer4_outputs(9229) <= a or b;
    layer4_outputs(9230) <= not b or a;
    layer4_outputs(9231) <= 1'b0;
    layer4_outputs(9232) <= not (a xor b);
    layer4_outputs(9233) <= not (a and b);
    layer4_outputs(9234) <= not (a and b);
    layer4_outputs(9235) <= a;
    layer4_outputs(9236) <= b;
    layer4_outputs(9237) <= not b;
    layer4_outputs(9238) <= a;
    layer4_outputs(9239) <= not (a or b);
    layer4_outputs(9240) <= not b or a;
    layer4_outputs(9241) <= a and b;
    layer4_outputs(9242) <= not a or b;
    layer4_outputs(9243) <= a or b;
    layer4_outputs(9244) <= not b;
    layer4_outputs(9245) <= a;
    layer4_outputs(9246) <= 1'b0;
    layer4_outputs(9247) <= b;
    layer4_outputs(9248) <= b;
    layer4_outputs(9249) <= not b;
    layer4_outputs(9250) <= 1'b1;
    layer4_outputs(9251) <= 1'b0;
    layer4_outputs(9252) <= not a or b;
    layer4_outputs(9253) <= not (a xor b);
    layer4_outputs(9254) <= not a;
    layer4_outputs(9255) <= not (a or b);
    layer4_outputs(9256) <= not (a or b);
    layer4_outputs(9257) <= not a or b;
    layer4_outputs(9258) <= not b;
    layer4_outputs(9259) <= b;
    layer4_outputs(9260) <= 1'b1;
    layer4_outputs(9261) <= not b;
    layer4_outputs(9262) <= a and not b;
    layer4_outputs(9263) <= b;
    layer4_outputs(9264) <= a;
    layer4_outputs(9265) <= not b;
    layer4_outputs(9266) <= not a;
    layer4_outputs(9267) <= a and b;
    layer4_outputs(9268) <= a;
    layer4_outputs(9269) <= not (a or b);
    layer4_outputs(9270) <= a xor b;
    layer4_outputs(9271) <= not a or b;
    layer4_outputs(9272) <= not b;
    layer4_outputs(9273) <= not (a and b);
    layer4_outputs(9274) <= a and b;
    layer4_outputs(9275) <= a and b;
    layer4_outputs(9276) <= not a;
    layer4_outputs(9277) <= a and not b;
    layer4_outputs(9278) <= not a;
    layer4_outputs(9279) <= a or b;
    layer4_outputs(9280) <= not (a and b);
    layer4_outputs(9281) <= a and not b;
    layer4_outputs(9282) <= a or b;
    layer4_outputs(9283) <= a and not b;
    layer4_outputs(9284) <= not a or b;
    layer4_outputs(9285) <= 1'b1;
    layer4_outputs(9286) <= not a or b;
    layer4_outputs(9287) <= a;
    layer4_outputs(9288) <= not b;
    layer4_outputs(9289) <= not a;
    layer4_outputs(9290) <= not b or a;
    layer4_outputs(9291) <= not b or a;
    layer4_outputs(9292) <= a or b;
    layer4_outputs(9293) <= b and not a;
    layer4_outputs(9294) <= b;
    layer4_outputs(9295) <= a or b;
    layer4_outputs(9296) <= b;
    layer4_outputs(9297) <= b;
    layer4_outputs(9298) <= 1'b1;
    layer4_outputs(9299) <= a or b;
    layer4_outputs(9300) <= b and not a;
    layer4_outputs(9301) <= a or b;
    layer4_outputs(9302) <= a;
    layer4_outputs(9303) <= a and b;
    layer4_outputs(9304) <= not a;
    layer4_outputs(9305) <= a and b;
    layer4_outputs(9306) <= a and not b;
    layer4_outputs(9307) <= not a;
    layer4_outputs(9308) <= not a or b;
    layer4_outputs(9309) <= not a;
    layer4_outputs(9310) <= a or b;
    layer4_outputs(9311) <= b;
    layer4_outputs(9312) <= not b;
    layer4_outputs(9313) <= a or b;
    layer4_outputs(9314) <= 1'b1;
    layer4_outputs(9315) <= not (a xor b);
    layer4_outputs(9316) <= not (a xor b);
    layer4_outputs(9317) <= not b;
    layer4_outputs(9318) <= b;
    layer4_outputs(9319) <= not (a and b);
    layer4_outputs(9320) <= not b or a;
    layer4_outputs(9321) <= not b;
    layer4_outputs(9322) <= not (a or b);
    layer4_outputs(9323) <= b;
    layer4_outputs(9324) <= a or b;
    layer4_outputs(9325) <= not (a and b);
    layer4_outputs(9326) <= not b or a;
    layer4_outputs(9327) <= not (a or b);
    layer4_outputs(9328) <= not b or a;
    layer4_outputs(9329) <= 1'b1;
    layer4_outputs(9330) <= not a;
    layer4_outputs(9331) <= not b or a;
    layer4_outputs(9332) <= not b or a;
    layer4_outputs(9333) <= a or b;
    layer4_outputs(9334) <= not (a or b);
    layer4_outputs(9335) <= a and not b;
    layer4_outputs(9336) <= a xor b;
    layer4_outputs(9337) <= not (a and b);
    layer4_outputs(9338) <= not (a and b);
    layer4_outputs(9339) <= not (a and b);
    layer4_outputs(9340) <= not (a and b);
    layer4_outputs(9341) <= not a;
    layer4_outputs(9342) <= not b or a;
    layer4_outputs(9343) <= b;
    layer4_outputs(9344) <= not (a and b);
    layer4_outputs(9345) <= a or b;
    layer4_outputs(9346) <= not a or b;
    layer4_outputs(9347) <= a xor b;
    layer4_outputs(9348) <= 1'b1;
    layer4_outputs(9349) <= a or b;
    layer4_outputs(9350) <= 1'b1;
    layer4_outputs(9351) <= a and not b;
    layer4_outputs(9352) <= a and b;
    layer4_outputs(9353) <= a xor b;
    layer4_outputs(9354) <= not (a and b);
    layer4_outputs(9355) <= 1'b1;
    layer4_outputs(9356) <= not a;
    layer4_outputs(9357) <= a and b;
    layer4_outputs(9358) <= not a;
    layer4_outputs(9359) <= not a;
    layer4_outputs(9360) <= a and b;
    layer4_outputs(9361) <= not (a and b);
    layer4_outputs(9362) <= not (a or b);
    layer4_outputs(9363) <= a;
    layer4_outputs(9364) <= a and not b;
    layer4_outputs(9365) <= b and not a;
    layer4_outputs(9366) <= not (a and b);
    layer4_outputs(9367) <= not (a or b);
    layer4_outputs(9368) <= a or b;
    layer4_outputs(9369) <= not a or b;
    layer4_outputs(9370) <= not (a or b);
    layer4_outputs(9371) <= 1'b0;
    layer4_outputs(9372) <= a and b;
    layer4_outputs(9373) <= a;
    layer4_outputs(9374) <= not a;
    layer4_outputs(9375) <= not (a or b);
    layer4_outputs(9376) <= a or b;
    layer4_outputs(9377) <= not (a and b);
    layer4_outputs(9378) <= b;
    layer4_outputs(9379) <= not b;
    layer4_outputs(9380) <= not a;
    layer4_outputs(9381) <= not (a or b);
    layer4_outputs(9382) <= a and b;
    layer4_outputs(9383) <= not b;
    layer4_outputs(9384) <= not b;
    layer4_outputs(9385) <= not a or b;
    layer4_outputs(9386) <= 1'b1;
    layer4_outputs(9387) <= a xor b;
    layer4_outputs(9388) <= a;
    layer4_outputs(9389) <= b;
    layer4_outputs(9390) <= a;
    layer4_outputs(9391) <= 1'b1;
    layer4_outputs(9392) <= not a;
    layer4_outputs(9393) <= not (a and b);
    layer4_outputs(9394) <= 1'b1;
    layer4_outputs(9395) <= 1'b1;
    layer4_outputs(9396) <= not b;
    layer4_outputs(9397) <= not (a or b);
    layer4_outputs(9398) <= not (a and b);
    layer4_outputs(9399) <= a and not b;
    layer4_outputs(9400) <= not (a or b);
    layer4_outputs(9401) <= a or b;
    layer4_outputs(9402) <= not (a or b);
    layer4_outputs(9403) <= b;
    layer4_outputs(9404) <= a;
    layer4_outputs(9405) <= not (a and b);
    layer4_outputs(9406) <= b;
    layer4_outputs(9407) <= b and not a;
    layer4_outputs(9408) <= not (a and b);
    layer4_outputs(9409) <= not a;
    layer4_outputs(9410) <= 1'b0;
    layer4_outputs(9411) <= a and b;
    layer4_outputs(9412) <= b;
    layer4_outputs(9413) <= a and b;
    layer4_outputs(9414) <= b;
    layer4_outputs(9415) <= a or b;
    layer4_outputs(9416) <= not a or b;
    layer4_outputs(9417) <= b and not a;
    layer4_outputs(9418) <= b and not a;
    layer4_outputs(9419) <= not b;
    layer4_outputs(9420) <= not (a and b);
    layer4_outputs(9421) <= not b;
    layer4_outputs(9422) <= a and not b;
    layer4_outputs(9423) <= 1'b1;
    layer4_outputs(9424) <= not (a xor b);
    layer4_outputs(9425) <= not a;
    layer4_outputs(9426) <= not b or a;
    layer4_outputs(9427) <= a and not b;
    layer4_outputs(9428) <= 1'b0;
    layer4_outputs(9429) <= not b or a;
    layer4_outputs(9430) <= not a or b;
    layer4_outputs(9431) <= a;
    layer4_outputs(9432) <= not (a and b);
    layer4_outputs(9433) <= 1'b1;
    layer4_outputs(9434) <= a;
    layer4_outputs(9435) <= not a;
    layer4_outputs(9436) <= not b or a;
    layer4_outputs(9437) <= a and not b;
    layer4_outputs(9438) <= not b;
    layer4_outputs(9439) <= 1'b0;
    layer4_outputs(9440) <= b;
    layer4_outputs(9441) <= not (a xor b);
    layer4_outputs(9442) <= b;
    layer4_outputs(9443) <= not a;
    layer4_outputs(9444) <= not b;
    layer4_outputs(9445) <= b and not a;
    layer4_outputs(9446) <= not (a or b);
    layer4_outputs(9447) <= b;
    layer4_outputs(9448) <= not a or b;
    layer4_outputs(9449) <= a and not b;
    layer4_outputs(9450) <= not b or a;
    layer4_outputs(9451) <= not (a or b);
    layer4_outputs(9452) <= not b or a;
    layer4_outputs(9453) <= a or b;
    layer4_outputs(9454) <= a;
    layer4_outputs(9455) <= 1'b0;
    layer4_outputs(9456) <= a xor b;
    layer4_outputs(9457) <= not (a xor b);
    layer4_outputs(9458) <= not (a and b);
    layer4_outputs(9459) <= not a;
    layer4_outputs(9460) <= 1'b0;
    layer4_outputs(9461) <= a or b;
    layer4_outputs(9462) <= a;
    layer4_outputs(9463) <= not b;
    layer4_outputs(9464) <= a and not b;
    layer4_outputs(9465) <= a and not b;
    layer4_outputs(9466) <= 1'b0;
    layer4_outputs(9467) <= a or b;
    layer4_outputs(9468) <= not (a or b);
    layer4_outputs(9469) <= a or b;
    layer4_outputs(9470) <= not a;
    layer4_outputs(9471) <= not (a and b);
    layer4_outputs(9472) <= b and not a;
    layer4_outputs(9473) <= b and not a;
    layer4_outputs(9474) <= a and not b;
    layer4_outputs(9475) <= not b or a;
    layer4_outputs(9476) <= not b or a;
    layer4_outputs(9477) <= not a or b;
    layer4_outputs(9478) <= b;
    layer4_outputs(9479) <= a;
    layer4_outputs(9480) <= not b;
    layer4_outputs(9481) <= 1'b1;
    layer4_outputs(9482) <= a xor b;
    layer4_outputs(9483) <= a and b;
    layer4_outputs(9484) <= not a or b;
    layer4_outputs(9485) <= not b;
    layer4_outputs(9486) <= 1'b0;
    layer4_outputs(9487) <= not (a xor b);
    layer4_outputs(9488) <= b and not a;
    layer4_outputs(9489) <= a;
    layer4_outputs(9490) <= not (a and b);
    layer4_outputs(9491) <= 1'b1;
    layer4_outputs(9492) <= not (a and b);
    layer4_outputs(9493) <= not (a and b);
    layer4_outputs(9494) <= not b or a;
    layer4_outputs(9495) <= not b;
    layer4_outputs(9496) <= 1'b1;
    layer4_outputs(9497) <= not b;
    layer4_outputs(9498) <= not b or a;
    layer4_outputs(9499) <= not b;
    layer4_outputs(9500) <= not b;
    layer4_outputs(9501) <= 1'b1;
    layer4_outputs(9502) <= b;
    layer4_outputs(9503) <= a and not b;
    layer4_outputs(9504) <= a and b;
    layer4_outputs(9505) <= b;
    layer4_outputs(9506) <= not (a or b);
    layer4_outputs(9507) <= not b;
    layer4_outputs(9508) <= not b;
    layer4_outputs(9509) <= not a;
    layer4_outputs(9510) <= 1'b0;
    layer4_outputs(9511) <= not (a and b);
    layer4_outputs(9512) <= not a;
    layer4_outputs(9513) <= 1'b1;
    layer4_outputs(9514) <= not a;
    layer4_outputs(9515) <= a and b;
    layer4_outputs(9516) <= b;
    layer4_outputs(9517) <= 1'b1;
    layer4_outputs(9518) <= a;
    layer4_outputs(9519) <= not (a and b);
    layer4_outputs(9520) <= not (a and b);
    layer4_outputs(9521) <= a or b;
    layer4_outputs(9522) <= a and b;
    layer4_outputs(9523) <= a;
    layer4_outputs(9524) <= a or b;
    layer4_outputs(9525) <= a or b;
    layer4_outputs(9526) <= a and b;
    layer4_outputs(9527) <= not (a or b);
    layer4_outputs(9528) <= a;
    layer4_outputs(9529) <= a;
    layer4_outputs(9530) <= not a or b;
    layer4_outputs(9531) <= 1'b0;
    layer4_outputs(9532) <= 1'b1;
    layer4_outputs(9533) <= not a;
    layer4_outputs(9534) <= not b or a;
    layer4_outputs(9535) <= not b or a;
    layer4_outputs(9536) <= not b;
    layer4_outputs(9537) <= a and not b;
    layer4_outputs(9538) <= a and b;
    layer4_outputs(9539) <= not a;
    layer4_outputs(9540) <= not (a xor b);
    layer4_outputs(9541) <= a and b;
    layer4_outputs(9542) <= a;
    layer4_outputs(9543) <= a;
    layer4_outputs(9544) <= a xor b;
    layer4_outputs(9545) <= a and b;
    layer4_outputs(9546) <= 1'b0;
    layer4_outputs(9547) <= b;
    layer4_outputs(9548) <= 1'b1;
    layer4_outputs(9549) <= not (a or b);
    layer4_outputs(9550) <= not b or a;
    layer4_outputs(9551) <= not a;
    layer4_outputs(9552) <= a;
    layer4_outputs(9553) <= not b or a;
    layer4_outputs(9554) <= not b;
    layer4_outputs(9555) <= b;
    layer4_outputs(9556) <= a and b;
    layer4_outputs(9557) <= a or b;
    layer4_outputs(9558) <= a or b;
    layer4_outputs(9559) <= 1'b0;
    layer4_outputs(9560) <= b;
    layer4_outputs(9561) <= a xor b;
    layer4_outputs(9562) <= not a or b;
    layer4_outputs(9563) <= 1'b0;
    layer4_outputs(9564) <= 1'b1;
    layer4_outputs(9565) <= 1'b0;
    layer4_outputs(9566) <= not (a and b);
    layer4_outputs(9567) <= a and not b;
    layer4_outputs(9568) <= b;
    layer4_outputs(9569) <= not a or b;
    layer4_outputs(9570) <= not a or b;
    layer4_outputs(9571) <= not (a or b);
    layer4_outputs(9572) <= a;
    layer4_outputs(9573) <= not b;
    layer4_outputs(9574) <= 1'b1;
    layer4_outputs(9575) <= not a;
    layer4_outputs(9576) <= 1'b1;
    layer4_outputs(9577) <= not a;
    layer4_outputs(9578) <= b;
    layer4_outputs(9579) <= 1'b1;
    layer4_outputs(9580) <= not a;
    layer4_outputs(9581) <= a and b;
    layer4_outputs(9582) <= not (a or b);
    layer4_outputs(9583) <= not a;
    layer4_outputs(9584) <= not a;
    layer4_outputs(9585) <= b and not a;
    layer4_outputs(9586) <= b and not a;
    layer4_outputs(9587) <= a;
    layer4_outputs(9588) <= not (a and b);
    layer4_outputs(9589) <= not b;
    layer4_outputs(9590) <= b and not a;
    layer4_outputs(9591) <= b and not a;
    layer4_outputs(9592) <= b and not a;
    layer4_outputs(9593) <= not (a xor b);
    layer4_outputs(9594) <= not a;
    layer4_outputs(9595) <= not a or b;
    layer4_outputs(9596) <= a xor b;
    layer4_outputs(9597) <= a and not b;
    layer4_outputs(9598) <= not a or b;
    layer4_outputs(9599) <= a;
    layer4_outputs(9600) <= a;
    layer4_outputs(9601) <= a or b;
    layer4_outputs(9602) <= a and not b;
    layer4_outputs(9603) <= b;
    layer4_outputs(9604) <= not b or a;
    layer4_outputs(9605) <= not a or b;
    layer4_outputs(9606) <= 1'b0;
    layer4_outputs(9607) <= not b or a;
    layer4_outputs(9608) <= a and b;
    layer4_outputs(9609) <= not a or b;
    layer4_outputs(9610) <= not (a and b);
    layer4_outputs(9611) <= a;
    layer4_outputs(9612) <= a;
    layer4_outputs(9613) <= b;
    layer4_outputs(9614) <= not a or b;
    layer4_outputs(9615) <= a;
    layer4_outputs(9616) <= a or b;
    layer4_outputs(9617) <= not b or a;
    layer4_outputs(9618) <= not a;
    layer4_outputs(9619) <= a and not b;
    layer4_outputs(9620) <= a and b;
    layer4_outputs(9621) <= a;
    layer4_outputs(9622) <= b;
    layer4_outputs(9623) <= not (a xor b);
    layer4_outputs(9624) <= not (a xor b);
    layer4_outputs(9625) <= a xor b;
    layer4_outputs(9626) <= a or b;
    layer4_outputs(9627) <= not (a and b);
    layer4_outputs(9628) <= not b;
    layer4_outputs(9629) <= a;
    layer4_outputs(9630) <= not b or a;
    layer4_outputs(9631) <= a xor b;
    layer4_outputs(9632) <= not b or a;
    layer4_outputs(9633) <= not a;
    layer4_outputs(9634) <= not a;
    layer4_outputs(9635) <= not (a and b);
    layer4_outputs(9636) <= not b;
    layer4_outputs(9637) <= not (a xor b);
    layer4_outputs(9638) <= not (a or b);
    layer4_outputs(9639) <= not b or a;
    layer4_outputs(9640) <= 1'b1;
    layer4_outputs(9641) <= not a;
    layer4_outputs(9642) <= a or b;
    layer4_outputs(9643) <= not (a and b);
    layer4_outputs(9644) <= b and not a;
    layer4_outputs(9645) <= not b;
    layer4_outputs(9646) <= a or b;
    layer4_outputs(9647) <= a or b;
    layer4_outputs(9648) <= a or b;
    layer4_outputs(9649) <= not b;
    layer4_outputs(9650) <= 1'b0;
    layer4_outputs(9651) <= a;
    layer4_outputs(9652) <= a;
    layer4_outputs(9653) <= a;
    layer4_outputs(9654) <= not (a and b);
    layer4_outputs(9655) <= b;
    layer4_outputs(9656) <= not (a or b);
    layer4_outputs(9657) <= 1'b0;
    layer4_outputs(9658) <= b and not a;
    layer4_outputs(9659) <= 1'b0;
    layer4_outputs(9660) <= 1'b0;
    layer4_outputs(9661) <= a and not b;
    layer4_outputs(9662) <= not a or b;
    layer4_outputs(9663) <= not b;
    layer4_outputs(9664) <= not a;
    layer4_outputs(9665) <= a and not b;
    layer4_outputs(9666) <= not a or b;
    layer4_outputs(9667) <= a or b;
    layer4_outputs(9668) <= not b or a;
    layer4_outputs(9669) <= b;
    layer4_outputs(9670) <= a xor b;
    layer4_outputs(9671) <= 1'b1;
    layer4_outputs(9672) <= not (a and b);
    layer4_outputs(9673) <= not (a xor b);
    layer4_outputs(9674) <= not b;
    layer4_outputs(9675) <= a and b;
    layer4_outputs(9676) <= a;
    layer4_outputs(9677) <= a and not b;
    layer4_outputs(9678) <= 1'b0;
    layer4_outputs(9679) <= not a or b;
    layer4_outputs(9680) <= b;
    layer4_outputs(9681) <= a;
    layer4_outputs(9682) <= a and b;
    layer4_outputs(9683) <= a;
    layer4_outputs(9684) <= a and b;
    layer4_outputs(9685) <= 1'b1;
    layer4_outputs(9686) <= not b or a;
    layer4_outputs(9687) <= not (a and b);
    layer4_outputs(9688) <= a and not b;
    layer4_outputs(9689) <= not a;
    layer4_outputs(9690) <= not (a and b);
    layer4_outputs(9691) <= not b;
    layer4_outputs(9692) <= not b or a;
    layer4_outputs(9693) <= not (a and b);
    layer4_outputs(9694) <= a;
    layer4_outputs(9695) <= 1'b0;
    layer4_outputs(9696) <= a and not b;
    layer4_outputs(9697) <= b;
    layer4_outputs(9698) <= a;
    layer4_outputs(9699) <= not b or a;
    layer4_outputs(9700) <= a or b;
    layer4_outputs(9701) <= a and not b;
    layer4_outputs(9702) <= not (a or b);
    layer4_outputs(9703) <= 1'b1;
    layer4_outputs(9704) <= not a;
    layer4_outputs(9705) <= 1'b1;
    layer4_outputs(9706) <= a;
    layer4_outputs(9707) <= b;
    layer4_outputs(9708) <= not a;
    layer4_outputs(9709) <= not (a or b);
    layer4_outputs(9710) <= 1'b1;
    layer4_outputs(9711) <= a and b;
    layer4_outputs(9712) <= a and not b;
    layer4_outputs(9713) <= b;
    layer4_outputs(9714) <= not b;
    layer4_outputs(9715) <= a;
    layer4_outputs(9716) <= not b;
    layer4_outputs(9717) <= not a;
    layer4_outputs(9718) <= a;
    layer4_outputs(9719) <= b and not a;
    layer4_outputs(9720) <= a;
    layer4_outputs(9721) <= a or b;
    layer4_outputs(9722) <= not (a or b);
    layer4_outputs(9723) <= not (a and b);
    layer4_outputs(9724) <= not b;
    layer4_outputs(9725) <= a and b;
    layer4_outputs(9726) <= 1'b1;
    layer4_outputs(9727) <= 1'b0;
    layer4_outputs(9728) <= not a or b;
    layer4_outputs(9729) <= a and not b;
    layer4_outputs(9730) <= not b;
    layer4_outputs(9731) <= a;
    layer4_outputs(9732) <= not a;
    layer4_outputs(9733) <= not b or a;
    layer4_outputs(9734) <= b;
    layer4_outputs(9735) <= a and not b;
    layer4_outputs(9736) <= not (a or b);
    layer4_outputs(9737) <= not (a and b);
    layer4_outputs(9738) <= not a;
    layer4_outputs(9739) <= not a or b;
    layer4_outputs(9740) <= a or b;
    layer4_outputs(9741) <= not (a or b);
    layer4_outputs(9742) <= not a;
    layer4_outputs(9743) <= not (a or b);
    layer4_outputs(9744) <= not (a and b);
    layer4_outputs(9745) <= a or b;
    layer4_outputs(9746) <= not (a or b);
    layer4_outputs(9747) <= not b or a;
    layer4_outputs(9748) <= a and b;
    layer4_outputs(9749) <= not (a and b);
    layer4_outputs(9750) <= a and not b;
    layer4_outputs(9751) <= not (a and b);
    layer4_outputs(9752) <= b;
    layer4_outputs(9753) <= not (a and b);
    layer4_outputs(9754) <= a and not b;
    layer4_outputs(9755) <= not a;
    layer4_outputs(9756) <= b;
    layer4_outputs(9757) <= b and not a;
    layer4_outputs(9758) <= 1'b1;
    layer4_outputs(9759) <= b and not a;
    layer4_outputs(9760) <= 1'b0;
    layer4_outputs(9761) <= not b;
    layer4_outputs(9762) <= not a;
    layer4_outputs(9763) <= not (a xor b);
    layer4_outputs(9764) <= not a or b;
    layer4_outputs(9765) <= a and not b;
    layer4_outputs(9766) <= a;
    layer4_outputs(9767) <= b and not a;
    layer4_outputs(9768) <= a and not b;
    layer4_outputs(9769) <= not a;
    layer4_outputs(9770) <= a;
    layer4_outputs(9771) <= a;
    layer4_outputs(9772) <= a;
    layer4_outputs(9773) <= not a;
    layer4_outputs(9774) <= 1'b0;
    layer4_outputs(9775) <= a and b;
    layer4_outputs(9776) <= a and not b;
    layer4_outputs(9777) <= b and not a;
    layer4_outputs(9778) <= a and not b;
    layer4_outputs(9779) <= not b or a;
    layer4_outputs(9780) <= not a;
    layer4_outputs(9781) <= not a or b;
    layer4_outputs(9782) <= b and not a;
    layer4_outputs(9783) <= not b;
    layer4_outputs(9784) <= not (a xor b);
    layer4_outputs(9785) <= not a or b;
    layer4_outputs(9786) <= not a or b;
    layer4_outputs(9787) <= not (a or b);
    layer4_outputs(9788) <= not a or b;
    layer4_outputs(9789) <= not b;
    layer4_outputs(9790) <= a;
    layer4_outputs(9791) <= b and not a;
    layer4_outputs(9792) <= a;
    layer4_outputs(9793) <= 1'b1;
    layer4_outputs(9794) <= a and not b;
    layer4_outputs(9795) <= not a or b;
    layer4_outputs(9796) <= a and not b;
    layer4_outputs(9797) <= b;
    layer4_outputs(9798) <= not b or a;
    layer4_outputs(9799) <= not b or a;
    layer4_outputs(9800) <= not a;
    layer4_outputs(9801) <= not a or b;
    layer4_outputs(9802) <= a xor b;
    layer4_outputs(9803) <= not a;
    layer4_outputs(9804) <= not a or b;
    layer4_outputs(9805) <= a or b;
    layer4_outputs(9806) <= not b;
    layer4_outputs(9807) <= not a;
    layer4_outputs(9808) <= 1'b1;
    layer4_outputs(9809) <= not a;
    layer4_outputs(9810) <= a and not b;
    layer4_outputs(9811) <= 1'b1;
    layer4_outputs(9812) <= b and not a;
    layer4_outputs(9813) <= a and not b;
    layer4_outputs(9814) <= not b;
    layer4_outputs(9815) <= a;
    layer4_outputs(9816) <= not b;
    layer4_outputs(9817) <= 1'b0;
    layer4_outputs(9818) <= not (a or b);
    layer4_outputs(9819) <= not a or b;
    layer4_outputs(9820) <= 1'b1;
    layer4_outputs(9821) <= a or b;
    layer4_outputs(9822) <= not a;
    layer4_outputs(9823) <= a or b;
    layer4_outputs(9824) <= a and not b;
    layer4_outputs(9825) <= a;
    layer4_outputs(9826) <= b and not a;
    layer4_outputs(9827) <= not a;
    layer4_outputs(9828) <= b and not a;
    layer4_outputs(9829) <= not b;
    layer4_outputs(9830) <= 1'b0;
    layer4_outputs(9831) <= a;
    layer4_outputs(9832) <= not b;
    layer4_outputs(9833) <= not a;
    layer4_outputs(9834) <= b and not a;
    layer4_outputs(9835) <= b and not a;
    layer4_outputs(9836) <= not b or a;
    layer4_outputs(9837) <= a or b;
    layer4_outputs(9838) <= not b;
    layer4_outputs(9839) <= not (a and b);
    layer4_outputs(9840) <= a or b;
    layer4_outputs(9841) <= not b or a;
    layer4_outputs(9842) <= a;
    layer4_outputs(9843) <= not a;
    layer4_outputs(9844) <= not (a xor b);
    layer4_outputs(9845) <= not b;
    layer4_outputs(9846) <= not (a or b);
    layer4_outputs(9847) <= a and b;
    layer4_outputs(9848) <= a;
    layer4_outputs(9849) <= a xor b;
    layer4_outputs(9850) <= b and not a;
    layer4_outputs(9851) <= a and not b;
    layer4_outputs(9852) <= not b or a;
    layer4_outputs(9853) <= b;
    layer4_outputs(9854) <= not b or a;
    layer4_outputs(9855) <= a and not b;
    layer4_outputs(9856) <= a xor b;
    layer4_outputs(9857) <= not b or a;
    layer4_outputs(9858) <= b and not a;
    layer4_outputs(9859) <= not a;
    layer4_outputs(9860) <= 1'b0;
    layer4_outputs(9861) <= b;
    layer4_outputs(9862) <= 1'b1;
    layer4_outputs(9863) <= 1'b1;
    layer4_outputs(9864) <= not (a or b);
    layer4_outputs(9865) <= a xor b;
    layer4_outputs(9866) <= a;
    layer4_outputs(9867) <= not (a or b);
    layer4_outputs(9868) <= b;
    layer4_outputs(9869) <= a or b;
    layer4_outputs(9870) <= not b or a;
    layer4_outputs(9871) <= not (a or b);
    layer4_outputs(9872) <= a;
    layer4_outputs(9873) <= a and b;
    layer4_outputs(9874) <= 1'b0;
    layer4_outputs(9875) <= b and not a;
    layer4_outputs(9876) <= a and b;
    layer4_outputs(9877) <= not b or a;
    layer4_outputs(9878) <= not b;
    layer4_outputs(9879) <= a and not b;
    layer4_outputs(9880) <= a and b;
    layer4_outputs(9881) <= a and not b;
    layer4_outputs(9882) <= a and b;
    layer4_outputs(9883) <= not a or b;
    layer4_outputs(9884) <= b;
    layer4_outputs(9885) <= a and b;
    layer4_outputs(9886) <= not (a xor b);
    layer4_outputs(9887) <= a;
    layer4_outputs(9888) <= b;
    layer4_outputs(9889) <= 1'b1;
    layer4_outputs(9890) <= not b;
    layer4_outputs(9891) <= 1'b1;
    layer4_outputs(9892) <= not b;
    layer4_outputs(9893) <= b;
    layer4_outputs(9894) <= a and b;
    layer4_outputs(9895) <= not (a or b);
    layer4_outputs(9896) <= a;
    layer4_outputs(9897) <= a xor b;
    layer4_outputs(9898) <= a and not b;
    layer4_outputs(9899) <= not b;
    layer4_outputs(9900) <= not b or a;
    layer4_outputs(9901) <= 1'b1;
    layer4_outputs(9902) <= a;
    layer4_outputs(9903) <= b and not a;
    layer4_outputs(9904) <= a;
    layer4_outputs(9905) <= not a or b;
    layer4_outputs(9906) <= a and not b;
    layer4_outputs(9907) <= not a;
    layer4_outputs(9908) <= b and not a;
    layer4_outputs(9909) <= b;
    layer4_outputs(9910) <= 1'b0;
    layer4_outputs(9911) <= a and b;
    layer4_outputs(9912) <= not a;
    layer4_outputs(9913) <= not b or a;
    layer4_outputs(9914) <= not (a or b);
    layer4_outputs(9915) <= not b;
    layer4_outputs(9916) <= not (a and b);
    layer4_outputs(9917) <= 1'b0;
    layer4_outputs(9918) <= 1'b0;
    layer4_outputs(9919) <= 1'b0;
    layer4_outputs(9920) <= not (a xor b);
    layer4_outputs(9921) <= not (a or b);
    layer4_outputs(9922) <= not b;
    layer4_outputs(9923) <= 1'b1;
    layer4_outputs(9924) <= not b;
    layer4_outputs(9925) <= a;
    layer4_outputs(9926) <= not (a or b);
    layer4_outputs(9927) <= 1'b1;
    layer4_outputs(9928) <= not a;
    layer4_outputs(9929) <= a and b;
    layer4_outputs(9930) <= not b;
    layer4_outputs(9931) <= not b;
    layer4_outputs(9932) <= a or b;
    layer4_outputs(9933) <= a and not b;
    layer4_outputs(9934) <= not (a and b);
    layer4_outputs(9935) <= not a or b;
    layer4_outputs(9936) <= a and b;
    layer4_outputs(9937) <= a;
    layer4_outputs(9938) <= b;
    layer4_outputs(9939) <= not (a or b);
    layer4_outputs(9940) <= b and not a;
    layer4_outputs(9941) <= b and not a;
    layer4_outputs(9942) <= b and not a;
    layer4_outputs(9943) <= a and b;
    layer4_outputs(9944) <= not (a and b);
    layer4_outputs(9945) <= b and not a;
    layer4_outputs(9946) <= not b;
    layer4_outputs(9947) <= a and not b;
    layer4_outputs(9948) <= 1'b1;
    layer4_outputs(9949) <= a or b;
    layer4_outputs(9950) <= b and not a;
    layer4_outputs(9951) <= a or b;
    layer4_outputs(9952) <= not b or a;
    layer4_outputs(9953) <= b;
    layer4_outputs(9954) <= a or b;
    layer4_outputs(9955) <= a or b;
    layer4_outputs(9956) <= not b or a;
    layer4_outputs(9957) <= a and b;
    layer4_outputs(9958) <= not a or b;
    layer4_outputs(9959) <= a and not b;
    layer4_outputs(9960) <= a;
    layer4_outputs(9961) <= not (a and b);
    layer4_outputs(9962) <= a xor b;
    layer4_outputs(9963) <= not (a and b);
    layer4_outputs(9964) <= not a or b;
    layer4_outputs(9965) <= b;
    layer4_outputs(9966) <= not b;
    layer4_outputs(9967) <= not b;
    layer4_outputs(9968) <= not b;
    layer4_outputs(9969) <= a and b;
    layer4_outputs(9970) <= not (a xor b);
    layer4_outputs(9971) <= not b;
    layer4_outputs(9972) <= b and not a;
    layer4_outputs(9973) <= 1'b1;
    layer4_outputs(9974) <= not a or b;
    layer4_outputs(9975) <= not (a xor b);
    layer4_outputs(9976) <= b;
    layer4_outputs(9977) <= not (a xor b);
    layer4_outputs(9978) <= not (a or b);
    layer4_outputs(9979) <= not a or b;
    layer4_outputs(9980) <= not b or a;
    layer4_outputs(9981) <= b;
    layer4_outputs(9982) <= 1'b0;
    layer4_outputs(9983) <= 1'b1;
    layer4_outputs(9984) <= not b;
    layer4_outputs(9985) <= a and b;
    layer4_outputs(9986) <= a;
    layer4_outputs(9987) <= not a;
    layer4_outputs(9988) <= a and b;
    layer4_outputs(9989) <= a or b;
    layer4_outputs(9990) <= not b;
    layer4_outputs(9991) <= not (a or b);
    layer4_outputs(9992) <= 1'b0;
    layer4_outputs(9993) <= not b or a;
    layer4_outputs(9994) <= not b;
    layer4_outputs(9995) <= b and not a;
    layer4_outputs(9996) <= 1'b1;
    layer4_outputs(9997) <= b;
    layer4_outputs(9998) <= 1'b0;
    layer4_outputs(9999) <= a and b;
    layer4_outputs(10000) <= 1'b0;
    layer4_outputs(10001) <= a and not b;
    layer4_outputs(10002) <= a;
    layer4_outputs(10003) <= b;
    layer4_outputs(10004) <= a or b;
    layer4_outputs(10005) <= b;
    layer4_outputs(10006) <= not b or a;
    layer4_outputs(10007) <= a and not b;
    layer4_outputs(10008) <= 1'b1;
    layer4_outputs(10009) <= b;
    layer4_outputs(10010) <= a;
    layer4_outputs(10011) <= a and not b;
    layer4_outputs(10012) <= b and not a;
    layer4_outputs(10013) <= b;
    layer4_outputs(10014) <= not a or b;
    layer4_outputs(10015) <= not (a or b);
    layer4_outputs(10016) <= b;
    layer4_outputs(10017) <= not b or a;
    layer4_outputs(10018) <= 1'b1;
    layer4_outputs(10019) <= not a;
    layer4_outputs(10020) <= not a or b;
    layer4_outputs(10021) <= a and b;
    layer4_outputs(10022) <= not a or b;
    layer4_outputs(10023) <= not a;
    layer4_outputs(10024) <= 1'b0;
    layer4_outputs(10025) <= not (a and b);
    layer4_outputs(10026) <= not b;
    layer4_outputs(10027) <= 1'b1;
    layer4_outputs(10028) <= a and b;
    layer4_outputs(10029) <= not a;
    layer4_outputs(10030) <= not a or b;
    layer4_outputs(10031) <= a xor b;
    layer4_outputs(10032) <= not b;
    layer4_outputs(10033) <= a and b;
    layer4_outputs(10034) <= not (a or b);
    layer4_outputs(10035) <= not (a or b);
    layer4_outputs(10036) <= not (a xor b);
    layer4_outputs(10037) <= a;
    layer4_outputs(10038) <= b;
    layer4_outputs(10039) <= not b;
    layer4_outputs(10040) <= 1'b0;
    layer4_outputs(10041) <= a and not b;
    layer4_outputs(10042) <= a;
    layer4_outputs(10043) <= not b;
    layer4_outputs(10044) <= a and b;
    layer4_outputs(10045) <= not a;
    layer4_outputs(10046) <= b and not a;
    layer4_outputs(10047) <= not (a and b);
    layer4_outputs(10048) <= not a or b;
    layer4_outputs(10049) <= not b or a;
    layer4_outputs(10050) <= not a;
    layer4_outputs(10051) <= not a or b;
    layer4_outputs(10052) <= b;
    layer4_outputs(10053) <= a and not b;
    layer4_outputs(10054) <= not a;
    layer4_outputs(10055) <= not b or a;
    layer4_outputs(10056) <= 1'b1;
    layer4_outputs(10057) <= b;
    layer4_outputs(10058) <= a xor b;
    layer4_outputs(10059) <= a and not b;
    layer4_outputs(10060) <= not b or a;
    layer4_outputs(10061) <= 1'b1;
    layer4_outputs(10062) <= not b or a;
    layer4_outputs(10063) <= not a;
    layer4_outputs(10064) <= a xor b;
    layer4_outputs(10065) <= a and not b;
    layer4_outputs(10066) <= a and not b;
    layer4_outputs(10067) <= not a;
    layer4_outputs(10068) <= not a;
    layer4_outputs(10069) <= a or b;
    layer4_outputs(10070) <= not b or a;
    layer4_outputs(10071) <= not a;
    layer4_outputs(10072) <= not (a xor b);
    layer4_outputs(10073) <= 1'b1;
    layer4_outputs(10074) <= a or b;
    layer4_outputs(10075) <= not (a xor b);
    layer4_outputs(10076) <= not (a or b);
    layer4_outputs(10077) <= a xor b;
    layer4_outputs(10078) <= not b;
    layer4_outputs(10079) <= not a;
    layer4_outputs(10080) <= b and not a;
    layer4_outputs(10081) <= 1'b1;
    layer4_outputs(10082) <= not b or a;
    layer4_outputs(10083) <= 1'b1;
    layer4_outputs(10084) <= not a;
    layer4_outputs(10085) <= a or b;
    layer4_outputs(10086) <= not (a xor b);
    layer4_outputs(10087) <= b and not a;
    layer4_outputs(10088) <= b and not a;
    layer4_outputs(10089) <= 1'b0;
    layer4_outputs(10090) <= not a;
    layer4_outputs(10091) <= a;
    layer4_outputs(10092) <= a and not b;
    layer4_outputs(10093) <= not a;
    layer4_outputs(10094) <= not a;
    layer4_outputs(10095) <= a xor b;
    layer4_outputs(10096) <= not b;
    layer4_outputs(10097) <= not a;
    layer4_outputs(10098) <= not b or a;
    layer4_outputs(10099) <= not a or b;
    layer4_outputs(10100) <= 1'b0;
    layer4_outputs(10101) <= not a;
    layer4_outputs(10102) <= b;
    layer4_outputs(10103) <= not (a or b);
    layer4_outputs(10104) <= a and not b;
    layer4_outputs(10105) <= not (a and b);
    layer4_outputs(10106) <= not b;
    layer4_outputs(10107) <= a and b;
    layer4_outputs(10108) <= a xor b;
    layer4_outputs(10109) <= not (a and b);
    layer4_outputs(10110) <= 1'b1;
    layer4_outputs(10111) <= 1'b0;
    layer4_outputs(10112) <= not a;
    layer4_outputs(10113) <= b;
    layer4_outputs(10114) <= a and not b;
    layer4_outputs(10115) <= not b;
    layer4_outputs(10116) <= not (a and b);
    layer4_outputs(10117) <= a and not b;
    layer4_outputs(10118) <= b;
    layer4_outputs(10119) <= not b or a;
    layer4_outputs(10120) <= not a;
    layer4_outputs(10121) <= a and b;
    layer4_outputs(10122) <= not b or a;
    layer4_outputs(10123) <= not b;
    layer4_outputs(10124) <= b and not a;
    layer4_outputs(10125) <= not a;
    layer4_outputs(10126) <= 1'b0;
    layer4_outputs(10127) <= 1'b1;
    layer4_outputs(10128) <= b and not a;
    layer4_outputs(10129) <= 1'b1;
    layer4_outputs(10130) <= not (a or b);
    layer4_outputs(10131) <= a and b;
    layer4_outputs(10132) <= not a or b;
    layer4_outputs(10133) <= a or b;
    layer4_outputs(10134) <= not (a or b);
    layer4_outputs(10135) <= b and not a;
    layer4_outputs(10136) <= a xor b;
    layer4_outputs(10137) <= not b;
    layer4_outputs(10138) <= not b;
    layer4_outputs(10139) <= not (a or b);
    layer4_outputs(10140) <= a;
    layer4_outputs(10141) <= not a or b;
    layer4_outputs(10142) <= not b or a;
    layer4_outputs(10143) <= a or b;
    layer4_outputs(10144) <= b;
    layer4_outputs(10145) <= not a;
    layer4_outputs(10146) <= 1'b0;
    layer4_outputs(10147) <= not b;
    layer4_outputs(10148) <= not b or a;
    layer4_outputs(10149) <= a;
    layer4_outputs(10150) <= not b;
    layer4_outputs(10151) <= a and not b;
    layer4_outputs(10152) <= not a;
    layer4_outputs(10153) <= a and not b;
    layer4_outputs(10154) <= not a;
    layer4_outputs(10155) <= not b;
    layer4_outputs(10156) <= 1'b1;
    layer4_outputs(10157) <= a or b;
    layer4_outputs(10158) <= a and b;
    layer4_outputs(10159) <= 1'b1;
    layer4_outputs(10160) <= b;
    layer4_outputs(10161) <= 1'b1;
    layer4_outputs(10162) <= not b;
    layer4_outputs(10163) <= not (a or b);
    layer4_outputs(10164) <= b;
    layer4_outputs(10165) <= b and not a;
    layer4_outputs(10166) <= not (a xor b);
    layer4_outputs(10167) <= not b or a;
    layer4_outputs(10168) <= a and b;
    layer4_outputs(10169) <= 1'b0;
    layer4_outputs(10170) <= 1'b0;
    layer4_outputs(10171) <= 1'b1;
    layer4_outputs(10172) <= not b or a;
    layer4_outputs(10173) <= 1'b1;
    layer4_outputs(10174) <= a;
    layer4_outputs(10175) <= b and not a;
    layer4_outputs(10176) <= 1'b1;
    layer4_outputs(10177) <= a xor b;
    layer4_outputs(10178) <= not a or b;
    layer4_outputs(10179) <= a or b;
    layer4_outputs(10180) <= b and not a;
    layer4_outputs(10181) <= a;
    layer4_outputs(10182) <= a;
    layer4_outputs(10183) <= not b;
    layer4_outputs(10184) <= not (a xor b);
    layer4_outputs(10185) <= 1'b1;
    layer4_outputs(10186) <= a and not b;
    layer4_outputs(10187) <= 1'b0;
    layer4_outputs(10188) <= a or b;
    layer4_outputs(10189) <= not (a and b);
    layer4_outputs(10190) <= a and b;
    layer4_outputs(10191) <= a and not b;
    layer4_outputs(10192) <= not a;
    layer4_outputs(10193) <= not a or b;
    layer4_outputs(10194) <= not b;
    layer4_outputs(10195) <= a and not b;
    layer4_outputs(10196) <= 1'b0;
    layer4_outputs(10197) <= not (a xor b);
    layer4_outputs(10198) <= a;
    layer4_outputs(10199) <= a and b;
    layer4_outputs(10200) <= not b;
    layer4_outputs(10201) <= not a or b;
    layer4_outputs(10202) <= not (a or b);
    layer4_outputs(10203) <= b;
    layer4_outputs(10204) <= a and b;
    layer4_outputs(10205) <= not (a or b);
    layer4_outputs(10206) <= a;
    layer4_outputs(10207) <= not a;
    layer4_outputs(10208) <= 1'b0;
    layer4_outputs(10209) <= not (a xor b);
    layer4_outputs(10210) <= b and not a;
    layer4_outputs(10211) <= a;
    layer4_outputs(10212) <= b;
    layer4_outputs(10213) <= a or b;
    layer4_outputs(10214) <= not a;
    layer4_outputs(10215) <= a or b;
    layer4_outputs(10216) <= a and b;
    layer4_outputs(10217) <= a and b;
    layer4_outputs(10218) <= not a or b;
    layer4_outputs(10219) <= 1'b1;
    layer4_outputs(10220) <= a or b;
    layer4_outputs(10221) <= a and not b;
    layer4_outputs(10222) <= 1'b0;
    layer4_outputs(10223) <= not (a xor b);
    layer4_outputs(10224) <= a and b;
    layer4_outputs(10225) <= a xor b;
    layer4_outputs(10226) <= b;
    layer4_outputs(10227) <= not a or b;
    layer4_outputs(10228) <= 1'b1;
    layer4_outputs(10229) <= not b;
    layer4_outputs(10230) <= a and b;
    layer4_outputs(10231) <= a xor b;
    layer4_outputs(10232) <= not (a or b);
    layer4_outputs(10233) <= not (a and b);
    layer4_outputs(10234) <= b;
    layer4_outputs(10235) <= not b;
    layer4_outputs(10236) <= a or b;
    layer4_outputs(10237) <= 1'b1;
    layer4_outputs(10238) <= not b;
    layer4_outputs(10239) <= a and not b;
    layer5_outputs(0) <= not a or b;
    layer5_outputs(1) <= a xor b;
    layer5_outputs(2) <= not b;
    layer5_outputs(3) <= not a or b;
    layer5_outputs(4) <= not a;
    layer5_outputs(5) <= not b or a;
    layer5_outputs(6) <= not a or b;
    layer5_outputs(7) <= 1'b0;
    layer5_outputs(8) <= not a or b;
    layer5_outputs(9) <= not a;
    layer5_outputs(10) <= a or b;
    layer5_outputs(11) <= a or b;
    layer5_outputs(12) <= not a;
    layer5_outputs(13) <= a;
    layer5_outputs(14) <= not (a and b);
    layer5_outputs(15) <= not a;
    layer5_outputs(16) <= a and b;
    layer5_outputs(17) <= a xor b;
    layer5_outputs(18) <= not b or a;
    layer5_outputs(19) <= not a;
    layer5_outputs(20) <= not (a and b);
    layer5_outputs(21) <= not a or b;
    layer5_outputs(22) <= not a;
    layer5_outputs(23) <= b;
    layer5_outputs(24) <= b;
    layer5_outputs(25) <= not b;
    layer5_outputs(26) <= not (a or b);
    layer5_outputs(27) <= not a;
    layer5_outputs(28) <= not a or b;
    layer5_outputs(29) <= not (a or b);
    layer5_outputs(30) <= not b;
    layer5_outputs(31) <= a;
    layer5_outputs(32) <= a or b;
    layer5_outputs(33) <= not b;
    layer5_outputs(34) <= a xor b;
    layer5_outputs(35) <= not a;
    layer5_outputs(36) <= not b;
    layer5_outputs(37) <= not a or b;
    layer5_outputs(38) <= b;
    layer5_outputs(39) <= a xor b;
    layer5_outputs(40) <= a and b;
    layer5_outputs(41) <= b;
    layer5_outputs(42) <= not (a and b);
    layer5_outputs(43) <= not b;
    layer5_outputs(44) <= not b;
    layer5_outputs(45) <= not b or a;
    layer5_outputs(46) <= a or b;
    layer5_outputs(47) <= not (a and b);
    layer5_outputs(48) <= a and b;
    layer5_outputs(49) <= a;
    layer5_outputs(50) <= a or b;
    layer5_outputs(51) <= not b;
    layer5_outputs(52) <= not a;
    layer5_outputs(53) <= 1'b1;
    layer5_outputs(54) <= b;
    layer5_outputs(55) <= not a or b;
    layer5_outputs(56) <= not a;
    layer5_outputs(57) <= b;
    layer5_outputs(58) <= not a;
    layer5_outputs(59) <= b and not a;
    layer5_outputs(60) <= a and not b;
    layer5_outputs(61) <= not (a xor b);
    layer5_outputs(62) <= a and not b;
    layer5_outputs(63) <= not b;
    layer5_outputs(64) <= a and b;
    layer5_outputs(65) <= not b or a;
    layer5_outputs(66) <= not a or b;
    layer5_outputs(67) <= not a or b;
    layer5_outputs(68) <= b;
    layer5_outputs(69) <= not (a or b);
    layer5_outputs(70) <= b;
    layer5_outputs(71) <= not (a and b);
    layer5_outputs(72) <= a and not b;
    layer5_outputs(73) <= not a or b;
    layer5_outputs(74) <= not a or b;
    layer5_outputs(75) <= b;
    layer5_outputs(76) <= a;
    layer5_outputs(77) <= a;
    layer5_outputs(78) <= not b;
    layer5_outputs(79) <= 1'b0;
    layer5_outputs(80) <= not b;
    layer5_outputs(81) <= 1'b0;
    layer5_outputs(82) <= b;
    layer5_outputs(83) <= not b;
    layer5_outputs(84) <= a;
    layer5_outputs(85) <= not b;
    layer5_outputs(86) <= not a;
    layer5_outputs(87) <= b;
    layer5_outputs(88) <= a or b;
    layer5_outputs(89) <= not b or a;
    layer5_outputs(90) <= 1'b0;
    layer5_outputs(91) <= not (a and b);
    layer5_outputs(92) <= a or b;
    layer5_outputs(93) <= not (a or b);
    layer5_outputs(94) <= a and b;
    layer5_outputs(95) <= b and not a;
    layer5_outputs(96) <= a and not b;
    layer5_outputs(97) <= b;
    layer5_outputs(98) <= a and b;
    layer5_outputs(99) <= not a or b;
    layer5_outputs(100) <= not b or a;
    layer5_outputs(101) <= not a;
    layer5_outputs(102) <= b and not a;
    layer5_outputs(103) <= a or b;
    layer5_outputs(104) <= not b;
    layer5_outputs(105) <= not b;
    layer5_outputs(106) <= not (a and b);
    layer5_outputs(107) <= not (a and b);
    layer5_outputs(108) <= a and not b;
    layer5_outputs(109) <= not b;
    layer5_outputs(110) <= a or b;
    layer5_outputs(111) <= not (a xor b);
    layer5_outputs(112) <= not a or b;
    layer5_outputs(113) <= not b or a;
    layer5_outputs(114) <= a or b;
    layer5_outputs(115) <= not a;
    layer5_outputs(116) <= b;
    layer5_outputs(117) <= b;
    layer5_outputs(118) <= a xor b;
    layer5_outputs(119) <= not b;
    layer5_outputs(120) <= not (a and b);
    layer5_outputs(121) <= not b;
    layer5_outputs(122) <= a and not b;
    layer5_outputs(123) <= a and b;
    layer5_outputs(124) <= not a;
    layer5_outputs(125) <= 1'b0;
    layer5_outputs(126) <= b;
    layer5_outputs(127) <= not b;
    layer5_outputs(128) <= not a;
    layer5_outputs(129) <= a;
    layer5_outputs(130) <= not b or a;
    layer5_outputs(131) <= a and not b;
    layer5_outputs(132) <= not a;
    layer5_outputs(133) <= a;
    layer5_outputs(134) <= not b or a;
    layer5_outputs(135) <= not b;
    layer5_outputs(136) <= a and b;
    layer5_outputs(137) <= not (a xor b);
    layer5_outputs(138) <= not b or a;
    layer5_outputs(139) <= b;
    layer5_outputs(140) <= 1'b1;
    layer5_outputs(141) <= not b;
    layer5_outputs(142) <= not a;
    layer5_outputs(143) <= not b or a;
    layer5_outputs(144) <= 1'b0;
    layer5_outputs(145) <= not a;
    layer5_outputs(146) <= 1'b1;
    layer5_outputs(147) <= a or b;
    layer5_outputs(148) <= not b;
    layer5_outputs(149) <= 1'b1;
    layer5_outputs(150) <= a;
    layer5_outputs(151) <= a or b;
    layer5_outputs(152) <= b and not a;
    layer5_outputs(153) <= not (a and b);
    layer5_outputs(154) <= a and b;
    layer5_outputs(155) <= not a;
    layer5_outputs(156) <= a or b;
    layer5_outputs(157) <= not a or b;
    layer5_outputs(158) <= not (a or b);
    layer5_outputs(159) <= not a;
    layer5_outputs(160) <= a or b;
    layer5_outputs(161) <= not b;
    layer5_outputs(162) <= not b;
    layer5_outputs(163) <= a xor b;
    layer5_outputs(164) <= a and not b;
    layer5_outputs(165) <= 1'b1;
    layer5_outputs(166) <= 1'b1;
    layer5_outputs(167) <= not (a and b);
    layer5_outputs(168) <= b and not a;
    layer5_outputs(169) <= not (a and b);
    layer5_outputs(170) <= not b or a;
    layer5_outputs(171) <= not a;
    layer5_outputs(172) <= not b;
    layer5_outputs(173) <= 1'b0;
    layer5_outputs(174) <= 1'b1;
    layer5_outputs(175) <= not a;
    layer5_outputs(176) <= not (a and b);
    layer5_outputs(177) <= b and not a;
    layer5_outputs(178) <= a xor b;
    layer5_outputs(179) <= not b or a;
    layer5_outputs(180) <= a or b;
    layer5_outputs(181) <= not (a xor b);
    layer5_outputs(182) <= b;
    layer5_outputs(183) <= not (a and b);
    layer5_outputs(184) <= not b or a;
    layer5_outputs(185) <= b;
    layer5_outputs(186) <= not (a or b);
    layer5_outputs(187) <= 1'b1;
    layer5_outputs(188) <= 1'b0;
    layer5_outputs(189) <= 1'b0;
    layer5_outputs(190) <= not b;
    layer5_outputs(191) <= a and b;
    layer5_outputs(192) <= a and b;
    layer5_outputs(193) <= not (a and b);
    layer5_outputs(194) <= not (a or b);
    layer5_outputs(195) <= not (a and b);
    layer5_outputs(196) <= not (a or b);
    layer5_outputs(197) <= not a;
    layer5_outputs(198) <= a or b;
    layer5_outputs(199) <= b;
    layer5_outputs(200) <= not b or a;
    layer5_outputs(201) <= not (a xor b);
    layer5_outputs(202) <= not (a and b);
    layer5_outputs(203) <= b;
    layer5_outputs(204) <= not b;
    layer5_outputs(205) <= a;
    layer5_outputs(206) <= not (a and b);
    layer5_outputs(207) <= a;
    layer5_outputs(208) <= not (a and b);
    layer5_outputs(209) <= not a;
    layer5_outputs(210) <= not (a xor b);
    layer5_outputs(211) <= not a;
    layer5_outputs(212) <= a;
    layer5_outputs(213) <= a;
    layer5_outputs(214) <= not b;
    layer5_outputs(215) <= a and not b;
    layer5_outputs(216) <= not (a and b);
    layer5_outputs(217) <= a;
    layer5_outputs(218) <= not b;
    layer5_outputs(219) <= b;
    layer5_outputs(220) <= not (a and b);
    layer5_outputs(221) <= b and not a;
    layer5_outputs(222) <= not b or a;
    layer5_outputs(223) <= b and not a;
    layer5_outputs(224) <= 1'b1;
    layer5_outputs(225) <= not b;
    layer5_outputs(226) <= b;
    layer5_outputs(227) <= not b;
    layer5_outputs(228) <= a and not b;
    layer5_outputs(229) <= a and b;
    layer5_outputs(230) <= a or b;
    layer5_outputs(231) <= 1'b0;
    layer5_outputs(232) <= b and not a;
    layer5_outputs(233) <= a and not b;
    layer5_outputs(234) <= not b;
    layer5_outputs(235) <= not (a or b);
    layer5_outputs(236) <= not b;
    layer5_outputs(237) <= not a or b;
    layer5_outputs(238) <= not a or b;
    layer5_outputs(239) <= not b;
    layer5_outputs(240) <= not a or b;
    layer5_outputs(241) <= a;
    layer5_outputs(242) <= not b or a;
    layer5_outputs(243) <= a and b;
    layer5_outputs(244) <= a and not b;
    layer5_outputs(245) <= not a;
    layer5_outputs(246) <= not b;
    layer5_outputs(247) <= not b;
    layer5_outputs(248) <= not a or b;
    layer5_outputs(249) <= not b;
    layer5_outputs(250) <= 1'b1;
    layer5_outputs(251) <= 1'b0;
    layer5_outputs(252) <= not b;
    layer5_outputs(253) <= a and b;
    layer5_outputs(254) <= a xor b;
    layer5_outputs(255) <= not a or b;
    layer5_outputs(256) <= not (a xor b);
    layer5_outputs(257) <= not b;
    layer5_outputs(258) <= 1'b0;
    layer5_outputs(259) <= 1'b1;
    layer5_outputs(260) <= a and b;
    layer5_outputs(261) <= b and not a;
    layer5_outputs(262) <= not b or a;
    layer5_outputs(263) <= not b or a;
    layer5_outputs(264) <= not b or a;
    layer5_outputs(265) <= not a;
    layer5_outputs(266) <= a and not b;
    layer5_outputs(267) <= a and b;
    layer5_outputs(268) <= b;
    layer5_outputs(269) <= not b or a;
    layer5_outputs(270) <= a xor b;
    layer5_outputs(271) <= not (a and b);
    layer5_outputs(272) <= not a;
    layer5_outputs(273) <= a xor b;
    layer5_outputs(274) <= 1'b1;
    layer5_outputs(275) <= not b or a;
    layer5_outputs(276) <= not (a and b);
    layer5_outputs(277) <= not a;
    layer5_outputs(278) <= not a or b;
    layer5_outputs(279) <= not a or b;
    layer5_outputs(280) <= a and b;
    layer5_outputs(281) <= not b or a;
    layer5_outputs(282) <= a and b;
    layer5_outputs(283) <= a or b;
    layer5_outputs(284) <= a or b;
    layer5_outputs(285) <= b and not a;
    layer5_outputs(286) <= b;
    layer5_outputs(287) <= not b or a;
    layer5_outputs(288) <= not a;
    layer5_outputs(289) <= not b;
    layer5_outputs(290) <= a and not b;
    layer5_outputs(291) <= not (a or b);
    layer5_outputs(292) <= not (a or b);
    layer5_outputs(293) <= not b or a;
    layer5_outputs(294) <= not (a or b);
    layer5_outputs(295) <= a xor b;
    layer5_outputs(296) <= a xor b;
    layer5_outputs(297) <= a;
    layer5_outputs(298) <= b;
    layer5_outputs(299) <= b and not a;
    layer5_outputs(300) <= not b;
    layer5_outputs(301) <= not b;
    layer5_outputs(302) <= not (a or b);
    layer5_outputs(303) <= a;
    layer5_outputs(304) <= not a;
    layer5_outputs(305) <= b;
    layer5_outputs(306) <= not b;
    layer5_outputs(307) <= a and not b;
    layer5_outputs(308) <= not b or a;
    layer5_outputs(309) <= b and not a;
    layer5_outputs(310) <= not a;
    layer5_outputs(311) <= not b;
    layer5_outputs(312) <= not b;
    layer5_outputs(313) <= not a;
    layer5_outputs(314) <= b;
    layer5_outputs(315) <= b and not a;
    layer5_outputs(316) <= a and b;
    layer5_outputs(317) <= 1'b0;
    layer5_outputs(318) <= not b;
    layer5_outputs(319) <= not a;
    layer5_outputs(320) <= a xor b;
    layer5_outputs(321) <= b;
    layer5_outputs(322) <= a;
    layer5_outputs(323) <= not b or a;
    layer5_outputs(324) <= not (a and b);
    layer5_outputs(325) <= not b;
    layer5_outputs(326) <= a and not b;
    layer5_outputs(327) <= not (a or b);
    layer5_outputs(328) <= a or b;
    layer5_outputs(329) <= a or b;
    layer5_outputs(330) <= b;
    layer5_outputs(331) <= not (a or b);
    layer5_outputs(332) <= not b;
    layer5_outputs(333) <= not a;
    layer5_outputs(334) <= a or b;
    layer5_outputs(335) <= not (a and b);
    layer5_outputs(336) <= b;
    layer5_outputs(337) <= a or b;
    layer5_outputs(338) <= not a or b;
    layer5_outputs(339) <= not (a xor b);
    layer5_outputs(340) <= not b;
    layer5_outputs(341) <= b;
    layer5_outputs(342) <= not a or b;
    layer5_outputs(343) <= b;
    layer5_outputs(344) <= a and b;
    layer5_outputs(345) <= a;
    layer5_outputs(346) <= a;
    layer5_outputs(347) <= b;
    layer5_outputs(348) <= 1'b0;
    layer5_outputs(349) <= a;
    layer5_outputs(350) <= 1'b1;
    layer5_outputs(351) <= a;
    layer5_outputs(352) <= not b or a;
    layer5_outputs(353) <= not (a xor b);
    layer5_outputs(354) <= a and b;
    layer5_outputs(355) <= not b;
    layer5_outputs(356) <= a;
    layer5_outputs(357) <= 1'b0;
    layer5_outputs(358) <= b and not a;
    layer5_outputs(359) <= b;
    layer5_outputs(360) <= b and not a;
    layer5_outputs(361) <= not (a and b);
    layer5_outputs(362) <= not (a and b);
    layer5_outputs(363) <= a or b;
    layer5_outputs(364) <= not a or b;
    layer5_outputs(365) <= not a;
    layer5_outputs(366) <= 1'b0;
    layer5_outputs(367) <= not (a and b);
    layer5_outputs(368) <= a and not b;
    layer5_outputs(369) <= not (a and b);
    layer5_outputs(370) <= b;
    layer5_outputs(371) <= not a or b;
    layer5_outputs(372) <= 1'b1;
    layer5_outputs(373) <= a xor b;
    layer5_outputs(374) <= b and not a;
    layer5_outputs(375) <= not (a xor b);
    layer5_outputs(376) <= a;
    layer5_outputs(377) <= not b;
    layer5_outputs(378) <= not a;
    layer5_outputs(379) <= a and b;
    layer5_outputs(380) <= a and not b;
    layer5_outputs(381) <= a and b;
    layer5_outputs(382) <= not b or a;
    layer5_outputs(383) <= b;
    layer5_outputs(384) <= not b or a;
    layer5_outputs(385) <= a;
    layer5_outputs(386) <= not a or b;
    layer5_outputs(387) <= not (a xor b);
    layer5_outputs(388) <= a and b;
    layer5_outputs(389) <= not b or a;
    layer5_outputs(390) <= not (a or b);
    layer5_outputs(391) <= not (a xor b);
    layer5_outputs(392) <= 1'b1;
    layer5_outputs(393) <= b;
    layer5_outputs(394) <= not a;
    layer5_outputs(395) <= a and b;
    layer5_outputs(396) <= not a or b;
    layer5_outputs(397) <= b;
    layer5_outputs(398) <= a;
    layer5_outputs(399) <= not (a xor b);
    layer5_outputs(400) <= not b;
    layer5_outputs(401) <= not b;
    layer5_outputs(402) <= a or b;
    layer5_outputs(403) <= a and not b;
    layer5_outputs(404) <= 1'b1;
    layer5_outputs(405) <= a and not b;
    layer5_outputs(406) <= a and not b;
    layer5_outputs(407) <= b;
    layer5_outputs(408) <= a or b;
    layer5_outputs(409) <= not b or a;
    layer5_outputs(410) <= not b or a;
    layer5_outputs(411) <= not (a and b);
    layer5_outputs(412) <= not a or b;
    layer5_outputs(413) <= not a;
    layer5_outputs(414) <= not (a or b);
    layer5_outputs(415) <= not a;
    layer5_outputs(416) <= not (a and b);
    layer5_outputs(417) <= 1'b0;
    layer5_outputs(418) <= 1'b0;
    layer5_outputs(419) <= not b;
    layer5_outputs(420) <= not b;
    layer5_outputs(421) <= not (a or b);
    layer5_outputs(422) <= b and not a;
    layer5_outputs(423) <= not (a and b);
    layer5_outputs(424) <= a;
    layer5_outputs(425) <= b;
    layer5_outputs(426) <= a and not b;
    layer5_outputs(427) <= not a or b;
    layer5_outputs(428) <= a and b;
    layer5_outputs(429) <= not b or a;
    layer5_outputs(430) <= not b;
    layer5_outputs(431) <= not a;
    layer5_outputs(432) <= a;
    layer5_outputs(433) <= a and b;
    layer5_outputs(434) <= not (a and b);
    layer5_outputs(435) <= 1'b1;
    layer5_outputs(436) <= a;
    layer5_outputs(437) <= 1'b1;
    layer5_outputs(438) <= b and not a;
    layer5_outputs(439) <= a and not b;
    layer5_outputs(440) <= 1'b0;
    layer5_outputs(441) <= a xor b;
    layer5_outputs(442) <= a;
    layer5_outputs(443) <= not (a xor b);
    layer5_outputs(444) <= not a;
    layer5_outputs(445) <= not a or b;
    layer5_outputs(446) <= a and not b;
    layer5_outputs(447) <= a xor b;
    layer5_outputs(448) <= not (a xor b);
    layer5_outputs(449) <= not a or b;
    layer5_outputs(450) <= b and not a;
    layer5_outputs(451) <= not b;
    layer5_outputs(452) <= not (a and b);
    layer5_outputs(453) <= a or b;
    layer5_outputs(454) <= b and not a;
    layer5_outputs(455) <= not (a and b);
    layer5_outputs(456) <= not (a and b);
    layer5_outputs(457) <= a and b;
    layer5_outputs(458) <= 1'b0;
    layer5_outputs(459) <= not b;
    layer5_outputs(460) <= a and b;
    layer5_outputs(461) <= a and not b;
    layer5_outputs(462) <= a;
    layer5_outputs(463) <= 1'b1;
    layer5_outputs(464) <= 1'b0;
    layer5_outputs(465) <= not a;
    layer5_outputs(466) <= a and b;
    layer5_outputs(467) <= a;
    layer5_outputs(468) <= not a;
    layer5_outputs(469) <= not (a and b);
    layer5_outputs(470) <= not (a xor b);
    layer5_outputs(471) <= b and not a;
    layer5_outputs(472) <= not b or a;
    layer5_outputs(473) <= not a or b;
    layer5_outputs(474) <= a;
    layer5_outputs(475) <= not a;
    layer5_outputs(476) <= not (a and b);
    layer5_outputs(477) <= not a or b;
    layer5_outputs(478) <= not a or b;
    layer5_outputs(479) <= not a or b;
    layer5_outputs(480) <= not (a and b);
    layer5_outputs(481) <= 1'b1;
    layer5_outputs(482) <= a and not b;
    layer5_outputs(483) <= not a or b;
    layer5_outputs(484) <= not a or b;
    layer5_outputs(485) <= a;
    layer5_outputs(486) <= b;
    layer5_outputs(487) <= b;
    layer5_outputs(488) <= not a;
    layer5_outputs(489) <= a;
    layer5_outputs(490) <= not (a or b);
    layer5_outputs(491) <= a or b;
    layer5_outputs(492) <= not a or b;
    layer5_outputs(493) <= not a;
    layer5_outputs(494) <= not a;
    layer5_outputs(495) <= not a or b;
    layer5_outputs(496) <= b;
    layer5_outputs(497) <= 1'b0;
    layer5_outputs(498) <= a;
    layer5_outputs(499) <= not b or a;
    layer5_outputs(500) <= not a or b;
    layer5_outputs(501) <= b;
    layer5_outputs(502) <= not b;
    layer5_outputs(503) <= not a;
    layer5_outputs(504) <= not a or b;
    layer5_outputs(505) <= 1'b1;
    layer5_outputs(506) <= a;
    layer5_outputs(507) <= not (a or b);
    layer5_outputs(508) <= not (a xor b);
    layer5_outputs(509) <= a xor b;
    layer5_outputs(510) <= 1'b0;
    layer5_outputs(511) <= not a;
    layer5_outputs(512) <= b;
    layer5_outputs(513) <= a and b;
    layer5_outputs(514) <= a;
    layer5_outputs(515) <= a;
    layer5_outputs(516) <= not (a and b);
    layer5_outputs(517) <= b;
    layer5_outputs(518) <= not a;
    layer5_outputs(519) <= a;
    layer5_outputs(520) <= not (a or b);
    layer5_outputs(521) <= 1'b1;
    layer5_outputs(522) <= b;
    layer5_outputs(523) <= b;
    layer5_outputs(524) <= 1'b1;
    layer5_outputs(525) <= a and not b;
    layer5_outputs(526) <= 1'b1;
    layer5_outputs(527) <= not (a or b);
    layer5_outputs(528) <= not (a or b);
    layer5_outputs(529) <= not (a and b);
    layer5_outputs(530) <= a and b;
    layer5_outputs(531) <= not (a or b);
    layer5_outputs(532) <= a and not b;
    layer5_outputs(533) <= 1'b1;
    layer5_outputs(534) <= b and not a;
    layer5_outputs(535) <= 1'b0;
    layer5_outputs(536) <= not a;
    layer5_outputs(537) <= not (a xor b);
    layer5_outputs(538) <= b and not a;
    layer5_outputs(539) <= not a or b;
    layer5_outputs(540) <= a or b;
    layer5_outputs(541) <= not (a and b);
    layer5_outputs(542) <= a or b;
    layer5_outputs(543) <= a or b;
    layer5_outputs(544) <= not (a or b);
    layer5_outputs(545) <= not b;
    layer5_outputs(546) <= not a;
    layer5_outputs(547) <= 1'b0;
    layer5_outputs(548) <= not (a xor b);
    layer5_outputs(549) <= not (a or b);
    layer5_outputs(550) <= not a;
    layer5_outputs(551) <= not (a and b);
    layer5_outputs(552) <= b;
    layer5_outputs(553) <= a or b;
    layer5_outputs(554) <= not (a or b);
    layer5_outputs(555) <= a or b;
    layer5_outputs(556) <= not a;
    layer5_outputs(557) <= a or b;
    layer5_outputs(558) <= a;
    layer5_outputs(559) <= not (a xor b);
    layer5_outputs(560) <= not a;
    layer5_outputs(561) <= a;
    layer5_outputs(562) <= b and not a;
    layer5_outputs(563) <= a;
    layer5_outputs(564) <= not (a or b);
    layer5_outputs(565) <= a and b;
    layer5_outputs(566) <= not a or b;
    layer5_outputs(567) <= not (a or b);
    layer5_outputs(568) <= 1'b1;
    layer5_outputs(569) <= not (a and b);
    layer5_outputs(570) <= a and not b;
    layer5_outputs(571) <= not b or a;
    layer5_outputs(572) <= b and not a;
    layer5_outputs(573) <= a;
    layer5_outputs(574) <= a and not b;
    layer5_outputs(575) <= not b or a;
    layer5_outputs(576) <= a or b;
    layer5_outputs(577) <= a xor b;
    layer5_outputs(578) <= b;
    layer5_outputs(579) <= not (a and b);
    layer5_outputs(580) <= a xor b;
    layer5_outputs(581) <= not a or b;
    layer5_outputs(582) <= a and b;
    layer5_outputs(583) <= not a or b;
    layer5_outputs(584) <= 1'b1;
    layer5_outputs(585) <= a;
    layer5_outputs(586) <= not b;
    layer5_outputs(587) <= 1'b1;
    layer5_outputs(588) <= a and b;
    layer5_outputs(589) <= a;
    layer5_outputs(590) <= not b or a;
    layer5_outputs(591) <= 1'b0;
    layer5_outputs(592) <= b and not a;
    layer5_outputs(593) <= a and b;
    layer5_outputs(594) <= not a;
    layer5_outputs(595) <= not (a and b);
    layer5_outputs(596) <= not (a or b);
    layer5_outputs(597) <= not a;
    layer5_outputs(598) <= not a;
    layer5_outputs(599) <= b;
    layer5_outputs(600) <= a;
    layer5_outputs(601) <= b;
    layer5_outputs(602) <= a;
    layer5_outputs(603) <= not a or b;
    layer5_outputs(604) <= not a;
    layer5_outputs(605) <= not b or a;
    layer5_outputs(606) <= not (a and b);
    layer5_outputs(607) <= a and not b;
    layer5_outputs(608) <= a;
    layer5_outputs(609) <= b;
    layer5_outputs(610) <= b and not a;
    layer5_outputs(611) <= a;
    layer5_outputs(612) <= a;
    layer5_outputs(613) <= a;
    layer5_outputs(614) <= a or b;
    layer5_outputs(615) <= a xor b;
    layer5_outputs(616) <= a and not b;
    layer5_outputs(617) <= 1'b0;
    layer5_outputs(618) <= b and not a;
    layer5_outputs(619) <= a and not b;
    layer5_outputs(620) <= a;
    layer5_outputs(621) <= not a;
    layer5_outputs(622) <= not b or a;
    layer5_outputs(623) <= b;
    layer5_outputs(624) <= a or b;
    layer5_outputs(625) <= not b;
    layer5_outputs(626) <= not a or b;
    layer5_outputs(627) <= a or b;
    layer5_outputs(628) <= not b;
    layer5_outputs(629) <= b;
    layer5_outputs(630) <= b and not a;
    layer5_outputs(631) <= not b;
    layer5_outputs(632) <= 1'b0;
    layer5_outputs(633) <= a;
    layer5_outputs(634) <= not a or b;
    layer5_outputs(635) <= not (a and b);
    layer5_outputs(636) <= b;
    layer5_outputs(637) <= not a;
    layer5_outputs(638) <= not b or a;
    layer5_outputs(639) <= b and not a;
    layer5_outputs(640) <= a;
    layer5_outputs(641) <= a or b;
    layer5_outputs(642) <= a or b;
    layer5_outputs(643) <= a and not b;
    layer5_outputs(644) <= a or b;
    layer5_outputs(645) <= not b or a;
    layer5_outputs(646) <= not a or b;
    layer5_outputs(647) <= not b or a;
    layer5_outputs(648) <= not b or a;
    layer5_outputs(649) <= not b or a;
    layer5_outputs(650) <= b;
    layer5_outputs(651) <= a;
    layer5_outputs(652) <= not a;
    layer5_outputs(653) <= not b;
    layer5_outputs(654) <= not (a and b);
    layer5_outputs(655) <= not (a and b);
    layer5_outputs(656) <= not (a xor b);
    layer5_outputs(657) <= not a;
    layer5_outputs(658) <= not b or a;
    layer5_outputs(659) <= not b;
    layer5_outputs(660) <= a and b;
    layer5_outputs(661) <= a;
    layer5_outputs(662) <= a or b;
    layer5_outputs(663) <= not a;
    layer5_outputs(664) <= not a or b;
    layer5_outputs(665) <= a or b;
    layer5_outputs(666) <= a;
    layer5_outputs(667) <= a and b;
    layer5_outputs(668) <= 1'b0;
    layer5_outputs(669) <= not b or a;
    layer5_outputs(670) <= not (a or b);
    layer5_outputs(671) <= a and b;
    layer5_outputs(672) <= 1'b1;
    layer5_outputs(673) <= b;
    layer5_outputs(674) <= not a;
    layer5_outputs(675) <= b and not a;
    layer5_outputs(676) <= not (a or b);
    layer5_outputs(677) <= not (a and b);
    layer5_outputs(678) <= not a or b;
    layer5_outputs(679) <= not a;
    layer5_outputs(680) <= a and not b;
    layer5_outputs(681) <= not b;
    layer5_outputs(682) <= a or b;
    layer5_outputs(683) <= not b;
    layer5_outputs(684) <= a and not b;
    layer5_outputs(685) <= b and not a;
    layer5_outputs(686) <= b;
    layer5_outputs(687) <= not (a xor b);
    layer5_outputs(688) <= not a or b;
    layer5_outputs(689) <= a;
    layer5_outputs(690) <= a or b;
    layer5_outputs(691) <= a and not b;
    layer5_outputs(692) <= not (a or b);
    layer5_outputs(693) <= b and not a;
    layer5_outputs(694) <= a;
    layer5_outputs(695) <= not b;
    layer5_outputs(696) <= not a;
    layer5_outputs(697) <= a;
    layer5_outputs(698) <= not a;
    layer5_outputs(699) <= not b;
    layer5_outputs(700) <= a;
    layer5_outputs(701) <= b and not a;
    layer5_outputs(702) <= b;
    layer5_outputs(703) <= b;
    layer5_outputs(704) <= not b;
    layer5_outputs(705) <= not a;
    layer5_outputs(706) <= b;
    layer5_outputs(707) <= 1'b0;
    layer5_outputs(708) <= 1'b0;
    layer5_outputs(709) <= not a;
    layer5_outputs(710) <= not a;
    layer5_outputs(711) <= 1'b0;
    layer5_outputs(712) <= a and b;
    layer5_outputs(713) <= not a;
    layer5_outputs(714) <= not a;
    layer5_outputs(715) <= not a;
    layer5_outputs(716) <= not a;
    layer5_outputs(717) <= a;
    layer5_outputs(718) <= a and b;
    layer5_outputs(719) <= not a;
    layer5_outputs(720) <= not a or b;
    layer5_outputs(721) <= not b;
    layer5_outputs(722) <= not a;
    layer5_outputs(723) <= a or b;
    layer5_outputs(724) <= b and not a;
    layer5_outputs(725) <= not b;
    layer5_outputs(726) <= a or b;
    layer5_outputs(727) <= not (a and b);
    layer5_outputs(728) <= a and not b;
    layer5_outputs(729) <= not (a and b);
    layer5_outputs(730) <= not a or b;
    layer5_outputs(731) <= 1'b1;
    layer5_outputs(732) <= not (a and b);
    layer5_outputs(733) <= not b or a;
    layer5_outputs(734) <= a;
    layer5_outputs(735) <= not b;
    layer5_outputs(736) <= not (a or b);
    layer5_outputs(737) <= not a;
    layer5_outputs(738) <= not a;
    layer5_outputs(739) <= a and b;
    layer5_outputs(740) <= a or b;
    layer5_outputs(741) <= 1'b0;
    layer5_outputs(742) <= not a;
    layer5_outputs(743) <= a or b;
    layer5_outputs(744) <= a or b;
    layer5_outputs(745) <= b and not a;
    layer5_outputs(746) <= a and not b;
    layer5_outputs(747) <= a;
    layer5_outputs(748) <= a and not b;
    layer5_outputs(749) <= a or b;
    layer5_outputs(750) <= a;
    layer5_outputs(751) <= a or b;
    layer5_outputs(752) <= a and not b;
    layer5_outputs(753) <= a;
    layer5_outputs(754) <= b;
    layer5_outputs(755) <= not (a or b);
    layer5_outputs(756) <= b;
    layer5_outputs(757) <= not a;
    layer5_outputs(758) <= not a or b;
    layer5_outputs(759) <= a and b;
    layer5_outputs(760) <= not a or b;
    layer5_outputs(761) <= b;
    layer5_outputs(762) <= not (a or b);
    layer5_outputs(763) <= not (a or b);
    layer5_outputs(764) <= a and not b;
    layer5_outputs(765) <= b;
    layer5_outputs(766) <= not b;
    layer5_outputs(767) <= a;
    layer5_outputs(768) <= not a;
    layer5_outputs(769) <= 1'b0;
    layer5_outputs(770) <= not b;
    layer5_outputs(771) <= a and b;
    layer5_outputs(772) <= b and not a;
    layer5_outputs(773) <= 1'b1;
    layer5_outputs(774) <= a and b;
    layer5_outputs(775) <= not b;
    layer5_outputs(776) <= b;
    layer5_outputs(777) <= not b;
    layer5_outputs(778) <= a;
    layer5_outputs(779) <= not b or a;
    layer5_outputs(780) <= not (a or b);
    layer5_outputs(781) <= not (a and b);
    layer5_outputs(782) <= a xor b;
    layer5_outputs(783) <= b and not a;
    layer5_outputs(784) <= not a;
    layer5_outputs(785) <= b and not a;
    layer5_outputs(786) <= a and b;
    layer5_outputs(787) <= a;
    layer5_outputs(788) <= a and not b;
    layer5_outputs(789) <= a xor b;
    layer5_outputs(790) <= b;
    layer5_outputs(791) <= not a;
    layer5_outputs(792) <= 1'b0;
    layer5_outputs(793) <= b and not a;
    layer5_outputs(794) <= b and not a;
    layer5_outputs(795) <= b and not a;
    layer5_outputs(796) <= not b or a;
    layer5_outputs(797) <= not b;
    layer5_outputs(798) <= a and not b;
    layer5_outputs(799) <= not a;
    layer5_outputs(800) <= b and not a;
    layer5_outputs(801) <= not b or a;
    layer5_outputs(802) <= a;
    layer5_outputs(803) <= not b;
    layer5_outputs(804) <= not b;
    layer5_outputs(805) <= a and b;
    layer5_outputs(806) <= a;
    layer5_outputs(807) <= not (a and b);
    layer5_outputs(808) <= 1'b1;
    layer5_outputs(809) <= a xor b;
    layer5_outputs(810) <= not b;
    layer5_outputs(811) <= not (a or b);
    layer5_outputs(812) <= 1'b0;
    layer5_outputs(813) <= not a or b;
    layer5_outputs(814) <= a and b;
    layer5_outputs(815) <= b;
    layer5_outputs(816) <= not b;
    layer5_outputs(817) <= b;
    layer5_outputs(818) <= not a;
    layer5_outputs(819) <= not (a xor b);
    layer5_outputs(820) <= a;
    layer5_outputs(821) <= b;
    layer5_outputs(822) <= 1'b1;
    layer5_outputs(823) <= 1'b0;
    layer5_outputs(824) <= b;
    layer5_outputs(825) <= a or b;
    layer5_outputs(826) <= b and not a;
    layer5_outputs(827) <= not b or a;
    layer5_outputs(828) <= b;
    layer5_outputs(829) <= not a;
    layer5_outputs(830) <= not a;
    layer5_outputs(831) <= a;
    layer5_outputs(832) <= b;
    layer5_outputs(833) <= a;
    layer5_outputs(834) <= not (a xor b);
    layer5_outputs(835) <= not b;
    layer5_outputs(836) <= a or b;
    layer5_outputs(837) <= a and not b;
    layer5_outputs(838) <= a xor b;
    layer5_outputs(839) <= not (a xor b);
    layer5_outputs(840) <= a or b;
    layer5_outputs(841) <= 1'b1;
    layer5_outputs(842) <= 1'b1;
    layer5_outputs(843) <= a xor b;
    layer5_outputs(844) <= a or b;
    layer5_outputs(845) <= not (a and b);
    layer5_outputs(846) <= a;
    layer5_outputs(847) <= not (a and b);
    layer5_outputs(848) <= not a;
    layer5_outputs(849) <= a xor b;
    layer5_outputs(850) <= a and not b;
    layer5_outputs(851) <= not a;
    layer5_outputs(852) <= a and not b;
    layer5_outputs(853) <= not (a and b);
    layer5_outputs(854) <= b and not a;
    layer5_outputs(855) <= a and b;
    layer5_outputs(856) <= 1'b0;
    layer5_outputs(857) <= a;
    layer5_outputs(858) <= a xor b;
    layer5_outputs(859) <= a and not b;
    layer5_outputs(860) <= a;
    layer5_outputs(861) <= b;
    layer5_outputs(862) <= not a;
    layer5_outputs(863) <= a and b;
    layer5_outputs(864) <= not b;
    layer5_outputs(865) <= not b;
    layer5_outputs(866) <= a or b;
    layer5_outputs(867) <= b;
    layer5_outputs(868) <= b;
    layer5_outputs(869) <= a and b;
    layer5_outputs(870) <= not b or a;
    layer5_outputs(871) <= not (a and b);
    layer5_outputs(872) <= b and not a;
    layer5_outputs(873) <= not b or a;
    layer5_outputs(874) <= not a or b;
    layer5_outputs(875) <= b and not a;
    layer5_outputs(876) <= a or b;
    layer5_outputs(877) <= not a or b;
    layer5_outputs(878) <= a or b;
    layer5_outputs(879) <= not (a xor b);
    layer5_outputs(880) <= a and not b;
    layer5_outputs(881) <= b and not a;
    layer5_outputs(882) <= not a or b;
    layer5_outputs(883) <= not (a xor b);
    layer5_outputs(884) <= not b;
    layer5_outputs(885) <= not a or b;
    layer5_outputs(886) <= 1'b0;
    layer5_outputs(887) <= not b;
    layer5_outputs(888) <= a xor b;
    layer5_outputs(889) <= a or b;
    layer5_outputs(890) <= not a or b;
    layer5_outputs(891) <= not a;
    layer5_outputs(892) <= a;
    layer5_outputs(893) <= b;
    layer5_outputs(894) <= a and not b;
    layer5_outputs(895) <= not b or a;
    layer5_outputs(896) <= not a;
    layer5_outputs(897) <= b;
    layer5_outputs(898) <= a or b;
    layer5_outputs(899) <= b;
    layer5_outputs(900) <= not (a and b);
    layer5_outputs(901) <= a and b;
    layer5_outputs(902) <= a and not b;
    layer5_outputs(903) <= a and not b;
    layer5_outputs(904) <= 1'b1;
    layer5_outputs(905) <= not b;
    layer5_outputs(906) <= not (a or b);
    layer5_outputs(907) <= not (a xor b);
    layer5_outputs(908) <= not b;
    layer5_outputs(909) <= not b;
    layer5_outputs(910) <= not (a xor b);
    layer5_outputs(911) <= not a;
    layer5_outputs(912) <= a;
    layer5_outputs(913) <= not (a xor b);
    layer5_outputs(914) <= a and not b;
    layer5_outputs(915) <= b and not a;
    layer5_outputs(916) <= not a or b;
    layer5_outputs(917) <= not a or b;
    layer5_outputs(918) <= b;
    layer5_outputs(919) <= not b or a;
    layer5_outputs(920) <= a and b;
    layer5_outputs(921) <= not b;
    layer5_outputs(922) <= a and b;
    layer5_outputs(923) <= a;
    layer5_outputs(924) <= b and not a;
    layer5_outputs(925) <= not a or b;
    layer5_outputs(926) <= b and not a;
    layer5_outputs(927) <= a or b;
    layer5_outputs(928) <= a and not b;
    layer5_outputs(929) <= 1'b1;
    layer5_outputs(930) <= not b or a;
    layer5_outputs(931) <= a or b;
    layer5_outputs(932) <= a or b;
    layer5_outputs(933) <= 1'b1;
    layer5_outputs(934) <= a;
    layer5_outputs(935) <= a;
    layer5_outputs(936) <= not b or a;
    layer5_outputs(937) <= b;
    layer5_outputs(938) <= not a or b;
    layer5_outputs(939) <= not b;
    layer5_outputs(940) <= not a;
    layer5_outputs(941) <= 1'b0;
    layer5_outputs(942) <= a or b;
    layer5_outputs(943) <= not b;
    layer5_outputs(944) <= not b or a;
    layer5_outputs(945) <= a xor b;
    layer5_outputs(946) <= not a or b;
    layer5_outputs(947) <= 1'b0;
    layer5_outputs(948) <= a or b;
    layer5_outputs(949) <= a and not b;
    layer5_outputs(950) <= b;
    layer5_outputs(951) <= not b;
    layer5_outputs(952) <= a;
    layer5_outputs(953) <= not (a and b);
    layer5_outputs(954) <= not b or a;
    layer5_outputs(955) <= b;
    layer5_outputs(956) <= not (a and b);
    layer5_outputs(957) <= a and b;
    layer5_outputs(958) <= not b;
    layer5_outputs(959) <= not b or a;
    layer5_outputs(960) <= not b;
    layer5_outputs(961) <= b and not a;
    layer5_outputs(962) <= not (a or b);
    layer5_outputs(963) <= not (a or b);
    layer5_outputs(964) <= not a or b;
    layer5_outputs(965) <= not b;
    layer5_outputs(966) <= not b or a;
    layer5_outputs(967) <= not b;
    layer5_outputs(968) <= not a or b;
    layer5_outputs(969) <= 1'b1;
    layer5_outputs(970) <= a or b;
    layer5_outputs(971) <= b and not a;
    layer5_outputs(972) <= not a or b;
    layer5_outputs(973) <= not (a or b);
    layer5_outputs(974) <= a and b;
    layer5_outputs(975) <= not (a or b);
    layer5_outputs(976) <= b;
    layer5_outputs(977) <= a and not b;
    layer5_outputs(978) <= a;
    layer5_outputs(979) <= a or b;
    layer5_outputs(980) <= a and not b;
    layer5_outputs(981) <= a and not b;
    layer5_outputs(982) <= a;
    layer5_outputs(983) <= not (a and b);
    layer5_outputs(984) <= 1'b0;
    layer5_outputs(985) <= a and b;
    layer5_outputs(986) <= a and b;
    layer5_outputs(987) <= b;
    layer5_outputs(988) <= 1'b1;
    layer5_outputs(989) <= not (a xor b);
    layer5_outputs(990) <= b and not a;
    layer5_outputs(991) <= not (a and b);
    layer5_outputs(992) <= a;
    layer5_outputs(993) <= b;
    layer5_outputs(994) <= not b or a;
    layer5_outputs(995) <= a;
    layer5_outputs(996) <= not (a or b);
    layer5_outputs(997) <= a;
    layer5_outputs(998) <= a xor b;
    layer5_outputs(999) <= not a or b;
    layer5_outputs(1000) <= a or b;
    layer5_outputs(1001) <= not (a or b);
    layer5_outputs(1002) <= a xor b;
    layer5_outputs(1003) <= not b;
    layer5_outputs(1004) <= not a;
    layer5_outputs(1005) <= a and b;
    layer5_outputs(1006) <= a and not b;
    layer5_outputs(1007) <= not b;
    layer5_outputs(1008) <= b and not a;
    layer5_outputs(1009) <= a xor b;
    layer5_outputs(1010) <= a and not b;
    layer5_outputs(1011) <= not (a or b);
    layer5_outputs(1012) <= not a or b;
    layer5_outputs(1013) <= a or b;
    layer5_outputs(1014) <= a or b;
    layer5_outputs(1015) <= not b;
    layer5_outputs(1016) <= not a or b;
    layer5_outputs(1017) <= a xor b;
    layer5_outputs(1018) <= b and not a;
    layer5_outputs(1019) <= a and not b;
    layer5_outputs(1020) <= a and not b;
    layer5_outputs(1021) <= a xor b;
    layer5_outputs(1022) <= not (a and b);
    layer5_outputs(1023) <= b and not a;
    layer5_outputs(1024) <= a and b;
    layer5_outputs(1025) <= 1'b0;
    layer5_outputs(1026) <= b;
    layer5_outputs(1027) <= a and not b;
    layer5_outputs(1028) <= not (a or b);
    layer5_outputs(1029) <= a and b;
    layer5_outputs(1030) <= a or b;
    layer5_outputs(1031) <= not a;
    layer5_outputs(1032) <= a;
    layer5_outputs(1033) <= a xor b;
    layer5_outputs(1034) <= a;
    layer5_outputs(1035) <= b;
    layer5_outputs(1036) <= not b;
    layer5_outputs(1037) <= not a or b;
    layer5_outputs(1038) <= a and not b;
    layer5_outputs(1039) <= b and not a;
    layer5_outputs(1040) <= not b;
    layer5_outputs(1041) <= a and not b;
    layer5_outputs(1042) <= a;
    layer5_outputs(1043) <= a or b;
    layer5_outputs(1044) <= 1'b0;
    layer5_outputs(1045) <= not b or a;
    layer5_outputs(1046) <= not a;
    layer5_outputs(1047) <= not b;
    layer5_outputs(1048) <= a and not b;
    layer5_outputs(1049) <= not a or b;
    layer5_outputs(1050) <= not (a or b);
    layer5_outputs(1051) <= not b;
    layer5_outputs(1052) <= not (a and b);
    layer5_outputs(1053) <= not b;
    layer5_outputs(1054) <= 1'b1;
    layer5_outputs(1055) <= not (a or b);
    layer5_outputs(1056) <= a and not b;
    layer5_outputs(1057) <= a;
    layer5_outputs(1058) <= not a;
    layer5_outputs(1059) <= a xor b;
    layer5_outputs(1060) <= not b or a;
    layer5_outputs(1061) <= a and b;
    layer5_outputs(1062) <= 1'b0;
    layer5_outputs(1063) <= not (a xor b);
    layer5_outputs(1064) <= a;
    layer5_outputs(1065) <= a and not b;
    layer5_outputs(1066) <= a and not b;
    layer5_outputs(1067) <= not b;
    layer5_outputs(1068) <= a and not b;
    layer5_outputs(1069) <= not a;
    layer5_outputs(1070) <= b;
    layer5_outputs(1071) <= not b or a;
    layer5_outputs(1072) <= b;
    layer5_outputs(1073) <= not (a and b);
    layer5_outputs(1074) <= 1'b1;
    layer5_outputs(1075) <= a and not b;
    layer5_outputs(1076) <= 1'b1;
    layer5_outputs(1077) <= a;
    layer5_outputs(1078) <= a and b;
    layer5_outputs(1079) <= not b;
    layer5_outputs(1080) <= not b;
    layer5_outputs(1081) <= b;
    layer5_outputs(1082) <= a and b;
    layer5_outputs(1083) <= b;
    layer5_outputs(1084) <= 1'b0;
    layer5_outputs(1085) <= b;
    layer5_outputs(1086) <= not (a and b);
    layer5_outputs(1087) <= not a;
    layer5_outputs(1088) <= a and b;
    layer5_outputs(1089) <= b;
    layer5_outputs(1090) <= not a or b;
    layer5_outputs(1091) <= not (a and b);
    layer5_outputs(1092) <= not a;
    layer5_outputs(1093) <= a;
    layer5_outputs(1094) <= b;
    layer5_outputs(1095) <= not a;
    layer5_outputs(1096) <= 1'b0;
    layer5_outputs(1097) <= a;
    layer5_outputs(1098) <= 1'b0;
    layer5_outputs(1099) <= not b;
    layer5_outputs(1100) <= not (a and b);
    layer5_outputs(1101) <= b;
    layer5_outputs(1102) <= a;
    layer5_outputs(1103) <= not (a and b);
    layer5_outputs(1104) <= b and not a;
    layer5_outputs(1105) <= a and b;
    layer5_outputs(1106) <= not (a and b);
    layer5_outputs(1107) <= a;
    layer5_outputs(1108) <= not b or a;
    layer5_outputs(1109) <= not b or a;
    layer5_outputs(1110) <= a;
    layer5_outputs(1111) <= b and not a;
    layer5_outputs(1112) <= not a;
    layer5_outputs(1113) <= 1'b1;
    layer5_outputs(1114) <= 1'b1;
    layer5_outputs(1115) <= b and not a;
    layer5_outputs(1116) <= not b;
    layer5_outputs(1117) <= not b;
    layer5_outputs(1118) <= not a;
    layer5_outputs(1119) <= 1'b1;
    layer5_outputs(1120) <= not (a and b);
    layer5_outputs(1121) <= not a;
    layer5_outputs(1122) <= b;
    layer5_outputs(1123) <= not a or b;
    layer5_outputs(1124) <= not a;
    layer5_outputs(1125) <= a or b;
    layer5_outputs(1126) <= a and b;
    layer5_outputs(1127) <= a;
    layer5_outputs(1128) <= a xor b;
    layer5_outputs(1129) <= b and not a;
    layer5_outputs(1130) <= not b or a;
    layer5_outputs(1131) <= a or b;
    layer5_outputs(1132) <= not b;
    layer5_outputs(1133) <= not b;
    layer5_outputs(1134) <= b;
    layer5_outputs(1135) <= not a;
    layer5_outputs(1136) <= not a or b;
    layer5_outputs(1137) <= b;
    layer5_outputs(1138) <= a and not b;
    layer5_outputs(1139) <= a;
    layer5_outputs(1140) <= not a;
    layer5_outputs(1141) <= not a;
    layer5_outputs(1142) <= not a;
    layer5_outputs(1143) <= not (a and b);
    layer5_outputs(1144) <= not b;
    layer5_outputs(1145) <= not a;
    layer5_outputs(1146) <= not (a or b);
    layer5_outputs(1147) <= a;
    layer5_outputs(1148) <= not (a and b);
    layer5_outputs(1149) <= b and not a;
    layer5_outputs(1150) <= not (a or b);
    layer5_outputs(1151) <= not b or a;
    layer5_outputs(1152) <= not a;
    layer5_outputs(1153) <= not b or a;
    layer5_outputs(1154) <= b;
    layer5_outputs(1155) <= b;
    layer5_outputs(1156) <= not a or b;
    layer5_outputs(1157) <= b and not a;
    layer5_outputs(1158) <= not (a or b);
    layer5_outputs(1159) <= a;
    layer5_outputs(1160) <= not (a xor b);
    layer5_outputs(1161) <= b and not a;
    layer5_outputs(1162) <= not b;
    layer5_outputs(1163) <= not (a xor b);
    layer5_outputs(1164) <= not b or a;
    layer5_outputs(1165) <= not b;
    layer5_outputs(1166) <= a or b;
    layer5_outputs(1167) <= not b;
    layer5_outputs(1168) <= a and b;
    layer5_outputs(1169) <= not b;
    layer5_outputs(1170) <= not a;
    layer5_outputs(1171) <= a;
    layer5_outputs(1172) <= b;
    layer5_outputs(1173) <= not a;
    layer5_outputs(1174) <= not (a and b);
    layer5_outputs(1175) <= not a;
    layer5_outputs(1176) <= 1'b0;
    layer5_outputs(1177) <= a;
    layer5_outputs(1178) <= not (a or b);
    layer5_outputs(1179) <= not (a or b);
    layer5_outputs(1180) <= b and not a;
    layer5_outputs(1181) <= not b;
    layer5_outputs(1182) <= not a;
    layer5_outputs(1183) <= not a or b;
    layer5_outputs(1184) <= b and not a;
    layer5_outputs(1185) <= b and not a;
    layer5_outputs(1186) <= b and not a;
    layer5_outputs(1187) <= not (a xor b);
    layer5_outputs(1188) <= b;
    layer5_outputs(1189) <= b and not a;
    layer5_outputs(1190) <= b and not a;
    layer5_outputs(1191) <= not (a xor b);
    layer5_outputs(1192) <= not a;
    layer5_outputs(1193) <= not a;
    layer5_outputs(1194) <= b and not a;
    layer5_outputs(1195) <= a and b;
    layer5_outputs(1196) <= b;
    layer5_outputs(1197) <= 1'b1;
    layer5_outputs(1198) <= not a;
    layer5_outputs(1199) <= not a or b;
    layer5_outputs(1200) <= a and not b;
    layer5_outputs(1201) <= not a;
    layer5_outputs(1202) <= not (a or b);
    layer5_outputs(1203) <= a or b;
    layer5_outputs(1204) <= not a;
    layer5_outputs(1205) <= a;
    layer5_outputs(1206) <= not b;
    layer5_outputs(1207) <= not (a and b);
    layer5_outputs(1208) <= not a;
    layer5_outputs(1209) <= 1'b1;
    layer5_outputs(1210) <= 1'b1;
    layer5_outputs(1211) <= b;
    layer5_outputs(1212) <= a;
    layer5_outputs(1213) <= not (a and b);
    layer5_outputs(1214) <= a;
    layer5_outputs(1215) <= not a;
    layer5_outputs(1216) <= a;
    layer5_outputs(1217) <= a;
    layer5_outputs(1218) <= a or b;
    layer5_outputs(1219) <= b;
    layer5_outputs(1220) <= a or b;
    layer5_outputs(1221) <= not (a xor b);
    layer5_outputs(1222) <= not b or a;
    layer5_outputs(1223) <= a;
    layer5_outputs(1224) <= a and b;
    layer5_outputs(1225) <= 1'b1;
    layer5_outputs(1226) <= not b or a;
    layer5_outputs(1227) <= not (a xor b);
    layer5_outputs(1228) <= 1'b1;
    layer5_outputs(1229) <= a or b;
    layer5_outputs(1230) <= 1'b0;
    layer5_outputs(1231) <= a;
    layer5_outputs(1232) <= not b;
    layer5_outputs(1233) <= b and not a;
    layer5_outputs(1234) <= not b;
    layer5_outputs(1235) <= not a;
    layer5_outputs(1236) <= b;
    layer5_outputs(1237) <= b;
    layer5_outputs(1238) <= a;
    layer5_outputs(1239) <= not b or a;
    layer5_outputs(1240) <= not (a xor b);
    layer5_outputs(1241) <= a;
    layer5_outputs(1242) <= not (a or b);
    layer5_outputs(1243) <= 1'b1;
    layer5_outputs(1244) <= 1'b0;
    layer5_outputs(1245) <= not a or b;
    layer5_outputs(1246) <= not a or b;
    layer5_outputs(1247) <= a and not b;
    layer5_outputs(1248) <= not a;
    layer5_outputs(1249) <= not a or b;
    layer5_outputs(1250) <= a or b;
    layer5_outputs(1251) <= b;
    layer5_outputs(1252) <= b;
    layer5_outputs(1253) <= not (a xor b);
    layer5_outputs(1254) <= not a;
    layer5_outputs(1255) <= not (a and b);
    layer5_outputs(1256) <= not a or b;
    layer5_outputs(1257) <= not a;
    layer5_outputs(1258) <= 1'b0;
    layer5_outputs(1259) <= b;
    layer5_outputs(1260) <= a and not b;
    layer5_outputs(1261) <= not b or a;
    layer5_outputs(1262) <= not a;
    layer5_outputs(1263) <= 1'b1;
    layer5_outputs(1264) <= a and not b;
    layer5_outputs(1265) <= a xor b;
    layer5_outputs(1266) <= not (a and b);
    layer5_outputs(1267) <= not a or b;
    layer5_outputs(1268) <= not (a and b);
    layer5_outputs(1269) <= not (a and b);
    layer5_outputs(1270) <= a or b;
    layer5_outputs(1271) <= b and not a;
    layer5_outputs(1272) <= a or b;
    layer5_outputs(1273) <= 1'b0;
    layer5_outputs(1274) <= a or b;
    layer5_outputs(1275) <= not b or a;
    layer5_outputs(1276) <= 1'b0;
    layer5_outputs(1277) <= a xor b;
    layer5_outputs(1278) <= a and b;
    layer5_outputs(1279) <= b and not a;
    layer5_outputs(1280) <= a xor b;
    layer5_outputs(1281) <= not a or b;
    layer5_outputs(1282) <= not a;
    layer5_outputs(1283) <= not a or b;
    layer5_outputs(1284) <= a and not b;
    layer5_outputs(1285) <= not a;
    layer5_outputs(1286) <= not (a or b);
    layer5_outputs(1287) <= not a or b;
    layer5_outputs(1288) <= not a or b;
    layer5_outputs(1289) <= 1'b0;
    layer5_outputs(1290) <= a or b;
    layer5_outputs(1291) <= a and b;
    layer5_outputs(1292) <= not (a or b);
    layer5_outputs(1293) <= not a or b;
    layer5_outputs(1294) <= a and not b;
    layer5_outputs(1295) <= a xor b;
    layer5_outputs(1296) <= b;
    layer5_outputs(1297) <= not b or a;
    layer5_outputs(1298) <= a xor b;
    layer5_outputs(1299) <= b;
    layer5_outputs(1300) <= not a;
    layer5_outputs(1301) <= a and b;
    layer5_outputs(1302) <= b and not a;
    layer5_outputs(1303) <= not a;
    layer5_outputs(1304) <= b and not a;
    layer5_outputs(1305) <= b;
    layer5_outputs(1306) <= b;
    layer5_outputs(1307) <= a and not b;
    layer5_outputs(1308) <= a;
    layer5_outputs(1309) <= 1'b1;
    layer5_outputs(1310) <= not (a or b);
    layer5_outputs(1311) <= a;
    layer5_outputs(1312) <= b and not a;
    layer5_outputs(1313) <= not a or b;
    layer5_outputs(1314) <= not (a or b);
    layer5_outputs(1315) <= not a or b;
    layer5_outputs(1316) <= not b;
    layer5_outputs(1317) <= b and not a;
    layer5_outputs(1318) <= 1'b1;
    layer5_outputs(1319) <= 1'b1;
    layer5_outputs(1320) <= 1'b0;
    layer5_outputs(1321) <= not a;
    layer5_outputs(1322) <= a or b;
    layer5_outputs(1323) <= not (a and b);
    layer5_outputs(1324) <= not b;
    layer5_outputs(1325) <= not (a or b);
    layer5_outputs(1326) <= 1'b1;
    layer5_outputs(1327) <= b;
    layer5_outputs(1328) <= not b or a;
    layer5_outputs(1329) <= not (a and b);
    layer5_outputs(1330) <= 1'b1;
    layer5_outputs(1331) <= b;
    layer5_outputs(1332) <= b;
    layer5_outputs(1333) <= not (a and b);
    layer5_outputs(1334) <= not b;
    layer5_outputs(1335) <= not a;
    layer5_outputs(1336) <= not a;
    layer5_outputs(1337) <= a and b;
    layer5_outputs(1338) <= not a or b;
    layer5_outputs(1339) <= b;
    layer5_outputs(1340) <= not (a and b);
    layer5_outputs(1341) <= not a;
    layer5_outputs(1342) <= not a;
    layer5_outputs(1343) <= not a;
    layer5_outputs(1344) <= not a or b;
    layer5_outputs(1345) <= a or b;
    layer5_outputs(1346) <= not b;
    layer5_outputs(1347) <= 1'b0;
    layer5_outputs(1348) <= a;
    layer5_outputs(1349) <= a and b;
    layer5_outputs(1350) <= not a;
    layer5_outputs(1351) <= a and not b;
    layer5_outputs(1352) <= not (a or b);
    layer5_outputs(1353) <= not (a and b);
    layer5_outputs(1354) <= not b;
    layer5_outputs(1355) <= not a;
    layer5_outputs(1356) <= not b or a;
    layer5_outputs(1357) <= b;
    layer5_outputs(1358) <= not a or b;
    layer5_outputs(1359) <= not (a or b);
    layer5_outputs(1360) <= not (a and b);
    layer5_outputs(1361) <= not b or a;
    layer5_outputs(1362) <= a;
    layer5_outputs(1363) <= a;
    layer5_outputs(1364) <= b;
    layer5_outputs(1365) <= not a or b;
    layer5_outputs(1366) <= not b;
    layer5_outputs(1367) <= a and b;
    layer5_outputs(1368) <= a;
    layer5_outputs(1369) <= a and not b;
    layer5_outputs(1370) <= a or b;
    layer5_outputs(1371) <= b and not a;
    layer5_outputs(1372) <= a and not b;
    layer5_outputs(1373) <= b and not a;
    layer5_outputs(1374) <= not a;
    layer5_outputs(1375) <= b and not a;
    layer5_outputs(1376) <= not b;
    layer5_outputs(1377) <= not b or a;
    layer5_outputs(1378) <= not a or b;
    layer5_outputs(1379) <= 1'b0;
    layer5_outputs(1380) <= a and not b;
    layer5_outputs(1381) <= a and not b;
    layer5_outputs(1382) <= a;
    layer5_outputs(1383) <= not a;
    layer5_outputs(1384) <= a and not b;
    layer5_outputs(1385) <= not b;
    layer5_outputs(1386) <= b and not a;
    layer5_outputs(1387) <= 1'b1;
    layer5_outputs(1388) <= not a;
    layer5_outputs(1389) <= a and b;
    layer5_outputs(1390) <= a or b;
    layer5_outputs(1391) <= b;
    layer5_outputs(1392) <= not (a and b);
    layer5_outputs(1393) <= not a;
    layer5_outputs(1394) <= a and b;
    layer5_outputs(1395) <= not b or a;
    layer5_outputs(1396) <= a xor b;
    layer5_outputs(1397) <= not b;
    layer5_outputs(1398) <= not (a or b);
    layer5_outputs(1399) <= a;
    layer5_outputs(1400) <= not a or b;
    layer5_outputs(1401) <= not (a xor b);
    layer5_outputs(1402) <= 1'b1;
    layer5_outputs(1403) <= b;
    layer5_outputs(1404) <= not a;
    layer5_outputs(1405) <= not (a xor b);
    layer5_outputs(1406) <= not (a xor b);
    layer5_outputs(1407) <= not a or b;
    layer5_outputs(1408) <= a xor b;
    layer5_outputs(1409) <= not b;
    layer5_outputs(1410) <= 1'b1;
    layer5_outputs(1411) <= not a;
    layer5_outputs(1412) <= not b or a;
    layer5_outputs(1413) <= not b or a;
    layer5_outputs(1414) <= not a;
    layer5_outputs(1415) <= b;
    layer5_outputs(1416) <= b;
    layer5_outputs(1417) <= not b or a;
    layer5_outputs(1418) <= not a or b;
    layer5_outputs(1419) <= a or b;
    layer5_outputs(1420) <= not a or b;
    layer5_outputs(1421) <= a and b;
    layer5_outputs(1422) <= b;
    layer5_outputs(1423) <= not b;
    layer5_outputs(1424) <= a;
    layer5_outputs(1425) <= not (a or b);
    layer5_outputs(1426) <= a or b;
    layer5_outputs(1427) <= not a or b;
    layer5_outputs(1428) <= 1'b1;
    layer5_outputs(1429) <= b;
    layer5_outputs(1430) <= a;
    layer5_outputs(1431) <= 1'b0;
    layer5_outputs(1432) <= not b;
    layer5_outputs(1433) <= a and not b;
    layer5_outputs(1434) <= not (a xor b);
    layer5_outputs(1435) <= a and not b;
    layer5_outputs(1436) <= not b;
    layer5_outputs(1437) <= a or b;
    layer5_outputs(1438) <= not a or b;
    layer5_outputs(1439) <= a or b;
    layer5_outputs(1440) <= b;
    layer5_outputs(1441) <= not b;
    layer5_outputs(1442) <= not b;
    layer5_outputs(1443) <= b and not a;
    layer5_outputs(1444) <= a xor b;
    layer5_outputs(1445) <= not b;
    layer5_outputs(1446) <= 1'b1;
    layer5_outputs(1447) <= not a;
    layer5_outputs(1448) <= not a or b;
    layer5_outputs(1449) <= a and b;
    layer5_outputs(1450) <= b;
    layer5_outputs(1451) <= not b or a;
    layer5_outputs(1452) <= a;
    layer5_outputs(1453) <= a;
    layer5_outputs(1454) <= not a;
    layer5_outputs(1455) <= not b or a;
    layer5_outputs(1456) <= not b or a;
    layer5_outputs(1457) <= 1'b0;
    layer5_outputs(1458) <= not a or b;
    layer5_outputs(1459) <= 1'b1;
    layer5_outputs(1460) <= not (a xor b);
    layer5_outputs(1461) <= not b;
    layer5_outputs(1462) <= b and not a;
    layer5_outputs(1463) <= not b;
    layer5_outputs(1464) <= b;
    layer5_outputs(1465) <= a xor b;
    layer5_outputs(1466) <= not a;
    layer5_outputs(1467) <= b;
    layer5_outputs(1468) <= not (a or b);
    layer5_outputs(1469) <= 1'b1;
    layer5_outputs(1470) <= not a;
    layer5_outputs(1471) <= not (a or b);
    layer5_outputs(1472) <= not b;
    layer5_outputs(1473) <= not (a and b);
    layer5_outputs(1474) <= not b;
    layer5_outputs(1475) <= not (a and b);
    layer5_outputs(1476) <= a and b;
    layer5_outputs(1477) <= not a;
    layer5_outputs(1478) <= not b;
    layer5_outputs(1479) <= not a or b;
    layer5_outputs(1480) <= not b or a;
    layer5_outputs(1481) <= not b;
    layer5_outputs(1482) <= a;
    layer5_outputs(1483) <= not a;
    layer5_outputs(1484) <= 1'b1;
    layer5_outputs(1485) <= not (a xor b);
    layer5_outputs(1486) <= a or b;
    layer5_outputs(1487) <= not b or a;
    layer5_outputs(1488) <= b;
    layer5_outputs(1489) <= 1'b0;
    layer5_outputs(1490) <= not (a and b);
    layer5_outputs(1491) <= not a;
    layer5_outputs(1492) <= not a;
    layer5_outputs(1493) <= not (a or b);
    layer5_outputs(1494) <= 1'b1;
    layer5_outputs(1495) <= a xor b;
    layer5_outputs(1496) <= a;
    layer5_outputs(1497) <= not (a or b);
    layer5_outputs(1498) <= a;
    layer5_outputs(1499) <= 1'b0;
    layer5_outputs(1500) <= not b or a;
    layer5_outputs(1501) <= a;
    layer5_outputs(1502) <= a or b;
    layer5_outputs(1503) <= b;
    layer5_outputs(1504) <= not (a and b);
    layer5_outputs(1505) <= not (a or b);
    layer5_outputs(1506) <= not b or a;
    layer5_outputs(1507) <= a and b;
    layer5_outputs(1508) <= not b;
    layer5_outputs(1509) <= a;
    layer5_outputs(1510) <= 1'b0;
    layer5_outputs(1511) <= b;
    layer5_outputs(1512) <= not (a xor b);
    layer5_outputs(1513) <= not (a or b);
    layer5_outputs(1514) <= a and not b;
    layer5_outputs(1515) <= a and not b;
    layer5_outputs(1516) <= a;
    layer5_outputs(1517) <= a or b;
    layer5_outputs(1518) <= 1'b0;
    layer5_outputs(1519) <= b;
    layer5_outputs(1520) <= b and not a;
    layer5_outputs(1521) <= b and not a;
    layer5_outputs(1522) <= not a;
    layer5_outputs(1523) <= a;
    layer5_outputs(1524) <= b;
    layer5_outputs(1525) <= a xor b;
    layer5_outputs(1526) <= a or b;
    layer5_outputs(1527) <= not b or a;
    layer5_outputs(1528) <= b and not a;
    layer5_outputs(1529) <= a;
    layer5_outputs(1530) <= not a or b;
    layer5_outputs(1531) <= b;
    layer5_outputs(1532) <= not (a and b);
    layer5_outputs(1533) <= a;
    layer5_outputs(1534) <= a and b;
    layer5_outputs(1535) <= a and b;
    layer5_outputs(1536) <= a;
    layer5_outputs(1537) <= 1'b0;
    layer5_outputs(1538) <= not a;
    layer5_outputs(1539) <= not (a xor b);
    layer5_outputs(1540) <= 1'b1;
    layer5_outputs(1541) <= not (a or b);
    layer5_outputs(1542) <= b;
    layer5_outputs(1543) <= b and not a;
    layer5_outputs(1544) <= b;
    layer5_outputs(1545) <= 1'b1;
    layer5_outputs(1546) <= not (a xor b);
    layer5_outputs(1547) <= not b;
    layer5_outputs(1548) <= b and not a;
    layer5_outputs(1549) <= not a or b;
    layer5_outputs(1550) <= a and not b;
    layer5_outputs(1551) <= b;
    layer5_outputs(1552) <= not b;
    layer5_outputs(1553) <= not b;
    layer5_outputs(1554) <= not (a or b);
    layer5_outputs(1555) <= a or b;
    layer5_outputs(1556) <= not b or a;
    layer5_outputs(1557) <= b and not a;
    layer5_outputs(1558) <= not a;
    layer5_outputs(1559) <= not a or b;
    layer5_outputs(1560) <= 1'b1;
    layer5_outputs(1561) <= not a or b;
    layer5_outputs(1562) <= not (a xor b);
    layer5_outputs(1563) <= 1'b1;
    layer5_outputs(1564) <= not b;
    layer5_outputs(1565) <= b and not a;
    layer5_outputs(1566) <= not a;
    layer5_outputs(1567) <= a;
    layer5_outputs(1568) <= not b or a;
    layer5_outputs(1569) <= a or b;
    layer5_outputs(1570) <= not a;
    layer5_outputs(1571) <= a;
    layer5_outputs(1572) <= b;
    layer5_outputs(1573) <= a and b;
    layer5_outputs(1574) <= a;
    layer5_outputs(1575) <= a;
    layer5_outputs(1576) <= not (a or b);
    layer5_outputs(1577) <= b;
    layer5_outputs(1578) <= a and b;
    layer5_outputs(1579) <= b;
    layer5_outputs(1580) <= not b;
    layer5_outputs(1581) <= 1'b1;
    layer5_outputs(1582) <= not a;
    layer5_outputs(1583) <= not b;
    layer5_outputs(1584) <= not b or a;
    layer5_outputs(1585) <= a or b;
    layer5_outputs(1586) <= not a;
    layer5_outputs(1587) <= not (a and b);
    layer5_outputs(1588) <= b;
    layer5_outputs(1589) <= not (a and b);
    layer5_outputs(1590) <= a and b;
    layer5_outputs(1591) <= not b or a;
    layer5_outputs(1592) <= b;
    layer5_outputs(1593) <= a and not b;
    layer5_outputs(1594) <= not a;
    layer5_outputs(1595) <= not b or a;
    layer5_outputs(1596) <= a or b;
    layer5_outputs(1597) <= a xor b;
    layer5_outputs(1598) <= a;
    layer5_outputs(1599) <= not b or a;
    layer5_outputs(1600) <= not a;
    layer5_outputs(1601) <= not a;
    layer5_outputs(1602) <= b;
    layer5_outputs(1603) <= not a;
    layer5_outputs(1604) <= not b or a;
    layer5_outputs(1605) <= a and not b;
    layer5_outputs(1606) <= b;
    layer5_outputs(1607) <= 1'b0;
    layer5_outputs(1608) <= not a;
    layer5_outputs(1609) <= not a;
    layer5_outputs(1610) <= not b;
    layer5_outputs(1611) <= a and not b;
    layer5_outputs(1612) <= 1'b1;
    layer5_outputs(1613) <= not b;
    layer5_outputs(1614) <= not a or b;
    layer5_outputs(1615) <= not b;
    layer5_outputs(1616) <= not (a and b);
    layer5_outputs(1617) <= not a;
    layer5_outputs(1618) <= not a;
    layer5_outputs(1619) <= b;
    layer5_outputs(1620) <= 1'b0;
    layer5_outputs(1621) <= a or b;
    layer5_outputs(1622) <= b;
    layer5_outputs(1623) <= 1'b1;
    layer5_outputs(1624) <= b;
    layer5_outputs(1625) <= a or b;
    layer5_outputs(1626) <= a xor b;
    layer5_outputs(1627) <= not (a xor b);
    layer5_outputs(1628) <= not b or a;
    layer5_outputs(1629) <= not (a or b);
    layer5_outputs(1630) <= a and not b;
    layer5_outputs(1631) <= not (a xor b);
    layer5_outputs(1632) <= not (a or b);
    layer5_outputs(1633) <= not a;
    layer5_outputs(1634) <= a;
    layer5_outputs(1635) <= a xor b;
    layer5_outputs(1636) <= b;
    layer5_outputs(1637) <= not (a or b);
    layer5_outputs(1638) <= not b or a;
    layer5_outputs(1639) <= a and not b;
    layer5_outputs(1640) <= a xor b;
    layer5_outputs(1641) <= b;
    layer5_outputs(1642) <= a or b;
    layer5_outputs(1643) <= a and b;
    layer5_outputs(1644) <= not (a or b);
    layer5_outputs(1645) <= not b;
    layer5_outputs(1646) <= not (a and b);
    layer5_outputs(1647) <= 1'b0;
    layer5_outputs(1648) <= a;
    layer5_outputs(1649) <= not (a xor b);
    layer5_outputs(1650) <= a or b;
    layer5_outputs(1651) <= a;
    layer5_outputs(1652) <= not a or b;
    layer5_outputs(1653) <= not (a and b);
    layer5_outputs(1654) <= not b;
    layer5_outputs(1655) <= not b;
    layer5_outputs(1656) <= a and b;
    layer5_outputs(1657) <= not (a and b);
    layer5_outputs(1658) <= a and b;
    layer5_outputs(1659) <= not a;
    layer5_outputs(1660) <= a;
    layer5_outputs(1661) <= not (a or b);
    layer5_outputs(1662) <= a;
    layer5_outputs(1663) <= not a;
    layer5_outputs(1664) <= a and b;
    layer5_outputs(1665) <= not (a or b);
    layer5_outputs(1666) <= not b or a;
    layer5_outputs(1667) <= not b;
    layer5_outputs(1668) <= not b;
    layer5_outputs(1669) <= 1'b0;
    layer5_outputs(1670) <= b;
    layer5_outputs(1671) <= not (a and b);
    layer5_outputs(1672) <= b and not a;
    layer5_outputs(1673) <= 1'b1;
    layer5_outputs(1674) <= not a;
    layer5_outputs(1675) <= a and b;
    layer5_outputs(1676) <= not (a xor b);
    layer5_outputs(1677) <= not (a and b);
    layer5_outputs(1678) <= not a;
    layer5_outputs(1679) <= a or b;
    layer5_outputs(1680) <= a or b;
    layer5_outputs(1681) <= b;
    layer5_outputs(1682) <= not a;
    layer5_outputs(1683) <= a or b;
    layer5_outputs(1684) <= not (a or b);
    layer5_outputs(1685) <= 1'b0;
    layer5_outputs(1686) <= not a;
    layer5_outputs(1687) <= not a or b;
    layer5_outputs(1688) <= a and not b;
    layer5_outputs(1689) <= b and not a;
    layer5_outputs(1690) <= not (a and b);
    layer5_outputs(1691) <= not b or a;
    layer5_outputs(1692) <= not (a and b);
    layer5_outputs(1693) <= a and b;
    layer5_outputs(1694) <= not b or a;
    layer5_outputs(1695) <= a xor b;
    layer5_outputs(1696) <= not b;
    layer5_outputs(1697) <= a or b;
    layer5_outputs(1698) <= not a;
    layer5_outputs(1699) <= not (a or b);
    layer5_outputs(1700) <= not b;
    layer5_outputs(1701) <= b;
    layer5_outputs(1702) <= not b or a;
    layer5_outputs(1703) <= a or b;
    layer5_outputs(1704) <= not (a or b);
    layer5_outputs(1705) <= not (a or b);
    layer5_outputs(1706) <= not a;
    layer5_outputs(1707) <= not b;
    layer5_outputs(1708) <= not b;
    layer5_outputs(1709) <= not a;
    layer5_outputs(1710) <= a;
    layer5_outputs(1711) <= not a or b;
    layer5_outputs(1712) <= not (a and b);
    layer5_outputs(1713) <= not a;
    layer5_outputs(1714) <= a and not b;
    layer5_outputs(1715) <= 1'b0;
    layer5_outputs(1716) <= not b;
    layer5_outputs(1717) <= a;
    layer5_outputs(1718) <= not a;
    layer5_outputs(1719) <= a;
    layer5_outputs(1720) <= not b or a;
    layer5_outputs(1721) <= not b;
    layer5_outputs(1722) <= not (a and b);
    layer5_outputs(1723) <= b;
    layer5_outputs(1724) <= not a;
    layer5_outputs(1725) <= not b;
    layer5_outputs(1726) <= not b;
    layer5_outputs(1727) <= not b or a;
    layer5_outputs(1728) <= not (a and b);
    layer5_outputs(1729) <= b;
    layer5_outputs(1730) <= b;
    layer5_outputs(1731) <= a and b;
    layer5_outputs(1732) <= a or b;
    layer5_outputs(1733) <= not a;
    layer5_outputs(1734) <= not a or b;
    layer5_outputs(1735) <= b;
    layer5_outputs(1736) <= a and not b;
    layer5_outputs(1737) <= b;
    layer5_outputs(1738) <= a and b;
    layer5_outputs(1739) <= b;
    layer5_outputs(1740) <= not a;
    layer5_outputs(1741) <= a xor b;
    layer5_outputs(1742) <= not (a xor b);
    layer5_outputs(1743) <= a and not b;
    layer5_outputs(1744) <= not a;
    layer5_outputs(1745) <= 1'b0;
    layer5_outputs(1746) <= not b;
    layer5_outputs(1747) <= not b or a;
    layer5_outputs(1748) <= a or b;
    layer5_outputs(1749) <= a;
    layer5_outputs(1750) <= a or b;
    layer5_outputs(1751) <= not a;
    layer5_outputs(1752) <= not a or b;
    layer5_outputs(1753) <= b and not a;
    layer5_outputs(1754) <= not b or a;
    layer5_outputs(1755) <= 1'b0;
    layer5_outputs(1756) <= not (a or b);
    layer5_outputs(1757) <= b;
    layer5_outputs(1758) <= not b;
    layer5_outputs(1759) <= not a or b;
    layer5_outputs(1760) <= a and b;
    layer5_outputs(1761) <= not a;
    layer5_outputs(1762) <= not a;
    layer5_outputs(1763) <= not (a xor b);
    layer5_outputs(1764) <= not a or b;
    layer5_outputs(1765) <= not b or a;
    layer5_outputs(1766) <= not b or a;
    layer5_outputs(1767) <= not (a xor b);
    layer5_outputs(1768) <= 1'b1;
    layer5_outputs(1769) <= not a;
    layer5_outputs(1770) <= 1'b1;
    layer5_outputs(1771) <= a xor b;
    layer5_outputs(1772) <= a and not b;
    layer5_outputs(1773) <= b and not a;
    layer5_outputs(1774) <= 1'b0;
    layer5_outputs(1775) <= not b;
    layer5_outputs(1776) <= a;
    layer5_outputs(1777) <= not (a xor b);
    layer5_outputs(1778) <= a;
    layer5_outputs(1779) <= a xor b;
    layer5_outputs(1780) <= a and b;
    layer5_outputs(1781) <= b;
    layer5_outputs(1782) <= a or b;
    layer5_outputs(1783) <= b;
    layer5_outputs(1784) <= not a;
    layer5_outputs(1785) <= a and not b;
    layer5_outputs(1786) <= 1'b1;
    layer5_outputs(1787) <= 1'b1;
    layer5_outputs(1788) <= b;
    layer5_outputs(1789) <= not (a xor b);
    layer5_outputs(1790) <= not (a and b);
    layer5_outputs(1791) <= b and not a;
    layer5_outputs(1792) <= a;
    layer5_outputs(1793) <= a and b;
    layer5_outputs(1794) <= not (a or b);
    layer5_outputs(1795) <= not b or a;
    layer5_outputs(1796) <= not b;
    layer5_outputs(1797) <= a;
    layer5_outputs(1798) <= a;
    layer5_outputs(1799) <= a or b;
    layer5_outputs(1800) <= b;
    layer5_outputs(1801) <= a and not b;
    layer5_outputs(1802) <= not b;
    layer5_outputs(1803) <= not a;
    layer5_outputs(1804) <= 1'b1;
    layer5_outputs(1805) <= a or b;
    layer5_outputs(1806) <= a;
    layer5_outputs(1807) <= b;
    layer5_outputs(1808) <= b;
    layer5_outputs(1809) <= a;
    layer5_outputs(1810) <= not a or b;
    layer5_outputs(1811) <= a and b;
    layer5_outputs(1812) <= not (a and b);
    layer5_outputs(1813) <= 1'b0;
    layer5_outputs(1814) <= a xor b;
    layer5_outputs(1815) <= a;
    layer5_outputs(1816) <= not (a or b);
    layer5_outputs(1817) <= a or b;
    layer5_outputs(1818) <= b;
    layer5_outputs(1819) <= not b;
    layer5_outputs(1820) <= a;
    layer5_outputs(1821) <= not b or a;
    layer5_outputs(1822) <= not a;
    layer5_outputs(1823) <= not b or a;
    layer5_outputs(1824) <= a or b;
    layer5_outputs(1825) <= a;
    layer5_outputs(1826) <= not a;
    layer5_outputs(1827) <= a and b;
    layer5_outputs(1828) <= not b;
    layer5_outputs(1829) <= 1'b1;
    layer5_outputs(1830) <= a;
    layer5_outputs(1831) <= a and b;
    layer5_outputs(1832) <= not b;
    layer5_outputs(1833) <= b and not a;
    layer5_outputs(1834) <= a or b;
    layer5_outputs(1835) <= not (a xor b);
    layer5_outputs(1836) <= not (a and b);
    layer5_outputs(1837) <= not b;
    layer5_outputs(1838) <= not b;
    layer5_outputs(1839) <= not (a and b);
    layer5_outputs(1840) <= b;
    layer5_outputs(1841) <= 1'b0;
    layer5_outputs(1842) <= not a;
    layer5_outputs(1843) <= not (a and b);
    layer5_outputs(1844) <= not (a xor b);
    layer5_outputs(1845) <= a or b;
    layer5_outputs(1846) <= not (a or b);
    layer5_outputs(1847) <= b and not a;
    layer5_outputs(1848) <= a or b;
    layer5_outputs(1849) <= a and not b;
    layer5_outputs(1850) <= not b;
    layer5_outputs(1851) <= a;
    layer5_outputs(1852) <= not (a and b);
    layer5_outputs(1853) <= a and not b;
    layer5_outputs(1854) <= not (a and b);
    layer5_outputs(1855) <= b;
    layer5_outputs(1856) <= 1'b0;
    layer5_outputs(1857) <= a and b;
    layer5_outputs(1858) <= not a;
    layer5_outputs(1859) <= a and b;
    layer5_outputs(1860) <= a and b;
    layer5_outputs(1861) <= a xor b;
    layer5_outputs(1862) <= not a or b;
    layer5_outputs(1863) <= not a or b;
    layer5_outputs(1864) <= not b;
    layer5_outputs(1865) <= a;
    layer5_outputs(1866) <= not (a xor b);
    layer5_outputs(1867) <= not a;
    layer5_outputs(1868) <= a;
    layer5_outputs(1869) <= b;
    layer5_outputs(1870) <= not (a xor b);
    layer5_outputs(1871) <= a;
    layer5_outputs(1872) <= a and not b;
    layer5_outputs(1873) <= b;
    layer5_outputs(1874) <= not (a xor b);
    layer5_outputs(1875) <= a and not b;
    layer5_outputs(1876) <= not a;
    layer5_outputs(1877) <= not b or a;
    layer5_outputs(1878) <= b;
    layer5_outputs(1879) <= b and not a;
    layer5_outputs(1880) <= not a;
    layer5_outputs(1881) <= a xor b;
    layer5_outputs(1882) <= not b;
    layer5_outputs(1883) <= not a or b;
    layer5_outputs(1884) <= not b;
    layer5_outputs(1885) <= a or b;
    layer5_outputs(1886) <= not b or a;
    layer5_outputs(1887) <= a;
    layer5_outputs(1888) <= 1'b0;
    layer5_outputs(1889) <= not (a xor b);
    layer5_outputs(1890) <= a and b;
    layer5_outputs(1891) <= a or b;
    layer5_outputs(1892) <= b and not a;
    layer5_outputs(1893) <= b;
    layer5_outputs(1894) <= a;
    layer5_outputs(1895) <= not b;
    layer5_outputs(1896) <= 1'b1;
    layer5_outputs(1897) <= a or b;
    layer5_outputs(1898) <= not a;
    layer5_outputs(1899) <= not a or b;
    layer5_outputs(1900) <= 1'b1;
    layer5_outputs(1901) <= not b;
    layer5_outputs(1902) <= b;
    layer5_outputs(1903) <= not b;
    layer5_outputs(1904) <= b and not a;
    layer5_outputs(1905) <= b;
    layer5_outputs(1906) <= a;
    layer5_outputs(1907) <= not a;
    layer5_outputs(1908) <= not b;
    layer5_outputs(1909) <= b;
    layer5_outputs(1910) <= b;
    layer5_outputs(1911) <= not b;
    layer5_outputs(1912) <= a;
    layer5_outputs(1913) <= 1'b0;
    layer5_outputs(1914) <= not b or a;
    layer5_outputs(1915) <= 1'b1;
    layer5_outputs(1916) <= b;
    layer5_outputs(1917) <= a or b;
    layer5_outputs(1918) <= b and not a;
    layer5_outputs(1919) <= not b;
    layer5_outputs(1920) <= 1'b1;
    layer5_outputs(1921) <= b;
    layer5_outputs(1922) <= not a;
    layer5_outputs(1923) <= not (a and b);
    layer5_outputs(1924) <= b and not a;
    layer5_outputs(1925) <= a xor b;
    layer5_outputs(1926) <= a or b;
    layer5_outputs(1927) <= 1'b1;
    layer5_outputs(1928) <= a and b;
    layer5_outputs(1929) <= not a or b;
    layer5_outputs(1930) <= not b;
    layer5_outputs(1931) <= 1'b1;
    layer5_outputs(1932) <= not (a or b);
    layer5_outputs(1933) <= a and b;
    layer5_outputs(1934) <= 1'b0;
    layer5_outputs(1935) <= a and not b;
    layer5_outputs(1936) <= a or b;
    layer5_outputs(1937) <= not (a or b);
    layer5_outputs(1938) <= not (a and b);
    layer5_outputs(1939) <= not b;
    layer5_outputs(1940) <= not a or b;
    layer5_outputs(1941) <= not b;
    layer5_outputs(1942) <= b;
    layer5_outputs(1943) <= not a;
    layer5_outputs(1944) <= not a or b;
    layer5_outputs(1945) <= a and not b;
    layer5_outputs(1946) <= not a;
    layer5_outputs(1947) <= b and not a;
    layer5_outputs(1948) <= not b or a;
    layer5_outputs(1949) <= a and b;
    layer5_outputs(1950) <= a or b;
    layer5_outputs(1951) <= not (a and b);
    layer5_outputs(1952) <= a and not b;
    layer5_outputs(1953) <= b;
    layer5_outputs(1954) <= not a;
    layer5_outputs(1955) <= not a;
    layer5_outputs(1956) <= a and not b;
    layer5_outputs(1957) <= not a or b;
    layer5_outputs(1958) <= b and not a;
    layer5_outputs(1959) <= not a or b;
    layer5_outputs(1960) <= not (a and b);
    layer5_outputs(1961) <= a and not b;
    layer5_outputs(1962) <= a and not b;
    layer5_outputs(1963) <= b;
    layer5_outputs(1964) <= a or b;
    layer5_outputs(1965) <= not a or b;
    layer5_outputs(1966) <= not (a and b);
    layer5_outputs(1967) <= not (a or b);
    layer5_outputs(1968) <= 1'b0;
    layer5_outputs(1969) <= a;
    layer5_outputs(1970) <= not a;
    layer5_outputs(1971) <= a;
    layer5_outputs(1972) <= b and not a;
    layer5_outputs(1973) <= not a;
    layer5_outputs(1974) <= a and not b;
    layer5_outputs(1975) <= not a;
    layer5_outputs(1976) <= not b;
    layer5_outputs(1977) <= a;
    layer5_outputs(1978) <= a or b;
    layer5_outputs(1979) <= a and b;
    layer5_outputs(1980) <= not a;
    layer5_outputs(1981) <= not (a and b);
    layer5_outputs(1982) <= not a;
    layer5_outputs(1983) <= a or b;
    layer5_outputs(1984) <= b;
    layer5_outputs(1985) <= not b or a;
    layer5_outputs(1986) <= not (a and b);
    layer5_outputs(1987) <= 1'b0;
    layer5_outputs(1988) <= 1'b1;
    layer5_outputs(1989) <= not b or a;
    layer5_outputs(1990) <= b;
    layer5_outputs(1991) <= not (a or b);
    layer5_outputs(1992) <= not a or b;
    layer5_outputs(1993) <= not (a or b);
    layer5_outputs(1994) <= not b or a;
    layer5_outputs(1995) <= b;
    layer5_outputs(1996) <= a or b;
    layer5_outputs(1997) <= not a or b;
    layer5_outputs(1998) <= not b;
    layer5_outputs(1999) <= 1'b0;
    layer5_outputs(2000) <= not b;
    layer5_outputs(2001) <= not b or a;
    layer5_outputs(2002) <= not a;
    layer5_outputs(2003) <= not (a and b);
    layer5_outputs(2004) <= a or b;
    layer5_outputs(2005) <= not (a xor b);
    layer5_outputs(2006) <= not (a and b);
    layer5_outputs(2007) <= a or b;
    layer5_outputs(2008) <= not (a or b);
    layer5_outputs(2009) <= b and not a;
    layer5_outputs(2010) <= a and b;
    layer5_outputs(2011) <= b;
    layer5_outputs(2012) <= a and b;
    layer5_outputs(2013) <= a or b;
    layer5_outputs(2014) <= a or b;
    layer5_outputs(2015) <= b;
    layer5_outputs(2016) <= a and b;
    layer5_outputs(2017) <= a or b;
    layer5_outputs(2018) <= b;
    layer5_outputs(2019) <= b;
    layer5_outputs(2020) <= not b;
    layer5_outputs(2021) <= a and not b;
    layer5_outputs(2022) <= not (a xor b);
    layer5_outputs(2023) <= b;
    layer5_outputs(2024) <= not b or a;
    layer5_outputs(2025) <= not b;
    layer5_outputs(2026) <= not a or b;
    layer5_outputs(2027) <= b;
    layer5_outputs(2028) <= not a or b;
    layer5_outputs(2029) <= not (a or b);
    layer5_outputs(2030) <= b and not a;
    layer5_outputs(2031) <= not b;
    layer5_outputs(2032) <= b;
    layer5_outputs(2033) <= not (a and b);
    layer5_outputs(2034) <= b;
    layer5_outputs(2035) <= not (a and b);
    layer5_outputs(2036) <= not a;
    layer5_outputs(2037) <= a;
    layer5_outputs(2038) <= not a;
    layer5_outputs(2039) <= a;
    layer5_outputs(2040) <= not (a and b);
    layer5_outputs(2041) <= not b;
    layer5_outputs(2042) <= not (a and b);
    layer5_outputs(2043) <= b;
    layer5_outputs(2044) <= not a;
    layer5_outputs(2045) <= a;
    layer5_outputs(2046) <= not b;
    layer5_outputs(2047) <= not b;
    layer5_outputs(2048) <= not a;
    layer5_outputs(2049) <= not b;
    layer5_outputs(2050) <= not b;
    layer5_outputs(2051) <= b and not a;
    layer5_outputs(2052) <= not b;
    layer5_outputs(2053) <= not b;
    layer5_outputs(2054) <= not b;
    layer5_outputs(2055) <= b;
    layer5_outputs(2056) <= a and not b;
    layer5_outputs(2057) <= not a;
    layer5_outputs(2058) <= not b;
    layer5_outputs(2059) <= not a;
    layer5_outputs(2060) <= a and b;
    layer5_outputs(2061) <= a;
    layer5_outputs(2062) <= not a;
    layer5_outputs(2063) <= not (a and b);
    layer5_outputs(2064) <= 1'b0;
    layer5_outputs(2065) <= a xor b;
    layer5_outputs(2066) <= not b;
    layer5_outputs(2067) <= a and not b;
    layer5_outputs(2068) <= b and not a;
    layer5_outputs(2069) <= 1'b0;
    layer5_outputs(2070) <= a or b;
    layer5_outputs(2071) <= not b or a;
    layer5_outputs(2072) <= b;
    layer5_outputs(2073) <= a or b;
    layer5_outputs(2074) <= b;
    layer5_outputs(2075) <= not a;
    layer5_outputs(2076) <= not (a and b);
    layer5_outputs(2077) <= 1'b0;
    layer5_outputs(2078) <= not a;
    layer5_outputs(2079) <= 1'b0;
    layer5_outputs(2080) <= b;
    layer5_outputs(2081) <= not (a xor b);
    layer5_outputs(2082) <= b;
    layer5_outputs(2083) <= a;
    layer5_outputs(2084) <= not b;
    layer5_outputs(2085) <= not b or a;
    layer5_outputs(2086) <= not a or b;
    layer5_outputs(2087) <= not b;
    layer5_outputs(2088) <= a xor b;
    layer5_outputs(2089) <= b;
    layer5_outputs(2090) <= a xor b;
    layer5_outputs(2091) <= not b;
    layer5_outputs(2092) <= a and not b;
    layer5_outputs(2093) <= not b or a;
    layer5_outputs(2094) <= b and not a;
    layer5_outputs(2095) <= not a;
    layer5_outputs(2096) <= 1'b0;
    layer5_outputs(2097) <= a and not b;
    layer5_outputs(2098) <= a and not b;
    layer5_outputs(2099) <= 1'b1;
    layer5_outputs(2100) <= not (a and b);
    layer5_outputs(2101) <= not (a xor b);
    layer5_outputs(2102) <= not b or a;
    layer5_outputs(2103) <= a;
    layer5_outputs(2104) <= not (a and b);
    layer5_outputs(2105) <= not b or a;
    layer5_outputs(2106) <= not (a xor b);
    layer5_outputs(2107) <= not a;
    layer5_outputs(2108) <= a and not b;
    layer5_outputs(2109) <= not (a or b);
    layer5_outputs(2110) <= a and not b;
    layer5_outputs(2111) <= a or b;
    layer5_outputs(2112) <= a or b;
    layer5_outputs(2113) <= not a or b;
    layer5_outputs(2114) <= not b or a;
    layer5_outputs(2115) <= a or b;
    layer5_outputs(2116) <= not (a and b);
    layer5_outputs(2117) <= a xor b;
    layer5_outputs(2118) <= not (a xor b);
    layer5_outputs(2119) <= a;
    layer5_outputs(2120) <= b and not a;
    layer5_outputs(2121) <= not b;
    layer5_outputs(2122) <= not b;
    layer5_outputs(2123) <= not b or a;
    layer5_outputs(2124) <= b;
    layer5_outputs(2125) <= not b;
    layer5_outputs(2126) <= not (a xor b);
    layer5_outputs(2127) <= not a;
    layer5_outputs(2128) <= a and b;
    layer5_outputs(2129) <= 1'b1;
    layer5_outputs(2130) <= not (a or b);
    layer5_outputs(2131) <= not b;
    layer5_outputs(2132) <= 1'b1;
    layer5_outputs(2133) <= a and b;
    layer5_outputs(2134) <= a or b;
    layer5_outputs(2135) <= not b or a;
    layer5_outputs(2136) <= a xor b;
    layer5_outputs(2137) <= not b;
    layer5_outputs(2138) <= not (a and b);
    layer5_outputs(2139) <= not b;
    layer5_outputs(2140) <= not b;
    layer5_outputs(2141) <= a or b;
    layer5_outputs(2142) <= a xor b;
    layer5_outputs(2143) <= a and b;
    layer5_outputs(2144) <= not a or b;
    layer5_outputs(2145) <= not (a and b);
    layer5_outputs(2146) <= not a or b;
    layer5_outputs(2147) <= a;
    layer5_outputs(2148) <= not a or b;
    layer5_outputs(2149) <= not a;
    layer5_outputs(2150) <= b;
    layer5_outputs(2151) <= 1'b1;
    layer5_outputs(2152) <= not b;
    layer5_outputs(2153) <= not a or b;
    layer5_outputs(2154) <= not b;
    layer5_outputs(2155) <= 1'b0;
    layer5_outputs(2156) <= not b;
    layer5_outputs(2157) <= not (a and b);
    layer5_outputs(2158) <= a and not b;
    layer5_outputs(2159) <= not a;
    layer5_outputs(2160) <= not b;
    layer5_outputs(2161) <= not b or a;
    layer5_outputs(2162) <= a;
    layer5_outputs(2163) <= not (a or b);
    layer5_outputs(2164) <= b;
    layer5_outputs(2165) <= a and b;
    layer5_outputs(2166) <= not (a or b);
    layer5_outputs(2167) <= not b;
    layer5_outputs(2168) <= b and not a;
    layer5_outputs(2169) <= not (a or b);
    layer5_outputs(2170) <= not a or b;
    layer5_outputs(2171) <= not b;
    layer5_outputs(2172) <= not b;
    layer5_outputs(2173) <= b;
    layer5_outputs(2174) <= not a;
    layer5_outputs(2175) <= not b;
    layer5_outputs(2176) <= not (a xor b);
    layer5_outputs(2177) <= not b or a;
    layer5_outputs(2178) <= not a;
    layer5_outputs(2179) <= not a;
    layer5_outputs(2180) <= a and b;
    layer5_outputs(2181) <= 1'b0;
    layer5_outputs(2182) <= not b;
    layer5_outputs(2183) <= not a;
    layer5_outputs(2184) <= a;
    layer5_outputs(2185) <= not a;
    layer5_outputs(2186) <= b;
    layer5_outputs(2187) <= a or b;
    layer5_outputs(2188) <= a and b;
    layer5_outputs(2189) <= not b or a;
    layer5_outputs(2190) <= a;
    layer5_outputs(2191) <= a and not b;
    layer5_outputs(2192) <= not a;
    layer5_outputs(2193) <= not b or a;
    layer5_outputs(2194) <= not b or a;
    layer5_outputs(2195) <= 1'b0;
    layer5_outputs(2196) <= not b;
    layer5_outputs(2197) <= not a;
    layer5_outputs(2198) <= b;
    layer5_outputs(2199) <= a and b;
    layer5_outputs(2200) <= b;
    layer5_outputs(2201) <= a or b;
    layer5_outputs(2202) <= not b;
    layer5_outputs(2203) <= 1'b0;
    layer5_outputs(2204) <= a xor b;
    layer5_outputs(2205) <= not b;
    layer5_outputs(2206) <= a;
    layer5_outputs(2207) <= 1'b0;
    layer5_outputs(2208) <= 1'b1;
    layer5_outputs(2209) <= not (a and b);
    layer5_outputs(2210) <= not (a and b);
    layer5_outputs(2211) <= not a;
    layer5_outputs(2212) <= b and not a;
    layer5_outputs(2213) <= b and not a;
    layer5_outputs(2214) <= not a;
    layer5_outputs(2215) <= not b;
    layer5_outputs(2216) <= not b;
    layer5_outputs(2217) <= not b;
    layer5_outputs(2218) <= a and not b;
    layer5_outputs(2219) <= not (a or b);
    layer5_outputs(2220) <= not (a and b);
    layer5_outputs(2221) <= not a or b;
    layer5_outputs(2222) <= not b;
    layer5_outputs(2223) <= a and b;
    layer5_outputs(2224) <= 1'b1;
    layer5_outputs(2225) <= not b;
    layer5_outputs(2226) <= not a or b;
    layer5_outputs(2227) <= a;
    layer5_outputs(2228) <= a xor b;
    layer5_outputs(2229) <= not b;
    layer5_outputs(2230) <= a xor b;
    layer5_outputs(2231) <= b;
    layer5_outputs(2232) <= not b or a;
    layer5_outputs(2233) <= not a;
    layer5_outputs(2234) <= not (a and b);
    layer5_outputs(2235) <= a and b;
    layer5_outputs(2236) <= not (a or b);
    layer5_outputs(2237) <= a xor b;
    layer5_outputs(2238) <= not a or b;
    layer5_outputs(2239) <= b;
    layer5_outputs(2240) <= not a;
    layer5_outputs(2241) <= 1'b0;
    layer5_outputs(2242) <= not a;
    layer5_outputs(2243) <= not b;
    layer5_outputs(2244) <= b and not a;
    layer5_outputs(2245) <= not (a xor b);
    layer5_outputs(2246) <= 1'b1;
    layer5_outputs(2247) <= not a;
    layer5_outputs(2248) <= 1'b1;
    layer5_outputs(2249) <= a or b;
    layer5_outputs(2250) <= not a or b;
    layer5_outputs(2251) <= not (a xor b);
    layer5_outputs(2252) <= not (a xor b);
    layer5_outputs(2253) <= not b;
    layer5_outputs(2254) <= not a;
    layer5_outputs(2255) <= not a;
    layer5_outputs(2256) <= b;
    layer5_outputs(2257) <= a and b;
    layer5_outputs(2258) <= b and not a;
    layer5_outputs(2259) <= not b;
    layer5_outputs(2260) <= not (a and b);
    layer5_outputs(2261) <= a and not b;
    layer5_outputs(2262) <= not b;
    layer5_outputs(2263) <= b and not a;
    layer5_outputs(2264) <= not a;
    layer5_outputs(2265) <= not (a and b);
    layer5_outputs(2266) <= not a;
    layer5_outputs(2267) <= b and not a;
    layer5_outputs(2268) <= a;
    layer5_outputs(2269) <= 1'b0;
    layer5_outputs(2270) <= b and not a;
    layer5_outputs(2271) <= not (a and b);
    layer5_outputs(2272) <= a or b;
    layer5_outputs(2273) <= 1'b0;
    layer5_outputs(2274) <= a and b;
    layer5_outputs(2275) <= b and not a;
    layer5_outputs(2276) <= not (a and b);
    layer5_outputs(2277) <= not b;
    layer5_outputs(2278) <= a or b;
    layer5_outputs(2279) <= a and b;
    layer5_outputs(2280) <= 1'b1;
    layer5_outputs(2281) <= a;
    layer5_outputs(2282) <= a and not b;
    layer5_outputs(2283) <= not b;
    layer5_outputs(2284) <= b;
    layer5_outputs(2285) <= not b;
    layer5_outputs(2286) <= b;
    layer5_outputs(2287) <= not (a xor b);
    layer5_outputs(2288) <= not b;
    layer5_outputs(2289) <= 1'b0;
    layer5_outputs(2290) <= a xor b;
    layer5_outputs(2291) <= a and not b;
    layer5_outputs(2292) <= not b or a;
    layer5_outputs(2293) <= not (a and b);
    layer5_outputs(2294) <= not b;
    layer5_outputs(2295) <= not a;
    layer5_outputs(2296) <= not b;
    layer5_outputs(2297) <= not a or b;
    layer5_outputs(2298) <= not b;
    layer5_outputs(2299) <= b;
    layer5_outputs(2300) <= not (a or b);
    layer5_outputs(2301) <= b;
    layer5_outputs(2302) <= a;
    layer5_outputs(2303) <= b and not a;
    layer5_outputs(2304) <= not (a and b);
    layer5_outputs(2305) <= a;
    layer5_outputs(2306) <= a;
    layer5_outputs(2307) <= b;
    layer5_outputs(2308) <= not a;
    layer5_outputs(2309) <= not b;
    layer5_outputs(2310) <= b and not a;
    layer5_outputs(2311) <= b and not a;
    layer5_outputs(2312) <= not b or a;
    layer5_outputs(2313) <= a xor b;
    layer5_outputs(2314) <= a and b;
    layer5_outputs(2315) <= a;
    layer5_outputs(2316) <= not b;
    layer5_outputs(2317) <= a or b;
    layer5_outputs(2318) <= a and not b;
    layer5_outputs(2319) <= 1'b1;
    layer5_outputs(2320) <= not (a or b);
    layer5_outputs(2321) <= not (a or b);
    layer5_outputs(2322) <= a and not b;
    layer5_outputs(2323) <= b and not a;
    layer5_outputs(2324) <= b;
    layer5_outputs(2325) <= not b or a;
    layer5_outputs(2326) <= a or b;
    layer5_outputs(2327) <= not b;
    layer5_outputs(2328) <= a xor b;
    layer5_outputs(2329) <= not a or b;
    layer5_outputs(2330) <= not (a or b);
    layer5_outputs(2331) <= 1'b0;
    layer5_outputs(2332) <= b;
    layer5_outputs(2333) <= a and b;
    layer5_outputs(2334) <= b;
    layer5_outputs(2335) <= b;
    layer5_outputs(2336) <= not b or a;
    layer5_outputs(2337) <= a and b;
    layer5_outputs(2338) <= not b or a;
    layer5_outputs(2339) <= not a;
    layer5_outputs(2340) <= a xor b;
    layer5_outputs(2341) <= a;
    layer5_outputs(2342) <= not (a xor b);
    layer5_outputs(2343) <= b and not a;
    layer5_outputs(2344) <= 1'b1;
    layer5_outputs(2345) <= not a or b;
    layer5_outputs(2346) <= not a or b;
    layer5_outputs(2347) <= not a or b;
    layer5_outputs(2348) <= a xor b;
    layer5_outputs(2349) <= not a;
    layer5_outputs(2350) <= a or b;
    layer5_outputs(2351) <= not a or b;
    layer5_outputs(2352) <= not (a or b);
    layer5_outputs(2353) <= a and not b;
    layer5_outputs(2354) <= a xor b;
    layer5_outputs(2355) <= a;
    layer5_outputs(2356) <= a;
    layer5_outputs(2357) <= not b or a;
    layer5_outputs(2358) <= 1'b1;
    layer5_outputs(2359) <= not a;
    layer5_outputs(2360) <= a and not b;
    layer5_outputs(2361) <= not b;
    layer5_outputs(2362) <= not (a and b);
    layer5_outputs(2363) <= not a;
    layer5_outputs(2364) <= not (a xor b);
    layer5_outputs(2365) <= a;
    layer5_outputs(2366) <= b and not a;
    layer5_outputs(2367) <= b;
    layer5_outputs(2368) <= a or b;
    layer5_outputs(2369) <= not (a and b);
    layer5_outputs(2370) <= not (a xor b);
    layer5_outputs(2371) <= b and not a;
    layer5_outputs(2372) <= b;
    layer5_outputs(2373) <= not a;
    layer5_outputs(2374) <= 1'b1;
    layer5_outputs(2375) <= a;
    layer5_outputs(2376) <= not (a or b);
    layer5_outputs(2377) <= 1'b0;
    layer5_outputs(2378) <= a xor b;
    layer5_outputs(2379) <= a and not b;
    layer5_outputs(2380) <= a xor b;
    layer5_outputs(2381) <= not a or b;
    layer5_outputs(2382) <= a and not b;
    layer5_outputs(2383) <= not (a or b);
    layer5_outputs(2384) <= b and not a;
    layer5_outputs(2385) <= a or b;
    layer5_outputs(2386) <= b;
    layer5_outputs(2387) <= not a;
    layer5_outputs(2388) <= not a or b;
    layer5_outputs(2389) <= a and b;
    layer5_outputs(2390) <= b;
    layer5_outputs(2391) <= b;
    layer5_outputs(2392) <= b;
    layer5_outputs(2393) <= a or b;
    layer5_outputs(2394) <= not b;
    layer5_outputs(2395) <= a;
    layer5_outputs(2396) <= a and not b;
    layer5_outputs(2397) <= 1'b1;
    layer5_outputs(2398) <= not (a and b);
    layer5_outputs(2399) <= b and not a;
    layer5_outputs(2400) <= not (a and b);
    layer5_outputs(2401) <= a and b;
    layer5_outputs(2402) <= not a;
    layer5_outputs(2403) <= not a;
    layer5_outputs(2404) <= not (a or b);
    layer5_outputs(2405) <= b;
    layer5_outputs(2406) <= not (a and b);
    layer5_outputs(2407) <= a and b;
    layer5_outputs(2408) <= not (a xor b);
    layer5_outputs(2409) <= b;
    layer5_outputs(2410) <= a and not b;
    layer5_outputs(2411) <= b;
    layer5_outputs(2412) <= not b;
    layer5_outputs(2413) <= 1'b0;
    layer5_outputs(2414) <= a;
    layer5_outputs(2415) <= a or b;
    layer5_outputs(2416) <= not a or b;
    layer5_outputs(2417) <= not b;
    layer5_outputs(2418) <= b and not a;
    layer5_outputs(2419) <= 1'b1;
    layer5_outputs(2420) <= not b;
    layer5_outputs(2421) <= not (a and b);
    layer5_outputs(2422) <= a and not b;
    layer5_outputs(2423) <= not b;
    layer5_outputs(2424) <= not a;
    layer5_outputs(2425) <= not (a xor b);
    layer5_outputs(2426) <= a or b;
    layer5_outputs(2427) <= not (a or b);
    layer5_outputs(2428) <= a and b;
    layer5_outputs(2429) <= not b;
    layer5_outputs(2430) <= not a or b;
    layer5_outputs(2431) <= not b or a;
    layer5_outputs(2432) <= not (a or b);
    layer5_outputs(2433) <= a or b;
    layer5_outputs(2434) <= not (a or b);
    layer5_outputs(2435) <= not (a and b);
    layer5_outputs(2436) <= not a;
    layer5_outputs(2437) <= not b or a;
    layer5_outputs(2438) <= a and b;
    layer5_outputs(2439) <= not (a and b);
    layer5_outputs(2440) <= a and b;
    layer5_outputs(2441) <= 1'b1;
    layer5_outputs(2442) <= a and b;
    layer5_outputs(2443) <= a or b;
    layer5_outputs(2444) <= b and not a;
    layer5_outputs(2445) <= a;
    layer5_outputs(2446) <= b;
    layer5_outputs(2447) <= a or b;
    layer5_outputs(2448) <= 1'b0;
    layer5_outputs(2449) <= not b;
    layer5_outputs(2450) <= a and not b;
    layer5_outputs(2451) <= not b;
    layer5_outputs(2452) <= b;
    layer5_outputs(2453) <= not a;
    layer5_outputs(2454) <= not a or b;
    layer5_outputs(2455) <= b;
    layer5_outputs(2456) <= not (a or b);
    layer5_outputs(2457) <= not a;
    layer5_outputs(2458) <= 1'b1;
    layer5_outputs(2459) <= not b;
    layer5_outputs(2460) <= not a;
    layer5_outputs(2461) <= a and b;
    layer5_outputs(2462) <= b and not a;
    layer5_outputs(2463) <= a and b;
    layer5_outputs(2464) <= not a or b;
    layer5_outputs(2465) <= b;
    layer5_outputs(2466) <= a and not b;
    layer5_outputs(2467) <= a xor b;
    layer5_outputs(2468) <= not b;
    layer5_outputs(2469) <= not (a xor b);
    layer5_outputs(2470) <= b;
    layer5_outputs(2471) <= b and not a;
    layer5_outputs(2472) <= a and b;
    layer5_outputs(2473) <= a and not b;
    layer5_outputs(2474) <= not b or a;
    layer5_outputs(2475) <= a and not b;
    layer5_outputs(2476) <= not (a and b);
    layer5_outputs(2477) <= not a;
    layer5_outputs(2478) <= not (a or b);
    layer5_outputs(2479) <= not b;
    layer5_outputs(2480) <= a;
    layer5_outputs(2481) <= a or b;
    layer5_outputs(2482) <= b;
    layer5_outputs(2483) <= 1'b0;
    layer5_outputs(2484) <= not a;
    layer5_outputs(2485) <= 1'b0;
    layer5_outputs(2486) <= 1'b0;
    layer5_outputs(2487) <= a and not b;
    layer5_outputs(2488) <= a and b;
    layer5_outputs(2489) <= not (a and b);
    layer5_outputs(2490) <= b and not a;
    layer5_outputs(2491) <= b and not a;
    layer5_outputs(2492) <= 1'b1;
    layer5_outputs(2493) <= a;
    layer5_outputs(2494) <= not (a and b);
    layer5_outputs(2495) <= not a or b;
    layer5_outputs(2496) <= b;
    layer5_outputs(2497) <= not a;
    layer5_outputs(2498) <= not b or a;
    layer5_outputs(2499) <= b;
    layer5_outputs(2500) <= not b or a;
    layer5_outputs(2501) <= not a or b;
    layer5_outputs(2502) <= not b;
    layer5_outputs(2503) <= b;
    layer5_outputs(2504) <= 1'b0;
    layer5_outputs(2505) <= 1'b0;
    layer5_outputs(2506) <= a and b;
    layer5_outputs(2507) <= a and b;
    layer5_outputs(2508) <= a;
    layer5_outputs(2509) <= not (a or b);
    layer5_outputs(2510) <= a and not b;
    layer5_outputs(2511) <= not a;
    layer5_outputs(2512) <= not a;
    layer5_outputs(2513) <= a xor b;
    layer5_outputs(2514) <= not b;
    layer5_outputs(2515) <= a and not b;
    layer5_outputs(2516) <= not (a and b);
    layer5_outputs(2517) <= a;
    layer5_outputs(2518) <= a;
    layer5_outputs(2519) <= not b or a;
    layer5_outputs(2520) <= b;
    layer5_outputs(2521) <= not (a and b);
    layer5_outputs(2522) <= a and not b;
    layer5_outputs(2523) <= not a or b;
    layer5_outputs(2524) <= not a;
    layer5_outputs(2525) <= a;
    layer5_outputs(2526) <= a xor b;
    layer5_outputs(2527) <= not b;
    layer5_outputs(2528) <= not (a and b);
    layer5_outputs(2529) <= b;
    layer5_outputs(2530) <= 1'b0;
    layer5_outputs(2531) <= not b or a;
    layer5_outputs(2532) <= a and not b;
    layer5_outputs(2533) <= 1'b1;
    layer5_outputs(2534) <= not (a or b);
    layer5_outputs(2535) <= a;
    layer5_outputs(2536) <= a xor b;
    layer5_outputs(2537) <= b;
    layer5_outputs(2538) <= not (a xor b);
    layer5_outputs(2539) <= not b;
    layer5_outputs(2540) <= a;
    layer5_outputs(2541) <= a and b;
    layer5_outputs(2542) <= a or b;
    layer5_outputs(2543) <= a and b;
    layer5_outputs(2544) <= not b or a;
    layer5_outputs(2545) <= not (a xor b);
    layer5_outputs(2546) <= a;
    layer5_outputs(2547) <= b;
    layer5_outputs(2548) <= not b or a;
    layer5_outputs(2549) <= not a;
    layer5_outputs(2550) <= a and not b;
    layer5_outputs(2551) <= not (a and b);
    layer5_outputs(2552) <= 1'b0;
    layer5_outputs(2553) <= a;
    layer5_outputs(2554) <= not (a and b);
    layer5_outputs(2555) <= not a or b;
    layer5_outputs(2556) <= a or b;
    layer5_outputs(2557) <= b and not a;
    layer5_outputs(2558) <= not a or b;
    layer5_outputs(2559) <= not b;
    layer5_outputs(2560) <= not (a or b);
    layer5_outputs(2561) <= a;
    layer5_outputs(2562) <= a xor b;
    layer5_outputs(2563) <= not (a xor b);
    layer5_outputs(2564) <= not b;
    layer5_outputs(2565) <= 1'b1;
    layer5_outputs(2566) <= 1'b0;
    layer5_outputs(2567) <= 1'b0;
    layer5_outputs(2568) <= a or b;
    layer5_outputs(2569) <= b;
    layer5_outputs(2570) <= not (a or b);
    layer5_outputs(2571) <= not (a xor b);
    layer5_outputs(2572) <= not b;
    layer5_outputs(2573) <= not b;
    layer5_outputs(2574) <= not a;
    layer5_outputs(2575) <= not (a or b);
    layer5_outputs(2576) <= a;
    layer5_outputs(2577) <= not a;
    layer5_outputs(2578) <= not b or a;
    layer5_outputs(2579) <= a and not b;
    layer5_outputs(2580) <= a xor b;
    layer5_outputs(2581) <= not (a or b);
    layer5_outputs(2582) <= a or b;
    layer5_outputs(2583) <= not (a and b);
    layer5_outputs(2584) <= a xor b;
    layer5_outputs(2585) <= not b;
    layer5_outputs(2586) <= a;
    layer5_outputs(2587) <= a or b;
    layer5_outputs(2588) <= not (a or b);
    layer5_outputs(2589) <= a and not b;
    layer5_outputs(2590) <= a and not b;
    layer5_outputs(2591) <= not b;
    layer5_outputs(2592) <= not (a and b);
    layer5_outputs(2593) <= a or b;
    layer5_outputs(2594) <= a and not b;
    layer5_outputs(2595) <= not (a or b);
    layer5_outputs(2596) <= 1'b1;
    layer5_outputs(2597) <= not b or a;
    layer5_outputs(2598) <= 1'b1;
    layer5_outputs(2599) <= not b;
    layer5_outputs(2600) <= not (a or b);
    layer5_outputs(2601) <= not a;
    layer5_outputs(2602) <= not a or b;
    layer5_outputs(2603) <= not b;
    layer5_outputs(2604) <= not (a and b);
    layer5_outputs(2605) <= b;
    layer5_outputs(2606) <= 1'b0;
    layer5_outputs(2607) <= a;
    layer5_outputs(2608) <= b;
    layer5_outputs(2609) <= not a;
    layer5_outputs(2610) <= b;
    layer5_outputs(2611) <= not (a and b);
    layer5_outputs(2612) <= not (a and b);
    layer5_outputs(2613) <= a;
    layer5_outputs(2614) <= not (a and b);
    layer5_outputs(2615) <= a and b;
    layer5_outputs(2616) <= a or b;
    layer5_outputs(2617) <= not a;
    layer5_outputs(2618) <= not (a or b);
    layer5_outputs(2619) <= a;
    layer5_outputs(2620) <= not (a xor b);
    layer5_outputs(2621) <= not b;
    layer5_outputs(2622) <= not b;
    layer5_outputs(2623) <= not a;
    layer5_outputs(2624) <= not a or b;
    layer5_outputs(2625) <= a and b;
    layer5_outputs(2626) <= 1'b1;
    layer5_outputs(2627) <= not a;
    layer5_outputs(2628) <= not a;
    layer5_outputs(2629) <= 1'b1;
    layer5_outputs(2630) <= b and not a;
    layer5_outputs(2631) <= 1'b0;
    layer5_outputs(2632) <= 1'b1;
    layer5_outputs(2633) <= b and not a;
    layer5_outputs(2634) <= not b;
    layer5_outputs(2635) <= a;
    layer5_outputs(2636) <= not a;
    layer5_outputs(2637) <= not (a xor b);
    layer5_outputs(2638) <= 1'b1;
    layer5_outputs(2639) <= b and not a;
    layer5_outputs(2640) <= not b;
    layer5_outputs(2641) <= a;
    layer5_outputs(2642) <= a and not b;
    layer5_outputs(2643) <= not (a or b);
    layer5_outputs(2644) <= not a;
    layer5_outputs(2645) <= not (a and b);
    layer5_outputs(2646) <= a or b;
    layer5_outputs(2647) <= not (a or b);
    layer5_outputs(2648) <= not a;
    layer5_outputs(2649) <= a or b;
    layer5_outputs(2650) <= not (a or b);
    layer5_outputs(2651) <= a;
    layer5_outputs(2652) <= 1'b1;
    layer5_outputs(2653) <= 1'b0;
    layer5_outputs(2654) <= not b or a;
    layer5_outputs(2655) <= a xor b;
    layer5_outputs(2656) <= not (a or b);
    layer5_outputs(2657) <= not (a and b);
    layer5_outputs(2658) <= b;
    layer5_outputs(2659) <= not a or b;
    layer5_outputs(2660) <= 1'b0;
    layer5_outputs(2661) <= not a;
    layer5_outputs(2662) <= not (a or b);
    layer5_outputs(2663) <= a xor b;
    layer5_outputs(2664) <= b;
    layer5_outputs(2665) <= a and not b;
    layer5_outputs(2666) <= not b;
    layer5_outputs(2667) <= not (a or b);
    layer5_outputs(2668) <= not (a and b);
    layer5_outputs(2669) <= b;
    layer5_outputs(2670) <= not a or b;
    layer5_outputs(2671) <= not (a xor b);
    layer5_outputs(2672) <= a;
    layer5_outputs(2673) <= not a;
    layer5_outputs(2674) <= not a;
    layer5_outputs(2675) <= a;
    layer5_outputs(2676) <= a;
    layer5_outputs(2677) <= a and b;
    layer5_outputs(2678) <= a and b;
    layer5_outputs(2679) <= a xor b;
    layer5_outputs(2680) <= not b;
    layer5_outputs(2681) <= a or b;
    layer5_outputs(2682) <= b;
    layer5_outputs(2683) <= a;
    layer5_outputs(2684) <= not a or b;
    layer5_outputs(2685) <= not a;
    layer5_outputs(2686) <= not b;
    layer5_outputs(2687) <= not b or a;
    layer5_outputs(2688) <= b and not a;
    layer5_outputs(2689) <= a and not b;
    layer5_outputs(2690) <= a and b;
    layer5_outputs(2691) <= a and not b;
    layer5_outputs(2692) <= not b;
    layer5_outputs(2693) <= not (a xor b);
    layer5_outputs(2694) <= not a;
    layer5_outputs(2695) <= a;
    layer5_outputs(2696) <= not a;
    layer5_outputs(2697) <= b;
    layer5_outputs(2698) <= b and not a;
    layer5_outputs(2699) <= not b;
    layer5_outputs(2700) <= a;
    layer5_outputs(2701) <= a and not b;
    layer5_outputs(2702) <= a and b;
    layer5_outputs(2703) <= not b or a;
    layer5_outputs(2704) <= 1'b0;
    layer5_outputs(2705) <= b and not a;
    layer5_outputs(2706) <= b and not a;
    layer5_outputs(2707) <= b and not a;
    layer5_outputs(2708) <= not (a and b);
    layer5_outputs(2709) <= b;
    layer5_outputs(2710) <= not (a xor b);
    layer5_outputs(2711) <= b;
    layer5_outputs(2712) <= not a;
    layer5_outputs(2713) <= a and not b;
    layer5_outputs(2714) <= a or b;
    layer5_outputs(2715) <= b;
    layer5_outputs(2716) <= not (a or b);
    layer5_outputs(2717) <= a and b;
    layer5_outputs(2718) <= a or b;
    layer5_outputs(2719) <= b and not a;
    layer5_outputs(2720) <= a and not b;
    layer5_outputs(2721) <= a and b;
    layer5_outputs(2722) <= b and not a;
    layer5_outputs(2723) <= b and not a;
    layer5_outputs(2724) <= not a;
    layer5_outputs(2725) <= b;
    layer5_outputs(2726) <= not (a and b);
    layer5_outputs(2727) <= a and b;
    layer5_outputs(2728) <= b;
    layer5_outputs(2729) <= a xor b;
    layer5_outputs(2730) <= not (a and b);
    layer5_outputs(2731) <= 1'b0;
    layer5_outputs(2732) <= b and not a;
    layer5_outputs(2733) <= b and not a;
    layer5_outputs(2734) <= a xor b;
    layer5_outputs(2735) <= not a or b;
    layer5_outputs(2736) <= not (a xor b);
    layer5_outputs(2737) <= a;
    layer5_outputs(2738) <= not (a and b);
    layer5_outputs(2739) <= 1'b0;
    layer5_outputs(2740) <= not a or b;
    layer5_outputs(2741) <= a;
    layer5_outputs(2742) <= b;
    layer5_outputs(2743) <= a and not b;
    layer5_outputs(2744) <= a and b;
    layer5_outputs(2745) <= not a;
    layer5_outputs(2746) <= not a;
    layer5_outputs(2747) <= not (a or b);
    layer5_outputs(2748) <= not b or a;
    layer5_outputs(2749) <= a xor b;
    layer5_outputs(2750) <= 1'b1;
    layer5_outputs(2751) <= b;
    layer5_outputs(2752) <= not b;
    layer5_outputs(2753) <= a and not b;
    layer5_outputs(2754) <= 1'b1;
    layer5_outputs(2755) <= not a or b;
    layer5_outputs(2756) <= 1'b0;
    layer5_outputs(2757) <= not b or a;
    layer5_outputs(2758) <= 1'b0;
    layer5_outputs(2759) <= not b;
    layer5_outputs(2760) <= not a;
    layer5_outputs(2761) <= not (a xor b);
    layer5_outputs(2762) <= a and b;
    layer5_outputs(2763) <= not a;
    layer5_outputs(2764) <= a and not b;
    layer5_outputs(2765) <= b and not a;
    layer5_outputs(2766) <= a or b;
    layer5_outputs(2767) <= a xor b;
    layer5_outputs(2768) <= a;
    layer5_outputs(2769) <= 1'b0;
    layer5_outputs(2770) <= b and not a;
    layer5_outputs(2771) <= 1'b0;
    layer5_outputs(2772) <= b;
    layer5_outputs(2773) <= a and not b;
    layer5_outputs(2774) <= not (a xor b);
    layer5_outputs(2775) <= b and not a;
    layer5_outputs(2776) <= a and b;
    layer5_outputs(2777) <= a;
    layer5_outputs(2778) <= not b;
    layer5_outputs(2779) <= not b;
    layer5_outputs(2780) <= not b;
    layer5_outputs(2781) <= not a or b;
    layer5_outputs(2782) <= not (a or b);
    layer5_outputs(2783) <= b and not a;
    layer5_outputs(2784) <= not a;
    layer5_outputs(2785) <= a;
    layer5_outputs(2786) <= 1'b0;
    layer5_outputs(2787) <= 1'b0;
    layer5_outputs(2788) <= not b;
    layer5_outputs(2789) <= b and not a;
    layer5_outputs(2790) <= a;
    layer5_outputs(2791) <= not (a or b);
    layer5_outputs(2792) <= a;
    layer5_outputs(2793) <= b;
    layer5_outputs(2794) <= not a;
    layer5_outputs(2795) <= a and b;
    layer5_outputs(2796) <= b and not a;
    layer5_outputs(2797) <= b;
    layer5_outputs(2798) <= not a;
    layer5_outputs(2799) <= 1'b0;
    layer5_outputs(2800) <= a and b;
    layer5_outputs(2801) <= 1'b0;
    layer5_outputs(2802) <= not a or b;
    layer5_outputs(2803) <= a;
    layer5_outputs(2804) <= not a;
    layer5_outputs(2805) <= a and b;
    layer5_outputs(2806) <= a or b;
    layer5_outputs(2807) <= not a or b;
    layer5_outputs(2808) <= not (a xor b);
    layer5_outputs(2809) <= b and not a;
    layer5_outputs(2810) <= not b;
    layer5_outputs(2811) <= 1'b1;
    layer5_outputs(2812) <= not (a and b);
    layer5_outputs(2813) <= a xor b;
    layer5_outputs(2814) <= a and not b;
    layer5_outputs(2815) <= b;
    layer5_outputs(2816) <= not b;
    layer5_outputs(2817) <= a or b;
    layer5_outputs(2818) <= a or b;
    layer5_outputs(2819) <= a xor b;
    layer5_outputs(2820) <= a and not b;
    layer5_outputs(2821) <= b;
    layer5_outputs(2822) <= not b;
    layer5_outputs(2823) <= b and not a;
    layer5_outputs(2824) <= a;
    layer5_outputs(2825) <= a and b;
    layer5_outputs(2826) <= 1'b1;
    layer5_outputs(2827) <= a xor b;
    layer5_outputs(2828) <= not b;
    layer5_outputs(2829) <= a;
    layer5_outputs(2830) <= not (a xor b);
    layer5_outputs(2831) <= not (a and b);
    layer5_outputs(2832) <= b;
    layer5_outputs(2833) <= a;
    layer5_outputs(2834) <= not b;
    layer5_outputs(2835) <= a;
    layer5_outputs(2836) <= not (a and b);
    layer5_outputs(2837) <= not (a xor b);
    layer5_outputs(2838) <= b and not a;
    layer5_outputs(2839) <= b;
    layer5_outputs(2840) <= 1'b1;
    layer5_outputs(2841) <= a and not b;
    layer5_outputs(2842) <= not a;
    layer5_outputs(2843) <= not a;
    layer5_outputs(2844) <= 1'b1;
    layer5_outputs(2845) <= not a;
    layer5_outputs(2846) <= 1'b0;
    layer5_outputs(2847) <= a xor b;
    layer5_outputs(2848) <= not b;
    layer5_outputs(2849) <= b;
    layer5_outputs(2850) <= not b or a;
    layer5_outputs(2851) <= b;
    layer5_outputs(2852) <= not a;
    layer5_outputs(2853) <= a and not b;
    layer5_outputs(2854) <= not (a and b);
    layer5_outputs(2855) <= a;
    layer5_outputs(2856) <= not a;
    layer5_outputs(2857) <= not a or b;
    layer5_outputs(2858) <= 1'b0;
    layer5_outputs(2859) <= not b or a;
    layer5_outputs(2860) <= a and not b;
    layer5_outputs(2861) <= a;
    layer5_outputs(2862) <= not (a or b);
    layer5_outputs(2863) <= b and not a;
    layer5_outputs(2864) <= 1'b1;
    layer5_outputs(2865) <= not b or a;
    layer5_outputs(2866) <= not a;
    layer5_outputs(2867) <= a;
    layer5_outputs(2868) <= b and not a;
    layer5_outputs(2869) <= not a or b;
    layer5_outputs(2870) <= a and not b;
    layer5_outputs(2871) <= 1'b1;
    layer5_outputs(2872) <= a;
    layer5_outputs(2873) <= not a or b;
    layer5_outputs(2874) <= b;
    layer5_outputs(2875) <= not (a and b);
    layer5_outputs(2876) <= 1'b1;
    layer5_outputs(2877) <= a or b;
    layer5_outputs(2878) <= not b or a;
    layer5_outputs(2879) <= b and not a;
    layer5_outputs(2880) <= not a;
    layer5_outputs(2881) <= not a;
    layer5_outputs(2882) <= b;
    layer5_outputs(2883) <= not (a and b);
    layer5_outputs(2884) <= a and b;
    layer5_outputs(2885) <= not a;
    layer5_outputs(2886) <= a or b;
    layer5_outputs(2887) <= b;
    layer5_outputs(2888) <= not a or b;
    layer5_outputs(2889) <= a or b;
    layer5_outputs(2890) <= b;
    layer5_outputs(2891) <= a and b;
    layer5_outputs(2892) <= not b;
    layer5_outputs(2893) <= b;
    layer5_outputs(2894) <= not b or a;
    layer5_outputs(2895) <= not (a or b);
    layer5_outputs(2896) <= a and b;
    layer5_outputs(2897) <= b and not a;
    layer5_outputs(2898) <= not a;
    layer5_outputs(2899) <= a and b;
    layer5_outputs(2900) <= b and not a;
    layer5_outputs(2901) <= a or b;
    layer5_outputs(2902) <= not (a or b);
    layer5_outputs(2903) <= not (a xor b);
    layer5_outputs(2904) <= a and not b;
    layer5_outputs(2905) <= not (a or b);
    layer5_outputs(2906) <= b and not a;
    layer5_outputs(2907) <= not b;
    layer5_outputs(2908) <= b and not a;
    layer5_outputs(2909) <= not b;
    layer5_outputs(2910) <= b and not a;
    layer5_outputs(2911) <= a and b;
    layer5_outputs(2912) <= a or b;
    layer5_outputs(2913) <= a and b;
    layer5_outputs(2914) <= b;
    layer5_outputs(2915) <= not b;
    layer5_outputs(2916) <= a;
    layer5_outputs(2917) <= a or b;
    layer5_outputs(2918) <= not b or a;
    layer5_outputs(2919) <= not b;
    layer5_outputs(2920) <= a;
    layer5_outputs(2921) <= a;
    layer5_outputs(2922) <= b;
    layer5_outputs(2923) <= b and not a;
    layer5_outputs(2924) <= b;
    layer5_outputs(2925) <= not (a or b);
    layer5_outputs(2926) <= a xor b;
    layer5_outputs(2927) <= not (a or b);
    layer5_outputs(2928) <= a and b;
    layer5_outputs(2929) <= not b;
    layer5_outputs(2930) <= not a;
    layer5_outputs(2931) <= not (a or b);
    layer5_outputs(2932) <= not b;
    layer5_outputs(2933) <= 1'b1;
    layer5_outputs(2934) <= b;
    layer5_outputs(2935) <= a and b;
    layer5_outputs(2936) <= b;
    layer5_outputs(2937) <= b and not a;
    layer5_outputs(2938) <= not (a and b);
    layer5_outputs(2939) <= not (a and b);
    layer5_outputs(2940) <= not b;
    layer5_outputs(2941) <= a;
    layer5_outputs(2942) <= not a;
    layer5_outputs(2943) <= a or b;
    layer5_outputs(2944) <= a and not b;
    layer5_outputs(2945) <= a and b;
    layer5_outputs(2946) <= a and not b;
    layer5_outputs(2947) <= 1'b1;
    layer5_outputs(2948) <= b;
    layer5_outputs(2949) <= b and not a;
    layer5_outputs(2950) <= not a;
    layer5_outputs(2951) <= a xor b;
    layer5_outputs(2952) <= not a;
    layer5_outputs(2953) <= not a;
    layer5_outputs(2954) <= not b;
    layer5_outputs(2955) <= a;
    layer5_outputs(2956) <= b and not a;
    layer5_outputs(2957) <= not (a xor b);
    layer5_outputs(2958) <= not b or a;
    layer5_outputs(2959) <= b and not a;
    layer5_outputs(2960) <= 1'b1;
    layer5_outputs(2961) <= b and not a;
    layer5_outputs(2962) <= not b;
    layer5_outputs(2963) <= a and not b;
    layer5_outputs(2964) <= a;
    layer5_outputs(2965) <= not (a or b);
    layer5_outputs(2966) <= not b;
    layer5_outputs(2967) <= not a or b;
    layer5_outputs(2968) <= a;
    layer5_outputs(2969) <= b;
    layer5_outputs(2970) <= a;
    layer5_outputs(2971) <= not (a or b);
    layer5_outputs(2972) <= not b or a;
    layer5_outputs(2973) <= not b or a;
    layer5_outputs(2974) <= b;
    layer5_outputs(2975) <= b and not a;
    layer5_outputs(2976) <= b;
    layer5_outputs(2977) <= a;
    layer5_outputs(2978) <= a;
    layer5_outputs(2979) <= a;
    layer5_outputs(2980) <= 1'b1;
    layer5_outputs(2981) <= a;
    layer5_outputs(2982) <= 1'b0;
    layer5_outputs(2983) <= a;
    layer5_outputs(2984) <= not b;
    layer5_outputs(2985) <= b and not a;
    layer5_outputs(2986) <= not a or b;
    layer5_outputs(2987) <= a or b;
    layer5_outputs(2988) <= not b;
    layer5_outputs(2989) <= a and b;
    layer5_outputs(2990) <= 1'b1;
    layer5_outputs(2991) <= not (a xor b);
    layer5_outputs(2992) <= not a;
    layer5_outputs(2993) <= not a or b;
    layer5_outputs(2994) <= not b or a;
    layer5_outputs(2995) <= b;
    layer5_outputs(2996) <= not a;
    layer5_outputs(2997) <= a;
    layer5_outputs(2998) <= 1'b0;
    layer5_outputs(2999) <= not (a and b);
    layer5_outputs(3000) <= a or b;
    layer5_outputs(3001) <= b;
    layer5_outputs(3002) <= a;
    layer5_outputs(3003) <= a xor b;
    layer5_outputs(3004) <= not a;
    layer5_outputs(3005) <= 1'b1;
    layer5_outputs(3006) <= not a or b;
    layer5_outputs(3007) <= b and not a;
    layer5_outputs(3008) <= 1'b1;
    layer5_outputs(3009) <= not (a or b);
    layer5_outputs(3010) <= not b;
    layer5_outputs(3011) <= not a or b;
    layer5_outputs(3012) <= not (a or b);
    layer5_outputs(3013) <= not b;
    layer5_outputs(3014) <= not b;
    layer5_outputs(3015) <= not b;
    layer5_outputs(3016) <= a or b;
    layer5_outputs(3017) <= 1'b0;
    layer5_outputs(3018) <= a and b;
    layer5_outputs(3019) <= not b;
    layer5_outputs(3020) <= not (a and b);
    layer5_outputs(3021) <= a and not b;
    layer5_outputs(3022) <= not a or b;
    layer5_outputs(3023) <= not (a xor b);
    layer5_outputs(3024) <= not (a and b);
    layer5_outputs(3025) <= not a or b;
    layer5_outputs(3026) <= 1'b1;
    layer5_outputs(3027) <= a or b;
    layer5_outputs(3028) <= not b;
    layer5_outputs(3029) <= not a or b;
    layer5_outputs(3030) <= b;
    layer5_outputs(3031) <= not (a or b);
    layer5_outputs(3032) <= not (a and b);
    layer5_outputs(3033) <= a;
    layer5_outputs(3034) <= a;
    layer5_outputs(3035) <= a and not b;
    layer5_outputs(3036) <= a and not b;
    layer5_outputs(3037) <= not a or b;
    layer5_outputs(3038) <= a or b;
    layer5_outputs(3039) <= not (a and b);
    layer5_outputs(3040) <= b;
    layer5_outputs(3041) <= a and not b;
    layer5_outputs(3042) <= not b;
    layer5_outputs(3043) <= a and b;
    layer5_outputs(3044) <= not (a or b);
    layer5_outputs(3045) <= b;
    layer5_outputs(3046) <= a and not b;
    layer5_outputs(3047) <= a and b;
    layer5_outputs(3048) <= a and b;
    layer5_outputs(3049) <= b;
    layer5_outputs(3050) <= not b;
    layer5_outputs(3051) <= not a or b;
    layer5_outputs(3052) <= a and b;
    layer5_outputs(3053) <= a and b;
    layer5_outputs(3054) <= b and not a;
    layer5_outputs(3055) <= not (a or b);
    layer5_outputs(3056) <= not (a and b);
    layer5_outputs(3057) <= b;
    layer5_outputs(3058) <= a and not b;
    layer5_outputs(3059) <= 1'b0;
    layer5_outputs(3060) <= 1'b1;
    layer5_outputs(3061) <= b;
    layer5_outputs(3062) <= not a or b;
    layer5_outputs(3063) <= not b;
    layer5_outputs(3064) <= not (a and b);
    layer5_outputs(3065) <= a and b;
    layer5_outputs(3066) <= not (a xor b);
    layer5_outputs(3067) <= not a or b;
    layer5_outputs(3068) <= not b or a;
    layer5_outputs(3069) <= 1'b1;
    layer5_outputs(3070) <= not (a xor b);
    layer5_outputs(3071) <= a;
    layer5_outputs(3072) <= a xor b;
    layer5_outputs(3073) <= b and not a;
    layer5_outputs(3074) <= not a or b;
    layer5_outputs(3075) <= b;
    layer5_outputs(3076) <= not a or b;
    layer5_outputs(3077) <= not (a and b);
    layer5_outputs(3078) <= a and not b;
    layer5_outputs(3079) <= not (a and b);
    layer5_outputs(3080) <= not b;
    layer5_outputs(3081) <= not (a xor b);
    layer5_outputs(3082) <= not (a xor b);
    layer5_outputs(3083) <= a;
    layer5_outputs(3084) <= not a;
    layer5_outputs(3085) <= b;
    layer5_outputs(3086) <= b;
    layer5_outputs(3087) <= a xor b;
    layer5_outputs(3088) <= a and b;
    layer5_outputs(3089) <= not (a and b);
    layer5_outputs(3090) <= not a;
    layer5_outputs(3091) <= a or b;
    layer5_outputs(3092) <= 1'b0;
    layer5_outputs(3093) <= b and not a;
    layer5_outputs(3094) <= not b or a;
    layer5_outputs(3095) <= not b or a;
    layer5_outputs(3096) <= not b or a;
    layer5_outputs(3097) <= not b;
    layer5_outputs(3098) <= b;
    layer5_outputs(3099) <= not (a or b);
    layer5_outputs(3100) <= a and b;
    layer5_outputs(3101) <= not (a and b);
    layer5_outputs(3102) <= b and not a;
    layer5_outputs(3103) <= not b or a;
    layer5_outputs(3104) <= a or b;
    layer5_outputs(3105) <= not a or b;
    layer5_outputs(3106) <= not (a or b);
    layer5_outputs(3107) <= a or b;
    layer5_outputs(3108) <= not b;
    layer5_outputs(3109) <= a xor b;
    layer5_outputs(3110) <= a and b;
    layer5_outputs(3111) <= a or b;
    layer5_outputs(3112) <= not (a and b);
    layer5_outputs(3113) <= b;
    layer5_outputs(3114) <= b;
    layer5_outputs(3115) <= not b;
    layer5_outputs(3116) <= b and not a;
    layer5_outputs(3117) <= a or b;
    layer5_outputs(3118) <= a and not b;
    layer5_outputs(3119) <= not b or a;
    layer5_outputs(3120) <= a;
    layer5_outputs(3121) <= a and b;
    layer5_outputs(3122) <= b;
    layer5_outputs(3123) <= a;
    layer5_outputs(3124) <= not (a or b);
    layer5_outputs(3125) <= a;
    layer5_outputs(3126) <= not (a and b);
    layer5_outputs(3127) <= a or b;
    layer5_outputs(3128) <= not b or a;
    layer5_outputs(3129) <= b and not a;
    layer5_outputs(3130) <= a or b;
    layer5_outputs(3131) <= b;
    layer5_outputs(3132) <= not (a and b);
    layer5_outputs(3133) <= not b;
    layer5_outputs(3134) <= b;
    layer5_outputs(3135) <= not b;
    layer5_outputs(3136) <= not b;
    layer5_outputs(3137) <= not (a xor b);
    layer5_outputs(3138) <= a;
    layer5_outputs(3139) <= b and not a;
    layer5_outputs(3140) <= not b;
    layer5_outputs(3141) <= not a or b;
    layer5_outputs(3142) <= 1'b0;
    layer5_outputs(3143) <= a and not b;
    layer5_outputs(3144) <= not a or b;
    layer5_outputs(3145) <= a xor b;
    layer5_outputs(3146) <= b;
    layer5_outputs(3147) <= a and not b;
    layer5_outputs(3148) <= not a;
    layer5_outputs(3149) <= not a or b;
    layer5_outputs(3150) <= b;
    layer5_outputs(3151) <= not a;
    layer5_outputs(3152) <= not (a or b);
    layer5_outputs(3153) <= not (a or b);
    layer5_outputs(3154) <= not a or b;
    layer5_outputs(3155) <= not a;
    layer5_outputs(3156) <= not (a and b);
    layer5_outputs(3157) <= a and b;
    layer5_outputs(3158) <= not (a xor b);
    layer5_outputs(3159) <= not a or b;
    layer5_outputs(3160) <= b;
    layer5_outputs(3161) <= 1'b1;
    layer5_outputs(3162) <= 1'b0;
    layer5_outputs(3163) <= a or b;
    layer5_outputs(3164) <= a xor b;
    layer5_outputs(3165) <= not a;
    layer5_outputs(3166) <= not b;
    layer5_outputs(3167) <= b;
    layer5_outputs(3168) <= not (a or b);
    layer5_outputs(3169) <= not a;
    layer5_outputs(3170) <= a or b;
    layer5_outputs(3171) <= 1'b0;
    layer5_outputs(3172) <= not (a or b);
    layer5_outputs(3173) <= not (a or b);
    layer5_outputs(3174) <= 1'b1;
    layer5_outputs(3175) <= not b;
    layer5_outputs(3176) <= a and not b;
    layer5_outputs(3177) <= a and b;
    layer5_outputs(3178) <= b;
    layer5_outputs(3179) <= not b;
    layer5_outputs(3180) <= 1'b0;
    layer5_outputs(3181) <= not (a or b);
    layer5_outputs(3182) <= not a or b;
    layer5_outputs(3183) <= not a or b;
    layer5_outputs(3184) <= not (a or b);
    layer5_outputs(3185) <= not b;
    layer5_outputs(3186) <= b and not a;
    layer5_outputs(3187) <= b;
    layer5_outputs(3188) <= 1'b1;
    layer5_outputs(3189) <= not (a and b);
    layer5_outputs(3190) <= a xor b;
    layer5_outputs(3191) <= b;
    layer5_outputs(3192) <= not a;
    layer5_outputs(3193) <= 1'b0;
    layer5_outputs(3194) <= not (a or b);
    layer5_outputs(3195) <= a and not b;
    layer5_outputs(3196) <= not a or b;
    layer5_outputs(3197) <= b;
    layer5_outputs(3198) <= a and not b;
    layer5_outputs(3199) <= a and not b;
    layer5_outputs(3200) <= b and not a;
    layer5_outputs(3201) <= not a;
    layer5_outputs(3202) <= not (a or b);
    layer5_outputs(3203) <= a;
    layer5_outputs(3204) <= not b;
    layer5_outputs(3205) <= not (a or b);
    layer5_outputs(3206) <= a or b;
    layer5_outputs(3207) <= a xor b;
    layer5_outputs(3208) <= a;
    layer5_outputs(3209) <= a;
    layer5_outputs(3210) <= not (a or b);
    layer5_outputs(3211) <= not a or b;
    layer5_outputs(3212) <= 1'b0;
    layer5_outputs(3213) <= a and not b;
    layer5_outputs(3214) <= not b or a;
    layer5_outputs(3215) <= not (a and b);
    layer5_outputs(3216) <= 1'b0;
    layer5_outputs(3217) <= not b;
    layer5_outputs(3218) <= a and b;
    layer5_outputs(3219) <= not a;
    layer5_outputs(3220) <= not (a xor b);
    layer5_outputs(3221) <= not (a xor b);
    layer5_outputs(3222) <= not b;
    layer5_outputs(3223) <= not (a xor b);
    layer5_outputs(3224) <= b;
    layer5_outputs(3225) <= b;
    layer5_outputs(3226) <= not a;
    layer5_outputs(3227) <= not a;
    layer5_outputs(3228) <= 1'b1;
    layer5_outputs(3229) <= a;
    layer5_outputs(3230) <= a and b;
    layer5_outputs(3231) <= a;
    layer5_outputs(3232) <= b and not a;
    layer5_outputs(3233) <= b;
    layer5_outputs(3234) <= a;
    layer5_outputs(3235) <= a and b;
    layer5_outputs(3236) <= not (a and b);
    layer5_outputs(3237) <= b;
    layer5_outputs(3238) <= not (a xor b);
    layer5_outputs(3239) <= a;
    layer5_outputs(3240) <= not (a xor b);
    layer5_outputs(3241) <= a;
    layer5_outputs(3242) <= not a or b;
    layer5_outputs(3243) <= not b;
    layer5_outputs(3244) <= not (a or b);
    layer5_outputs(3245) <= 1'b0;
    layer5_outputs(3246) <= not b;
    layer5_outputs(3247) <= not b or a;
    layer5_outputs(3248) <= 1'b0;
    layer5_outputs(3249) <= a;
    layer5_outputs(3250) <= not a or b;
    layer5_outputs(3251) <= a and b;
    layer5_outputs(3252) <= a or b;
    layer5_outputs(3253) <= a and not b;
    layer5_outputs(3254) <= 1'b1;
    layer5_outputs(3255) <= not b or a;
    layer5_outputs(3256) <= not b;
    layer5_outputs(3257) <= not b;
    layer5_outputs(3258) <= not a;
    layer5_outputs(3259) <= a or b;
    layer5_outputs(3260) <= a and not b;
    layer5_outputs(3261) <= a;
    layer5_outputs(3262) <= not b;
    layer5_outputs(3263) <= a and not b;
    layer5_outputs(3264) <= a;
    layer5_outputs(3265) <= a;
    layer5_outputs(3266) <= a;
    layer5_outputs(3267) <= not a;
    layer5_outputs(3268) <= a;
    layer5_outputs(3269) <= a or b;
    layer5_outputs(3270) <= a and b;
    layer5_outputs(3271) <= b;
    layer5_outputs(3272) <= a;
    layer5_outputs(3273) <= b and not a;
    layer5_outputs(3274) <= not a;
    layer5_outputs(3275) <= a or b;
    layer5_outputs(3276) <= 1'b0;
    layer5_outputs(3277) <= 1'b0;
    layer5_outputs(3278) <= not (a and b);
    layer5_outputs(3279) <= a or b;
    layer5_outputs(3280) <= a xor b;
    layer5_outputs(3281) <= b and not a;
    layer5_outputs(3282) <= a and b;
    layer5_outputs(3283) <= not b or a;
    layer5_outputs(3284) <= a and b;
    layer5_outputs(3285) <= 1'b0;
    layer5_outputs(3286) <= b;
    layer5_outputs(3287) <= a and b;
    layer5_outputs(3288) <= b and not a;
    layer5_outputs(3289) <= a or b;
    layer5_outputs(3290) <= a;
    layer5_outputs(3291) <= a and not b;
    layer5_outputs(3292) <= not b;
    layer5_outputs(3293) <= b and not a;
    layer5_outputs(3294) <= not (a or b);
    layer5_outputs(3295) <= not b;
    layer5_outputs(3296) <= not a;
    layer5_outputs(3297) <= 1'b0;
    layer5_outputs(3298) <= a or b;
    layer5_outputs(3299) <= not a;
    layer5_outputs(3300) <= 1'b1;
    layer5_outputs(3301) <= a or b;
    layer5_outputs(3302) <= 1'b1;
    layer5_outputs(3303) <= not b;
    layer5_outputs(3304) <= not a;
    layer5_outputs(3305) <= not b;
    layer5_outputs(3306) <= not b;
    layer5_outputs(3307) <= not b or a;
    layer5_outputs(3308) <= not a or b;
    layer5_outputs(3309) <= a and not b;
    layer5_outputs(3310) <= a;
    layer5_outputs(3311) <= not b;
    layer5_outputs(3312) <= a xor b;
    layer5_outputs(3313) <= a or b;
    layer5_outputs(3314) <= not (a and b);
    layer5_outputs(3315) <= not (a xor b);
    layer5_outputs(3316) <= a;
    layer5_outputs(3317) <= not (a and b);
    layer5_outputs(3318) <= a;
    layer5_outputs(3319) <= a and not b;
    layer5_outputs(3320) <= not (a or b);
    layer5_outputs(3321) <= a;
    layer5_outputs(3322) <= not b;
    layer5_outputs(3323) <= not b;
    layer5_outputs(3324) <= b;
    layer5_outputs(3325) <= a;
    layer5_outputs(3326) <= b and not a;
    layer5_outputs(3327) <= b and not a;
    layer5_outputs(3328) <= a and b;
    layer5_outputs(3329) <= not a;
    layer5_outputs(3330) <= not b;
    layer5_outputs(3331) <= not a;
    layer5_outputs(3332) <= b and not a;
    layer5_outputs(3333) <= not (a or b);
    layer5_outputs(3334) <= 1'b1;
    layer5_outputs(3335) <= not (a xor b);
    layer5_outputs(3336) <= a xor b;
    layer5_outputs(3337) <= not b or a;
    layer5_outputs(3338) <= a and b;
    layer5_outputs(3339) <= not (a or b);
    layer5_outputs(3340) <= a and b;
    layer5_outputs(3341) <= not a;
    layer5_outputs(3342) <= b;
    layer5_outputs(3343) <= a and b;
    layer5_outputs(3344) <= a and b;
    layer5_outputs(3345) <= a or b;
    layer5_outputs(3346) <= not a;
    layer5_outputs(3347) <= not a;
    layer5_outputs(3348) <= 1'b0;
    layer5_outputs(3349) <= a and not b;
    layer5_outputs(3350) <= 1'b1;
    layer5_outputs(3351) <= a;
    layer5_outputs(3352) <= a and b;
    layer5_outputs(3353) <= not a;
    layer5_outputs(3354) <= 1'b1;
    layer5_outputs(3355) <= not a or b;
    layer5_outputs(3356) <= not a;
    layer5_outputs(3357) <= not b;
    layer5_outputs(3358) <= b and not a;
    layer5_outputs(3359) <= not a;
    layer5_outputs(3360) <= b and not a;
    layer5_outputs(3361) <= b;
    layer5_outputs(3362) <= a;
    layer5_outputs(3363) <= not b;
    layer5_outputs(3364) <= a and b;
    layer5_outputs(3365) <= a xor b;
    layer5_outputs(3366) <= b;
    layer5_outputs(3367) <= not (a xor b);
    layer5_outputs(3368) <= b;
    layer5_outputs(3369) <= b and not a;
    layer5_outputs(3370) <= b;
    layer5_outputs(3371) <= a xor b;
    layer5_outputs(3372) <= not a or b;
    layer5_outputs(3373) <= not a;
    layer5_outputs(3374) <= not (a and b);
    layer5_outputs(3375) <= a xor b;
    layer5_outputs(3376) <= 1'b1;
    layer5_outputs(3377) <= a or b;
    layer5_outputs(3378) <= a;
    layer5_outputs(3379) <= not b;
    layer5_outputs(3380) <= a and b;
    layer5_outputs(3381) <= b;
    layer5_outputs(3382) <= not a;
    layer5_outputs(3383) <= not a or b;
    layer5_outputs(3384) <= a and not b;
    layer5_outputs(3385) <= a and b;
    layer5_outputs(3386) <= not b;
    layer5_outputs(3387) <= a and not b;
    layer5_outputs(3388) <= not a;
    layer5_outputs(3389) <= a or b;
    layer5_outputs(3390) <= a and not b;
    layer5_outputs(3391) <= a and b;
    layer5_outputs(3392) <= a;
    layer5_outputs(3393) <= 1'b1;
    layer5_outputs(3394) <= b;
    layer5_outputs(3395) <= a and b;
    layer5_outputs(3396) <= 1'b0;
    layer5_outputs(3397) <= not b or a;
    layer5_outputs(3398) <= not b;
    layer5_outputs(3399) <= a and not b;
    layer5_outputs(3400) <= 1'b0;
    layer5_outputs(3401) <= not (a and b);
    layer5_outputs(3402) <= a and b;
    layer5_outputs(3403) <= a or b;
    layer5_outputs(3404) <= a and not b;
    layer5_outputs(3405) <= not (a and b);
    layer5_outputs(3406) <= not (a xor b);
    layer5_outputs(3407) <= not (a xor b);
    layer5_outputs(3408) <= not b;
    layer5_outputs(3409) <= not a or b;
    layer5_outputs(3410) <= a;
    layer5_outputs(3411) <= 1'b0;
    layer5_outputs(3412) <= b;
    layer5_outputs(3413) <= not a;
    layer5_outputs(3414) <= b and not a;
    layer5_outputs(3415) <= a or b;
    layer5_outputs(3416) <= a xor b;
    layer5_outputs(3417) <= not (a xor b);
    layer5_outputs(3418) <= b;
    layer5_outputs(3419) <= not (a xor b);
    layer5_outputs(3420) <= not a;
    layer5_outputs(3421) <= not b;
    layer5_outputs(3422) <= b;
    layer5_outputs(3423) <= 1'b1;
    layer5_outputs(3424) <= not b or a;
    layer5_outputs(3425) <= not (a or b);
    layer5_outputs(3426) <= not (a or b);
    layer5_outputs(3427) <= a;
    layer5_outputs(3428) <= not (a or b);
    layer5_outputs(3429) <= a xor b;
    layer5_outputs(3430) <= a and b;
    layer5_outputs(3431) <= not (a and b);
    layer5_outputs(3432) <= a or b;
    layer5_outputs(3433) <= not a or b;
    layer5_outputs(3434) <= 1'b1;
    layer5_outputs(3435) <= not (a and b);
    layer5_outputs(3436) <= not (a and b);
    layer5_outputs(3437) <= 1'b0;
    layer5_outputs(3438) <= 1'b0;
    layer5_outputs(3439) <= b;
    layer5_outputs(3440) <= not b;
    layer5_outputs(3441) <= not b or a;
    layer5_outputs(3442) <= a or b;
    layer5_outputs(3443) <= a and not b;
    layer5_outputs(3444) <= a and b;
    layer5_outputs(3445) <= not b or a;
    layer5_outputs(3446) <= b;
    layer5_outputs(3447) <= not b;
    layer5_outputs(3448) <= not a;
    layer5_outputs(3449) <= 1'b0;
    layer5_outputs(3450) <= b;
    layer5_outputs(3451) <= b;
    layer5_outputs(3452) <= a;
    layer5_outputs(3453) <= not b;
    layer5_outputs(3454) <= 1'b0;
    layer5_outputs(3455) <= 1'b0;
    layer5_outputs(3456) <= not (a and b);
    layer5_outputs(3457) <= a;
    layer5_outputs(3458) <= b and not a;
    layer5_outputs(3459) <= b and not a;
    layer5_outputs(3460) <= 1'b0;
    layer5_outputs(3461) <= 1'b0;
    layer5_outputs(3462) <= a or b;
    layer5_outputs(3463) <= not (a and b);
    layer5_outputs(3464) <= b and not a;
    layer5_outputs(3465) <= not (a and b);
    layer5_outputs(3466) <= not a or b;
    layer5_outputs(3467) <= not b;
    layer5_outputs(3468) <= not (a or b);
    layer5_outputs(3469) <= not (a or b);
    layer5_outputs(3470) <= not a;
    layer5_outputs(3471) <= b;
    layer5_outputs(3472) <= not (a or b);
    layer5_outputs(3473) <= a xor b;
    layer5_outputs(3474) <= b;
    layer5_outputs(3475) <= b;
    layer5_outputs(3476) <= not b;
    layer5_outputs(3477) <= not (a and b);
    layer5_outputs(3478) <= 1'b1;
    layer5_outputs(3479) <= a and not b;
    layer5_outputs(3480) <= not a or b;
    layer5_outputs(3481) <= a or b;
    layer5_outputs(3482) <= not a;
    layer5_outputs(3483) <= 1'b1;
    layer5_outputs(3484) <= not (a and b);
    layer5_outputs(3485) <= not b or a;
    layer5_outputs(3486) <= a and not b;
    layer5_outputs(3487) <= a and not b;
    layer5_outputs(3488) <= b and not a;
    layer5_outputs(3489) <= a and not b;
    layer5_outputs(3490) <= a;
    layer5_outputs(3491) <= a and not b;
    layer5_outputs(3492) <= not (a or b);
    layer5_outputs(3493) <= not (a and b);
    layer5_outputs(3494) <= not b;
    layer5_outputs(3495) <= not (a or b);
    layer5_outputs(3496) <= 1'b0;
    layer5_outputs(3497) <= b;
    layer5_outputs(3498) <= not a;
    layer5_outputs(3499) <= not a;
    layer5_outputs(3500) <= not (a and b);
    layer5_outputs(3501) <= a and b;
    layer5_outputs(3502) <= not (a and b);
    layer5_outputs(3503) <= not (a xor b);
    layer5_outputs(3504) <= a or b;
    layer5_outputs(3505) <= not b;
    layer5_outputs(3506) <= not (a xor b);
    layer5_outputs(3507) <= not (a and b);
    layer5_outputs(3508) <= not (a and b);
    layer5_outputs(3509) <= a and b;
    layer5_outputs(3510) <= not (a and b);
    layer5_outputs(3511) <= not a or b;
    layer5_outputs(3512) <= not (a and b);
    layer5_outputs(3513) <= 1'b1;
    layer5_outputs(3514) <= a xor b;
    layer5_outputs(3515) <= b and not a;
    layer5_outputs(3516) <= a;
    layer5_outputs(3517) <= not (a and b);
    layer5_outputs(3518) <= not a;
    layer5_outputs(3519) <= not (a xor b);
    layer5_outputs(3520) <= not (a or b);
    layer5_outputs(3521) <= b;
    layer5_outputs(3522) <= b;
    layer5_outputs(3523) <= not (a or b);
    layer5_outputs(3524) <= not b or a;
    layer5_outputs(3525) <= not a or b;
    layer5_outputs(3526) <= a xor b;
    layer5_outputs(3527) <= not b or a;
    layer5_outputs(3528) <= a;
    layer5_outputs(3529) <= a;
    layer5_outputs(3530) <= not a;
    layer5_outputs(3531) <= b;
    layer5_outputs(3532) <= not b;
    layer5_outputs(3533) <= not b or a;
    layer5_outputs(3534) <= b and not a;
    layer5_outputs(3535) <= b;
    layer5_outputs(3536) <= not a;
    layer5_outputs(3537) <= a and b;
    layer5_outputs(3538) <= a and b;
    layer5_outputs(3539) <= a or b;
    layer5_outputs(3540) <= 1'b0;
    layer5_outputs(3541) <= 1'b0;
    layer5_outputs(3542) <= a xor b;
    layer5_outputs(3543) <= not a or b;
    layer5_outputs(3544) <= b and not a;
    layer5_outputs(3545) <= b;
    layer5_outputs(3546) <= not (a or b);
    layer5_outputs(3547) <= 1'b0;
    layer5_outputs(3548) <= a xor b;
    layer5_outputs(3549) <= not b;
    layer5_outputs(3550) <= 1'b1;
    layer5_outputs(3551) <= a and not b;
    layer5_outputs(3552) <= not a;
    layer5_outputs(3553) <= not b;
    layer5_outputs(3554) <= 1'b0;
    layer5_outputs(3555) <= 1'b0;
    layer5_outputs(3556) <= b;
    layer5_outputs(3557) <= not (a or b);
    layer5_outputs(3558) <= b;
    layer5_outputs(3559) <= not (a or b);
    layer5_outputs(3560) <= a and b;
    layer5_outputs(3561) <= not a or b;
    layer5_outputs(3562) <= not a or b;
    layer5_outputs(3563) <= not (a or b);
    layer5_outputs(3564) <= not (a xor b);
    layer5_outputs(3565) <= not b or a;
    layer5_outputs(3566) <= a and b;
    layer5_outputs(3567) <= a and not b;
    layer5_outputs(3568) <= a xor b;
    layer5_outputs(3569) <= not a or b;
    layer5_outputs(3570) <= a and not b;
    layer5_outputs(3571) <= not b or a;
    layer5_outputs(3572) <= a and b;
    layer5_outputs(3573) <= not b;
    layer5_outputs(3574) <= a or b;
    layer5_outputs(3575) <= not b;
    layer5_outputs(3576) <= 1'b0;
    layer5_outputs(3577) <= not a;
    layer5_outputs(3578) <= a;
    layer5_outputs(3579) <= not b;
    layer5_outputs(3580) <= a;
    layer5_outputs(3581) <= a or b;
    layer5_outputs(3582) <= not b or a;
    layer5_outputs(3583) <= a or b;
    layer5_outputs(3584) <= not b or a;
    layer5_outputs(3585) <= not b;
    layer5_outputs(3586) <= not b;
    layer5_outputs(3587) <= not b or a;
    layer5_outputs(3588) <= not b;
    layer5_outputs(3589) <= b and not a;
    layer5_outputs(3590) <= b and not a;
    layer5_outputs(3591) <= not (a xor b);
    layer5_outputs(3592) <= not a or b;
    layer5_outputs(3593) <= not a or b;
    layer5_outputs(3594) <= not b;
    layer5_outputs(3595) <= b;
    layer5_outputs(3596) <= a or b;
    layer5_outputs(3597) <= b and not a;
    layer5_outputs(3598) <= not b or a;
    layer5_outputs(3599) <= a;
    layer5_outputs(3600) <= not b or a;
    layer5_outputs(3601) <= not (a and b);
    layer5_outputs(3602) <= not a or b;
    layer5_outputs(3603) <= not b;
    layer5_outputs(3604) <= a;
    layer5_outputs(3605) <= b;
    layer5_outputs(3606) <= not (a or b);
    layer5_outputs(3607) <= not a or b;
    layer5_outputs(3608) <= not b;
    layer5_outputs(3609) <= a;
    layer5_outputs(3610) <= 1'b1;
    layer5_outputs(3611) <= b;
    layer5_outputs(3612) <= 1'b1;
    layer5_outputs(3613) <= b and not a;
    layer5_outputs(3614) <= b and not a;
    layer5_outputs(3615) <= 1'b1;
    layer5_outputs(3616) <= not (a xor b);
    layer5_outputs(3617) <= not b or a;
    layer5_outputs(3618) <= a xor b;
    layer5_outputs(3619) <= a;
    layer5_outputs(3620) <= not b;
    layer5_outputs(3621) <= not a or b;
    layer5_outputs(3622) <= not b or a;
    layer5_outputs(3623) <= not a;
    layer5_outputs(3624) <= not b or a;
    layer5_outputs(3625) <= not b;
    layer5_outputs(3626) <= a and b;
    layer5_outputs(3627) <= not (a xor b);
    layer5_outputs(3628) <= not (a xor b);
    layer5_outputs(3629) <= a and b;
    layer5_outputs(3630) <= a;
    layer5_outputs(3631) <= 1'b0;
    layer5_outputs(3632) <= not a;
    layer5_outputs(3633) <= 1'b0;
    layer5_outputs(3634) <= not (a or b);
    layer5_outputs(3635) <= b;
    layer5_outputs(3636) <= b and not a;
    layer5_outputs(3637) <= not (a and b);
    layer5_outputs(3638) <= a and not b;
    layer5_outputs(3639) <= a and not b;
    layer5_outputs(3640) <= not (a and b);
    layer5_outputs(3641) <= b and not a;
    layer5_outputs(3642) <= 1'b1;
    layer5_outputs(3643) <= not (a or b);
    layer5_outputs(3644) <= b;
    layer5_outputs(3645) <= not a;
    layer5_outputs(3646) <= a or b;
    layer5_outputs(3647) <= not (a xor b);
    layer5_outputs(3648) <= b and not a;
    layer5_outputs(3649) <= b and not a;
    layer5_outputs(3650) <= b;
    layer5_outputs(3651) <= a and not b;
    layer5_outputs(3652) <= b and not a;
    layer5_outputs(3653) <= a and b;
    layer5_outputs(3654) <= a and not b;
    layer5_outputs(3655) <= not a or b;
    layer5_outputs(3656) <= not a;
    layer5_outputs(3657) <= not a;
    layer5_outputs(3658) <= a and b;
    layer5_outputs(3659) <= 1'b0;
    layer5_outputs(3660) <= a;
    layer5_outputs(3661) <= not a;
    layer5_outputs(3662) <= a;
    layer5_outputs(3663) <= not b or a;
    layer5_outputs(3664) <= not b or a;
    layer5_outputs(3665) <= a;
    layer5_outputs(3666) <= not a;
    layer5_outputs(3667) <= not (a or b);
    layer5_outputs(3668) <= a and b;
    layer5_outputs(3669) <= not b;
    layer5_outputs(3670) <= b;
    layer5_outputs(3671) <= b;
    layer5_outputs(3672) <= a and not b;
    layer5_outputs(3673) <= not a or b;
    layer5_outputs(3674) <= not (a and b);
    layer5_outputs(3675) <= not a;
    layer5_outputs(3676) <= a and not b;
    layer5_outputs(3677) <= not b or a;
    layer5_outputs(3678) <= a or b;
    layer5_outputs(3679) <= not (a or b);
    layer5_outputs(3680) <= not b;
    layer5_outputs(3681) <= not b;
    layer5_outputs(3682) <= not b or a;
    layer5_outputs(3683) <= not (a and b);
    layer5_outputs(3684) <= 1'b1;
    layer5_outputs(3685) <= not b;
    layer5_outputs(3686) <= b and not a;
    layer5_outputs(3687) <= 1'b1;
    layer5_outputs(3688) <= a and not b;
    layer5_outputs(3689) <= not a or b;
    layer5_outputs(3690) <= b and not a;
    layer5_outputs(3691) <= not (a xor b);
    layer5_outputs(3692) <= a;
    layer5_outputs(3693) <= not (a and b);
    layer5_outputs(3694) <= 1'b1;
    layer5_outputs(3695) <= b and not a;
    layer5_outputs(3696) <= a and b;
    layer5_outputs(3697) <= a or b;
    layer5_outputs(3698) <= a and not b;
    layer5_outputs(3699) <= not a;
    layer5_outputs(3700) <= not a;
    layer5_outputs(3701) <= not a;
    layer5_outputs(3702) <= not (a and b);
    layer5_outputs(3703) <= a and not b;
    layer5_outputs(3704) <= a or b;
    layer5_outputs(3705) <= not b or a;
    layer5_outputs(3706) <= not a;
    layer5_outputs(3707) <= 1'b1;
    layer5_outputs(3708) <= b;
    layer5_outputs(3709) <= not a;
    layer5_outputs(3710) <= not b or a;
    layer5_outputs(3711) <= b;
    layer5_outputs(3712) <= a and not b;
    layer5_outputs(3713) <= not (a and b);
    layer5_outputs(3714) <= not (a or b);
    layer5_outputs(3715) <= a xor b;
    layer5_outputs(3716) <= 1'b0;
    layer5_outputs(3717) <= not b;
    layer5_outputs(3718) <= a;
    layer5_outputs(3719) <= not a or b;
    layer5_outputs(3720) <= a and not b;
    layer5_outputs(3721) <= b and not a;
    layer5_outputs(3722) <= b;
    layer5_outputs(3723) <= not (a xor b);
    layer5_outputs(3724) <= a and not b;
    layer5_outputs(3725) <= not a;
    layer5_outputs(3726) <= not (a or b);
    layer5_outputs(3727) <= a and not b;
    layer5_outputs(3728) <= 1'b1;
    layer5_outputs(3729) <= a;
    layer5_outputs(3730) <= a and not b;
    layer5_outputs(3731) <= not (a xor b);
    layer5_outputs(3732) <= not (a xor b);
    layer5_outputs(3733) <= not b or a;
    layer5_outputs(3734) <= not (a and b);
    layer5_outputs(3735) <= not (a or b);
    layer5_outputs(3736) <= 1'b1;
    layer5_outputs(3737) <= not a;
    layer5_outputs(3738) <= not a or b;
    layer5_outputs(3739) <= not b;
    layer5_outputs(3740) <= b;
    layer5_outputs(3741) <= not a or b;
    layer5_outputs(3742) <= b and not a;
    layer5_outputs(3743) <= not (a and b);
    layer5_outputs(3744) <= a;
    layer5_outputs(3745) <= not (a xor b);
    layer5_outputs(3746) <= not (a or b);
    layer5_outputs(3747) <= not b;
    layer5_outputs(3748) <= a;
    layer5_outputs(3749) <= not b;
    layer5_outputs(3750) <= a and b;
    layer5_outputs(3751) <= not b;
    layer5_outputs(3752) <= a and b;
    layer5_outputs(3753) <= b and not a;
    layer5_outputs(3754) <= a and not b;
    layer5_outputs(3755) <= not b;
    layer5_outputs(3756) <= b and not a;
    layer5_outputs(3757) <= 1'b0;
    layer5_outputs(3758) <= a;
    layer5_outputs(3759) <= not a or b;
    layer5_outputs(3760) <= b and not a;
    layer5_outputs(3761) <= not (a or b);
    layer5_outputs(3762) <= not a;
    layer5_outputs(3763) <= 1'b1;
    layer5_outputs(3764) <= a and b;
    layer5_outputs(3765) <= a or b;
    layer5_outputs(3766) <= a xor b;
    layer5_outputs(3767) <= not a;
    layer5_outputs(3768) <= not (a or b);
    layer5_outputs(3769) <= not a;
    layer5_outputs(3770) <= a and not b;
    layer5_outputs(3771) <= a and b;
    layer5_outputs(3772) <= b;
    layer5_outputs(3773) <= b and not a;
    layer5_outputs(3774) <= 1'b0;
    layer5_outputs(3775) <= not b;
    layer5_outputs(3776) <= a or b;
    layer5_outputs(3777) <= not a or b;
    layer5_outputs(3778) <= b;
    layer5_outputs(3779) <= a or b;
    layer5_outputs(3780) <= not a;
    layer5_outputs(3781) <= not a or b;
    layer5_outputs(3782) <= not (a or b);
    layer5_outputs(3783) <= not a or b;
    layer5_outputs(3784) <= not b or a;
    layer5_outputs(3785) <= not (a and b);
    layer5_outputs(3786) <= a and not b;
    layer5_outputs(3787) <= not b or a;
    layer5_outputs(3788) <= not (a xor b);
    layer5_outputs(3789) <= not (a xor b);
    layer5_outputs(3790) <= a or b;
    layer5_outputs(3791) <= a and b;
    layer5_outputs(3792) <= a xor b;
    layer5_outputs(3793) <= not (a and b);
    layer5_outputs(3794) <= a;
    layer5_outputs(3795) <= a xor b;
    layer5_outputs(3796) <= a xor b;
    layer5_outputs(3797) <= 1'b1;
    layer5_outputs(3798) <= not a;
    layer5_outputs(3799) <= b and not a;
    layer5_outputs(3800) <= not a;
    layer5_outputs(3801) <= a;
    layer5_outputs(3802) <= b and not a;
    layer5_outputs(3803) <= not b or a;
    layer5_outputs(3804) <= not b;
    layer5_outputs(3805) <= a or b;
    layer5_outputs(3806) <= b and not a;
    layer5_outputs(3807) <= a xor b;
    layer5_outputs(3808) <= not b;
    layer5_outputs(3809) <= b;
    layer5_outputs(3810) <= b;
    layer5_outputs(3811) <= a;
    layer5_outputs(3812) <= 1'b0;
    layer5_outputs(3813) <= not a;
    layer5_outputs(3814) <= b;
    layer5_outputs(3815) <= not a or b;
    layer5_outputs(3816) <= a and b;
    layer5_outputs(3817) <= b and not a;
    layer5_outputs(3818) <= not a or b;
    layer5_outputs(3819) <= a;
    layer5_outputs(3820) <= not a or b;
    layer5_outputs(3821) <= not a;
    layer5_outputs(3822) <= a;
    layer5_outputs(3823) <= not a or b;
    layer5_outputs(3824) <= not (a or b);
    layer5_outputs(3825) <= a;
    layer5_outputs(3826) <= not a;
    layer5_outputs(3827) <= not (a and b);
    layer5_outputs(3828) <= not (a and b);
    layer5_outputs(3829) <= a and not b;
    layer5_outputs(3830) <= not (a and b);
    layer5_outputs(3831) <= a;
    layer5_outputs(3832) <= not b;
    layer5_outputs(3833) <= not b or a;
    layer5_outputs(3834) <= a;
    layer5_outputs(3835) <= 1'b1;
    layer5_outputs(3836) <= b;
    layer5_outputs(3837) <= not (a or b);
    layer5_outputs(3838) <= not (a xor b);
    layer5_outputs(3839) <= not (a xor b);
    layer5_outputs(3840) <= not b;
    layer5_outputs(3841) <= not b;
    layer5_outputs(3842) <= not b;
    layer5_outputs(3843) <= not a or b;
    layer5_outputs(3844) <= b;
    layer5_outputs(3845) <= not (a or b);
    layer5_outputs(3846) <= 1'b1;
    layer5_outputs(3847) <= b;
    layer5_outputs(3848) <= b and not a;
    layer5_outputs(3849) <= a or b;
    layer5_outputs(3850) <= not b;
    layer5_outputs(3851) <= a or b;
    layer5_outputs(3852) <= a;
    layer5_outputs(3853) <= b and not a;
    layer5_outputs(3854) <= not a;
    layer5_outputs(3855) <= b;
    layer5_outputs(3856) <= not b;
    layer5_outputs(3857) <= not (a or b);
    layer5_outputs(3858) <= not a or b;
    layer5_outputs(3859) <= not a or b;
    layer5_outputs(3860) <= not (a and b);
    layer5_outputs(3861) <= a and not b;
    layer5_outputs(3862) <= not a;
    layer5_outputs(3863) <= b and not a;
    layer5_outputs(3864) <= b;
    layer5_outputs(3865) <= a;
    layer5_outputs(3866) <= not b;
    layer5_outputs(3867) <= a;
    layer5_outputs(3868) <= not (a xor b);
    layer5_outputs(3869) <= b;
    layer5_outputs(3870) <= a and not b;
    layer5_outputs(3871) <= a or b;
    layer5_outputs(3872) <= not b;
    layer5_outputs(3873) <= a and b;
    layer5_outputs(3874) <= not a or b;
    layer5_outputs(3875) <= b;
    layer5_outputs(3876) <= not (a or b);
    layer5_outputs(3877) <= a and not b;
    layer5_outputs(3878) <= b and not a;
    layer5_outputs(3879) <= a;
    layer5_outputs(3880) <= not b;
    layer5_outputs(3881) <= 1'b1;
    layer5_outputs(3882) <= not (a and b);
    layer5_outputs(3883) <= not (a and b);
    layer5_outputs(3884) <= a and b;
    layer5_outputs(3885) <= b and not a;
    layer5_outputs(3886) <= b;
    layer5_outputs(3887) <= a;
    layer5_outputs(3888) <= a;
    layer5_outputs(3889) <= not a or b;
    layer5_outputs(3890) <= b and not a;
    layer5_outputs(3891) <= b;
    layer5_outputs(3892) <= not b or a;
    layer5_outputs(3893) <= b and not a;
    layer5_outputs(3894) <= b and not a;
    layer5_outputs(3895) <= not a;
    layer5_outputs(3896) <= 1'b1;
    layer5_outputs(3897) <= a and b;
    layer5_outputs(3898) <= a and b;
    layer5_outputs(3899) <= not b;
    layer5_outputs(3900) <= not b or a;
    layer5_outputs(3901) <= b;
    layer5_outputs(3902) <= a and not b;
    layer5_outputs(3903) <= not a or b;
    layer5_outputs(3904) <= not (a and b);
    layer5_outputs(3905) <= not b or a;
    layer5_outputs(3906) <= a or b;
    layer5_outputs(3907) <= a and b;
    layer5_outputs(3908) <= a and b;
    layer5_outputs(3909) <= a;
    layer5_outputs(3910) <= 1'b1;
    layer5_outputs(3911) <= a;
    layer5_outputs(3912) <= not a or b;
    layer5_outputs(3913) <= b;
    layer5_outputs(3914) <= not a;
    layer5_outputs(3915) <= not (a and b);
    layer5_outputs(3916) <= not b or a;
    layer5_outputs(3917) <= a;
    layer5_outputs(3918) <= not (a and b);
    layer5_outputs(3919) <= not a or b;
    layer5_outputs(3920) <= b;
    layer5_outputs(3921) <= b and not a;
    layer5_outputs(3922) <= not a or b;
    layer5_outputs(3923) <= not a;
    layer5_outputs(3924) <= not b or a;
    layer5_outputs(3925) <= a or b;
    layer5_outputs(3926) <= 1'b0;
    layer5_outputs(3927) <= not (a and b);
    layer5_outputs(3928) <= a;
    layer5_outputs(3929) <= a and not b;
    layer5_outputs(3930) <= not a or b;
    layer5_outputs(3931) <= not a or b;
    layer5_outputs(3932) <= not (a or b);
    layer5_outputs(3933) <= a;
    layer5_outputs(3934) <= not b or a;
    layer5_outputs(3935) <= not a or b;
    layer5_outputs(3936) <= not (a or b);
    layer5_outputs(3937) <= not b or a;
    layer5_outputs(3938) <= a or b;
    layer5_outputs(3939) <= b;
    layer5_outputs(3940) <= not b or a;
    layer5_outputs(3941) <= a and b;
    layer5_outputs(3942) <= 1'b1;
    layer5_outputs(3943) <= not b;
    layer5_outputs(3944) <= a and not b;
    layer5_outputs(3945) <= a or b;
    layer5_outputs(3946) <= not a or b;
    layer5_outputs(3947) <= b and not a;
    layer5_outputs(3948) <= not b or a;
    layer5_outputs(3949) <= 1'b0;
    layer5_outputs(3950) <= 1'b0;
    layer5_outputs(3951) <= a and not b;
    layer5_outputs(3952) <= not a;
    layer5_outputs(3953) <= not b or a;
    layer5_outputs(3954) <= a and b;
    layer5_outputs(3955) <= not a;
    layer5_outputs(3956) <= a xor b;
    layer5_outputs(3957) <= a and not b;
    layer5_outputs(3958) <= a;
    layer5_outputs(3959) <= not b;
    layer5_outputs(3960) <= a and not b;
    layer5_outputs(3961) <= not b or a;
    layer5_outputs(3962) <= a xor b;
    layer5_outputs(3963) <= a and b;
    layer5_outputs(3964) <= a and b;
    layer5_outputs(3965) <= not a or b;
    layer5_outputs(3966) <= a;
    layer5_outputs(3967) <= 1'b0;
    layer5_outputs(3968) <= a and not b;
    layer5_outputs(3969) <= b;
    layer5_outputs(3970) <= b;
    layer5_outputs(3971) <= not b or a;
    layer5_outputs(3972) <= not a;
    layer5_outputs(3973) <= b and not a;
    layer5_outputs(3974) <= a;
    layer5_outputs(3975) <= not a;
    layer5_outputs(3976) <= b;
    layer5_outputs(3977) <= not b or a;
    layer5_outputs(3978) <= a;
    layer5_outputs(3979) <= not (a or b);
    layer5_outputs(3980) <= 1'b0;
    layer5_outputs(3981) <= a;
    layer5_outputs(3982) <= a;
    layer5_outputs(3983) <= not a;
    layer5_outputs(3984) <= not (a and b);
    layer5_outputs(3985) <= a;
    layer5_outputs(3986) <= b and not a;
    layer5_outputs(3987) <= a and b;
    layer5_outputs(3988) <= not a or b;
    layer5_outputs(3989) <= not a;
    layer5_outputs(3990) <= a and b;
    layer5_outputs(3991) <= a or b;
    layer5_outputs(3992) <= 1'b1;
    layer5_outputs(3993) <= not (a or b);
    layer5_outputs(3994) <= a xor b;
    layer5_outputs(3995) <= a and not b;
    layer5_outputs(3996) <= not b or a;
    layer5_outputs(3997) <= a;
    layer5_outputs(3998) <= a xor b;
    layer5_outputs(3999) <= not b or a;
    layer5_outputs(4000) <= not (a or b);
    layer5_outputs(4001) <= a;
    layer5_outputs(4002) <= b and not a;
    layer5_outputs(4003) <= b;
    layer5_outputs(4004) <= b;
    layer5_outputs(4005) <= not a;
    layer5_outputs(4006) <= 1'b1;
    layer5_outputs(4007) <= b;
    layer5_outputs(4008) <= a and b;
    layer5_outputs(4009) <= not b;
    layer5_outputs(4010) <= b;
    layer5_outputs(4011) <= b;
    layer5_outputs(4012) <= not b;
    layer5_outputs(4013) <= 1'b0;
    layer5_outputs(4014) <= not (a and b);
    layer5_outputs(4015) <= not b;
    layer5_outputs(4016) <= not a or b;
    layer5_outputs(4017) <= not b;
    layer5_outputs(4018) <= a;
    layer5_outputs(4019) <= b;
    layer5_outputs(4020) <= a or b;
    layer5_outputs(4021) <= b;
    layer5_outputs(4022) <= not b;
    layer5_outputs(4023) <= 1'b1;
    layer5_outputs(4024) <= a xor b;
    layer5_outputs(4025) <= b;
    layer5_outputs(4026) <= not b or a;
    layer5_outputs(4027) <= b;
    layer5_outputs(4028) <= not b;
    layer5_outputs(4029) <= not b or a;
    layer5_outputs(4030) <= b;
    layer5_outputs(4031) <= 1'b0;
    layer5_outputs(4032) <= b and not a;
    layer5_outputs(4033) <= b;
    layer5_outputs(4034) <= not a or b;
    layer5_outputs(4035) <= b;
    layer5_outputs(4036) <= not (a or b);
    layer5_outputs(4037) <= not a;
    layer5_outputs(4038) <= not b;
    layer5_outputs(4039) <= not a or b;
    layer5_outputs(4040) <= a and not b;
    layer5_outputs(4041) <= a and not b;
    layer5_outputs(4042) <= a or b;
    layer5_outputs(4043) <= a and b;
    layer5_outputs(4044) <= a or b;
    layer5_outputs(4045) <= a xor b;
    layer5_outputs(4046) <= not a or b;
    layer5_outputs(4047) <= not b;
    layer5_outputs(4048) <= a and b;
    layer5_outputs(4049) <= not (a xor b);
    layer5_outputs(4050) <= a;
    layer5_outputs(4051) <= a or b;
    layer5_outputs(4052) <= a and not b;
    layer5_outputs(4053) <= not a or b;
    layer5_outputs(4054) <= a and b;
    layer5_outputs(4055) <= not b;
    layer5_outputs(4056) <= a;
    layer5_outputs(4057) <= not a;
    layer5_outputs(4058) <= a and b;
    layer5_outputs(4059) <= a;
    layer5_outputs(4060) <= a;
    layer5_outputs(4061) <= not a;
    layer5_outputs(4062) <= 1'b1;
    layer5_outputs(4063) <= b;
    layer5_outputs(4064) <= not b;
    layer5_outputs(4065) <= a;
    layer5_outputs(4066) <= a and b;
    layer5_outputs(4067) <= a;
    layer5_outputs(4068) <= not a or b;
    layer5_outputs(4069) <= not b or a;
    layer5_outputs(4070) <= b;
    layer5_outputs(4071) <= not b or a;
    layer5_outputs(4072) <= not b;
    layer5_outputs(4073) <= not a;
    layer5_outputs(4074) <= not (a and b);
    layer5_outputs(4075) <= a and not b;
    layer5_outputs(4076) <= b and not a;
    layer5_outputs(4077) <= b and not a;
    layer5_outputs(4078) <= a and not b;
    layer5_outputs(4079) <= not a or b;
    layer5_outputs(4080) <= not (a and b);
    layer5_outputs(4081) <= a and b;
    layer5_outputs(4082) <= not b or a;
    layer5_outputs(4083) <= not b;
    layer5_outputs(4084) <= not b;
    layer5_outputs(4085) <= not b or a;
    layer5_outputs(4086) <= not b;
    layer5_outputs(4087) <= a and not b;
    layer5_outputs(4088) <= not b or a;
    layer5_outputs(4089) <= b and not a;
    layer5_outputs(4090) <= not (a and b);
    layer5_outputs(4091) <= a or b;
    layer5_outputs(4092) <= not b or a;
    layer5_outputs(4093) <= not b;
    layer5_outputs(4094) <= not b or a;
    layer5_outputs(4095) <= b;
    layer5_outputs(4096) <= 1'b1;
    layer5_outputs(4097) <= not a;
    layer5_outputs(4098) <= a and b;
    layer5_outputs(4099) <= 1'b0;
    layer5_outputs(4100) <= not a;
    layer5_outputs(4101) <= 1'b0;
    layer5_outputs(4102) <= not a;
    layer5_outputs(4103) <= not (a and b);
    layer5_outputs(4104) <= not (a or b);
    layer5_outputs(4105) <= not a;
    layer5_outputs(4106) <= not (a or b);
    layer5_outputs(4107) <= not (a or b);
    layer5_outputs(4108) <= not b;
    layer5_outputs(4109) <= not a or b;
    layer5_outputs(4110) <= not a;
    layer5_outputs(4111) <= a xor b;
    layer5_outputs(4112) <= not b or a;
    layer5_outputs(4113) <= b;
    layer5_outputs(4114) <= a and b;
    layer5_outputs(4115) <= b and not a;
    layer5_outputs(4116) <= not a;
    layer5_outputs(4117) <= not b;
    layer5_outputs(4118) <= a or b;
    layer5_outputs(4119) <= not b;
    layer5_outputs(4120) <= not b;
    layer5_outputs(4121) <= a;
    layer5_outputs(4122) <= a or b;
    layer5_outputs(4123) <= not b;
    layer5_outputs(4124) <= not b or a;
    layer5_outputs(4125) <= a and not b;
    layer5_outputs(4126) <= not (a or b);
    layer5_outputs(4127) <= a;
    layer5_outputs(4128) <= not a or b;
    layer5_outputs(4129) <= not a;
    layer5_outputs(4130) <= not b;
    layer5_outputs(4131) <= a xor b;
    layer5_outputs(4132) <= not (a or b);
    layer5_outputs(4133) <= a or b;
    layer5_outputs(4134) <= not (a and b);
    layer5_outputs(4135) <= not b;
    layer5_outputs(4136) <= a or b;
    layer5_outputs(4137) <= a or b;
    layer5_outputs(4138) <= a and b;
    layer5_outputs(4139) <= b;
    layer5_outputs(4140) <= not a or b;
    layer5_outputs(4141) <= not a or b;
    layer5_outputs(4142) <= not a or b;
    layer5_outputs(4143) <= a and b;
    layer5_outputs(4144) <= b;
    layer5_outputs(4145) <= not a;
    layer5_outputs(4146) <= not b;
    layer5_outputs(4147) <= 1'b1;
    layer5_outputs(4148) <= a and b;
    layer5_outputs(4149) <= a;
    layer5_outputs(4150) <= not a;
    layer5_outputs(4151) <= not (a xor b);
    layer5_outputs(4152) <= not a;
    layer5_outputs(4153) <= a;
    layer5_outputs(4154) <= not (a xor b);
    layer5_outputs(4155) <= a;
    layer5_outputs(4156) <= b and not a;
    layer5_outputs(4157) <= not a;
    layer5_outputs(4158) <= not a;
    layer5_outputs(4159) <= b;
    layer5_outputs(4160) <= a or b;
    layer5_outputs(4161) <= not a;
    layer5_outputs(4162) <= b;
    layer5_outputs(4163) <= a and not b;
    layer5_outputs(4164) <= not a or b;
    layer5_outputs(4165) <= b;
    layer5_outputs(4166) <= not b;
    layer5_outputs(4167) <= a xor b;
    layer5_outputs(4168) <= not a or b;
    layer5_outputs(4169) <= a xor b;
    layer5_outputs(4170) <= a;
    layer5_outputs(4171) <= 1'b1;
    layer5_outputs(4172) <= 1'b1;
    layer5_outputs(4173) <= not a;
    layer5_outputs(4174) <= not a or b;
    layer5_outputs(4175) <= not a;
    layer5_outputs(4176) <= not (a and b);
    layer5_outputs(4177) <= b;
    layer5_outputs(4178) <= not a;
    layer5_outputs(4179) <= not (a and b);
    layer5_outputs(4180) <= not b or a;
    layer5_outputs(4181) <= a or b;
    layer5_outputs(4182) <= not b or a;
    layer5_outputs(4183) <= a;
    layer5_outputs(4184) <= 1'b0;
    layer5_outputs(4185) <= b and not a;
    layer5_outputs(4186) <= a;
    layer5_outputs(4187) <= not (a or b);
    layer5_outputs(4188) <= not a or b;
    layer5_outputs(4189) <= not (a or b);
    layer5_outputs(4190) <= b;
    layer5_outputs(4191) <= b;
    layer5_outputs(4192) <= not b;
    layer5_outputs(4193) <= 1'b1;
    layer5_outputs(4194) <= b and not a;
    layer5_outputs(4195) <= 1'b0;
    layer5_outputs(4196) <= not b;
    layer5_outputs(4197) <= 1'b1;
    layer5_outputs(4198) <= not (a and b);
    layer5_outputs(4199) <= b and not a;
    layer5_outputs(4200) <= a xor b;
    layer5_outputs(4201) <= a;
    layer5_outputs(4202) <= not b or a;
    layer5_outputs(4203) <= b;
    layer5_outputs(4204) <= b;
    layer5_outputs(4205) <= not (a and b);
    layer5_outputs(4206) <= a;
    layer5_outputs(4207) <= not a;
    layer5_outputs(4208) <= b;
    layer5_outputs(4209) <= a or b;
    layer5_outputs(4210) <= not a or b;
    layer5_outputs(4211) <= a;
    layer5_outputs(4212) <= a or b;
    layer5_outputs(4213) <= b;
    layer5_outputs(4214) <= a xor b;
    layer5_outputs(4215) <= not (a or b);
    layer5_outputs(4216) <= not b;
    layer5_outputs(4217) <= a;
    layer5_outputs(4218) <= not b;
    layer5_outputs(4219) <= not b;
    layer5_outputs(4220) <= not a;
    layer5_outputs(4221) <= a or b;
    layer5_outputs(4222) <= not a;
    layer5_outputs(4223) <= 1'b1;
    layer5_outputs(4224) <= 1'b0;
    layer5_outputs(4225) <= b and not a;
    layer5_outputs(4226) <= 1'b1;
    layer5_outputs(4227) <= not b;
    layer5_outputs(4228) <= not a or b;
    layer5_outputs(4229) <= a or b;
    layer5_outputs(4230) <= not (a or b);
    layer5_outputs(4231) <= 1'b0;
    layer5_outputs(4232) <= a or b;
    layer5_outputs(4233) <= a;
    layer5_outputs(4234) <= b;
    layer5_outputs(4235) <= b;
    layer5_outputs(4236) <= b;
    layer5_outputs(4237) <= a;
    layer5_outputs(4238) <= not b or a;
    layer5_outputs(4239) <= b;
    layer5_outputs(4240) <= not (a xor b);
    layer5_outputs(4241) <= a and b;
    layer5_outputs(4242) <= not a or b;
    layer5_outputs(4243) <= a and not b;
    layer5_outputs(4244) <= a and b;
    layer5_outputs(4245) <= not (a or b);
    layer5_outputs(4246) <= b and not a;
    layer5_outputs(4247) <= not b;
    layer5_outputs(4248) <= a xor b;
    layer5_outputs(4249) <= b;
    layer5_outputs(4250) <= a and not b;
    layer5_outputs(4251) <= a or b;
    layer5_outputs(4252) <= b;
    layer5_outputs(4253) <= a;
    layer5_outputs(4254) <= b;
    layer5_outputs(4255) <= 1'b0;
    layer5_outputs(4256) <= not b or a;
    layer5_outputs(4257) <= not (a xor b);
    layer5_outputs(4258) <= a;
    layer5_outputs(4259) <= not b;
    layer5_outputs(4260) <= b and not a;
    layer5_outputs(4261) <= not (a or b);
    layer5_outputs(4262) <= not a or b;
    layer5_outputs(4263) <= a;
    layer5_outputs(4264) <= a and not b;
    layer5_outputs(4265) <= not (a and b);
    layer5_outputs(4266) <= a and not b;
    layer5_outputs(4267) <= b and not a;
    layer5_outputs(4268) <= not a or b;
    layer5_outputs(4269) <= b;
    layer5_outputs(4270) <= b;
    layer5_outputs(4271) <= 1'b0;
    layer5_outputs(4272) <= a;
    layer5_outputs(4273) <= not a;
    layer5_outputs(4274) <= a;
    layer5_outputs(4275) <= b and not a;
    layer5_outputs(4276) <= not a;
    layer5_outputs(4277) <= not (a xor b);
    layer5_outputs(4278) <= not b;
    layer5_outputs(4279) <= not (a and b);
    layer5_outputs(4280) <= 1'b1;
    layer5_outputs(4281) <= not b;
    layer5_outputs(4282) <= a or b;
    layer5_outputs(4283) <= b;
    layer5_outputs(4284) <= not b or a;
    layer5_outputs(4285) <= a;
    layer5_outputs(4286) <= a;
    layer5_outputs(4287) <= b;
    layer5_outputs(4288) <= a;
    layer5_outputs(4289) <= a and not b;
    layer5_outputs(4290) <= a and not b;
    layer5_outputs(4291) <= not (a or b);
    layer5_outputs(4292) <= a and b;
    layer5_outputs(4293) <= not (a or b);
    layer5_outputs(4294) <= not a;
    layer5_outputs(4295) <= a;
    layer5_outputs(4296) <= b;
    layer5_outputs(4297) <= not (a or b);
    layer5_outputs(4298) <= b;
    layer5_outputs(4299) <= not a or b;
    layer5_outputs(4300) <= not b;
    layer5_outputs(4301) <= a or b;
    layer5_outputs(4302) <= a;
    layer5_outputs(4303) <= not (a and b);
    layer5_outputs(4304) <= not b or a;
    layer5_outputs(4305) <= not a;
    layer5_outputs(4306) <= not (a and b);
    layer5_outputs(4307) <= not a or b;
    layer5_outputs(4308) <= 1'b0;
    layer5_outputs(4309) <= a and b;
    layer5_outputs(4310) <= a and not b;
    layer5_outputs(4311) <= a xor b;
    layer5_outputs(4312) <= not b;
    layer5_outputs(4313) <= not b or a;
    layer5_outputs(4314) <= not (a xor b);
    layer5_outputs(4315) <= b and not a;
    layer5_outputs(4316) <= b and not a;
    layer5_outputs(4317) <= a;
    layer5_outputs(4318) <= b;
    layer5_outputs(4319) <= a;
    layer5_outputs(4320) <= not (a xor b);
    layer5_outputs(4321) <= b;
    layer5_outputs(4322) <= a and b;
    layer5_outputs(4323) <= 1'b0;
    layer5_outputs(4324) <= 1'b0;
    layer5_outputs(4325) <= a;
    layer5_outputs(4326) <= b and not a;
    layer5_outputs(4327) <= b;
    layer5_outputs(4328) <= a xor b;
    layer5_outputs(4329) <= not b;
    layer5_outputs(4330) <= b and not a;
    layer5_outputs(4331) <= a and b;
    layer5_outputs(4332) <= a;
    layer5_outputs(4333) <= a;
    layer5_outputs(4334) <= not b;
    layer5_outputs(4335) <= not a or b;
    layer5_outputs(4336) <= not a;
    layer5_outputs(4337) <= b;
    layer5_outputs(4338) <= a or b;
    layer5_outputs(4339) <= b;
    layer5_outputs(4340) <= b and not a;
    layer5_outputs(4341) <= a and b;
    layer5_outputs(4342) <= a and b;
    layer5_outputs(4343) <= not (a or b);
    layer5_outputs(4344) <= 1'b1;
    layer5_outputs(4345) <= not b;
    layer5_outputs(4346) <= not b or a;
    layer5_outputs(4347) <= not b;
    layer5_outputs(4348) <= not b or a;
    layer5_outputs(4349) <= not b;
    layer5_outputs(4350) <= not (a xor b);
    layer5_outputs(4351) <= not a;
    layer5_outputs(4352) <= not a or b;
    layer5_outputs(4353) <= not b;
    layer5_outputs(4354) <= not b or a;
    layer5_outputs(4355) <= a and b;
    layer5_outputs(4356) <= not (a and b);
    layer5_outputs(4357) <= a or b;
    layer5_outputs(4358) <= not a;
    layer5_outputs(4359) <= b and not a;
    layer5_outputs(4360) <= 1'b1;
    layer5_outputs(4361) <= b and not a;
    layer5_outputs(4362) <= a and not b;
    layer5_outputs(4363) <= b and not a;
    layer5_outputs(4364) <= not (a xor b);
    layer5_outputs(4365) <= not (a xor b);
    layer5_outputs(4366) <= 1'b0;
    layer5_outputs(4367) <= not b;
    layer5_outputs(4368) <= a and b;
    layer5_outputs(4369) <= not (a xor b);
    layer5_outputs(4370) <= not a or b;
    layer5_outputs(4371) <= not (a or b);
    layer5_outputs(4372) <= b and not a;
    layer5_outputs(4373) <= a xor b;
    layer5_outputs(4374) <= b;
    layer5_outputs(4375) <= b;
    layer5_outputs(4376) <= a;
    layer5_outputs(4377) <= a and not b;
    layer5_outputs(4378) <= not b;
    layer5_outputs(4379) <= a and not b;
    layer5_outputs(4380) <= not a;
    layer5_outputs(4381) <= a and b;
    layer5_outputs(4382) <= a or b;
    layer5_outputs(4383) <= not b or a;
    layer5_outputs(4384) <= not (a or b);
    layer5_outputs(4385) <= not (a or b);
    layer5_outputs(4386) <= a and b;
    layer5_outputs(4387) <= b;
    layer5_outputs(4388) <= a or b;
    layer5_outputs(4389) <= 1'b0;
    layer5_outputs(4390) <= 1'b1;
    layer5_outputs(4391) <= 1'b0;
    layer5_outputs(4392) <= a and b;
    layer5_outputs(4393) <= 1'b0;
    layer5_outputs(4394) <= not (a xor b);
    layer5_outputs(4395) <= not b;
    layer5_outputs(4396) <= not b;
    layer5_outputs(4397) <= a and b;
    layer5_outputs(4398) <= not a;
    layer5_outputs(4399) <= a;
    layer5_outputs(4400) <= not b;
    layer5_outputs(4401) <= not a or b;
    layer5_outputs(4402) <= a;
    layer5_outputs(4403) <= not b;
    layer5_outputs(4404) <= not b or a;
    layer5_outputs(4405) <= not a or b;
    layer5_outputs(4406) <= not (a and b);
    layer5_outputs(4407) <= b;
    layer5_outputs(4408) <= not a;
    layer5_outputs(4409) <= not (a and b);
    layer5_outputs(4410) <= not a or b;
    layer5_outputs(4411) <= not a;
    layer5_outputs(4412) <= b and not a;
    layer5_outputs(4413) <= not (a and b);
    layer5_outputs(4414) <= not a;
    layer5_outputs(4415) <= b;
    layer5_outputs(4416) <= not (a xor b);
    layer5_outputs(4417) <= a or b;
    layer5_outputs(4418) <= not a;
    layer5_outputs(4419) <= not (a xor b);
    layer5_outputs(4420) <= a and not b;
    layer5_outputs(4421) <= a;
    layer5_outputs(4422) <= a or b;
    layer5_outputs(4423) <= not b or a;
    layer5_outputs(4424) <= not b;
    layer5_outputs(4425) <= a xor b;
    layer5_outputs(4426) <= not b;
    layer5_outputs(4427) <= not a or b;
    layer5_outputs(4428) <= a;
    layer5_outputs(4429) <= a;
    layer5_outputs(4430) <= not b;
    layer5_outputs(4431) <= 1'b1;
    layer5_outputs(4432) <= a or b;
    layer5_outputs(4433) <= not (a and b);
    layer5_outputs(4434) <= a or b;
    layer5_outputs(4435) <= a and not b;
    layer5_outputs(4436) <= a;
    layer5_outputs(4437) <= a and b;
    layer5_outputs(4438) <= not a;
    layer5_outputs(4439) <= not (a and b);
    layer5_outputs(4440) <= 1'b0;
    layer5_outputs(4441) <= not (a or b);
    layer5_outputs(4442) <= not b or a;
    layer5_outputs(4443) <= b and not a;
    layer5_outputs(4444) <= b and not a;
    layer5_outputs(4445) <= not a or b;
    layer5_outputs(4446) <= a and b;
    layer5_outputs(4447) <= not a or b;
    layer5_outputs(4448) <= not a;
    layer5_outputs(4449) <= b;
    layer5_outputs(4450) <= not a or b;
    layer5_outputs(4451) <= not (a or b);
    layer5_outputs(4452) <= not a or b;
    layer5_outputs(4453) <= a;
    layer5_outputs(4454) <= a and not b;
    layer5_outputs(4455) <= not (a xor b);
    layer5_outputs(4456) <= not (a and b);
    layer5_outputs(4457) <= not (a or b);
    layer5_outputs(4458) <= not (a or b);
    layer5_outputs(4459) <= not a;
    layer5_outputs(4460) <= not a;
    layer5_outputs(4461) <= not b;
    layer5_outputs(4462) <= b and not a;
    layer5_outputs(4463) <= a;
    layer5_outputs(4464) <= not (a xor b);
    layer5_outputs(4465) <= not b or a;
    layer5_outputs(4466) <= b and not a;
    layer5_outputs(4467) <= a or b;
    layer5_outputs(4468) <= a or b;
    layer5_outputs(4469) <= a;
    layer5_outputs(4470) <= not a;
    layer5_outputs(4471) <= not b or a;
    layer5_outputs(4472) <= a and not b;
    layer5_outputs(4473) <= a;
    layer5_outputs(4474) <= a and b;
    layer5_outputs(4475) <= not a;
    layer5_outputs(4476) <= not (a or b);
    layer5_outputs(4477) <= a;
    layer5_outputs(4478) <= a and b;
    layer5_outputs(4479) <= b;
    layer5_outputs(4480) <= b and not a;
    layer5_outputs(4481) <= not (a xor b);
    layer5_outputs(4482) <= not b;
    layer5_outputs(4483) <= not (a and b);
    layer5_outputs(4484) <= not b;
    layer5_outputs(4485) <= not b;
    layer5_outputs(4486) <= not a;
    layer5_outputs(4487) <= b and not a;
    layer5_outputs(4488) <= b;
    layer5_outputs(4489) <= not (a and b);
    layer5_outputs(4490) <= not (a or b);
    layer5_outputs(4491) <= a and not b;
    layer5_outputs(4492) <= 1'b0;
    layer5_outputs(4493) <= not (a and b);
    layer5_outputs(4494) <= b;
    layer5_outputs(4495) <= not a;
    layer5_outputs(4496) <= a and b;
    layer5_outputs(4497) <= b and not a;
    layer5_outputs(4498) <= a or b;
    layer5_outputs(4499) <= a and not b;
    layer5_outputs(4500) <= a;
    layer5_outputs(4501) <= 1'b1;
    layer5_outputs(4502) <= not (a or b);
    layer5_outputs(4503) <= not b or a;
    layer5_outputs(4504) <= a or b;
    layer5_outputs(4505) <= b;
    layer5_outputs(4506) <= a and b;
    layer5_outputs(4507) <= not (a or b);
    layer5_outputs(4508) <= not b;
    layer5_outputs(4509) <= not b or a;
    layer5_outputs(4510) <= a or b;
    layer5_outputs(4511) <= b;
    layer5_outputs(4512) <= a;
    layer5_outputs(4513) <= a;
    layer5_outputs(4514) <= not b;
    layer5_outputs(4515) <= a;
    layer5_outputs(4516) <= not a or b;
    layer5_outputs(4517) <= not b;
    layer5_outputs(4518) <= a and b;
    layer5_outputs(4519) <= b;
    layer5_outputs(4520) <= a;
    layer5_outputs(4521) <= not b;
    layer5_outputs(4522) <= a or b;
    layer5_outputs(4523) <= not b or a;
    layer5_outputs(4524) <= not b;
    layer5_outputs(4525) <= not a or b;
    layer5_outputs(4526) <= a and not b;
    layer5_outputs(4527) <= not a;
    layer5_outputs(4528) <= a;
    layer5_outputs(4529) <= a and b;
    layer5_outputs(4530) <= not a or b;
    layer5_outputs(4531) <= 1'b0;
    layer5_outputs(4532) <= not (a or b);
    layer5_outputs(4533) <= not (a and b);
    layer5_outputs(4534) <= 1'b1;
    layer5_outputs(4535) <= a and not b;
    layer5_outputs(4536) <= 1'b1;
    layer5_outputs(4537) <= not (a and b);
    layer5_outputs(4538) <= a;
    layer5_outputs(4539) <= not (a and b);
    layer5_outputs(4540) <= 1'b0;
    layer5_outputs(4541) <= a and not b;
    layer5_outputs(4542) <= not a;
    layer5_outputs(4543) <= b;
    layer5_outputs(4544) <= not (a and b);
    layer5_outputs(4545) <= a or b;
    layer5_outputs(4546) <= a xor b;
    layer5_outputs(4547) <= a xor b;
    layer5_outputs(4548) <= not a or b;
    layer5_outputs(4549) <= b;
    layer5_outputs(4550) <= not (a and b);
    layer5_outputs(4551) <= a and not b;
    layer5_outputs(4552) <= b;
    layer5_outputs(4553) <= a or b;
    layer5_outputs(4554) <= b and not a;
    layer5_outputs(4555) <= b;
    layer5_outputs(4556) <= not b;
    layer5_outputs(4557) <= not a;
    layer5_outputs(4558) <= not (a or b);
    layer5_outputs(4559) <= a xor b;
    layer5_outputs(4560) <= a and not b;
    layer5_outputs(4561) <= not b or a;
    layer5_outputs(4562) <= a xor b;
    layer5_outputs(4563) <= not b;
    layer5_outputs(4564) <= 1'b0;
    layer5_outputs(4565) <= a and not b;
    layer5_outputs(4566) <= not (a or b);
    layer5_outputs(4567) <= a xor b;
    layer5_outputs(4568) <= a;
    layer5_outputs(4569) <= not (a or b);
    layer5_outputs(4570) <= not a;
    layer5_outputs(4571) <= a or b;
    layer5_outputs(4572) <= b;
    layer5_outputs(4573) <= a or b;
    layer5_outputs(4574) <= a;
    layer5_outputs(4575) <= not (a and b);
    layer5_outputs(4576) <= 1'b0;
    layer5_outputs(4577) <= a or b;
    layer5_outputs(4578) <= b;
    layer5_outputs(4579) <= not a or b;
    layer5_outputs(4580) <= a and b;
    layer5_outputs(4581) <= a and not b;
    layer5_outputs(4582) <= a and b;
    layer5_outputs(4583) <= b and not a;
    layer5_outputs(4584) <= a;
    layer5_outputs(4585) <= 1'b1;
    layer5_outputs(4586) <= b and not a;
    layer5_outputs(4587) <= a and b;
    layer5_outputs(4588) <= b and not a;
    layer5_outputs(4589) <= b;
    layer5_outputs(4590) <= a xor b;
    layer5_outputs(4591) <= not (a or b);
    layer5_outputs(4592) <= not a;
    layer5_outputs(4593) <= b;
    layer5_outputs(4594) <= not b or a;
    layer5_outputs(4595) <= b;
    layer5_outputs(4596) <= a or b;
    layer5_outputs(4597) <= not a;
    layer5_outputs(4598) <= not a or b;
    layer5_outputs(4599) <= not a;
    layer5_outputs(4600) <= a;
    layer5_outputs(4601) <= not a;
    layer5_outputs(4602) <= not a;
    layer5_outputs(4603) <= not (a or b);
    layer5_outputs(4604) <= a;
    layer5_outputs(4605) <= a;
    layer5_outputs(4606) <= b;
    layer5_outputs(4607) <= not a or b;
    layer5_outputs(4608) <= not (a or b);
    layer5_outputs(4609) <= a and b;
    layer5_outputs(4610) <= not a;
    layer5_outputs(4611) <= 1'b1;
    layer5_outputs(4612) <= not a;
    layer5_outputs(4613) <= b and not a;
    layer5_outputs(4614) <= a and not b;
    layer5_outputs(4615) <= b;
    layer5_outputs(4616) <= a xor b;
    layer5_outputs(4617) <= b and not a;
    layer5_outputs(4618) <= a and not b;
    layer5_outputs(4619) <= a and not b;
    layer5_outputs(4620) <= b and not a;
    layer5_outputs(4621) <= a;
    layer5_outputs(4622) <= not a;
    layer5_outputs(4623) <= not a or b;
    layer5_outputs(4624) <= a;
    layer5_outputs(4625) <= not b or a;
    layer5_outputs(4626) <= b and not a;
    layer5_outputs(4627) <= a and not b;
    layer5_outputs(4628) <= 1'b1;
    layer5_outputs(4629) <= not a;
    layer5_outputs(4630) <= not a or b;
    layer5_outputs(4631) <= not (a and b);
    layer5_outputs(4632) <= a or b;
    layer5_outputs(4633) <= a xor b;
    layer5_outputs(4634) <= not (a or b);
    layer5_outputs(4635) <= not a;
    layer5_outputs(4636) <= a and b;
    layer5_outputs(4637) <= a and b;
    layer5_outputs(4638) <= a;
    layer5_outputs(4639) <= b;
    layer5_outputs(4640) <= a and b;
    layer5_outputs(4641) <= not b;
    layer5_outputs(4642) <= not b;
    layer5_outputs(4643) <= not b;
    layer5_outputs(4644) <= not a;
    layer5_outputs(4645) <= 1'b1;
    layer5_outputs(4646) <= not a;
    layer5_outputs(4647) <= not (a and b);
    layer5_outputs(4648) <= not b or a;
    layer5_outputs(4649) <= a or b;
    layer5_outputs(4650) <= not (a or b);
    layer5_outputs(4651) <= 1'b0;
    layer5_outputs(4652) <= b;
    layer5_outputs(4653) <= not (a or b);
    layer5_outputs(4654) <= a or b;
    layer5_outputs(4655) <= a and b;
    layer5_outputs(4656) <= 1'b1;
    layer5_outputs(4657) <= not b;
    layer5_outputs(4658) <= a;
    layer5_outputs(4659) <= not (a or b);
    layer5_outputs(4660) <= b;
    layer5_outputs(4661) <= not a or b;
    layer5_outputs(4662) <= not b;
    layer5_outputs(4663) <= b and not a;
    layer5_outputs(4664) <= not b;
    layer5_outputs(4665) <= a and not b;
    layer5_outputs(4666) <= a and not b;
    layer5_outputs(4667) <= not a or b;
    layer5_outputs(4668) <= not b;
    layer5_outputs(4669) <= not b;
    layer5_outputs(4670) <= not b;
    layer5_outputs(4671) <= not a or b;
    layer5_outputs(4672) <= 1'b1;
    layer5_outputs(4673) <= a and not b;
    layer5_outputs(4674) <= b and not a;
    layer5_outputs(4675) <= not (a and b);
    layer5_outputs(4676) <= not b;
    layer5_outputs(4677) <= b;
    layer5_outputs(4678) <= b and not a;
    layer5_outputs(4679) <= not (a and b);
    layer5_outputs(4680) <= b;
    layer5_outputs(4681) <= a;
    layer5_outputs(4682) <= a;
    layer5_outputs(4683) <= a and not b;
    layer5_outputs(4684) <= b;
    layer5_outputs(4685) <= a or b;
    layer5_outputs(4686) <= not (a or b);
    layer5_outputs(4687) <= a xor b;
    layer5_outputs(4688) <= not a;
    layer5_outputs(4689) <= not a or b;
    layer5_outputs(4690) <= b;
    layer5_outputs(4691) <= not b;
    layer5_outputs(4692) <= a and not b;
    layer5_outputs(4693) <= 1'b0;
    layer5_outputs(4694) <= a and b;
    layer5_outputs(4695) <= a;
    layer5_outputs(4696) <= a;
    layer5_outputs(4697) <= a and not b;
    layer5_outputs(4698) <= a;
    layer5_outputs(4699) <= b;
    layer5_outputs(4700) <= a or b;
    layer5_outputs(4701) <= not a;
    layer5_outputs(4702) <= not b or a;
    layer5_outputs(4703) <= b and not a;
    layer5_outputs(4704) <= not b;
    layer5_outputs(4705) <= not a or b;
    layer5_outputs(4706) <= a or b;
    layer5_outputs(4707) <= not a;
    layer5_outputs(4708) <= 1'b1;
    layer5_outputs(4709) <= not a or b;
    layer5_outputs(4710) <= a and b;
    layer5_outputs(4711) <= b;
    layer5_outputs(4712) <= not (a or b);
    layer5_outputs(4713) <= a xor b;
    layer5_outputs(4714) <= not b or a;
    layer5_outputs(4715) <= b and not a;
    layer5_outputs(4716) <= not (a xor b);
    layer5_outputs(4717) <= a xor b;
    layer5_outputs(4718) <= not a;
    layer5_outputs(4719) <= not b or a;
    layer5_outputs(4720) <= a or b;
    layer5_outputs(4721) <= b;
    layer5_outputs(4722) <= not a;
    layer5_outputs(4723) <= a;
    layer5_outputs(4724) <= b and not a;
    layer5_outputs(4725) <= not a;
    layer5_outputs(4726) <= a or b;
    layer5_outputs(4727) <= not a;
    layer5_outputs(4728) <= 1'b0;
    layer5_outputs(4729) <= not a;
    layer5_outputs(4730) <= not (a and b);
    layer5_outputs(4731) <= b and not a;
    layer5_outputs(4732) <= not (a xor b);
    layer5_outputs(4733) <= b and not a;
    layer5_outputs(4734) <= b;
    layer5_outputs(4735) <= a xor b;
    layer5_outputs(4736) <= not (a and b);
    layer5_outputs(4737) <= a or b;
    layer5_outputs(4738) <= not (a or b);
    layer5_outputs(4739) <= not (a or b);
    layer5_outputs(4740) <= not (a or b);
    layer5_outputs(4741) <= b and not a;
    layer5_outputs(4742) <= a and b;
    layer5_outputs(4743) <= not a or b;
    layer5_outputs(4744) <= b and not a;
    layer5_outputs(4745) <= b and not a;
    layer5_outputs(4746) <= not a;
    layer5_outputs(4747) <= a;
    layer5_outputs(4748) <= b and not a;
    layer5_outputs(4749) <= not (a and b);
    layer5_outputs(4750) <= b and not a;
    layer5_outputs(4751) <= not a;
    layer5_outputs(4752) <= not a;
    layer5_outputs(4753) <= b;
    layer5_outputs(4754) <= b and not a;
    layer5_outputs(4755) <= not a;
    layer5_outputs(4756) <= not (a xor b);
    layer5_outputs(4757) <= b;
    layer5_outputs(4758) <= b;
    layer5_outputs(4759) <= not b;
    layer5_outputs(4760) <= not (a xor b);
    layer5_outputs(4761) <= a or b;
    layer5_outputs(4762) <= not (a and b);
    layer5_outputs(4763) <= a xor b;
    layer5_outputs(4764) <= not a;
    layer5_outputs(4765) <= a or b;
    layer5_outputs(4766) <= a;
    layer5_outputs(4767) <= not b;
    layer5_outputs(4768) <= a;
    layer5_outputs(4769) <= a or b;
    layer5_outputs(4770) <= b;
    layer5_outputs(4771) <= not b or a;
    layer5_outputs(4772) <= 1'b0;
    layer5_outputs(4773) <= b;
    layer5_outputs(4774) <= 1'b0;
    layer5_outputs(4775) <= not b;
    layer5_outputs(4776) <= not b;
    layer5_outputs(4777) <= a;
    layer5_outputs(4778) <= not b or a;
    layer5_outputs(4779) <= not a;
    layer5_outputs(4780) <= not (a and b);
    layer5_outputs(4781) <= a and b;
    layer5_outputs(4782) <= not b;
    layer5_outputs(4783) <= b;
    layer5_outputs(4784) <= b;
    layer5_outputs(4785) <= not (a or b);
    layer5_outputs(4786) <= not b or a;
    layer5_outputs(4787) <= not (a and b);
    layer5_outputs(4788) <= not (a xor b);
    layer5_outputs(4789) <= 1'b0;
    layer5_outputs(4790) <= 1'b0;
    layer5_outputs(4791) <= not b;
    layer5_outputs(4792) <= b;
    layer5_outputs(4793) <= not a;
    layer5_outputs(4794) <= not (a and b);
    layer5_outputs(4795) <= not a or b;
    layer5_outputs(4796) <= not (a or b);
    layer5_outputs(4797) <= not a;
    layer5_outputs(4798) <= not a;
    layer5_outputs(4799) <= a;
    layer5_outputs(4800) <= not b;
    layer5_outputs(4801) <= b;
    layer5_outputs(4802) <= not a or b;
    layer5_outputs(4803) <= 1'b0;
    layer5_outputs(4804) <= not (a and b);
    layer5_outputs(4805) <= b and not a;
    layer5_outputs(4806) <= b and not a;
    layer5_outputs(4807) <= not (a xor b);
    layer5_outputs(4808) <= not b;
    layer5_outputs(4809) <= not (a and b);
    layer5_outputs(4810) <= a;
    layer5_outputs(4811) <= not a;
    layer5_outputs(4812) <= not b;
    layer5_outputs(4813) <= a and not b;
    layer5_outputs(4814) <= not b or a;
    layer5_outputs(4815) <= a xor b;
    layer5_outputs(4816) <= b and not a;
    layer5_outputs(4817) <= 1'b1;
    layer5_outputs(4818) <= b and not a;
    layer5_outputs(4819) <= a and not b;
    layer5_outputs(4820) <= not b;
    layer5_outputs(4821) <= b;
    layer5_outputs(4822) <= not (a xor b);
    layer5_outputs(4823) <= not b;
    layer5_outputs(4824) <= not (a or b);
    layer5_outputs(4825) <= a xor b;
    layer5_outputs(4826) <= not a or b;
    layer5_outputs(4827) <= not a or b;
    layer5_outputs(4828) <= not a;
    layer5_outputs(4829) <= a;
    layer5_outputs(4830) <= not (a xor b);
    layer5_outputs(4831) <= not (a and b);
    layer5_outputs(4832) <= not (a and b);
    layer5_outputs(4833) <= not (a and b);
    layer5_outputs(4834) <= a and b;
    layer5_outputs(4835) <= a;
    layer5_outputs(4836) <= b;
    layer5_outputs(4837) <= 1'b0;
    layer5_outputs(4838) <= not (a xor b);
    layer5_outputs(4839) <= a or b;
    layer5_outputs(4840) <= a and not b;
    layer5_outputs(4841) <= a;
    layer5_outputs(4842) <= not (a xor b);
    layer5_outputs(4843) <= a;
    layer5_outputs(4844) <= b and not a;
    layer5_outputs(4845) <= not b;
    layer5_outputs(4846) <= not a;
    layer5_outputs(4847) <= 1'b1;
    layer5_outputs(4848) <= a;
    layer5_outputs(4849) <= not b or a;
    layer5_outputs(4850) <= a and not b;
    layer5_outputs(4851) <= a xor b;
    layer5_outputs(4852) <= not (a or b);
    layer5_outputs(4853) <= not (a xor b);
    layer5_outputs(4854) <= not b;
    layer5_outputs(4855) <= not a;
    layer5_outputs(4856) <= not b or a;
    layer5_outputs(4857) <= not b or a;
    layer5_outputs(4858) <= not b;
    layer5_outputs(4859) <= a;
    layer5_outputs(4860) <= a and b;
    layer5_outputs(4861) <= a and b;
    layer5_outputs(4862) <= a and not b;
    layer5_outputs(4863) <= b and not a;
    layer5_outputs(4864) <= b and not a;
    layer5_outputs(4865) <= not a or b;
    layer5_outputs(4866) <= not a;
    layer5_outputs(4867) <= 1'b0;
    layer5_outputs(4868) <= a or b;
    layer5_outputs(4869) <= not b or a;
    layer5_outputs(4870) <= 1'b0;
    layer5_outputs(4871) <= a and b;
    layer5_outputs(4872) <= not b;
    layer5_outputs(4873) <= b;
    layer5_outputs(4874) <= a or b;
    layer5_outputs(4875) <= a xor b;
    layer5_outputs(4876) <= not a;
    layer5_outputs(4877) <= b;
    layer5_outputs(4878) <= not b;
    layer5_outputs(4879) <= not (a and b);
    layer5_outputs(4880) <= not (a and b);
    layer5_outputs(4881) <= not (a xor b);
    layer5_outputs(4882) <= not (a xor b);
    layer5_outputs(4883) <= 1'b0;
    layer5_outputs(4884) <= not (a and b);
    layer5_outputs(4885) <= a or b;
    layer5_outputs(4886) <= not b or a;
    layer5_outputs(4887) <= not (a or b);
    layer5_outputs(4888) <= not (a xor b);
    layer5_outputs(4889) <= not b or a;
    layer5_outputs(4890) <= b;
    layer5_outputs(4891) <= not b;
    layer5_outputs(4892) <= a;
    layer5_outputs(4893) <= 1'b1;
    layer5_outputs(4894) <= b;
    layer5_outputs(4895) <= b and not a;
    layer5_outputs(4896) <= not a or b;
    layer5_outputs(4897) <= b;
    layer5_outputs(4898) <= not a;
    layer5_outputs(4899) <= not (a and b);
    layer5_outputs(4900) <= a;
    layer5_outputs(4901) <= b and not a;
    layer5_outputs(4902) <= not (a or b);
    layer5_outputs(4903) <= 1'b0;
    layer5_outputs(4904) <= not a;
    layer5_outputs(4905) <= not a;
    layer5_outputs(4906) <= a and not b;
    layer5_outputs(4907) <= a or b;
    layer5_outputs(4908) <= 1'b1;
    layer5_outputs(4909) <= b and not a;
    layer5_outputs(4910) <= not a;
    layer5_outputs(4911) <= not a or b;
    layer5_outputs(4912) <= b and not a;
    layer5_outputs(4913) <= 1'b0;
    layer5_outputs(4914) <= a;
    layer5_outputs(4915) <= not (a or b);
    layer5_outputs(4916) <= not a;
    layer5_outputs(4917) <= b and not a;
    layer5_outputs(4918) <= not a or b;
    layer5_outputs(4919) <= not a or b;
    layer5_outputs(4920) <= a;
    layer5_outputs(4921) <= a or b;
    layer5_outputs(4922) <= not b;
    layer5_outputs(4923) <= not a;
    layer5_outputs(4924) <= not a;
    layer5_outputs(4925) <= b and not a;
    layer5_outputs(4926) <= a and b;
    layer5_outputs(4927) <= b;
    layer5_outputs(4928) <= not b;
    layer5_outputs(4929) <= not a or b;
    layer5_outputs(4930) <= a and b;
    layer5_outputs(4931) <= b;
    layer5_outputs(4932) <= b;
    layer5_outputs(4933) <= b;
    layer5_outputs(4934) <= not (a and b);
    layer5_outputs(4935) <= not b;
    layer5_outputs(4936) <= b;
    layer5_outputs(4937) <= a;
    layer5_outputs(4938) <= a and not b;
    layer5_outputs(4939) <= not (a xor b);
    layer5_outputs(4940) <= not (a or b);
    layer5_outputs(4941) <= not (a or b);
    layer5_outputs(4942) <= not a;
    layer5_outputs(4943) <= b;
    layer5_outputs(4944) <= not a or b;
    layer5_outputs(4945) <= not a;
    layer5_outputs(4946) <= a and not b;
    layer5_outputs(4947) <= not a or b;
    layer5_outputs(4948) <= not b;
    layer5_outputs(4949) <= not (a or b);
    layer5_outputs(4950) <= a xor b;
    layer5_outputs(4951) <= not b;
    layer5_outputs(4952) <= a;
    layer5_outputs(4953) <= b and not a;
    layer5_outputs(4954) <= not b;
    layer5_outputs(4955) <= not a or b;
    layer5_outputs(4956) <= a;
    layer5_outputs(4957) <= a and not b;
    layer5_outputs(4958) <= 1'b0;
    layer5_outputs(4959) <= a;
    layer5_outputs(4960) <= not (a xor b);
    layer5_outputs(4961) <= not a;
    layer5_outputs(4962) <= not (a and b);
    layer5_outputs(4963) <= not a;
    layer5_outputs(4964) <= not (a and b);
    layer5_outputs(4965) <= b;
    layer5_outputs(4966) <= b and not a;
    layer5_outputs(4967) <= not a;
    layer5_outputs(4968) <= a;
    layer5_outputs(4969) <= not a;
    layer5_outputs(4970) <= a;
    layer5_outputs(4971) <= not b;
    layer5_outputs(4972) <= b and not a;
    layer5_outputs(4973) <= not (a or b);
    layer5_outputs(4974) <= b;
    layer5_outputs(4975) <= b and not a;
    layer5_outputs(4976) <= not (a xor b);
    layer5_outputs(4977) <= not a;
    layer5_outputs(4978) <= b and not a;
    layer5_outputs(4979) <= b and not a;
    layer5_outputs(4980) <= not (a and b);
    layer5_outputs(4981) <= b;
    layer5_outputs(4982) <= 1'b0;
    layer5_outputs(4983) <= not a or b;
    layer5_outputs(4984) <= a and not b;
    layer5_outputs(4985) <= a;
    layer5_outputs(4986) <= b;
    layer5_outputs(4987) <= a;
    layer5_outputs(4988) <= a or b;
    layer5_outputs(4989) <= a;
    layer5_outputs(4990) <= a xor b;
    layer5_outputs(4991) <= not (a and b);
    layer5_outputs(4992) <= a;
    layer5_outputs(4993) <= not (a and b);
    layer5_outputs(4994) <= not (a or b);
    layer5_outputs(4995) <= a;
    layer5_outputs(4996) <= not b;
    layer5_outputs(4997) <= a and not b;
    layer5_outputs(4998) <= a;
    layer5_outputs(4999) <= not b or a;
    layer5_outputs(5000) <= a;
    layer5_outputs(5001) <= b;
    layer5_outputs(5002) <= not b or a;
    layer5_outputs(5003) <= 1'b1;
    layer5_outputs(5004) <= not a;
    layer5_outputs(5005) <= a xor b;
    layer5_outputs(5006) <= 1'b1;
    layer5_outputs(5007) <= a xor b;
    layer5_outputs(5008) <= not b or a;
    layer5_outputs(5009) <= 1'b1;
    layer5_outputs(5010) <= not (a and b);
    layer5_outputs(5011) <= a xor b;
    layer5_outputs(5012) <= not a or b;
    layer5_outputs(5013) <= b and not a;
    layer5_outputs(5014) <= not a;
    layer5_outputs(5015) <= not a or b;
    layer5_outputs(5016) <= not a or b;
    layer5_outputs(5017) <= not a;
    layer5_outputs(5018) <= a xor b;
    layer5_outputs(5019) <= not (a and b);
    layer5_outputs(5020) <= not (a or b);
    layer5_outputs(5021) <= b;
    layer5_outputs(5022) <= not b;
    layer5_outputs(5023) <= a;
    layer5_outputs(5024) <= not b;
    layer5_outputs(5025) <= not b;
    layer5_outputs(5026) <= not (a or b);
    layer5_outputs(5027) <= not b;
    layer5_outputs(5028) <= b;
    layer5_outputs(5029) <= not (a and b);
    layer5_outputs(5030) <= a;
    layer5_outputs(5031) <= not (a xor b);
    layer5_outputs(5032) <= not a or b;
    layer5_outputs(5033) <= not (a or b);
    layer5_outputs(5034) <= a and b;
    layer5_outputs(5035) <= b;
    layer5_outputs(5036) <= b and not a;
    layer5_outputs(5037) <= b;
    layer5_outputs(5038) <= a or b;
    layer5_outputs(5039) <= a xor b;
    layer5_outputs(5040) <= a and b;
    layer5_outputs(5041) <= 1'b0;
    layer5_outputs(5042) <= a and not b;
    layer5_outputs(5043) <= a or b;
    layer5_outputs(5044) <= 1'b1;
    layer5_outputs(5045) <= a and not b;
    layer5_outputs(5046) <= not (a or b);
    layer5_outputs(5047) <= not (a and b);
    layer5_outputs(5048) <= a and not b;
    layer5_outputs(5049) <= a or b;
    layer5_outputs(5050) <= not (a xor b);
    layer5_outputs(5051) <= not (a xor b);
    layer5_outputs(5052) <= not a;
    layer5_outputs(5053) <= a;
    layer5_outputs(5054) <= a xor b;
    layer5_outputs(5055) <= not a;
    layer5_outputs(5056) <= b and not a;
    layer5_outputs(5057) <= not (a xor b);
    layer5_outputs(5058) <= not (a or b);
    layer5_outputs(5059) <= not a;
    layer5_outputs(5060) <= b;
    layer5_outputs(5061) <= not b or a;
    layer5_outputs(5062) <= not a;
    layer5_outputs(5063) <= 1'b0;
    layer5_outputs(5064) <= b;
    layer5_outputs(5065) <= not a or b;
    layer5_outputs(5066) <= a or b;
    layer5_outputs(5067) <= b;
    layer5_outputs(5068) <= b;
    layer5_outputs(5069) <= not (a or b);
    layer5_outputs(5070) <= not a;
    layer5_outputs(5071) <= not a;
    layer5_outputs(5072) <= not a or b;
    layer5_outputs(5073) <= not a;
    layer5_outputs(5074) <= a or b;
    layer5_outputs(5075) <= 1'b0;
    layer5_outputs(5076) <= b and not a;
    layer5_outputs(5077) <= a xor b;
    layer5_outputs(5078) <= a;
    layer5_outputs(5079) <= 1'b0;
    layer5_outputs(5080) <= not (a xor b);
    layer5_outputs(5081) <= b;
    layer5_outputs(5082) <= a or b;
    layer5_outputs(5083) <= b and not a;
    layer5_outputs(5084) <= not b or a;
    layer5_outputs(5085) <= b and not a;
    layer5_outputs(5086) <= not a;
    layer5_outputs(5087) <= not (a xor b);
    layer5_outputs(5088) <= b;
    layer5_outputs(5089) <= not (a or b);
    layer5_outputs(5090) <= b;
    layer5_outputs(5091) <= a;
    layer5_outputs(5092) <= not b or a;
    layer5_outputs(5093) <= 1'b0;
    layer5_outputs(5094) <= not (a xor b);
    layer5_outputs(5095) <= not a;
    layer5_outputs(5096) <= not b or a;
    layer5_outputs(5097) <= 1'b1;
    layer5_outputs(5098) <= a;
    layer5_outputs(5099) <= b and not a;
    layer5_outputs(5100) <= b and not a;
    layer5_outputs(5101) <= not (a or b);
    layer5_outputs(5102) <= b;
    layer5_outputs(5103) <= b and not a;
    layer5_outputs(5104) <= a xor b;
    layer5_outputs(5105) <= not b;
    layer5_outputs(5106) <= a and not b;
    layer5_outputs(5107) <= 1'b1;
    layer5_outputs(5108) <= not a;
    layer5_outputs(5109) <= b and not a;
    layer5_outputs(5110) <= not b;
    layer5_outputs(5111) <= a;
    layer5_outputs(5112) <= a and b;
    layer5_outputs(5113) <= not a;
    layer5_outputs(5114) <= a or b;
    layer5_outputs(5115) <= a and b;
    layer5_outputs(5116) <= a and b;
    layer5_outputs(5117) <= not b or a;
    layer5_outputs(5118) <= 1'b0;
    layer5_outputs(5119) <= a and b;
    layer5_outputs(5120) <= not a;
    layer5_outputs(5121) <= b;
    layer5_outputs(5122) <= not a;
    layer5_outputs(5123) <= a and b;
    layer5_outputs(5124) <= not a;
    layer5_outputs(5125) <= 1'b0;
    layer5_outputs(5126) <= not a;
    layer5_outputs(5127) <= a and b;
    layer5_outputs(5128) <= not b;
    layer5_outputs(5129) <= 1'b1;
    layer5_outputs(5130) <= not a or b;
    layer5_outputs(5131) <= a and not b;
    layer5_outputs(5132) <= a;
    layer5_outputs(5133) <= a or b;
    layer5_outputs(5134) <= b;
    layer5_outputs(5135) <= a and not b;
    layer5_outputs(5136) <= not b;
    layer5_outputs(5137) <= not b;
    layer5_outputs(5138) <= b;
    layer5_outputs(5139) <= b;
    layer5_outputs(5140) <= not a or b;
    layer5_outputs(5141) <= not (a or b);
    layer5_outputs(5142) <= not b or a;
    layer5_outputs(5143) <= a;
    layer5_outputs(5144) <= b;
    layer5_outputs(5145) <= b and not a;
    layer5_outputs(5146) <= not (a and b);
    layer5_outputs(5147) <= not (a and b);
    layer5_outputs(5148) <= a;
    layer5_outputs(5149) <= not a;
    layer5_outputs(5150) <= not a or b;
    layer5_outputs(5151) <= not (a or b);
    layer5_outputs(5152) <= not a;
    layer5_outputs(5153) <= not (a or b);
    layer5_outputs(5154) <= a or b;
    layer5_outputs(5155) <= not a;
    layer5_outputs(5156) <= not a or b;
    layer5_outputs(5157) <= a;
    layer5_outputs(5158) <= not b;
    layer5_outputs(5159) <= a and not b;
    layer5_outputs(5160) <= a or b;
    layer5_outputs(5161) <= b;
    layer5_outputs(5162) <= a;
    layer5_outputs(5163) <= a and b;
    layer5_outputs(5164) <= not a or b;
    layer5_outputs(5165) <= not a or b;
    layer5_outputs(5166) <= a and not b;
    layer5_outputs(5167) <= not a;
    layer5_outputs(5168) <= not a;
    layer5_outputs(5169) <= a;
    layer5_outputs(5170) <= a and not b;
    layer5_outputs(5171) <= a and b;
    layer5_outputs(5172) <= b and not a;
    layer5_outputs(5173) <= not a or b;
    layer5_outputs(5174) <= not a;
    layer5_outputs(5175) <= not (a or b);
    layer5_outputs(5176) <= a or b;
    layer5_outputs(5177) <= a and not b;
    layer5_outputs(5178) <= not (a xor b);
    layer5_outputs(5179) <= not b or a;
    layer5_outputs(5180) <= b;
    layer5_outputs(5181) <= a and not b;
    layer5_outputs(5182) <= a and not b;
    layer5_outputs(5183) <= not (a xor b);
    layer5_outputs(5184) <= not (a xor b);
    layer5_outputs(5185) <= a or b;
    layer5_outputs(5186) <= not b;
    layer5_outputs(5187) <= a;
    layer5_outputs(5188) <= 1'b1;
    layer5_outputs(5189) <= not a;
    layer5_outputs(5190) <= not (a or b);
    layer5_outputs(5191) <= not a;
    layer5_outputs(5192) <= 1'b1;
    layer5_outputs(5193) <= not b;
    layer5_outputs(5194) <= b and not a;
    layer5_outputs(5195) <= not b or a;
    layer5_outputs(5196) <= 1'b0;
    layer5_outputs(5197) <= not a or b;
    layer5_outputs(5198) <= not b;
    layer5_outputs(5199) <= a and b;
    layer5_outputs(5200) <= a;
    layer5_outputs(5201) <= not (a xor b);
    layer5_outputs(5202) <= not a;
    layer5_outputs(5203) <= a xor b;
    layer5_outputs(5204) <= not b;
    layer5_outputs(5205) <= not a or b;
    layer5_outputs(5206) <= b;
    layer5_outputs(5207) <= b and not a;
    layer5_outputs(5208) <= b;
    layer5_outputs(5209) <= b;
    layer5_outputs(5210) <= not a;
    layer5_outputs(5211) <= not (a or b);
    layer5_outputs(5212) <= b;
    layer5_outputs(5213) <= a or b;
    layer5_outputs(5214) <= not a;
    layer5_outputs(5215) <= b;
    layer5_outputs(5216) <= not (a xor b);
    layer5_outputs(5217) <= not a or b;
    layer5_outputs(5218) <= a xor b;
    layer5_outputs(5219) <= not (a and b);
    layer5_outputs(5220) <= a and not b;
    layer5_outputs(5221) <= 1'b0;
    layer5_outputs(5222) <= b and not a;
    layer5_outputs(5223) <= b;
    layer5_outputs(5224) <= a;
    layer5_outputs(5225) <= a xor b;
    layer5_outputs(5226) <= a;
    layer5_outputs(5227) <= not (a and b);
    layer5_outputs(5228) <= not b;
    layer5_outputs(5229) <= not (a or b);
    layer5_outputs(5230) <= a;
    layer5_outputs(5231) <= not b or a;
    layer5_outputs(5232) <= b and not a;
    layer5_outputs(5233) <= not a or b;
    layer5_outputs(5234) <= not a;
    layer5_outputs(5235) <= not a or b;
    layer5_outputs(5236) <= not (a and b);
    layer5_outputs(5237) <= b;
    layer5_outputs(5238) <= b and not a;
    layer5_outputs(5239) <= b;
    layer5_outputs(5240) <= a and b;
    layer5_outputs(5241) <= not b;
    layer5_outputs(5242) <= b;
    layer5_outputs(5243) <= not (a or b);
    layer5_outputs(5244) <= not b;
    layer5_outputs(5245) <= a and not b;
    layer5_outputs(5246) <= not b;
    layer5_outputs(5247) <= a;
    layer5_outputs(5248) <= not (a and b);
    layer5_outputs(5249) <= not b;
    layer5_outputs(5250) <= not a;
    layer5_outputs(5251) <= not (a or b);
    layer5_outputs(5252) <= a and not b;
    layer5_outputs(5253) <= b;
    layer5_outputs(5254) <= a xor b;
    layer5_outputs(5255) <= a;
    layer5_outputs(5256) <= b;
    layer5_outputs(5257) <= not a;
    layer5_outputs(5258) <= a or b;
    layer5_outputs(5259) <= not a;
    layer5_outputs(5260) <= not (a xor b);
    layer5_outputs(5261) <= not (a and b);
    layer5_outputs(5262) <= a and b;
    layer5_outputs(5263) <= a or b;
    layer5_outputs(5264) <= not a;
    layer5_outputs(5265) <= a and not b;
    layer5_outputs(5266) <= not (a or b);
    layer5_outputs(5267) <= a and b;
    layer5_outputs(5268) <= 1'b0;
    layer5_outputs(5269) <= not (a or b);
    layer5_outputs(5270) <= b and not a;
    layer5_outputs(5271) <= not b or a;
    layer5_outputs(5272) <= a and not b;
    layer5_outputs(5273) <= 1'b0;
    layer5_outputs(5274) <= a;
    layer5_outputs(5275) <= not (a or b);
    layer5_outputs(5276) <= b;
    layer5_outputs(5277) <= not (a and b);
    layer5_outputs(5278) <= a and not b;
    layer5_outputs(5279) <= not (a and b);
    layer5_outputs(5280) <= not a or b;
    layer5_outputs(5281) <= not a;
    layer5_outputs(5282) <= not b or a;
    layer5_outputs(5283) <= not a or b;
    layer5_outputs(5284) <= a and not b;
    layer5_outputs(5285) <= not b;
    layer5_outputs(5286) <= 1'b1;
    layer5_outputs(5287) <= a or b;
    layer5_outputs(5288) <= not a or b;
    layer5_outputs(5289) <= not b;
    layer5_outputs(5290) <= not b or a;
    layer5_outputs(5291) <= not b;
    layer5_outputs(5292) <= a and not b;
    layer5_outputs(5293) <= a;
    layer5_outputs(5294) <= a xor b;
    layer5_outputs(5295) <= not a or b;
    layer5_outputs(5296) <= not b;
    layer5_outputs(5297) <= not (a xor b);
    layer5_outputs(5298) <= a;
    layer5_outputs(5299) <= not (a xor b);
    layer5_outputs(5300) <= a and b;
    layer5_outputs(5301) <= not (a or b);
    layer5_outputs(5302) <= not b;
    layer5_outputs(5303) <= not (a or b);
    layer5_outputs(5304) <= 1'b1;
    layer5_outputs(5305) <= not b;
    layer5_outputs(5306) <= a and not b;
    layer5_outputs(5307) <= a and not b;
    layer5_outputs(5308) <= a and not b;
    layer5_outputs(5309) <= not (a or b);
    layer5_outputs(5310) <= 1'b1;
    layer5_outputs(5311) <= not b;
    layer5_outputs(5312) <= 1'b0;
    layer5_outputs(5313) <= not a;
    layer5_outputs(5314) <= a or b;
    layer5_outputs(5315) <= a xor b;
    layer5_outputs(5316) <= a;
    layer5_outputs(5317) <= a and b;
    layer5_outputs(5318) <= a and b;
    layer5_outputs(5319) <= 1'b1;
    layer5_outputs(5320) <= b;
    layer5_outputs(5321) <= not (a xor b);
    layer5_outputs(5322) <= a;
    layer5_outputs(5323) <= a and not b;
    layer5_outputs(5324) <= b;
    layer5_outputs(5325) <= a and not b;
    layer5_outputs(5326) <= a and b;
    layer5_outputs(5327) <= a and not b;
    layer5_outputs(5328) <= not (a or b);
    layer5_outputs(5329) <= 1'b0;
    layer5_outputs(5330) <= not b or a;
    layer5_outputs(5331) <= not (a or b);
    layer5_outputs(5332) <= a and not b;
    layer5_outputs(5333) <= a;
    layer5_outputs(5334) <= a;
    layer5_outputs(5335) <= not a or b;
    layer5_outputs(5336) <= a and b;
    layer5_outputs(5337) <= a;
    layer5_outputs(5338) <= a or b;
    layer5_outputs(5339) <= not (a or b);
    layer5_outputs(5340) <= b;
    layer5_outputs(5341) <= a or b;
    layer5_outputs(5342) <= not a;
    layer5_outputs(5343) <= a;
    layer5_outputs(5344) <= not a;
    layer5_outputs(5345) <= a;
    layer5_outputs(5346) <= a and b;
    layer5_outputs(5347) <= b and not a;
    layer5_outputs(5348) <= a;
    layer5_outputs(5349) <= not a or b;
    layer5_outputs(5350) <= not (a or b);
    layer5_outputs(5351) <= a xor b;
    layer5_outputs(5352) <= not a;
    layer5_outputs(5353) <= not a or b;
    layer5_outputs(5354) <= not (a or b);
    layer5_outputs(5355) <= a or b;
    layer5_outputs(5356) <= b and not a;
    layer5_outputs(5357) <= a or b;
    layer5_outputs(5358) <= 1'b1;
    layer5_outputs(5359) <= 1'b0;
    layer5_outputs(5360) <= b;
    layer5_outputs(5361) <= not a;
    layer5_outputs(5362) <= b and not a;
    layer5_outputs(5363) <= not b;
    layer5_outputs(5364) <= b;
    layer5_outputs(5365) <= b and not a;
    layer5_outputs(5366) <= a and not b;
    layer5_outputs(5367) <= a xor b;
    layer5_outputs(5368) <= b;
    layer5_outputs(5369) <= b;
    layer5_outputs(5370) <= not a;
    layer5_outputs(5371) <= not b;
    layer5_outputs(5372) <= not (a or b);
    layer5_outputs(5373) <= not b;
    layer5_outputs(5374) <= not (a and b);
    layer5_outputs(5375) <= not b or a;
    layer5_outputs(5376) <= b;
    layer5_outputs(5377) <= a;
    layer5_outputs(5378) <= not (a xor b);
    layer5_outputs(5379) <= a or b;
    layer5_outputs(5380) <= b and not a;
    layer5_outputs(5381) <= 1'b0;
    layer5_outputs(5382) <= a;
    layer5_outputs(5383) <= 1'b0;
    layer5_outputs(5384) <= a;
    layer5_outputs(5385) <= a or b;
    layer5_outputs(5386) <= a or b;
    layer5_outputs(5387) <= not (a xor b);
    layer5_outputs(5388) <= b and not a;
    layer5_outputs(5389) <= not b;
    layer5_outputs(5390) <= not (a or b);
    layer5_outputs(5391) <= not (a and b);
    layer5_outputs(5392) <= not b;
    layer5_outputs(5393) <= a and not b;
    layer5_outputs(5394) <= a;
    layer5_outputs(5395) <= a and not b;
    layer5_outputs(5396) <= a or b;
    layer5_outputs(5397) <= b and not a;
    layer5_outputs(5398) <= b;
    layer5_outputs(5399) <= not (a or b);
    layer5_outputs(5400) <= a and not b;
    layer5_outputs(5401) <= not b or a;
    layer5_outputs(5402) <= not (a xor b);
    layer5_outputs(5403) <= not b;
    layer5_outputs(5404) <= not (a and b);
    layer5_outputs(5405) <= a;
    layer5_outputs(5406) <= a;
    layer5_outputs(5407) <= a and b;
    layer5_outputs(5408) <= b;
    layer5_outputs(5409) <= not (a and b);
    layer5_outputs(5410) <= a or b;
    layer5_outputs(5411) <= 1'b0;
    layer5_outputs(5412) <= not a or b;
    layer5_outputs(5413) <= not a;
    layer5_outputs(5414) <= b and not a;
    layer5_outputs(5415) <= not a;
    layer5_outputs(5416) <= not b;
    layer5_outputs(5417) <= not (a and b);
    layer5_outputs(5418) <= b;
    layer5_outputs(5419) <= b and not a;
    layer5_outputs(5420) <= b;
    layer5_outputs(5421) <= not (a and b);
    layer5_outputs(5422) <= not b;
    layer5_outputs(5423) <= not (a and b);
    layer5_outputs(5424) <= 1'b1;
    layer5_outputs(5425) <= not (a or b);
    layer5_outputs(5426) <= a and not b;
    layer5_outputs(5427) <= not b;
    layer5_outputs(5428) <= b and not a;
    layer5_outputs(5429) <= 1'b1;
    layer5_outputs(5430) <= not b;
    layer5_outputs(5431) <= a xor b;
    layer5_outputs(5432) <= b;
    layer5_outputs(5433) <= a and b;
    layer5_outputs(5434) <= not a or b;
    layer5_outputs(5435) <= b and not a;
    layer5_outputs(5436) <= not a;
    layer5_outputs(5437) <= not b or a;
    layer5_outputs(5438) <= not (a or b);
    layer5_outputs(5439) <= not b;
    layer5_outputs(5440) <= a and b;
    layer5_outputs(5441) <= a and not b;
    layer5_outputs(5442) <= a;
    layer5_outputs(5443) <= a or b;
    layer5_outputs(5444) <= a and b;
    layer5_outputs(5445) <= not a or b;
    layer5_outputs(5446) <= not b;
    layer5_outputs(5447) <= not a;
    layer5_outputs(5448) <= a and b;
    layer5_outputs(5449) <= not b or a;
    layer5_outputs(5450) <= not b or a;
    layer5_outputs(5451) <= not a;
    layer5_outputs(5452) <= not b;
    layer5_outputs(5453) <= not a;
    layer5_outputs(5454) <= not a;
    layer5_outputs(5455) <= a;
    layer5_outputs(5456) <= b and not a;
    layer5_outputs(5457) <= a;
    layer5_outputs(5458) <= b;
    layer5_outputs(5459) <= not b;
    layer5_outputs(5460) <= a and not b;
    layer5_outputs(5461) <= a;
    layer5_outputs(5462) <= 1'b0;
    layer5_outputs(5463) <= not a;
    layer5_outputs(5464) <= a;
    layer5_outputs(5465) <= a and b;
    layer5_outputs(5466) <= a xor b;
    layer5_outputs(5467) <= not a;
    layer5_outputs(5468) <= a or b;
    layer5_outputs(5469) <= not b;
    layer5_outputs(5470) <= not a;
    layer5_outputs(5471) <= not a;
    layer5_outputs(5472) <= a;
    layer5_outputs(5473) <= not (a xor b);
    layer5_outputs(5474) <= not a or b;
    layer5_outputs(5475) <= b and not a;
    layer5_outputs(5476) <= not (a or b);
    layer5_outputs(5477) <= not (a and b);
    layer5_outputs(5478) <= a xor b;
    layer5_outputs(5479) <= not b;
    layer5_outputs(5480) <= not a;
    layer5_outputs(5481) <= not b or a;
    layer5_outputs(5482) <= not a;
    layer5_outputs(5483) <= a xor b;
    layer5_outputs(5484) <= not a;
    layer5_outputs(5485) <= not (a or b);
    layer5_outputs(5486) <= not a;
    layer5_outputs(5487) <= not (a or b);
    layer5_outputs(5488) <= not b;
    layer5_outputs(5489) <= b;
    layer5_outputs(5490) <= 1'b1;
    layer5_outputs(5491) <= not a;
    layer5_outputs(5492) <= a;
    layer5_outputs(5493) <= not b;
    layer5_outputs(5494) <= not b;
    layer5_outputs(5495) <= not b or a;
    layer5_outputs(5496) <= a and not b;
    layer5_outputs(5497) <= not (a or b);
    layer5_outputs(5498) <= a and b;
    layer5_outputs(5499) <= not a;
    layer5_outputs(5500) <= b and not a;
    layer5_outputs(5501) <= a xor b;
    layer5_outputs(5502) <= not a or b;
    layer5_outputs(5503) <= b;
    layer5_outputs(5504) <= a and not b;
    layer5_outputs(5505) <= not (a or b);
    layer5_outputs(5506) <= not a or b;
    layer5_outputs(5507) <= a;
    layer5_outputs(5508) <= b;
    layer5_outputs(5509) <= a xor b;
    layer5_outputs(5510) <= 1'b0;
    layer5_outputs(5511) <= not b;
    layer5_outputs(5512) <= a or b;
    layer5_outputs(5513) <= b;
    layer5_outputs(5514) <= not (a and b);
    layer5_outputs(5515) <= a;
    layer5_outputs(5516) <= a or b;
    layer5_outputs(5517) <= a and b;
    layer5_outputs(5518) <= a;
    layer5_outputs(5519) <= 1'b0;
    layer5_outputs(5520) <= not (a and b);
    layer5_outputs(5521) <= not (a and b);
    layer5_outputs(5522) <= not a or b;
    layer5_outputs(5523) <= b and not a;
    layer5_outputs(5524) <= b and not a;
    layer5_outputs(5525) <= a or b;
    layer5_outputs(5526) <= a and b;
    layer5_outputs(5527) <= a or b;
    layer5_outputs(5528) <= not a;
    layer5_outputs(5529) <= not b;
    layer5_outputs(5530) <= not (a or b);
    layer5_outputs(5531) <= a or b;
    layer5_outputs(5532) <= not (a xor b);
    layer5_outputs(5533) <= a xor b;
    layer5_outputs(5534) <= not a;
    layer5_outputs(5535) <= a or b;
    layer5_outputs(5536) <= not (a or b);
    layer5_outputs(5537) <= not b or a;
    layer5_outputs(5538) <= 1'b0;
    layer5_outputs(5539) <= b and not a;
    layer5_outputs(5540) <= a;
    layer5_outputs(5541) <= b and not a;
    layer5_outputs(5542) <= not (a or b);
    layer5_outputs(5543) <= not b;
    layer5_outputs(5544) <= 1'b0;
    layer5_outputs(5545) <= a xor b;
    layer5_outputs(5546) <= 1'b0;
    layer5_outputs(5547) <= a and not b;
    layer5_outputs(5548) <= a xor b;
    layer5_outputs(5549) <= b;
    layer5_outputs(5550) <= a;
    layer5_outputs(5551) <= a and b;
    layer5_outputs(5552) <= not b;
    layer5_outputs(5553) <= not b;
    layer5_outputs(5554) <= not (a or b);
    layer5_outputs(5555) <= b and not a;
    layer5_outputs(5556) <= a and not b;
    layer5_outputs(5557) <= b;
    layer5_outputs(5558) <= a or b;
    layer5_outputs(5559) <= 1'b0;
    layer5_outputs(5560) <= not b;
    layer5_outputs(5561) <= a;
    layer5_outputs(5562) <= not b;
    layer5_outputs(5563) <= a or b;
    layer5_outputs(5564) <= a and b;
    layer5_outputs(5565) <= not b;
    layer5_outputs(5566) <= a or b;
    layer5_outputs(5567) <= a and b;
    layer5_outputs(5568) <= not b;
    layer5_outputs(5569) <= a and b;
    layer5_outputs(5570) <= a or b;
    layer5_outputs(5571) <= b and not a;
    layer5_outputs(5572) <= b and not a;
    layer5_outputs(5573) <= not (a or b);
    layer5_outputs(5574) <= b;
    layer5_outputs(5575) <= not (a and b);
    layer5_outputs(5576) <= not a;
    layer5_outputs(5577) <= not (a xor b);
    layer5_outputs(5578) <= b;
    layer5_outputs(5579) <= not b;
    layer5_outputs(5580) <= a and not b;
    layer5_outputs(5581) <= b and not a;
    layer5_outputs(5582) <= b;
    layer5_outputs(5583) <= not b;
    layer5_outputs(5584) <= not (a or b);
    layer5_outputs(5585) <= not (a and b);
    layer5_outputs(5586) <= a or b;
    layer5_outputs(5587) <= b;
    layer5_outputs(5588) <= not a or b;
    layer5_outputs(5589) <= not b or a;
    layer5_outputs(5590) <= b;
    layer5_outputs(5591) <= a and not b;
    layer5_outputs(5592) <= a;
    layer5_outputs(5593) <= b;
    layer5_outputs(5594) <= a xor b;
    layer5_outputs(5595) <= a or b;
    layer5_outputs(5596) <= b;
    layer5_outputs(5597) <= a and b;
    layer5_outputs(5598) <= b;
    layer5_outputs(5599) <= b and not a;
    layer5_outputs(5600) <= not a;
    layer5_outputs(5601) <= a or b;
    layer5_outputs(5602) <= a;
    layer5_outputs(5603) <= b;
    layer5_outputs(5604) <= a and b;
    layer5_outputs(5605) <= not b or a;
    layer5_outputs(5606) <= not (a and b);
    layer5_outputs(5607) <= a xor b;
    layer5_outputs(5608) <= 1'b0;
    layer5_outputs(5609) <= not (a and b);
    layer5_outputs(5610) <= not (a xor b);
    layer5_outputs(5611) <= b;
    layer5_outputs(5612) <= not a;
    layer5_outputs(5613) <= b and not a;
    layer5_outputs(5614) <= not b or a;
    layer5_outputs(5615) <= a or b;
    layer5_outputs(5616) <= not (a xor b);
    layer5_outputs(5617) <= a and b;
    layer5_outputs(5618) <= b;
    layer5_outputs(5619) <= 1'b1;
    layer5_outputs(5620) <= not a;
    layer5_outputs(5621) <= not (a or b);
    layer5_outputs(5622) <= a and b;
    layer5_outputs(5623) <= not b;
    layer5_outputs(5624) <= not b;
    layer5_outputs(5625) <= not a;
    layer5_outputs(5626) <= not (a or b);
    layer5_outputs(5627) <= not a or b;
    layer5_outputs(5628) <= b;
    layer5_outputs(5629) <= a and b;
    layer5_outputs(5630) <= 1'b1;
    layer5_outputs(5631) <= not a;
    layer5_outputs(5632) <= not (a and b);
    layer5_outputs(5633) <= a xor b;
    layer5_outputs(5634) <= 1'b0;
    layer5_outputs(5635) <= b and not a;
    layer5_outputs(5636) <= a and not b;
    layer5_outputs(5637) <= b;
    layer5_outputs(5638) <= a and b;
    layer5_outputs(5639) <= 1'b0;
    layer5_outputs(5640) <= b;
    layer5_outputs(5641) <= b and not a;
    layer5_outputs(5642) <= a;
    layer5_outputs(5643) <= not a;
    layer5_outputs(5644) <= a and not b;
    layer5_outputs(5645) <= not (a and b);
    layer5_outputs(5646) <= a xor b;
    layer5_outputs(5647) <= not (a and b);
    layer5_outputs(5648) <= a or b;
    layer5_outputs(5649) <= b;
    layer5_outputs(5650) <= not (a and b);
    layer5_outputs(5651) <= b;
    layer5_outputs(5652) <= not b or a;
    layer5_outputs(5653) <= not b;
    layer5_outputs(5654) <= not a or b;
    layer5_outputs(5655) <= 1'b1;
    layer5_outputs(5656) <= a and not b;
    layer5_outputs(5657) <= not b or a;
    layer5_outputs(5658) <= not a;
    layer5_outputs(5659) <= not a;
    layer5_outputs(5660) <= b;
    layer5_outputs(5661) <= a or b;
    layer5_outputs(5662) <= not b or a;
    layer5_outputs(5663) <= not (a xor b);
    layer5_outputs(5664) <= not a;
    layer5_outputs(5665) <= a or b;
    layer5_outputs(5666) <= not (a xor b);
    layer5_outputs(5667) <= not (a and b);
    layer5_outputs(5668) <= a and not b;
    layer5_outputs(5669) <= not a or b;
    layer5_outputs(5670) <= a;
    layer5_outputs(5671) <= b and not a;
    layer5_outputs(5672) <= not (a or b);
    layer5_outputs(5673) <= a and not b;
    layer5_outputs(5674) <= a or b;
    layer5_outputs(5675) <= 1'b0;
    layer5_outputs(5676) <= b and not a;
    layer5_outputs(5677) <= not b;
    layer5_outputs(5678) <= a and b;
    layer5_outputs(5679) <= a;
    layer5_outputs(5680) <= b;
    layer5_outputs(5681) <= 1'b1;
    layer5_outputs(5682) <= not a;
    layer5_outputs(5683) <= b;
    layer5_outputs(5684) <= not (a and b);
    layer5_outputs(5685) <= not (a and b);
    layer5_outputs(5686) <= b;
    layer5_outputs(5687) <= b;
    layer5_outputs(5688) <= b and not a;
    layer5_outputs(5689) <= not a;
    layer5_outputs(5690) <= not a or b;
    layer5_outputs(5691) <= a and b;
    layer5_outputs(5692) <= b and not a;
    layer5_outputs(5693) <= not (a and b);
    layer5_outputs(5694) <= a;
    layer5_outputs(5695) <= a or b;
    layer5_outputs(5696) <= not a;
    layer5_outputs(5697) <= b and not a;
    layer5_outputs(5698) <= 1'b1;
    layer5_outputs(5699) <= 1'b1;
    layer5_outputs(5700) <= not b or a;
    layer5_outputs(5701) <= a and b;
    layer5_outputs(5702) <= a and b;
    layer5_outputs(5703) <= a or b;
    layer5_outputs(5704) <= a xor b;
    layer5_outputs(5705) <= 1'b1;
    layer5_outputs(5706) <= not a;
    layer5_outputs(5707) <= not (a and b);
    layer5_outputs(5708) <= not b;
    layer5_outputs(5709) <= a and b;
    layer5_outputs(5710) <= 1'b1;
    layer5_outputs(5711) <= a and not b;
    layer5_outputs(5712) <= b and not a;
    layer5_outputs(5713) <= not b;
    layer5_outputs(5714) <= not b;
    layer5_outputs(5715) <= not b;
    layer5_outputs(5716) <= a and not b;
    layer5_outputs(5717) <= b;
    layer5_outputs(5718) <= not (a or b);
    layer5_outputs(5719) <= not (a xor b);
    layer5_outputs(5720) <= 1'b1;
    layer5_outputs(5721) <= b and not a;
    layer5_outputs(5722) <= not b;
    layer5_outputs(5723) <= a and not b;
    layer5_outputs(5724) <= a;
    layer5_outputs(5725) <= b and not a;
    layer5_outputs(5726) <= 1'b1;
    layer5_outputs(5727) <= a;
    layer5_outputs(5728) <= not b;
    layer5_outputs(5729) <= b;
    layer5_outputs(5730) <= not b or a;
    layer5_outputs(5731) <= not b;
    layer5_outputs(5732) <= not b;
    layer5_outputs(5733) <= not b or a;
    layer5_outputs(5734) <= not a;
    layer5_outputs(5735) <= not b;
    layer5_outputs(5736) <= b and not a;
    layer5_outputs(5737) <= not b or a;
    layer5_outputs(5738) <= b;
    layer5_outputs(5739) <= a;
    layer5_outputs(5740) <= b;
    layer5_outputs(5741) <= not a;
    layer5_outputs(5742) <= b;
    layer5_outputs(5743) <= not (a or b);
    layer5_outputs(5744) <= not a;
    layer5_outputs(5745) <= not b or a;
    layer5_outputs(5746) <= not b;
    layer5_outputs(5747) <= b;
    layer5_outputs(5748) <= b;
    layer5_outputs(5749) <= 1'b0;
    layer5_outputs(5750) <= b;
    layer5_outputs(5751) <= not (a or b);
    layer5_outputs(5752) <= not (a and b);
    layer5_outputs(5753) <= a xor b;
    layer5_outputs(5754) <= not a or b;
    layer5_outputs(5755) <= a;
    layer5_outputs(5756) <= a and b;
    layer5_outputs(5757) <= not b;
    layer5_outputs(5758) <= not a or b;
    layer5_outputs(5759) <= b and not a;
    layer5_outputs(5760) <= b;
    layer5_outputs(5761) <= not b;
    layer5_outputs(5762) <= a;
    layer5_outputs(5763) <= not b;
    layer5_outputs(5764) <= b and not a;
    layer5_outputs(5765) <= a and b;
    layer5_outputs(5766) <= not a;
    layer5_outputs(5767) <= not (a and b);
    layer5_outputs(5768) <= not a;
    layer5_outputs(5769) <= a;
    layer5_outputs(5770) <= not a;
    layer5_outputs(5771) <= b;
    layer5_outputs(5772) <= b and not a;
    layer5_outputs(5773) <= not (a or b);
    layer5_outputs(5774) <= b;
    layer5_outputs(5775) <= not (a or b);
    layer5_outputs(5776) <= not a or b;
    layer5_outputs(5777) <= b and not a;
    layer5_outputs(5778) <= a and not b;
    layer5_outputs(5779) <= not (a or b);
    layer5_outputs(5780) <= not a or b;
    layer5_outputs(5781) <= not a;
    layer5_outputs(5782) <= b;
    layer5_outputs(5783) <= not b;
    layer5_outputs(5784) <= a xor b;
    layer5_outputs(5785) <= b and not a;
    layer5_outputs(5786) <= not a;
    layer5_outputs(5787) <= not a;
    layer5_outputs(5788) <= not a or b;
    layer5_outputs(5789) <= a;
    layer5_outputs(5790) <= a or b;
    layer5_outputs(5791) <= 1'b1;
    layer5_outputs(5792) <= b;
    layer5_outputs(5793) <= not b;
    layer5_outputs(5794) <= a;
    layer5_outputs(5795) <= b and not a;
    layer5_outputs(5796) <= not (a and b);
    layer5_outputs(5797) <= a and b;
    layer5_outputs(5798) <= a and not b;
    layer5_outputs(5799) <= 1'b1;
    layer5_outputs(5800) <= a and not b;
    layer5_outputs(5801) <= a or b;
    layer5_outputs(5802) <= a and b;
    layer5_outputs(5803) <= b and not a;
    layer5_outputs(5804) <= a;
    layer5_outputs(5805) <= a or b;
    layer5_outputs(5806) <= not a;
    layer5_outputs(5807) <= not b or a;
    layer5_outputs(5808) <= not b or a;
    layer5_outputs(5809) <= a or b;
    layer5_outputs(5810) <= not a or b;
    layer5_outputs(5811) <= a and not b;
    layer5_outputs(5812) <= 1'b1;
    layer5_outputs(5813) <= 1'b1;
    layer5_outputs(5814) <= not (a and b);
    layer5_outputs(5815) <= not a or b;
    layer5_outputs(5816) <= not (a and b);
    layer5_outputs(5817) <= a;
    layer5_outputs(5818) <= a and b;
    layer5_outputs(5819) <= not b;
    layer5_outputs(5820) <= 1'b0;
    layer5_outputs(5821) <= b;
    layer5_outputs(5822) <= not a or b;
    layer5_outputs(5823) <= not a or b;
    layer5_outputs(5824) <= not b;
    layer5_outputs(5825) <= a and not b;
    layer5_outputs(5826) <= a and b;
    layer5_outputs(5827) <= not b or a;
    layer5_outputs(5828) <= b;
    layer5_outputs(5829) <= not (a or b);
    layer5_outputs(5830) <= not b;
    layer5_outputs(5831) <= not a;
    layer5_outputs(5832) <= not b;
    layer5_outputs(5833) <= a and not b;
    layer5_outputs(5834) <= not b;
    layer5_outputs(5835) <= b and not a;
    layer5_outputs(5836) <= a xor b;
    layer5_outputs(5837) <= not a or b;
    layer5_outputs(5838) <= a xor b;
    layer5_outputs(5839) <= not a or b;
    layer5_outputs(5840) <= b and not a;
    layer5_outputs(5841) <= not (a or b);
    layer5_outputs(5842) <= a;
    layer5_outputs(5843) <= b;
    layer5_outputs(5844) <= not b;
    layer5_outputs(5845) <= not a or b;
    layer5_outputs(5846) <= not a or b;
    layer5_outputs(5847) <= not (a and b);
    layer5_outputs(5848) <= 1'b0;
    layer5_outputs(5849) <= 1'b1;
    layer5_outputs(5850) <= not a;
    layer5_outputs(5851) <= not a or b;
    layer5_outputs(5852) <= not (a and b);
    layer5_outputs(5853) <= not b;
    layer5_outputs(5854) <= a and b;
    layer5_outputs(5855) <= a and b;
    layer5_outputs(5856) <= not a;
    layer5_outputs(5857) <= a;
    layer5_outputs(5858) <= 1'b1;
    layer5_outputs(5859) <= b and not a;
    layer5_outputs(5860) <= not a or b;
    layer5_outputs(5861) <= not b or a;
    layer5_outputs(5862) <= a;
    layer5_outputs(5863) <= not (a xor b);
    layer5_outputs(5864) <= not b or a;
    layer5_outputs(5865) <= not b or a;
    layer5_outputs(5866) <= not b or a;
    layer5_outputs(5867) <= b and not a;
    layer5_outputs(5868) <= b;
    layer5_outputs(5869) <= a;
    layer5_outputs(5870) <= a;
    layer5_outputs(5871) <= b;
    layer5_outputs(5872) <= a;
    layer5_outputs(5873) <= 1'b0;
    layer5_outputs(5874) <= not b or a;
    layer5_outputs(5875) <= a and b;
    layer5_outputs(5876) <= a xor b;
    layer5_outputs(5877) <= not a or b;
    layer5_outputs(5878) <= not b;
    layer5_outputs(5879) <= b;
    layer5_outputs(5880) <= not a or b;
    layer5_outputs(5881) <= 1'b0;
    layer5_outputs(5882) <= not a;
    layer5_outputs(5883) <= not (a and b);
    layer5_outputs(5884) <= not a;
    layer5_outputs(5885) <= a;
    layer5_outputs(5886) <= not a;
    layer5_outputs(5887) <= not b;
    layer5_outputs(5888) <= not (a and b);
    layer5_outputs(5889) <= a;
    layer5_outputs(5890) <= a and b;
    layer5_outputs(5891) <= not (a and b);
    layer5_outputs(5892) <= not (a or b);
    layer5_outputs(5893) <= not (a or b);
    layer5_outputs(5894) <= a or b;
    layer5_outputs(5895) <= not (a or b);
    layer5_outputs(5896) <= not b;
    layer5_outputs(5897) <= a;
    layer5_outputs(5898) <= a;
    layer5_outputs(5899) <= not b;
    layer5_outputs(5900) <= a and b;
    layer5_outputs(5901) <= 1'b1;
    layer5_outputs(5902) <= a and not b;
    layer5_outputs(5903) <= not b;
    layer5_outputs(5904) <= not a;
    layer5_outputs(5905) <= a or b;
    layer5_outputs(5906) <= b and not a;
    layer5_outputs(5907) <= not a or b;
    layer5_outputs(5908) <= a;
    layer5_outputs(5909) <= not (a or b);
    layer5_outputs(5910) <= not a;
    layer5_outputs(5911) <= not (a or b);
    layer5_outputs(5912) <= not (a or b);
    layer5_outputs(5913) <= not a;
    layer5_outputs(5914) <= not a;
    layer5_outputs(5915) <= 1'b0;
    layer5_outputs(5916) <= not b or a;
    layer5_outputs(5917) <= not b or a;
    layer5_outputs(5918) <= not (a or b);
    layer5_outputs(5919) <= a;
    layer5_outputs(5920) <= not (a and b);
    layer5_outputs(5921) <= a;
    layer5_outputs(5922) <= not (a and b);
    layer5_outputs(5923) <= a or b;
    layer5_outputs(5924) <= not b;
    layer5_outputs(5925) <= a or b;
    layer5_outputs(5926) <= a xor b;
    layer5_outputs(5927) <= b;
    layer5_outputs(5928) <= b;
    layer5_outputs(5929) <= not a;
    layer5_outputs(5930) <= b;
    layer5_outputs(5931) <= not b;
    layer5_outputs(5932) <= not b;
    layer5_outputs(5933) <= a;
    layer5_outputs(5934) <= 1'b0;
    layer5_outputs(5935) <= not a or b;
    layer5_outputs(5936) <= a;
    layer5_outputs(5937) <= a and b;
    layer5_outputs(5938) <= not a;
    layer5_outputs(5939) <= a and b;
    layer5_outputs(5940) <= a and not b;
    layer5_outputs(5941) <= not (a or b);
    layer5_outputs(5942) <= 1'b1;
    layer5_outputs(5943) <= a and not b;
    layer5_outputs(5944) <= a;
    layer5_outputs(5945) <= not a;
    layer5_outputs(5946) <= b;
    layer5_outputs(5947) <= not (a or b);
    layer5_outputs(5948) <= 1'b1;
    layer5_outputs(5949) <= a;
    layer5_outputs(5950) <= not a;
    layer5_outputs(5951) <= a;
    layer5_outputs(5952) <= a xor b;
    layer5_outputs(5953) <= not a;
    layer5_outputs(5954) <= a and not b;
    layer5_outputs(5955) <= b and not a;
    layer5_outputs(5956) <= not (a and b);
    layer5_outputs(5957) <= b;
    layer5_outputs(5958) <= not b or a;
    layer5_outputs(5959) <= a;
    layer5_outputs(5960) <= a and b;
    layer5_outputs(5961) <= not b;
    layer5_outputs(5962) <= not b;
    layer5_outputs(5963) <= not a;
    layer5_outputs(5964) <= b and not a;
    layer5_outputs(5965) <= 1'b0;
    layer5_outputs(5966) <= not a;
    layer5_outputs(5967) <= a;
    layer5_outputs(5968) <= 1'b0;
    layer5_outputs(5969) <= not a or b;
    layer5_outputs(5970) <= b and not a;
    layer5_outputs(5971) <= a xor b;
    layer5_outputs(5972) <= not a;
    layer5_outputs(5973) <= not a or b;
    layer5_outputs(5974) <= b;
    layer5_outputs(5975) <= a;
    layer5_outputs(5976) <= a and not b;
    layer5_outputs(5977) <= a and not b;
    layer5_outputs(5978) <= not a;
    layer5_outputs(5979) <= not a;
    layer5_outputs(5980) <= not b;
    layer5_outputs(5981) <= a and not b;
    layer5_outputs(5982) <= a xor b;
    layer5_outputs(5983) <= 1'b0;
    layer5_outputs(5984) <= not (a or b);
    layer5_outputs(5985) <= a;
    layer5_outputs(5986) <= not (a or b);
    layer5_outputs(5987) <= not a;
    layer5_outputs(5988) <= a or b;
    layer5_outputs(5989) <= not b;
    layer5_outputs(5990) <= not b;
    layer5_outputs(5991) <= a and not b;
    layer5_outputs(5992) <= not (a and b);
    layer5_outputs(5993) <= b and not a;
    layer5_outputs(5994) <= not a;
    layer5_outputs(5995) <= not b;
    layer5_outputs(5996) <= b and not a;
    layer5_outputs(5997) <= not a or b;
    layer5_outputs(5998) <= b;
    layer5_outputs(5999) <= 1'b1;
    layer5_outputs(6000) <= a xor b;
    layer5_outputs(6001) <= a or b;
    layer5_outputs(6002) <= 1'b0;
    layer5_outputs(6003) <= not a or b;
    layer5_outputs(6004) <= a;
    layer5_outputs(6005) <= a and b;
    layer5_outputs(6006) <= not a;
    layer5_outputs(6007) <= not a or b;
    layer5_outputs(6008) <= not a or b;
    layer5_outputs(6009) <= not b;
    layer5_outputs(6010) <= a and b;
    layer5_outputs(6011) <= a and not b;
    layer5_outputs(6012) <= not a;
    layer5_outputs(6013) <= not a;
    layer5_outputs(6014) <= not b;
    layer5_outputs(6015) <= not a;
    layer5_outputs(6016) <= a and not b;
    layer5_outputs(6017) <= a xor b;
    layer5_outputs(6018) <= a;
    layer5_outputs(6019) <= a;
    layer5_outputs(6020) <= not (a or b);
    layer5_outputs(6021) <= b and not a;
    layer5_outputs(6022) <= a and b;
    layer5_outputs(6023) <= not a or b;
    layer5_outputs(6024) <= not (a or b);
    layer5_outputs(6025) <= a;
    layer5_outputs(6026) <= not (a xor b);
    layer5_outputs(6027) <= not b or a;
    layer5_outputs(6028) <= not a;
    layer5_outputs(6029) <= b;
    layer5_outputs(6030) <= 1'b0;
    layer5_outputs(6031) <= b;
    layer5_outputs(6032) <= not a or b;
    layer5_outputs(6033) <= b;
    layer5_outputs(6034) <= not (a xor b);
    layer5_outputs(6035) <= not b;
    layer5_outputs(6036) <= a xor b;
    layer5_outputs(6037) <= a xor b;
    layer5_outputs(6038) <= 1'b0;
    layer5_outputs(6039) <= a;
    layer5_outputs(6040) <= not (a and b);
    layer5_outputs(6041) <= not (a xor b);
    layer5_outputs(6042) <= a or b;
    layer5_outputs(6043) <= 1'b0;
    layer5_outputs(6044) <= not (a xor b);
    layer5_outputs(6045) <= b;
    layer5_outputs(6046) <= not (a or b);
    layer5_outputs(6047) <= b;
    layer5_outputs(6048) <= not b;
    layer5_outputs(6049) <= not (a and b);
    layer5_outputs(6050) <= a or b;
    layer5_outputs(6051) <= b and not a;
    layer5_outputs(6052) <= a;
    layer5_outputs(6053) <= not (a and b);
    layer5_outputs(6054) <= not (a or b);
    layer5_outputs(6055) <= 1'b0;
    layer5_outputs(6056) <= not b;
    layer5_outputs(6057) <= not b or a;
    layer5_outputs(6058) <= not a;
    layer5_outputs(6059) <= not a;
    layer5_outputs(6060) <= b and not a;
    layer5_outputs(6061) <= 1'b1;
    layer5_outputs(6062) <= not (a xor b);
    layer5_outputs(6063) <= not b or a;
    layer5_outputs(6064) <= a or b;
    layer5_outputs(6065) <= a xor b;
    layer5_outputs(6066) <= not a;
    layer5_outputs(6067) <= a or b;
    layer5_outputs(6068) <= not (a xor b);
    layer5_outputs(6069) <= not (a or b);
    layer5_outputs(6070) <= not (a and b);
    layer5_outputs(6071) <= b and not a;
    layer5_outputs(6072) <= not a;
    layer5_outputs(6073) <= not a or b;
    layer5_outputs(6074) <= not b or a;
    layer5_outputs(6075) <= not b;
    layer5_outputs(6076) <= not (a and b);
    layer5_outputs(6077) <= a;
    layer5_outputs(6078) <= a and not b;
    layer5_outputs(6079) <= not (a and b);
    layer5_outputs(6080) <= a;
    layer5_outputs(6081) <= not (a and b);
    layer5_outputs(6082) <= b and not a;
    layer5_outputs(6083) <= b;
    layer5_outputs(6084) <= a and b;
    layer5_outputs(6085) <= not a;
    layer5_outputs(6086) <= a;
    layer5_outputs(6087) <= b;
    layer5_outputs(6088) <= b;
    layer5_outputs(6089) <= a and b;
    layer5_outputs(6090) <= a or b;
    layer5_outputs(6091) <= not b;
    layer5_outputs(6092) <= a;
    layer5_outputs(6093) <= a;
    layer5_outputs(6094) <= a;
    layer5_outputs(6095) <= not b;
    layer5_outputs(6096) <= not (a xor b);
    layer5_outputs(6097) <= 1'b0;
    layer5_outputs(6098) <= not b;
    layer5_outputs(6099) <= a and not b;
    layer5_outputs(6100) <= not b;
    layer5_outputs(6101) <= not a;
    layer5_outputs(6102) <= a or b;
    layer5_outputs(6103) <= a and b;
    layer5_outputs(6104) <= not (a xor b);
    layer5_outputs(6105) <= not b or a;
    layer5_outputs(6106) <= a and not b;
    layer5_outputs(6107) <= b and not a;
    layer5_outputs(6108) <= a or b;
    layer5_outputs(6109) <= 1'b1;
    layer5_outputs(6110) <= not (a and b);
    layer5_outputs(6111) <= a or b;
    layer5_outputs(6112) <= not b;
    layer5_outputs(6113) <= a;
    layer5_outputs(6114) <= not (a xor b);
    layer5_outputs(6115) <= not b or a;
    layer5_outputs(6116) <= not a;
    layer5_outputs(6117) <= not a;
    layer5_outputs(6118) <= 1'b0;
    layer5_outputs(6119) <= a or b;
    layer5_outputs(6120) <= not b;
    layer5_outputs(6121) <= not b;
    layer5_outputs(6122) <= a or b;
    layer5_outputs(6123) <= not (a or b);
    layer5_outputs(6124) <= b;
    layer5_outputs(6125) <= not (a xor b);
    layer5_outputs(6126) <= a or b;
    layer5_outputs(6127) <= a and b;
    layer5_outputs(6128) <= a xor b;
    layer5_outputs(6129) <= not b;
    layer5_outputs(6130) <= not a;
    layer5_outputs(6131) <= a and not b;
    layer5_outputs(6132) <= not b;
    layer5_outputs(6133) <= a or b;
    layer5_outputs(6134) <= not (a xor b);
    layer5_outputs(6135) <= not a or b;
    layer5_outputs(6136) <= not a;
    layer5_outputs(6137) <= a and b;
    layer5_outputs(6138) <= not b or a;
    layer5_outputs(6139) <= a and not b;
    layer5_outputs(6140) <= not (a xor b);
    layer5_outputs(6141) <= a;
    layer5_outputs(6142) <= not (a or b);
    layer5_outputs(6143) <= a xor b;
    layer5_outputs(6144) <= a xor b;
    layer5_outputs(6145) <= not b;
    layer5_outputs(6146) <= not a;
    layer5_outputs(6147) <= not b;
    layer5_outputs(6148) <= not (a xor b);
    layer5_outputs(6149) <= a and b;
    layer5_outputs(6150) <= not b;
    layer5_outputs(6151) <= b;
    layer5_outputs(6152) <= not a;
    layer5_outputs(6153) <= a and b;
    layer5_outputs(6154) <= a and b;
    layer5_outputs(6155) <= a;
    layer5_outputs(6156) <= b;
    layer5_outputs(6157) <= not a or b;
    layer5_outputs(6158) <= not b;
    layer5_outputs(6159) <= a and b;
    layer5_outputs(6160) <= a or b;
    layer5_outputs(6161) <= not a;
    layer5_outputs(6162) <= a or b;
    layer5_outputs(6163) <= a and not b;
    layer5_outputs(6164) <= a or b;
    layer5_outputs(6165) <= not a;
    layer5_outputs(6166) <= not a;
    layer5_outputs(6167) <= not a;
    layer5_outputs(6168) <= not a or b;
    layer5_outputs(6169) <= not b;
    layer5_outputs(6170) <= a or b;
    layer5_outputs(6171) <= a xor b;
    layer5_outputs(6172) <= not b;
    layer5_outputs(6173) <= 1'b0;
    layer5_outputs(6174) <= not (a or b);
    layer5_outputs(6175) <= not b or a;
    layer5_outputs(6176) <= not (a and b);
    layer5_outputs(6177) <= not (a xor b);
    layer5_outputs(6178) <= not b;
    layer5_outputs(6179) <= not b;
    layer5_outputs(6180) <= not a or b;
    layer5_outputs(6181) <= a and b;
    layer5_outputs(6182) <= not b;
    layer5_outputs(6183) <= not (a or b);
    layer5_outputs(6184) <= not (a and b);
    layer5_outputs(6185) <= not b or a;
    layer5_outputs(6186) <= a;
    layer5_outputs(6187) <= not a;
    layer5_outputs(6188) <= a and not b;
    layer5_outputs(6189) <= not (a or b);
    layer5_outputs(6190) <= not b or a;
    layer5_outputs(6191) <= a;
    layer5_outputs(6192) <= not b or a;
    layer5_outputs(6193) <= a and not b;
    layer5_outputs(6194) <= not a;
    layer5_outputs(6195) <= not a;
    layer5_outputs(6196) <= a;
    layer5_outputs(6197) <= not b or a;
    layer5_outputs(6198) <= a or b;
    layer5_outputs(6199) <= not a or b;
    layer5_outputs(6200) <= a or b;
    layer5_outputs(6201) <= not b;
    layer5_outputs(6202) <= not a;
    layer5_outputs(6203) <= a and not b;
    layer5_outputs(6204) <= 1'b1;
    layer5_outputs(6205) <= 1'b1;
    layer5_outputs(6206) <= a;
    layer5_outputs(6207) <= not (a or b);
    layer5_outputs(6208) <= not a or b;
    layer5_outputs(6209) <= not a;
    layer5_outputs(6210) <= a;
    layer5_outputs(6211) <= not b or a;
    layer5_outputs(6212) <= a and not b;
    layer5_outputs(6213) <= not (a and b);
    layer5_outputs(6214) <= not b or a;
    layer5_outputs(6215) <= not a;
    layer5_outputs(6216) <= not (a and b);
    layer5_outputs(6217) <= not (a or b);
    layer5_outputs(6218) <= not a or b;
    layer5_outputs(6219) <= a;
    layer5_outputs(6220) <= b and not a;
    layer5_outputs(6221) <= not (a or b);
    layer5_outputs(6222) <= not a;
    layer5_outputs(6223) <= 1'b0;
    layer5_outputs(6224) <= a;
    layer5_outputs(6225) <= a and b;
    layer5_outputs(6226) <= not (a and b);
    layer5_outputs(6227) <= not b;
    layer5_outputs(6228) <= b and not a;
    layer5_outputs(6229) <= not b;
    layer5_outputs(6230) <= b and not a;
    layer5_outputs(6231) <= a or b;
    layer5_outputs(6232) <= b;
    layer5_outputs(6233) <= 1'b0;
    layer5_outputs(6234) <= a and not b;
    layer5_outputs(6235) <= not a;
    layer5_outputs(6236) <= not b;
    layer5_outputs(6237) <= 1'b1;
    layer5_outputs(6238) <= not (a xor b);
    layer5_outputs(6239) <= a and not b;
    layer5_outputs(6240) <= not a;
    layer5_outputs(6241) <= b;
    layer5_outputs(6242) <= not b;
    layer5_outputs(6243) <= a and b;
    layer5_outputs(6244) <= 1'b0;
    layer5_outputs(6245) <= not b;
    layer5_outputs(6246) <= 1'b0;
    layer5_outputs(6247) <= not b;
    layer5_outputs(6248) <= a and not b;
    layer5_outputs(6249) <= not (a xor b);
    layer5_outputs(6250) <= not b;
    layer5_outputs(6251) <= not (a xor b);
    layer5_outputs(6252) <= a xor b;
    layer5_outputs(6253) <= a and b;
    layer5_outputs(6254) <= not (a or b);
    layer5_outputs(6255) <= not (a and b);
    layer5_outputs(6256) <= b;
    layer5_outputs(6257) <= not a or b;
    layer5_outputs(6258) <= not b;
    layer5_outputs(6259) <= not b or a;
    layer5_outputs(6260) <= a xor b;
    layer5_outputs(6261) <= 1'b0;
    layer5_outputs(6262) <= not a or b;
    layer5_outputs(6263) <= 1'b1;
    layer5_outputs(6264) <= a;
    layer5_outputs(6265) <= not a;
    layer5_outputs(6266) <= not (a or b);
    layer5_outputs(6267) <= a and b;
    layer5_outputs(6268) <= a or b;
    layer5_outputs(6269) <= a;
    layer5_outputs(6270) <= not (a xor b);
    layer5_outputs(6271) <= 1'b0;
    layer5_outputs(6272) <= b;
    layer5_outputs(6273) <= b and not a;
    layer5_outputs(6274) <= not a or b;
    layer5_outputs(6275) <= 1'b1;
    layer5_outputs(6276) <= a xor b;
    layer5_outputs(6277) <= not a or b;
    layer5_outputs(6278) <= not a or b;
    layer5_outputs(6279) <= b and not a;
    layer5_outputs(6280) <= a or b;
    layer5_outputs(6281) <= a and b;
    layer5_outputs(6282) <= not a or b;
    layer5_outputs(6283) <= not (a and b);
    layer5_outputs(6284) <= a;
    layer5_outputs(6285) <= not b or a;
    layer5_outputs(6286) <= not b;
    layer5_outputs(6287) <= not (a and b);
    layer5_outputs(6288) <= b and not a;
    layer5_outputs(6289) <= not a or b;
    layer5_outputs(6290) <= not a;
    layer5_outputs(6291) <= not (a and b);
    layer5_outputs(6292) <= b;
    layer5_outputs(6293) <= not a;
    layer5_outputs(6294) <= not a or b;
    layer5_outputs(6295) <= a and not b;
    layer5_outputs(6296) <= a xor b;
    layer5_outputs(6297) <= a and b;
    layer5_outputs(6298) <= a or b;
    layer5_outputs(6299) <= not b or a;
    layer5_outputs(6300) <= not a;
    layer5_outputs(6301) <= not a or b;
    layer5_outputs(6302) <= a or b;
    layer5_outputs(6303) <= not b;
    layer5_outputs(6304) <= a xor b;
    layer5_outputs(6305) <= not a or b;
    layer5_outputs(6306) <= a xor b;
    layer5_outputs(6307) <= a and b;
    layer5_outputs(6308) <= a and b;
    layer5_outputs(6309) <= a xor b;
    layer5_outputs(6310) <= a;
    layer5_outputs(6311) <= a or b;
    layer5_outputs(6312) <= not (a or b);
    layer5_outputs(6313) <= not (a xor b);
    layer5_outputs(6314) <= a or b;
    layer5_outputs(6315) <= b and not a;
    layer5_outputs(6316) <= 1'b1;
    layer5_outputs(6317) <= b and not a;
    layer5_outputs(6318) <= 1'b0;
    layer5_outputs(6319) <= not a;
    layer5_outputs(6320) <= 1'b0;
    layer5_outputs(6321) <= not a or b;
    layer5_outputs(6322) <= not (a and b);
    layer5_outputs(6323) <= not a or b;
    layer5_outputs(6324) <= 1'b1;
    layer5_outputs(6325) <= not a or b;
    layer5_outputs(6326) <= not a or b;
    layer5_outputs(6327) <= b;
    layer5_outputs(6328) <= not b or a;
    layer5_outputs(6329) <= b;
    layer5_outputs(6330) <= a or b;
    layer5_outputs(6331) <= not b;
    layer5_outputs(6332) <= b and not a;
    layer5_outputs(6333) <= a and not b;
    layer5_outputs(6334) <= b;
    layer5_outputs(6335) <= not (a xor b);
    layer5_outputs(6336) <= a xor b;
    layer5_outputs(6337) <= a xor b;
    layer5_outputs(6338) <= 1'b0;
    layer5_outputs(6339) <= not b;
    layer5_outputs(6340) <= not a;
    layer5_outputs(6341) <= a and not b;
    layer5_outputs(6342) <= not (a and b);
    layer5_outputs(6343) <= not b or a;
    layer5_outputs(6344) <= b and not a;
    layer5_outputs(6345) <= 1'b1;
    layer5_outputs(6346) <= b;
    layer5_outputs(6347) <= b and not a;
    layer5_outputs(6348) <= not b;
    layer5_outputs(6349) <= not b;
    layer5_outputs(6350) <= not a;
    layer5_outputs(6351) <= not a;
    layer5_outputs(6352) <= not b;
    layer5_outputs(6353) <= not b or a;
    layer5_outputs(6354) <= not (a xor b);
    layer5_outputs(6355) <= not a;
    layer5_outputs(6356) <= not (a and b);
    layer5_outputs(6357) <= a and not b;
    layer5_outputs(6358) <= b;
    layer5_outputs(6359) <= a and b;
    layer5_outputs(6360) <= a xor b;
    layer5_outputs(6361) <= a;
    layer5_outputs(6362) <= 1'b1;
    layer5_outputs(6363) <= not a or b;
    layer5_outputs(6364) <= b;
    layer5_outputs(6365) <= b and not a;
    layer5_outputs(6366) <= b;
    layer5_outputs(6367) <= b and not a;
    layer5_outputs(6368) <= b and not a;
    layer5_outputs(6369) <= not (a and b);
    layer5_outputs(6370) <= a xor b;
    layer5_outputs(6371) <= not a or b;
    layer5_outputs(6372) <= not b;
    layer5_outputs(6373) <= b;
    layer5_outputs(6374) <= not a;
    layer5_outputs(6375) <= not b;
    layer5_outputs(6376) <= not a;
    layer5_outputs(6377) <= a;
    layer5_outputs(6378) <= a and b;
    layer5_outputs(6379) <= not b;
    layer5_outputs(6380) <= not b;
    layer5_outputs(6381) <= not (a and b);
    layer5_outputs(6382) <= 1'b0;
    layer5_outputs(6383) <= not b or a;
    layer5_outputs(6384) <= not (a xor b);
    layer5_outputs(6385) <= a;
    layer5_outputs(6386) <= not a;
    layer5_outputs(6387) <= 1'b1;
    layer5_outputs(6388) <= not a or b;
    layer5_outputs(6389) <= not (a and b);
    layer5_outputs(6390) <= 1'b1;
    layer5_outputs(6391) <= not (a xor b);
    layer5_outputs(6392) <= a xor b;
    layer5_outputs(6393) <= 1'b1;
    layer5_outputs(6394) <= 1'b1;
    layer5_outputs(6395) <= not (a xor b);
    layer5_outputs(6396) <= not a;
    layer5_outputs(6397) <= not a;
    layer5_outputs(6398) <= not a or b;
    layer5_outputs(6399) <= not b or a;
    layer5_outputs(6400) <= a or b;
    layer5_outputs(6401) <= not b;
    layer5_outputs(6402) <= b and not a;
    layer5_outputs(6403) <= not (a and b);
    layer5_outputs(6404) <= b and not a;
    layer5_outputs(6405) <= b and not a;
    layer5_outputs(6406) <= a xor b;
    layer5_outputs(6407) <= not a;
    layer5_outputs(6408) <= a or b;
    layer5_outputs(6409) <= b;
    layer5_outputs(6410) <= not b;
    layer5_outputs(6411) <= a or b;
    layer5_outputs(6412) <= a or b;
    layer5_outputs(6413) <= b and not a;
    layer5_outputs(6414) <= not b;
    layer5_outputs(6415) <= not b;
    layer5_outputs(6416) <= a and b;
    layer5_outputs(6417) <= not (a xor b);
    layer5_outputs(6418) <= b and not a;
    layer5_outputs(6419) <= not a or b;
    layer5_outputs(6420) <= not a or b;
    layer5_outputs(6421) <= b;
    layer5_outputs(6422) <= a and b;
    layer5_outputs(6423) <= b;
    layer5_outputs(6424) <= a and b;
    layer5_outputs(6425) <= b and not a;
    layer5_outputs(6426) <= not a;
    layer5_outputs(6427) <= a;
    layer5_outputs(6428) <= b;
    layer5_outputs(6429) <= not (a and b);
    layer5_outputs(6430) <= not (a and b);
    layer5_outputs(6431) <= not (a and b);
    layer5_outputs(6432) <= not (a and b);
    layer5_outputs(6433) <= not a or b;
    layer5_outputs(6434) <= 1'b0;
    layer5_outputs(6435) <= b and not a;
    layer5_outputs(6436) <= 1'b1;
    layer5_outputs(6437) <= b and not a;
    layer5_outputs(6438) <= a and not b;
    layer5_outputs(6439) <= a;
    layer5_outputs(6440) <= a or b;
    layer5_outputs(6441) <= a and b;
    layer5_outputs(6442) <= not (a and b);
    layer5_outputs(6443) <= a or b;
    layer5_outputs(6444) <= not a;
    layer5_outputs(6445) <= a or b;
    layer5_outputs(6446) <= 1'b1;
    layer5_outputs(6447) <= not b;
    layer5_outputs(6448) <= 1'b1;
    layer5_outputs(6449) <= a and b;
    layer5_outputs(6450) <= b;
    layer5_outputs(6451) <= 1'b1;
    layer5_outputs(6452) <= 1'b1;
    layer5_outputs(6453) <= not (a or b);
    layer5_outputs(6454) <= b;
    layer5_outputs(6455) <= not (a or b);
    layer5_outputs(6456) <= b;
    layer5_outputs(6457) <= not (a and b);
    layer5_outputs(6458) <= not b;
    layer5_outputs(6459) <= not (a xor b);
    layer5_outputs(6460) <= not a;
    layer5_outputs(6461) <= a xor b;
    layer5_outputs(6462) <= not (a and b);
    layer5_outputs(6463) <= not (a or b);
    layer5_outputs(6464) <= not a or b;
    layer5_outputs(6465) <= not b;
    layer5_outputs(6466) <= b and not a;
    layer5_outputs(6467) <= not b or a;
    layer5_outputs(6468) <= a and b;
    layer5_outputs(6469) <= b;
    layer5_outputs(6470) <= b and not a;
    layer5_outputs(6471) <= not (a or b);
    layer5_outputs(6472) <= a or b;
    layer5_outputs(6473) <= 1'b0;
    layer5_outputs(6474) <= a;
    layer5_outputs(6475) <= not b or a;
    layer5_outputs(6476) <= not (a or b);
    layer5_outputs(6477) <= not b;
    layer5_outputs(6478) <= 1'b1;
    layer5_outputs(6479) <= not (a and b);
    layer5_outputs(6480) <= a;
    layer5_outputs(6481) <= a or b;
    layer5_outputs(6482) <= not a;
    layer5_outputs(6483) <= 1'b0;
    layer5_outputs(6484) <= not a;
    layer5_outputs(6485) <= b;
    layer5_outputs(6486) <= not a or b;
    layer5_outputs(6487) <= not (a or b);
    layer5_outputs(6488) <= a and b;
    layer5_outputs(6489) <= a and b;
    layer5_outputs(6490) <= a and not b;
    layer5_outputs(6491) <= not (a or b);
    layer5_outputs(6492) <= not (a or b);
    layer5_outputs(6493) <= not (a or b);
    layer5_outputs(6494) <= 1'b1;
    layer5_outputs(6495) <= a xor b;
    layer5_outputs(6496) <= b and not a;
    layer5_outputs(6497) <= a or b;
    layer5_outputs(6498) <= a;
    layer5_outputs(6499) <= b;
    layer5_outputs(6500) <= not a or b;
    layer5_outputs(6501) <= b and not a;
    layer5_outputs(6502) <= a and b;
    layer5_outputs(6503) <= a or b;
    layer5_outputs(6504) <= not (a and b);
    layer5_outputs(6505) <= a or b;
    layer5_outputs(6506) <= a xor b;
    layer5_outputs(6507) <= a and b;
    layer5_outputs(6508) <= not (a and b);
    layer5_outputs(6509) <= not b or a;
    layer5_outputs(6510) <= not a;
    layer5_outputs(6511) <= not a or b;
    layer5_outputs(6512) <= b;
    layer5_outputs(6513) <= not a;
    layer5_outputs(6514) <= a;
    layer5_outputs(6515) <= not a or b;
    layer5_outputs(6516) <= not b;
    layer5_outputs(6517) <= b;
    layer5_outputs(6518) <= not b;
    layer5_outputs(6519) <= b;
    layer5_outputs(6520) <= not a or b;
    layer5_outputs(6521) <= not a;
    layer5_outputs(6522) <= b;
    layer5_outputs(6523) <= a;
    layer5_outputs(6524) <= b;
    layer5_outputs(6525) <= not a;
    layer5_outputs(6526) <= 1'b1;
    layer5_outputs(6527) <= a;
    layer5_outputs(6528) <= a and b;
    layer5_outputs(6529) <= a;
    layer5_outputs(6530) <= b and not a;
    layer5_outputs(6531) <= b;
    layer5_outputs(6532) <= not (a or b);
    layer5_outputs(6533) <= a or b;
    layer5_outputs(6534) <= 1'b0;
    layer5_outputs(6535) <= not a or b;
    layer5_outputs(6536) <= 1'b1;
    layer5_outputs(6537) <= not b or a;
    layer5_outputs(6538) <= not (a xor b);
    layer5_outputs(6539) <= a;
    layer5_outputs(6540) <= b and not a;
    layer5_outputs(6541) <= not b;
    layer5_outputs(6542) <= b;
    layer5_outputs(6543) <= not b or a;
    layer5_outputs(6544) <= a and b;
    layer5_outputs(6545) <= b;
    layer5_outputs(6546) <= not a;
    layer5_outputs(6547) <= not a;
    layer5_outputs(6548) <= not a;
    layer5_outputs(6549) <= not (a and b);
    layer5_outputs(6550) <= a;
    layer5_outputs(6551) <= not (a and b);
    layer5_outputs(6552) <= a and b;
    layer5_outputs(6553) <= a and b;
    layer5_outputs(6554) <= not b;
    layer5_outputs(6555) <= a;
    layer5_outputs(6556) <= a and not b;
    layer5_outputs(6557) <= a;
    layer5_outputs(6558) <= b and not a;
    layer5_outputs(6559) <= not b;
    layer5_outputs(6560) <= not a;
    layer5_outputs(6561) <= a;
    layer5_outputs(6562) <= not a;
    layer5_outputs(6563) <= not b or a;
    layer5_outputs(6564) <= not (a and b);
    layer5_outputs(6565) <= not a;
    layer5_outputs(6566) <= not (a or b);
    layer5_outputs(6567) <= not a;
    layer5_outputs(6568) <= a or b;
    layer5_outputs(6569) <= not (a xor b);
    layer5_outputs(6570) <= 1'b1;
    layer5_outputs(6571) <= b;
    layer5_outputs(6572) <= not b;
    layer5_outputs(6573) <= b and not a;
    layer5_outputs(6574) <= a and b;
    layer5_outputs(6575) <= a xor b;
    layer5_outputs(6576) <= 1'b1;
    layer5_outputs(6577) <= a;
    layer5_outputs(6578) <= not b or a;
    layer5_outputs(6579) <= a;
    layer5_outputs(6580) <= a and b;
    layer5_outputs(6581) <= not b;
    layer5_outputs(6582) <= a and not b;
    layer5_outputs(6583) <= a;
    layer5_outputs(6584) <= not (a xor b);
    layer5_outputs(6585) <= not (a xor b);
    layer5_outputs(6586) <= not b or a;
    layer5_outputs(6587) <= b and not a;
    layer5_outputs(6588) <= not (a or b);
    layer5_outputs(6589) <= b;
    layer5_outputs(6590) <= not b;
    layer5_outputs(6591) <= not (a xor b);
    layer5_outputs(6592) <= a;
    layer5_outputs(6593) <= a and b;
    layer5_outputs(6594) <= a;
    layer5_outputs(6595) <= not a;
    layer5_outputs(6596) <= not a or b;
    layer5_outputs(6597) <= not a;
    layer5_outputs(6598) <= b and not a;
    layer5_outputs(6599) <= b;
    layer5_outputs(6600) <= b and not a;
    layer5_outputs(6601) <= not b or a;
    layer5_outputs(6602) <= a and b;
    layer5_outputs(6603) <= a or b;
    layer5_outputs(6604) <= not b or a;
    layer5_outputs(6605) <= a and not b;
    layer5_outputs(6606) <= a and b;
    layer5_outputs(6607) <= not (a and b);
    layer5_outputs(6608) <= not (a and b);
    layer5_outputs(6609) <= not a;
    layer5_outputs(6610) <= b;
    layer5_outputs(6611) <= not a;
    layer5_outputs(6612) <= b and not a;
    layer5_outputs(6613) <= a and b;
    layer5_outputs(6614) <= not a or b;
    layer5_outputs(6615) <= a;
    layer5_outputs(6616) <= not (a or b);
    layer5_outputs(6617) <= 1'b0;
    layer5_outputs(6618) <= not a;
    layer5_outputs(6619) <= b;
    layer5_outputs(6620) <= a and b;
    layer5_outputs(6621) <= a and not b;
    layer5_outputs(6622) <= a and b;
    layer5_outputs(6623) <= a or b;
    layer5_outputs(6624) <= a or b;
    layer5_outputs(6625) <= 1'b0;
    layer5_outputs(6626) <= b;
    layer5_outputs(6627) <= not b;
    layer5_outputs(6628) <= 1'b1;
    layer5_outputs(6629) <= b and not a;
    layer5_outputs(6630) <= not (a or b);
    layer5_outputs(6631) <= a or b;
    layer5_outputs(6632) <= not a;
    layer5_outputs(6633) <= not a;
    layer5_outputs(6634) <= not b;
    layer5_outputs(6635) <= a;
    layer5_outputs(6636) <= b and not a;
    layer5_outputs(6637) <= b and not a;
    layer5_outputs(6638) <= not (a xor b);
    layer5_outputs(6639) <= not (a or b);
    layer5_outputs(6640) <= b;
    layer5_outputs(6641) <= b;
    layer5_outputs(6642) <= not b;
    layer5_outputs(6643) <= not a;
    layer5_outputs(6644) <= b;
    layer5_outputs(6645) <= a;
    layer5_outputs(6646) <= a;
    layer5_outputs(6647) <= not a or b;
    layer5_outputs(6648) <= not a;
    layer5_outputs(6649) <= a xor b;
    layer5_outputs(6650) <= b;
    layer5_outputs(6651) <= b;
    layer5_outputs(6652) <= b and not a;
    layer5_outputs(6653) <= b;
    layer5_outputs(6654) <= not a;
    layer5_outputs(6655) <= b and not a;
    layer5_outputs(6656) <= b;
    layer5_outputs(6657) <= a and not b;
    layer5_outputs(6658) <= not (a xor b);
    layer5_outputs(6659) <= b;
    layer5_outputs(6660) <= a and not b;
    layer5_outputs(6661) <= not b or a;
    layer5_outputs(6662) <= a and b;
    layer5_outputs(6663) <= not b;
    layer5_outputs(6664) <= a;
    layer5_outputs(6665) <= not a;
    layer5_outputs(6666) <= b and not a;
    layer5_outputs(6667) <= b and not a;
    layer5_outputs(6668) <= b and not a;
    layer5_outputs(6669) <= b;
    layer5_outputs(6670) <= a xor b;
    layer5_outputs(6671) <= not b or a;
    layer5_outputs(6672) <= not (a xor b);
    layer5_outputs(6673) <= not a or b;
    layer5_outputs(6674) <= b;
    layer5_outputs(6675) <= not a;
    layer5_outputs(6676) <= not (a xor b);
    layer5_outputs(6677) <= not b or a;
    layer5_outputs(6678) <= not b;
    layer5_outputs(6679) <= not b;
    layer5_outputs(6680) <= 1'b1;
    layer5_outputs(6681) <= b and not a;
    layer5_outputs(6682) <= a;
    layer5_outputs(6683) <= not (a or b);
    layer5_outputs(6684) <= not a;
    layer5_outputs(6685) <= a and b;
    layer5_outputs(6686) <= a and not b;
    layer5_outputs(6687) <= b;
    layer5_outputs(6688) <= a and b;
    layer5_outputs(6689) <= b and not a;
    layer5_outputs(6690) <= not b or a;
    layer5_outputs(6691) <= b;
    layer5_outputs(6692) <= a;
    layer5_outputs(6693) <= not b;
    layer5_outputs(6694) <= not (a and b);
    layer5_outputs(6695) <= a and b;
    layer5_outputs(6696) <= not a;
    layer5_outputs(6697) <= not (a or b);
    layer5_outputs(6698) <= 1'b1;
    layer5_outputs(6699) <= a and b;
    layer5_outputs(6700) <= b;
    layer5_outputs(6701) <= not a or b;
    layer5_outputs(6702) <= not b;
    layer5_outputs(6703) <= b;
    layer5_outputs(6704) <= a or b;
    layer5_outputs(6705) <= not a or b;
    layer5_outputs(6706) <= b;
    layer5_outputs(6707) <= a;
    layer5_outputs(6708) <= b and not a;
    layer5_outputs(6709) <= not b or a;
    layer5_outputs(6710) <= 1'b0;
    layer5_outputs(6711) <= not b;
    layer5_outputs(6712) <= a and b;
    layer5_outputs(6713) <= not (a xor b);
    layer5_outputs(6714) <= a and not b;
    layer5_outputs(6715) <= a;
    layer5_outputs(6716) <= a;
    layer5_outputs(6717) <= not a;
    layer5_outputs(6718) <= a xor b;
    layer5_outputs(6719) <= not a or b;
    layer5_outputs(6720) <= not b;
    layer5_outputs(6721) <= a;
    layer5_outputs(6722) <= a xor b;
    layer5_outputs(6723) <= not b;
    layer5_outputs(6724) <= not b;
    layer5_outputs(6725) <= a;
    layer5_outputs(6726) <= a;
    layer5_outputs(6727) <= not a;
    layer5_outputs(6728) <= not a or b;
    layer5_outputs(6729) <= a and b;
    layer5_outputs(6730) <= not a or b;
    layer5_outputs(6731) <= a;
    layer5_outputs(6732) <= a;
    layer5_outputs(6733) <= not (a or b);
    layer5_outputs(6734) <= not a or b;
    layer5_outputs(6735) <= not (a and b);
    layer5_outputs(6736) <= not a or b;
    layer5_outputs(6737) <= a and b;
    layer5_outputs(6738) <= a or b;
    layer5_outputs(6739) <= not b;
    layer5_outputs(6740) <= not (a xor b);
    layer5_outputs(6741) <= not b;
    layer5_outputs(6742) <= not a or b;
    layer5_outputs(6743) <= b;
    layer5_outputs(6744) <= a and b;
    layer5_outputs(6745) <= not a;
    layer5_outputs(6746) <= not b or a;
    layer5_outputs(6747) <= b and not a;
    layer5_outputs(6748) <= not (a or b);
    layer5_outputs(6749) <= 1'b1;
    layer5_outputs(6750) <= a xor b;
    layer5_outputs(6751) <= not (a or b);
    layer5_outputs(6752) <= not b;
    layer5_outputs(6753) <= b;
    layer5_outputs(6754) <= b and not a;
    layer5_outputs(6755) <= a and b;
    layer5_outputs(6756) <= not a or b;
    layer5_outputs(6757) <= b;
    layer5_outputs(6758) <= not (a or b);
    layer5_outputs(6759) <= 1'b0;
    layer5_outputs(6760) <= a xor b;
    layer5_outputs(6761) <= not a or b;
    layer5_outputs(6762) <= b and not a;
    layer5_outputs(6763) <= not b;
    layer5_outputs(6764) <= not a;
    layer5_outputs(6765) <= a or b;
    layer5_outputs(6766) <= not (a and b);
    layer5_outputs(6767) <= not (a xor b);
    layer5_outputs(6768) <= not b;
    layer5_outputs(6769) <= a or b;
    layer5_outputs(6770) <= not (a and b);
    layer5_outputs(6771) <= not (a and b);
    layer5_outputs(6772) <= not b or a;
    layer5_outputs(6773) <= not (a or b);
    layer5_outputs(6774) <= a;
    layer5_outputs(6775) <= not a;
    layer5_outputs(6776) <= not (a and b);
    layer5_outputs(6777) <= a;
    layer5_outputs(6778) <= a and b;
    layer5_outputs(6779) <= a xor b;
    layer5_outputs(6780) <= not (a or b);
    layer5_outputs(6781) <= 1'b0;
    layer5_outputs(6782) <= a;
    layer5_outputs(6783) <= not a;
    layer5_outputs(6784) <= not a or b;
    layer5_outputs(6785) <= not (a or b);
    layer5_outputs(6786) <= not b;
    layer5_outputs(6787) <= a or b;
    layer5_outputs(6788) <= not (a and b);
    layer5_outputs(6789) <= a and not b;
    layer5_outputs(6790) <= not b;
    layer5_outputs(6791) <= not (a xor b);
    layer5_outputs(6792) <= not b;
    layer5_outputs(6793) <= not b;
    layer5_outputs(6794) <= b;
    layer5_outputs(6795) <= a and b;
    layer5_outputs(6796) <= a or b;
    layer5_outputs(6797) <= b;
    layer5_outputs(6798) <= not b;
    layer5_outputs(6799) <= a and not b;
    layer5_outputs(6800) <= not b;
    layer5_outputs(6801) <= a;
    layer5_outputs(6802) <= not (a or b);
    layer5_outputs(6803) <= not a;
    layer5_outputs(6804) <= b;
    layer5_outputs(6805) <= a and not b;
    layer5_outputs(6806) <= a;
    layer5_outputs(6807) <= a;
    layer5_outputs(6808) <= a and not b;
    layer5_outputs(6809) <= a;
    layer5_outputs(6810) <= not b;
    layer5_outputs(6811) <= a and b;
    layer5_outputs(6812) <= not a;
    layer5_outputs(6813) <= a or b;
    layer5_outputs(6814) <= not b;
    layer5_outputs(6815) <= 1'b0;
    layer5_outputs(6816) <= a xor b;
    layer5_outputs(6817) <= not (a or b);
    layer5_outputs(6818) <= not a;
    layer5_outputs(6819) <= not (a and b);
    layer5_outputs(6820) <= not (a and b);
    layer5_outputs(6821) <= not b;
    layer5_outputs(6822) <= b and not a;
    layer5_outputs(6823) <= a or b;
    layer5_outputs(6824) <= a and not b;
    layer5_outputs(6825) <= a;
    layer5_outputs(6826) <= not a;
    layer5_outputs(6827) <= a and not b;
    layer5_outputs(6828) <= a;
    layer5_outputs(6829) <= not b or a;
    layer5_outputs(6830) <= a;
    layer5_outputs(6831) <= not b;
    layer5_outputs(6832) <= not a or b;
    layer5_outputs(6833) <= a and not b;
    layer5_outputs(6834) <= a and not b;
    layer5_outputs(6835) <= not b or a;
    layer5_outputs(6836) <= not a or b;
    layer5_outputs(6837) <= 1'b0;
    layer5_outputs(6838) <= not b;
    layer5_outputs(6839) <= not a;
    layer5_outputs(6840) <= not b;
    layer5_outputs(6841) <= not (a and b);
    layer5_outputs(6842) <= not b;
    layer5_outputs(6843) <= not a or b;
    layer5_outputs(6844) <= not (a and b);
    layer5_outputs(6845) <= a;
    layer5_outputs(6846) <= 1'b1;
    layer5_outputs(6847) <= a or b;
    layer5_outputs(6848) <= not b or a;
    layer5_outputs(6849) <= not a;
    layer5_outputs(6850) <= not (a xor b);
    layer5_outputs(6851) <= a;
    layer5_outputs(6852) <= not a;
    layer5_outputs(6853) <= b;
    layer5_outputs(6854) <= not (a xor b);
    layer5_outputs(6855) <= not b;
    layer5_outputs(6856) <= not a;
    layer5_outputs(6857) <= a or b;
    layer5_outputs(6858) <= not a;
    layer5_outputs(6859) <= not a;
    layer5_outputs(6860) <= not b;
    layer5_outputs(6861) <= not (a or b);
    layer5_outputs(6862) <= a xor b;
    layer5_outputs(6863) <= not b;
    layer5_outputs(6864) <= a and b;
    layer5_outputs(6865) <= 1'b1;
    layer5_outputs(6866) <= b and not a;
    layer5_outputs(6867) <= 1'b1;
    layer5_outputs(6868) <= a and b;
    layer5_outputs(6869) <= a;
    layer5_outputs(6870) <= not a;
    layer5_outputs(6871) <= a xor b;
    layer5_outputs(6872) <= a;
    layer5_outputs(6873) <= a and not b;
    layer5_outputs(6874) <= a or b;
    layer5_outputs(6875) <= 1'b1;
    layer5_outputs(6876) <= not (a or b);
    layer5_outputs(6877) <= not (a xor b);
    layer5_outputs(6878) <= 1'b1;
    layer5_outputs(6879) <= a;
    layer5_outputs(6880) <= not a or b;
    layer5_outputs(6881) <= not (a and b);
    layer5_outputs(6882) <= not (a or b);
    layer5_outputs(6883) <= a and b;
    layer5_outputs(6884) <= a and not b;
    layer5_outputs(6885) <= not b;
    layer5_outputs(6886) <= a or b;
    layer5_outputs(6887) <= not (a xor b);
    layer5_outputs(6888) <= 1'b0;
    layer5_outputs(6889) <= not a;
    layer5_outputs(6890) <= b;
    layer5_outputs(6891) <= not a;
    layer5_outputs(6892) <= b;
    layer5_outputs(6893) <= not (a and b);
    layer5_outputs(6894) <= a or b;
    layer5_outputs(6895) <= a or b;
    layer5_outputs(6896) <= a and not b;
    layer5_outputs(6897) <= not a;
    layer5_outputs(6898) <= a or b;
    layer5_outputs(6899) <= not b or a;
    layer5_outputs(6900) <= b;
    layer5_outputs(6901) <= not (a and b);
    layer5_outputs(6902) <= b;
    layer5_outputs(6903) <= a;
    layer5_outputs(6904) <= not b;
    layer5_outputs(6905) <= a and not b;
    layer5_outputs(6906) <= b;
    layer5_outputs(6907) <= b;
    layer5_outputs(6908) <= a;
    layer5_outputs(6909) <= not (a xor b);
    layer5_outputs(6910) <= not (a or b);
    layer5_outputs(6911) <= not a or b;
    layer5_outputs(6912) <= not b;
    layer5_outputs(6913) <= a and b;
    layer5_outputs(6914) <= not a;
    layer5_outputs(6915) <= a;
    layer5_outputs(6916) <= b;
    layer5_outputs(6917) <= a;
    layer5_outputs(6918) <= b and not a;
    layer5_outputs(6919) <= a xor b;
    layer5_outputs(6920) <= not (a or b);
    layer5_outputs(6921) <= not b;
    layer5_outputs(6922) <= a and not b;
    layer5_outputs(6923) <= not a or b;
    layer5_outputs(6924) <= not b or a;
    layer5_outputs(6925) <= a and not b;
    layer5_outputs(6926) <= not b;
    layer5_outputs(6927) <= 1'b0;
    layer5_outputs(6928) <= not a or b;
    layer5_outputs(6929) <= b;
    layer5_outputs(6930) <= not b;
    layer5_outputs(6931) <= b;
    layer5_outputs(6932) <= not (a or b);
    layer5_outputs(6933) <= a;
    layer5_outputs(6934) <= not (a and b);
    layer5_outputs(6935) <= not a;
    layer5_outputs(6936) <= not a;
    layer5_outputs(6937) <= a xor b;
    layer5_outputs(6938) <= not a;
    layer5_outputs(6939) <= b and not a;
    layer5_outputs(6940) <= not (a or b);
    layer5_outputs(6941) <= not b;
    layer5_outputs(6942) <= a and b;
    layer5_outputs(6943) <= not (a and b);
    layer5_outputs(6944) <= not a;
    layer5_outputs(6945) <= not b or a;
    layer5_outputs(6946) <= b;
    layer5_outputs(6947) <= a and not b;
    layer5_outputs(6948) <= 1'b1;
    layer5_outputs(6949) <= b and not a;
    layer5_outputs(6950) <= b;
    layer5_outputs(6951) <= a and b;
    layer5_outputs(6952) <= b;
    layer5_outputs(6953) <= not b;
    layer5_outputs(6954) <= a and b;
    layer5_outputs(6955) <= not a;
    layer5_outputs(6956) <= a and b;
    layer5_outputs(6957) <= not a or b;
    layer5_outputs(6958) <= not (a and b);
    layer5_outputs(6959) <= b;
    layer5_outputs(6960) <= a;
    layer5_outputs(6961) <= not b or a;
    layer5_outputs(6962) <= a or b;
    layer5_outputs(6963) <= 1'b1;
    layer5_outputs(6964) <= 1'b0;
    layer5_outputs(6965) <= b;
    layer5_outputs(6966) <= b;
    layer5_outputs(6967) <= b;
    layer5_outputs(6968) <= b;
    layer5_outputs(6969) <= not a;
    layer5_outputs(6970) <= not (a and b);
    layer5_outputs(6971) <= not (a or b);
    layer5_outputs(6972) <= not b;
    layer5_outputs(6973) <= not b or a;
    layer5_outputs(6974) <= a or b;
    layer5_outputs(6975) <= 1'b1;
    layer5_outputs(6976) <= not a;
    layer5_outputs(6977) <= not (a or b);
    layer5_outputs(6978) <= not b or a;
    layer5_outputs(6979) <= not a or b;
    layer5_outputs(6980) <= 1'b1;
    layer5_outputs(6981) <= not b;
    layer5_outputs(6982) <= not b;
    layer5_outputs(6983) <= not b;
    layer5_outputs(6984) <= 1'b0;
    layer5_outputs(6985) <= not b;
    layer5_outputs(6986) <= a or b;
    layer5_outputs(6987) <= 1'b1;
    layer5_outputs(6988) <= not b;
    layer5_outputs(6989) <= not b;
    layer5_outputs(6990) <= a or b;
    layer5_outputs(6991) <= not b or a;
    layer5_outputs(6992) <= not a;
    layer5_outputs(6993) <= a or b;
    layer5_outputs(6994) <= not (a or b);
    layer5_outputs(6995) <= a or b;
    layer5_outputs(6996) <= b;
    layer5_outputs(6997) <= b;
    layer5_outputs(6998) <= not (a xor b);
    layer5_outputs(6999) <= a and b;
    layer5_outputs(7000) <= not (a or b);
    layer5_outputs(7001) <= b;
    layer5_outputs(7002) <= 1'b1;
    layer5_outputs(7003) <= not a or b;
    layer5_outputs(7004) <= not b;
    layer5_outputs(7005) <= 1'b1;
    layer5_outputs(7006) <= b and not a;
    layer5_outputs(7007) <= a;
    layer5_outputs(7008) <= a or b;
    layer5_outputs(7009) <= a or b;
    layer5_outputs(7010) <= not b or a;
    layer5_outputs(7011) <= b;
    layer5_outputs(7012) <= not a;
    layer5_outputs(7013) <= not (a xor b);
    layer5_outputs(7014) <= b and not a;
    layer5_outputs(7015) <= not a or b;
    layer5_outputs(7016) <= 1'b0;
    layer5_outputs(7017) <= b and not a;
    layer5_outputs(7018) <= not a;
    layer5_outputs(7019) <= 1'b1;
    layer5_outputs(7020) <= a and b;
    layer5_outputs(7021) <= a;
    layer5_outputs(7022) <= a or b;
    layer5_outputs(7023) <= not b;
    layer5_outputs(7024) <= 1'b0;
    layer5_outputs(7025) <= 1'b1;
    layer5_outputs(7026) <= b and not a;
    layer5_outputs(7027) <= not b;
    layer5_outputs(7028) <= a xor b;
    layer5_outputs(7029) <= a and not b;
    layer5_outputs(7030) <= a;
    layer5_outputs(7031) <= b and not a;
    layer5_outputs(7032) <= not a;
    layer5_outputs(7033) <= not a;
    layer5_outputs(7034) <= not a;
    layer5_outputs(7035) <= not a;
    layer5_outputs(7036) <= not b;
    layer5_outputs(7037) <= 1'b1;
    layer5_outputs(7038) <= a xor b;
    layer5_outputs(7039) <= not a;
    layer5_outputs(7040) <= not b or a;
    layer5_outputs(7041) <= not a or b;
    layer5_outputs(7042) <= a and not b;
    layer5_outputs(7043) <= not (a and b);
    layer5_outputs(7044) <= not b;
    layer5_outputs(7045) <= not (a and b);
    layer5_outputs(7046) <= b;
    layer5_outputs(7047) <= not b;
    layer5_outputs(7048) <= a or b;
    layer5_outputs(7049) <= b;
    layer5_outputs(7050) <= a;
    layer5_outputs(7051) <= a and b;
    layer5_outputs(7052) <= not (a or b);
    layer5_outputs(7053) <= not a;
    layer5_outputs(7054) <= not (a or b);
    layer5_outputs(7055) <= b;
    layer5_outputs(7056) <= a and b;
    layer5_outputs(7057) <= a and b;
    layer5_outputs(7058) <= b;
    layer5_outputs(7059) <= a and b;
    layer5_outputs(7060) <= not (a or b);
    layer5_outputs(7061) <= 1'b0;
    layer5_outputs(7062) <= a or b;
    layer5_outputs(7063) <= not a;
    layer5_outputs(7064) <= a;
    layer5_outputs(7065) <= a or b;
    layer5_outputs(7066) <= b;
    layer5_outputs(7067) <= a and not b;
    layer5_outputs(7068) <= a or b;
    layer5_outputs(7069) <= not a or b;
    layer5_outputs(7070) <= not a;
    layer5_outputs(7071) <= not b;
    layer5_outputs(7072) <= not b;
    layer5_outputs(7073) <= not a;
    layer5_outputs(7074) <= 1'b1;
    layer5_outputs(7075) <= a and b;
    layer5_outputs(7076) <= not (a or b);
    layer5_outputs(7077) <= b;
    layer5_outputs(7078) <= 1'b0;
    layer5_outputs(7079) <= not b;
    layer5_outputs(7080) <= not b;
    layer5_outputs(7081) <= b and not a;
    layer5_outputs(7082) <= not (a or b);
    layer5_outputs(7083) <= b;
    layer5_outputs(7084) <= not b or a;
    layer5_outputs(7085) <= not a;
    layer5_outputs(7086) <= b;
    layer5_outputs(7087) <= b and not a;
    layer5_outputs(7088) <= not b or a;
    layer5_outputs(7089) <= not (a xor b);
    layer5_outputs(7090) <= not b or a;
    layer5_outputs(7091) <= b;
    layer5_outputs(7092) <= a and b;
    layer5_outputs(7093) <= not (a or b);
    layer5_outputs(7094) <= b;
    layer5_outputs(7095) <= b;
    layer5_outputs(7096) <= b;
    layer5_outputs(7097) <= not a or b;
    layer5_outputs(7098) <= a or b;
    layer5_outputs(7099) <= a xor b;
    layer5_outputs(7100) <= a or b;
    layer5_outputs(7101) <= not b;
    layer5_outputs(7102) <= 1'b1;
    layer5_outputs(7103) <= not a;
    layer5_outputs(7104) <= a and not b;
    layer5_outputs(7105) <= a and not b;
    layer5_outputs(7106) <= not (a and b);
    layer5_outputs(7107) <= a;
    layer5_outputs(7108) <= not b or a;
    layer5_outputs(7109) <= not a or b;
    layer5_outputs(7110) <= not b or a;
    layer5_outputs(7111) <= not a or b;
    layer5_outputs(7112) <= b and not a;
    layer5_outputs(7113) <= a and not b;
    layer5_outputs(7114) <= not (a or b);
    layer5_outputs(7115) <= a xor b;
    layer5_outputs(7116) <= not (a or b);
    layer5_outputs(7117) <= b;
    layer5_outputs(7118) <= not (a or b);
    layer5_outputs(7119) <= not b;
    layer5_outputs(7120) <= a or b;
    layer5_outputs(7121) <= 1'b1;
    layer5_outputs(7122) <= 1'b1;
    layer5_outputs(7123) <= a and b;
    layer5_outputs(7124) <= not a or b;
    layer5_outputs(7125) <= not b or a;
    layer5_outputs(7126) <= 1'b1;
    layer5_outputs(7127) <= not (a xor b);
    layer5_outputs(7128) <= a and b;
    layer5_outputs(7129) <= not a;
    layer5_outputs(7130) <= not a;
    layer5_outputs(7131) <= not a;
    layer5_outputs(7132) <= not b or a;
    layer5_outputs(7133) <= b and not a;
    layer5_outputs(7134) <= not b or a;
    layer5_outputs(7135) <= not a;
    layer5_outputs(7136) <= 1'b0;
    layer5_outputs(7137) <= not a;
    layer5_outputs(7138) <= not b or a;
    layer5_outputs(7139) <= not b;
    layer5_outputs(7140) <= not b or a;
    layer5_outputs(7141) <= not (a xor b);
    layer5_outputs(7142) <= not (a or b);
    layer5_outputs(7143) <= 1'b0;
    layer5_outputs(7144) <= not a or b;
    layer5_outputs(7145) <= b;
    layer5_outputs(7146) <= a and not b;
    layer5_outputs(7147) <= not b or a;
    layer5_outputs(7148) <= not b or a;
    layer5_outputs(7149) <= not b or a;
    layer5_outputs(7150) <= a;
    layer5_outputs(7151) <= not b;
    layer5_outputs(7152) <= b;
    layer5_outputs(7153) <= not (a and b);
    layer5_outputs(7154) <= not b;
    layer5_outputs(7155) <= a xor b;
    layer5_outputs(7156) <= not b;
    layer5_outputs(7157) <= a or b;
    layer5_outputs(7158) <= a or b;
    layer5_outputs(7159) <= not a or b;
    layer5_outputs(7160) <= not b or a;
    layer5_outputs(7161) <= not (a xor b);
    layer5_outputs(7162) <= a or b;
    layer5_outputs(7163) <= a and b;
    layer5_outputs(7164) <= not a;
    layer5_outputs(7165) <= not b;
    layer5_outputs(7166) <= not (a or b);
    layer5_outputs(7167) <= b and not a;
    layer5_outputs(7168) <= b;
    layer5_outputs(7169) <= not (a xor b);
    layer5_outputs(7170) <= 1'b1;
    layer5_outputs(7171) <= a;
    layer5_outputs(7172) <= not (a xor b);
    layer5_outputs(7173) <= not a;
    layer5_outputs(7174) <= 1'b1;
    layer5_outputs(7175) <= a or b;
    layer5_outputs(7176) <= a;
    layer5_outputs(7177) <= not b;
    layer5_outputs(7178) <= a xor b;
    layer5_outputs(7179) <= b;
    layer5_outputs(7180) <= not b;
    layer5_outputs(7181) <= not (a or b);
    layer5_outputs(7182) <= not (a and b);
    layer5_outputs(7183) <= not (a or b);
    layer5_outputs(7184) <= not (a and b);
    layer5_outputs(7185) <= not a;
    layer5_outputs(7186) <= not a or b;
    layer5_outputs(7187) <= not (a and b);
    layer5_outputs(7188) <= not (a or b);
    layer5_outputs(7189) <= a and b;
    layer5_outputs(7190) <= a;
    layer5_outputs(7191) <= not b or a;
    layer5_outputs(7192) <= 1'b1;
    layer5_outputs(7193) <= not (a xor b);
    layer5_outputs(7194) <= b;
    layer5_outputs(7195) <= b and not a;
    layer5_outputs(7196) <= not b;
    layer5_outputs(7197) <= b;
    layer5_outputs(7198) <= not a;
    layer5_outputs(7199) <= not a;
    layer5_outputs(7200) <= not (a or b);
    layer5_outputs(7201) <= not a or b;
    layer5_outputs(7202) <= not a;
    layer5_outputs(7203) <= a and not b;
    layer5_outputs(7204) <= not a;
    layer5_outputs(7205) <= not b;
    layer5_outputs(7206) <= not a;
    layer5_outputs(7207) <= b;
    layer5_outputs(7208) <= not (a or b);
    layer5_outputs(7209) <= a or b;
    layer5_outputs(7210) <= a and b;
    layer5_outputs(7211) <= 1'b0;
    layer5_outputs(7212) <= b;
    layer5_outputs(7213) <= a or b;
    layer5_outputs(7214) <= not a;
    layer5_outputs(7215) <= b;
    layer5_outputs(7216) <= a xor b;
    layer5_outputs(7217) <= 1'b0;
    layer5_outputs(7218) <= not a;
    layer5_outputs(7219) <= not b or a;
    layer5_outputs(7220) <= b;
    layer5_outputs(7221) <= b;
    layer5_outputs(7222) <= not a;
    layer5_outputs(7223) <= 1'b0;
    layer5_outputs(7224) <= not b;
    layer5_outputs(7225) <= b and not a;
    layer5_outputs(7226) <= a;
    layer5_outputs(7227) <= 1'b1;
    layer5_outputs(7228) <= b;
    layer5_outputs(7229) <= not (a or b);
    layer5_outputs(7230) <= not (a xor b);
    layer5_outputs(7231) <= a and not b;
    layer5_outputs(7232) <= not a;
    layer5_outputs(7233) <= not b;
    layer5_outputs(7234) <= not (a xor b);
    layer5_outputs(7235) <= not (a xor b);
    layer5_outputs(7236) <= b and not a;
    layer5_outputs(7237) <= a;
    layer5_outputs(7238) <= not (a and b);
    layer5_outputs(7239) <= a xor b;
    layer5_outputs(7240) <= a and b;
    layer5_outputs(7241) <= b;
    layer5_outputs(7242) <= a;
    layer5_outputs(7243) <= not b;
    layer5_outputs(7244) <= a xor b;
    layer5_outputs(7245) <= not a;
    layer5_outputs(7246) <= 1'b0;
    layer5_outputs(7247) <= a;
    layer5_outputs(7248) <= 1'b0;
    layer5_outputs(7249) <= not (a or b);
    layer5_outputs(7250) <= not a;
    layer5_outputs(7251) <= a xor b;
    layer5_outputs(7252) <= 1'b0;
    layer5_outputs(7253) <= not a or b;
    layer5_outputs(7254) <= a or b;
    layer5_outputs(7255) <= 1'b1;
    layer5_outputs(7256) <= a;
    layer5_outputs(7257) <= a or b;
    layer5_outputs(7258) <= not (a and b);
    layer5_outputs(7259) <= b and not a;
    layer5_outputs(7260) <= b;
    layer5_outputs(7261) <= b;
    layer5_outputs(7262) <= not b;
    layer5_outputs(7263) <= a;
    layer5_outputs(7264) <= not b or a;
    layer5_outputs(7265) <= not b or a;
    layer5_outputs(7266) <= not b;
    layer5_outputs(7267) <= not b;
    layer5_outputs(7268) <= a;
    layer5_outputs(7269) <= b;
    layer5_outputs(7270) <= not a or b;
    layer5_outputs(7271) <= a xor b;
    layer5_outputs(7272) <= not (a or b);
    layer5_outputs(7273) <= b and not a;
    layer5_outputs(7274) <= not (a and b);
    layer5_outputs(7275) <= a xor b;
    layer5_outputs(7276) <= not b;
    layer5_outputs(7277) <= 1'b0;
    layer5_outputs(7278) <= 1'b1;
    layer5_outputs(7279) <= not b;
    layer5_outputs(7280) <= a or b;
    layer5_outputs(7281) <= a xor b;
    layer5_outputs(7282) <= not b or a;
    layer5_outputs(7283) <= a and b;
    layer5_outputs(7284) <= a and b;
    layer5_outputs(7285) <= b;
    layer5_outputs(7286) <= not (a and b);
    layer5_outputs(7287) <= not a or b;
    layer5_outputs(7288) <= a;
    layer5_outputs(7289) <= not (a and b);
    layer5_outputs(7290) <= not (a xor b);
    layer5_outputs(7291) <= not (a and b);
    layer5_outputs(7292) <= b;
    layer5_outputs(7293) <= not (a xor b);
    layer5_outputs(7294) <= 1'b0;
    layer5_outputs(7295) <= not b or a;
    layer5_outputs(7296) <= 1'b1;
    layer5_outputs(7297) <= b;
    layer5_outputs(7298) <= a;
    layer5_outputs(7299) <= a or b;
    layer5_outputs(7300) <= 1'b1;
    layer5_outputs(7301) <= not b or a;
    layer5_outputs(7302) <= not b;
    layer5_outputs(7303) <= not (a and b);
    layer5_outputs(7304) <= not b;
    layer5_outputs(7305) <= not b or a;
    layer5_outputs(7306) <= a and not b;
    layer5_outputs(7307) <= 1'b0;
    layer5_outputs(7308) <= b;
    layer5_outputs(7309) <= not (a and b);
    layer5_outputs(7310) <= 1'b0;
    layer5_outputs(7311) <= a and b;
    layer5_outputs(7312) <= a;
    layer5_outputs(7313) <= b;
    layer5_outputs(7314) <= not b;
    layer5_outputs(7315) <= 1'b1;
    layer5_outputs(7316) <= a xor b;
    layer5_outputs(7317) <= b and not a;
    layer5_outputs(7318) <= not b;
    layer5_outputs(7319) <= 1'b0;
    layer5_outputs(7320) <= not (a or b);
    layer5_outputs(7321) <= not b or a;
    layer5_outputs(7322) <= not (a or b);
    layer5_outputs(7323) <= 1'b1;
    layer5_outputs(7324) <= a or b;
    layer5_outputs(7325) <= a xor b;
    layer5_outputs(7326) <= not (a xor b);
    layer5_outputs(7327) <= a and not b;
    layer5_outputs(7328) <= not b or a;
    layer5_outputs(7329) <= a or b;
    layer5_outputs(7330) <= a;
    layer5_outputs(7331) <= a and b;
    layer5_outputs(7332) <= not b;
    layer5_outputs(7333) <= a and not b;
    layer5_outputs(7334) <= a;
    layer5_outputs(7335) <= 1'b0;
    layer5_outputs(7336) <= a;
    layer5_outputs(7337) <= not a or b;
    layer5_outputs(7338) <= a or b;
    layer5_outputs(7339) <= b;
    layer5_outputs(7340) <= b and not a;
    layer5_outputs(7341) <= not a or b;
    layer5_outputs(7342) <= 1'b0;
    layer5_outputs(7343) <= not a or b;
    layer5_outputs(7344) <= not (a and b);
    layer5_outputs(7345) <= a and not b;
    layer5_outputs(7346) <= not b or a;
    layer5_outputs(7347) <= not (a and b);
    layer5_outputs(7348) <= not b or a;
    layer5_outputs(7349) <= not a or b;
    layer5_outputs(7350) <= 1'b0;
    layer5_outputs(7351) <= a;
    layer5_outputs(7352) <= a;
    layer5_outputs(7353) <= not a or b;
    layer5_outputs(7354) <= b;
    layer5_outputs(7355) <= 1'b0;
    layer5_outputs(7356) <= a;
    layer5_outputs(7357) <= a and b;
    layer5_outputs(7358) <= not (a or b);
    layer5_outputs(7359) <= not b;
    layer5_outputs(7360) <= not (a and b);
    layer5_outputs(7361) <= not b;
    layer5_outputs(7362) <= b;
    layer5_outputs(7363) <= a;
    layer5_outputs(7364) <= not b;
    layer5_outputs(7365) <= not (a or b);
    layer5_outputs(7366) <= a xor b;
    layer5_outputs(7367) <= b;
    layer5_outputs(7368) <= a xor b;
    layer5_outputs(7369) <= a and not b;
    layer5_outputs(7370) <= b;
    layer5_outputs(7371) <= not b;
    layer5_outputs(7372) <= not a or b;
    layer5_outputs(7373) <= not b;
    layer5_outputs(7374) <= not b;
    layer5_outputs(7375) <= not a or b;
    layer5_outputs(7376) <= a and b;
    layer5_outputs(7377) <= a or b;
    layer5_outputs(7378) <= b;
    layer5_outputs(7379) <= b and not a;
    layer5_outputs(7380) <= not (a or b);
    layer5_outputs(7381) <= not (a xor b);
    layer5_outputs(7382) <= not a;
    layer5_outputs(7383) <= b;
    layer5_outputs(7384) <= b;
    layer5_outputs(7385) <= a xor b;
    layer5_outputs(7386) <= not (a or b);
    layer5_outputs(7387) <= not a;
    layer5_outputs(7388) <= a and not b;
    layer5_outputs(7389) <= b;
    layer5_outputs(7390) <= b and not a;
    layer5_outputs(7391) <= not a or b;
    layer5_outputs(7392) <= not b;
    layer5_outputs(7393) <= not (a or b);
    layer5_outputs(7394) <= not b;
    layer5_outputs(7395) <= not (a and b);
    layer5_outputs(7396) <= not a;
    layer5_outputs(7397) <= not b or a;
    layer5_outputs(7398) <= not a;
    layer5_outputs(7399) <= b;
    layer5_outputs(7400) <= a xor b;
    layer5_outputs(7401) <= not (a and b);
    layer5_outputs(7402) <= b;
    layer5_outputs(7403) <= not b or a;
    layer5_outputs(7404) <= a;
    layer5_outputs(7405) <= a and not b;
    layer5_outputs(7406) <= 1'b1;
    layer5_outputs(7407) <= not (a or b);
    layer5_outputs(7408) <= not b;
    layer5_outputs(7409) <= a;
    layer5_outputs(7410) <= not b;
    layer5_outputs(7411) <= not a or b;
    layer5_outputs(7412) <= b;
    layer5_outputs(7413) <= 1'b1;
    layer5_outputs(7414) <= not (a and b);
    layer5_outputs(7415) <= b;
    layer5_outputs(7416) <= a or b;
    layer5_outputs(7417) <= a and b;
    layer5_outputs(7418) <= not a;
    layer5_outputs(7419) <= b and not a;
    layer5_outputs(7420) <= a and not b;
    layer5_outputs(7421) <= b;
    layer5_outputs(7422) <= a xor b;
    layer5_outputs(7423) <= b;
    layer5_outputs(7424) <= not a;
    layer5_outputs(7425) <= not b or a;
    layer5_outputs(7426) <= not b;
    layer5_outputs(7427) <= not (a or b);
    layer5_outputs(7428) <= not a or b;
    layer5_outputs(7429) <= a;
    layer5_outputs(7430) <= not b or a;
    layer5_outputs(7431) <= a or b;
    layer5_outputs(7432) <= b;
    layer5_outputs(7433) <= a and not b;
    layer5_outputs(7434) <= not a;
    layer5_outputs(7435) <= 1'b1;
    layer5_outputs(7436) <= a xor b;
    layer5_outputs(7437) <= a xor b;
    layer5_outputs(7438) <= not b or a;
    layer5_outputs(7439) <= a and b;
    layer5_outputs(7440) <= not (a and b);
    layer5_outputs(7441) <= a;
    layer5_outputs(7442) <= not b;
    layer5_outputs(7443) <= a and not b;
    layer5_outputs(7444) <= not (a or b);
    layer5_outputs(7445) <= b and not a;
    layer5_outputs(7446) <= not a;
    layer5_outputs(7447) <= not a;
    layer5_outputs(7448) <= not a or b;
    layer5_outputs(7449) <= a;
    layer5_outputs(7450) <= 1'b0;
    layer5_outputs(7451) <= a and not b;
    layer5_outputs(7452) <= a xor b;
    layer5_outputs(7453) <= b;
    layer5_outputs(7454) <= not (a xor b);
    layer5_outputs(7455) <= not (a xor b);
    layer5_outputs(7456) <= b;
    layer5_outputs(7457) <= a or b;
    layer5_outputs(7458) <= not (a or b);
    layer5_outputs(7459) <= a or b;
    layer5_outputs(7460) <= not a or b;
    layer5_outputs(7461) <= not a;
    layer5_outputs(7462) <= not b;
    layer5_outputs(7463) <= b;
    layer5_outputs(7464) <= 1'b0;
    layer5_outputs(7465) <= not (a or b);
    layer5_outputs(7466) <= not a;
    layer5_outputs(7467) <= not b;
    layer5_outputs(7468) <= not b;
    layer5_outputs(7469) <= not b;
    layer5_outputs(7470) <= not b or a;
    layer5_outputs(7471) <= not (a and b);
    layer5_outputs(7472) <= a or b;
    layer5_outputs(7473) <= not a or b;
    layer5_outputs(7474) <= b;
    layer5_outputs(7475) <= b and not a;
    layer5_outputs(7476) <= not b;
    layer5_outputs(7477) <= not (a xor b);
    layer5_outputs(7478) <= a;
    layer5_outputs(7479) <= not a or b;
    layer5_outputs(7480) <= not a;
    layer5_outputs(7481) <= not b;
    layer5_outputs(7482) <= a xor b;
    layer5_outputs(7483) <= not b or a;
    layer5_outputs(7484) <= a;
    layer5_outputs(7485) <= b;
    layer5_outputs(7486) <= not b or a;
    layer5_outputs(7487) <= a;
    layer5_outputs(7488) <= not b;
    layer5_outputs(7489) <= 1'b0;
    layer5_outputs(7490) <= a;
    layer5_outputs(7491) <= not (a and b);
    layer5_outputs(7492) <= not a;
    layer5_outputs(7493) <= a;
    layer5_outputs(7494) <= a;
    layer5_outputs(7495) <= not (a or b);
    layer5_outputs(7496) <= 1'b0;
    layer5_outputs(7497) <= not a or b;
    layer5_outputs(7498) <= not b;
    layer5_outputs(7499) <= not (a and b);
    layer5_outputs(7500) <= 1'b1;
    layer5_outputs(7501) <= a and not b;
    layer5_outputs(7502) <= a and not b;
    layer5_outputs(7503) <= b and not a;
    layer5_outputs(7504) <= 1'b1;
    layer5_outputs(7505) <= not a;
    layer5_outputs(7506) <= a and not b;
    layer5_outputs(7507) <= not (a or b);
    layer5_outputs(7508) <= b and not a;
    layer5_outputs(7509) <= b and not a;
    layer5_outputs(7510) <= 1'b1;
    layer5_outputs(7511) <= not (a or b);
    layer5_outputs(7512) <= not a;
    layer5_outputs(7513) <= a and not b;
    layer5_outputs(7514) <= b and not a;
    layer5_outputs(7515) <= b;
    layer5_outputs(7516) <= a and not b;
    layer5_outputs(7517) <= not (a or b);
    layer5_outputs(7518) <= a and not b;
    layer5_outputs(7519) <= not (a and b);
    layer5_outputs(7520) <= not b;
    layer5_outputs(7521) <= not b;
    layer5_outputs(7522) <= not (a and b);
    layer5_outputs(7523) <= not b or a;
    layer5_outputs(7524) <= not (a or b);
    layer5_outputs(7525) <= not b;
    layer5_outputs(7526) <= not b;
    layer5_outputs(7527) <= 1'b1;
    layer5_outputs(7528) <= not (a or b);
    layer5_outputs(7529) <= b;
    layer5_outputs(7530) <= a and b;
    layer5_outputs(7531) <= not b;
    layer5_outputs(7532) <= a;
    layer5_outputs(7533) <= a or b;
    layer5_outputs(7534) <= a and b;
    layer5_outputs(7535) <= b and not a;
    layer5_outputs(7536) <= not (a or b);
    layer5_outputs(7537) <= not b;
    layer5_outputs(7538) <= 1'b1;
    layer5_outputs(7539) <= a;
    layer5_outputs(7540) <= not (a and b);
    layer5_outputs(7541) <= a and not b;
    layer5_outputs(7542) <= not b or a;
    layer5_outputs(7543) <= a or b;
    layer5_outputs(7544) <= a and not b;
    layer5_outputs(7545) <= not a or b;
    layer5_outputs(7546) <= a and not b;
    layer5_outputs(7547) <= not b or a;
    layer5_outputs(7548) <= not (a or b);
    layer5_outputs(7549) <= not b;
    layer5_outputs(7550) <= a or b;
    layer5_outputs(7551) <= not a or b;
    layer5_outputs(7552) <= b and not a;
    layer5_outputs(7553) <= a or b;
    layer5_outputs(7554) <= a and not b;
    layer5_outputs(7555) <= b;
    layer5_outputs(7556) <= b;
    layer5_outputs(7557) <= a;
    layer5_outputs(7558) <= not a or b;
    layer5_outputs(7559) <= not a;
    layer5_outputs(7560) <= b;
    layer5_outputs(7561) <= a and b;
    layer5_outputs(7562) <= a and b;
    layer5_outputs(7563) <= a and b;
    layer5_outputs(7564) <= not b or a;
    layer5_outputs(7565) <= b;
    layer5_outputs(7566) <= not a;
    layer5_outputs(7567) <= not a;
    layer5_outputs(7568) <= not b or a;
    layer5_outputs(7569) <= 1'b1;
    layer5_outputs(7570) <= a or b;
    layer5_outputs(7571) <= not (a or b);
    layer5_outputs(7572) <= 1'b1;
    layer5_outputs(7573) <= a or b;
    layer5_outputs(7574) <= 1'b0;
    layer5_outputs(7575) <= 1'b0;
    layer5_outputs(7576) <= not b or a;
    layer5_outputs(7577) <= 1'b1;
    layer5_outputs(7578) <= not a or b;
    layer5_outputs(7579) <= not (a xor b);
    layer5_outputs(7580) <= b and not a;
    layer5_outputs(7581) <= b;
    layer5_outputs(7582) <= 1'b1;
    layer5_outputs(7583) <= not a or b;
    layer5_outputs(7584) <= b;
    layer5_outputs(7585) <= not b or a;
    layer5_outputs(7586) <= a xor b;
    layer5_outputs(7587) <= not a;
    layer5_outputs(7588) <= b;
    layer5_outputs(7589) <= a xor b;
    layer5_outputs(7590) <= a or b;
    layer5_outputs(7591) <= not (a or b);
    layer5_outputs(7592) <= not (a or b);
    layer5_outputs(7593) <= not a;
    layer5_outputs(7594) <= not (a xor b);
    layer5_outputs(7595) <= a or b;
    layer5_outputs(7596) <= not b;
    layer5_outputs(7597) <= a or b;
    layer5_outputs(7598) <= not a;
    layer5_outputs(7599) <= 1'b1;
    layer5_outputs(7600) <= b;
    layer5_outputs(7601) <= not b or a;
    layer5_outputs(7602) <= not a or b;
    layer5_outputs(7603) <= a;
    layer5_outputs(7604) <= 1'b0;
    layer5_outputs(7605) <= not b;
    layer5_outputs(7606) <= b and not a;
    layer5_outputs(7607) <= b;
    layer5_outputs(7608) <= not a;
    layer5_outputs(7609) <= not a or b;
    layer5_outputs(7610) <= a and not b;
    layer5_outputs(7611) <= not (a and b);
    layer5_outputs(7612) <= a;
    layer5_outputs(7613) <= b and not a;
    layer5_outputs(7614) <= not b or a;
    layer5_outputs(7615) <= a or b;
    layer5_outputs(7616) <= not a;
    layer5_outputs(7617) <= a;
    layer5_outputs(7618) <= not (a xor b);
    layer5_outputs(7619) <= not a;
    layer5_outputs(7620) <= b;
    layer5_outputs(7621) <= a and not b;
    layer5_outputs(7622) <= a and not b;
    layer5_outputs(7623) <= not b or a;
    layer5_outputs(7624) <= a;
    layer5_outputs(7625) <= a;
    layer5_outputs(7626) <= a or b;
    layer5_outputs(7627) <= a and b;
    layer5_outputs(7628) <= a;
    layer5_outputs(7629) <= not b or a;
    layer5_outputs(7630) <= a and not b;
    layer5_outputs(7631) <= not b;
    layer5_outputs(7632) <= not a or b;
    layer5_outputs(7633) <= b and not a;
    layer5_outputs(7634) <= a or b;
    layer5_outputs(7635) <= a;
    layer5_outputs(7636) <= a and b;
    layer5_outputs(7637) <= b and not a;
    layer5_outputs(7638) <= not (a and b);
    layer5_outputs(7639) <= 1'b0;
    layer5_outputs(7640) <= not a;
    layer5_outputs(7641) <= a;
    layer5_outputs(7642) <= not a;
    layer5_outputs(7643) <= b and not a;
    layer5_outputs(7644) <= a and b;
    layer5_outputs(7645) <= 1'b0;
    layer5_outputs(7646) <= a and b;
    layer5_outputs(7647) <= a or b;
    layer5_outputs(7648) <= a and b;
    layer5_outputs(7649) <= 1'b0;
    layer5_outputs(7650) <= not a;
    layer5_outputs(7651) <= not a;
    layer5_outputs(7652) <= a and not b;
    layer5_outputs(7653) <= not b;
    layer5_outputs(7654) <= not b or a;
    layer5_outputs(7655) <= 1'b0;
    layer5_outputs(7656) <= not b;
    layer5_outputs(7657) <= not (a or b);
    layer5_outputs(7658) <= 1'b0;
    layer5_outputs(7659) <= not b;
    layer5_outputs(7660) <= not a or b;
    layer5_outputs(7661) <= a or b;
    layer5_outputs(7662) <= not (a or b);
    layer5_outputs(7663) <= not a;
    layer5_outputs(7664) <= a and not b;
    layer5_outputs(7665) <= not (a or b);
    layer5_outputs(7666) <= not a;
    layer5_outputs(7667) <= 1'b1;
    layer5_outputs(7668) <= a;
    layer5_outputs(7669) <= a;
    layer5_outputs(7670) <= b;
    layer5_outputs(7671) <= a and b;
    layer5_outputs(7672) <= a and not b;
    layer5_outputs(7673) <= not b or a;
    layer5_outputs(7674) <= a;
    layer5_outputs(7675) <= a xor b;
    layer5_outputs(7676) <= not b;
    layer5_outputs(7677) <= not a;
    layer5_outputs(7678) <= a;
    layer5_outputs(7679) <= a or b;
    layer5_outputs(7680) <= not b or a;
    layer5_outputs(7681) <= not a;
    layer5_outputs(7682) <= not a;
    layer5_outputs(7683) <= a and b;
    layer5_outputs(7684) <= a and b;
    layer5_outputs(7685) <= not (a or b);
    layer5_outputs(7686) <= not b;
    layer5_outputs(7687) <= b;
    layer5_outputs(7688) <= not b or a;
    layer5_outputs(7689) <= b and not a;
    layer5_outputs(7690) <= not (a and b);
    layer5_outputs(7691) <= not (a or b);
    layer5_outputs(7692) <= a xor b;
    layer5_outputs(7693) <= not a or b;
    layer5_outputs(7694) <= b;
    layer5_outputs(7695) <= 1'b0;
    layer5_outputs(7696) <= a xor b;
    layer5_outputs(7697) <= a and not b;
    layer5_outputs(7698) <= not b;
    layer5_outputs(7699) <= a and not b;
    layer5_outputs(7700) <= not (a and b);
    layer5_outputs(7701) <= not (a and b);
    layer5_outputs(7702) <= b and not a;
    layer5_outputs(7703) <= not a;
    layer5_outputs(7704) <= a and not b;
    layer5_outputs(7705) <= not a or b;
    layer5_outputs(7706) <= a and b;
    layer5_outputs(7707) <= b;
    layer5_outputs(7708) <= not a or b;
    layer5_outputs(7709) <= not (a or b);
    layer5_outputs(7710) <= 1'b0;
    layer5_outputs(7711) <= a xor b;
    layer5_outputs(7712) <= a and b;
    layer5_outputs(7713) <= not (a xor b);
    layer5_outputs(7714) <= 1'b1;
    layer5_outputs(7715) <= not (a or b);
    layer5_outputs(7716) <= b and not a;
    layer5_outputs(7717) <= b and not a;
    layer5_outputs(7718) <= b and not a;
    layer5_outputs(7719) <= 1'b0;
    layer5_outputs(7720) <= not a or b;
    layer5_outputs(7721) <= a and not b;
    layer5_outputs(7722) <= b and not a;
    layer5_outputs(7723) <= a;
    layer5_outputs(7724) <= b and not a;
    layer5_outputs(7725) <= not (a and b);
    layer5_outputs(7726) <= b;
    layer5_outputs(7727) <= not (a or b);
    layer5_outputs(7728) <= not a or b;
    layer5_outputs(7729) <= a and not b;
    layer5_outputs(7730) <= 1'b0;
    layer5_outputs(7731) <= a and not b;
    layer5_outputs(7732) <= not (a or b);
    layer5_outputs(7733) <= a and b;
    layer5_outputs(7734) <= a or b;
    layer5_outputs(7735) <= not b;
    layer5_outputs(7736) <= 1'b1;
    layer5_outputs(7737) <= b and not a;
    layer5_outputs(7738) <= not (a or b);
    layer5_outputs(7739) <= a and not b;
    layer5_outputs(7740) <= a;
    layer5_outputs(7741) <= a xor b;
    layer5_outputs(7742) <= not b;
    layer5_outputs(7743) <= a;
    layer5_outputs(7744) <= not a;
    layer5_outputs(7745) <= not b;
    layer5_outputs(7746) <= not (a or b);
    layer5_outputs(7747) <= not b;
    layer5_outputs(7748) <= a or b;
    layer5_outputs(7749) <= not a;
    layer5_outputs(7750) <= a;
    layer5_outputs(7751) <= not a;
    layer5_outputs(7752) <= a;
    layer5_outputs(7753) <= 1'b0;
    layer5_outputs(7754) <= not b or a;
    layer5_outputs(7755) <= a;
    layer5_outputs(7756) <= a;
    layer5_outputs(7757) <= a and b;
    layer5_outputs(7758) <= a or b;
    layer5_outputs(7759) <= not a or b;
    layer5_outputs(7760) <= b;
    layer5_outputs(7761) <= a xor b;
    layer5_outputs(7762) <= b;
    layer5_outputs(7763) <= not a;
    layer5_outputs(7764) <= 1'b1;
    layer5_outputs(7765) <= not (a xor b);
    layer5_outputs(7766) <= not a or b;
    layer5_outputs(7767) <= not a;
    layer5_outputs(7768) <= a and not b;
    layer5_outputs(7769) <= not a;
    layer5_outputs(7770) <= not (a or b);
    layer5_outputs(7771) <= b;
    layer5_outputs(7772) <= not a;
    layer5_outputs(7773) <= b and not a;
    layer5_outputs(7774) <= not a;
    layer5_outputs(7775) <= not a or b;
    layer5_outputs(7776) <= b and not a;
    layer5_outputs(7777) <= not b;
    layer5_outputs(7778) <= b and not a;
    layer5_outputs(7779) <= a and b;
    layer5_outputs(7780) <= not (a or b);
    layer5_outputs(7781) <= not a;
    layer5_outputs(7782) <= a and b;
    layer5_outputs(7783) <= not a or b;
    layer5_outputs(7784) <= a xor b;
    layer5_outputs(7785) <= a and b;
    layer5_outputs(7786) <= not (a xor b);
    layer5_outputs(7787) <= b;
    layer5_outputs(7788) <= not (a or b);
    layer5_outputs(7789) <= a xor b;
    layer5_outputs(7790) <= a xor b;
    layer5_outputs(7791) <= 1'b0;
    layer5_outputs(7792) <= b and not a;
    layer5_outputs(7793) <= b;
    layer5_outputs(7794) <= a and not b;
    layer5_outputs(7795) <= not a;
    layer5_outputs(7796) <= not (a xor b);
    layer5_outputs(7797) <= not (a and b);
    layer5_outputs(7798) <= not (a and b);
    layer5_outputs(7799) <= not a;
    layer5_outputs(7800) <= b and not a;
    layer5_outputs(7801) <= not (a and b);
    layer5_outputs(7802) <= b;
    layer5_outputs(7803) <= not a or b;
    layer5_outputs(7804) <= 1'b0;
    layer5_outputs(7805) <= not (a xor b);
    layer5_outputs(7806) <= b and not a;
    layer5_outputs(7807) <= b;
    layer5_outputs(7808) <= b and not a;
    layer5_outputs(7809) <= not b;
    layer5_outputs(7810) <= b;
    layer5_outputs(7811) <= not a;
    layer5_outputs(7812) <= a;
    layer5_outputs(7813) <= a;
    layer5_outputs(7814) <= a;
    layer5_outputs(7815) <= a or b;
    layer5_outputs(7816) <= not b or a;
    layer5_outputs(7817) <= not b;
    layer5_outputs(7818) <= a or b;
    layer5_outputs(7819) <= not (a or b);
    layer5_outputs(7820) <= not (a or b);
    layer5_outputs(7821) <= b;
    layer5_outputs(7822) <= b;
    layer5_outputs(7823) <= a or b;
    layer5_outputs(7824) <= not (a and b);
    layer5_outputs(7825) <= a and not b;
    layer5_outputs(7826) <= a and b;
    layer5_outputs(7827) <= a or b;
    layer5_outputs(7828) <= a and b;
    layer5_outputs(7829) <= a and not b;
    layer5_outputs(7830) <= not (a or b);
    layer5_outputs(7831) <= not (a or b);
    layer5_outputs(7832) <= b and not a;
    layer5_outputs(7833) <= b;
    layer5_outputs(7834) <= a;
    layer5_outputs(7835) <= b and not a;
    layer5_outputs(7836) <= a;
    layer5_outputs(7837) <= not b;
    layer5_outputs(7838) <= 1'b0;
    layer5_outputs(7839) <= b and not a;
    layer5_outputs(7840) <= a xor b;
    layer5_outputs(7841) <= 1'b1;
    layer5_outputs(7842) <= a;
    layer5_outputs(7843) <= b and not a;
    layer5_outputs(7844) <= a;
    layer5_outputs(7845) <= not a or b;
    layer5_outputs(7846) <= 1'b0;
    layer5_outputs(7847) <= b;
    layer5_outputs(7848) <= not (a and b);
    layer5_outputs(7849) <= not b or a;
    layer5_outputs(7850) <= b;
    layer5_outputs(7851) <= not a or b;
    layer5_outputs(7852) <= not b;
    layer5_outputs(7853) <= not a or b;
    layer5_outputs(7854) <= a xor b;
    layer5_outputs(7855) <= not (a xor b);
    layer5_outputs(7856) <= not a;
    layer5_outputs(7857) <= not a or b;
    layer5_outputs(7858) <= not (a and b);
    layer5_outputs(7859) <= a and not b;
    layer5_outputs(7860) <= b and not a;
    layer5_outputs(7861) <= b;
    layer5_outputs(7862) <= not b;
    layer5_outputs(7863) <= not (a and b);
    layer5_outputs(7864) <= 1'b0;
    layer5_outputs(7865) <= a and not b;
    layer5_outputs(7866) <= 1'b1;
    layer5_outputs(7867) <= a;
    layer5_outputs(7868) <= not b;
    layer5_outputs(7869) <= not b;
    layer5_outputs(7870) <= not a or b;
    layer5_outputs(7871) <= a;
    layer5_outputs(7872) <= not (a or b);
    layer5_outputs(7873) <= not b or a;
    layer5_outputs(7874) <= b;
    layer5_outputs(7875) <= a;
    layer5_outputs(7876) <= a xor b;
    layer5_outputs(7877) <= b and not a;
    layer5_outputs(7878) <= not (a or b);
    layer5_outputs(7879) <= not b or a;
    layer5_outputs(7880) <= not a or b;
    layer5_outputs(7881) <= b;
    layer5_outputs(7882) <= not b;
    layer5_outputs(7883) <= not b or a;
    layer5_outputs(7884) <= b;
    layer5_outputs(7885) <= 1'b1;
    layer5_outputs(7886) <= not a or b;
    layer5_outputs(7887) <= not (a and b);
    layer5_outputs(7888) <= not b or a;
    layer5_outputs(7889) <= a or b;
    layer5_outputs(7890) <= 1'b0;
    layer5_outputs(7891) <= a;
    layer5_outputs(7892) <= not (a and b);
    layer5_outputs(7893) <= a or b;
    layer5_outputs(7894) <= 1'b0;
    layer5_outputs(7895) <= not a;
    layer5_outputs(7896) <= b;
    layer5_outputs(7897) <= a and not b;
    layer5_outputs(7898) <= a xor b;
    layer5_outputs(7899) <= b;
    layer5_outputs(7900) <= not a or b;
    layer5_outputs(7901) <= not b or a;
    layer5_outputs(7902) <= b;
    layer5_outputs(7903) <= not b or a;
    layer5_outputs(7904) <= not b;
    layer5_outputs(7905) <= not (a and b);
    layer5_outputs(7906) <= a and b;
    layer5_outputs(7907) <= a;
    layer5_outputs(7908) <= b and not a;
    layer5_outputs(7909) <= a;
    layer5_outputs(7910) <= not (a and b);
    layer5_outputs(7911) <= b and not a;
    layer5_outputs(7912) <= not (a and b);
    layer5_outputs(7913) <= not a or b;
    layer5_outputs(7914) <= b and not a;
    layer5_outputs(7915) <= b and not a;
    layer5_outputs(7916) <= not (a and b);
    layer5_outputs(7917) <= not b;
    layer5_outputs(7918) <= not b or a;
    layer5_outputs(7919) <= b;
    layer5_outputs(7920) <= a;
    layer5_outputs(7921) <= a and not b;
    layer5_outputs(7922) <= b;
    layer5_outputs(7923) <= not b;
    layer5_outputs(7924) <= not (a and b);
    layer5_outputs(7925) <= not (a and b);
    layer5_outputs(7926) <= not (a or b);
    layer5_outputs(7927) <= not a;
    layer5_outputs(7928) <= not a;
    layer5_outputs(7929) <= not b;
    layer5_outputs(7930) <= 1'b1;
    layer5_outputs(7931) <= not b;
    layer5_outputs(7932) <= a or b;
    layer5_outputs(7933) <= b and not a;
    layer5_outputs(7934) <= a or b;
    layer5_outputs(7935) <= not a or b;
    layer5_outputs(7936) <= not b;
    layer5_outputs(7937) <= b;
    layer5_outputs(7938) <= a xor b;
    layer5_outputs(7939) <= a and not b;
    layer5_outputs(7940) <= 1'b1;
    layer5_outputs(7941) <= a;
    layer5_outputs(7942) <= not b;
    layer5_outputs(7943) <= not (a and b);
    layer5_outputs(7944) <= not (a xor b);
    layer5_outputs(7945) <= a xor b;
    layer5_outputs(7946) <= not a;
    layer5_outputs(7947) <= a xor b;
    layer5_outputs(7948) <= not (a and b);
    layer5_outputs(7949) <= not a;
    layer5_outputs(7950) <= a;
    layer5_outputs(7951) <= a;
    layer5_outputs(7952) <= 1'b1;
    layer5_outputs(7953) <= not (a xor b);
    layer5_outputs(7954) <= a;
    layer5_outputs(7955) <= a xor b;
    layer5_outputs(7956) <= a xor b;
    layer5_outputs(7957) <= not a;
    layer5_outputs(7958) <= not a;
    layer5_outputs(7959) <= b and not a;
    layer5_outputs(7960) <= a and not b;
    layer5_outputs(7961) <= not b;
    layer5_outputs(7962) <= not (a xor b);
    layer5_outputs(7963) <= not a or b;
    layer5_outputs(7964) <= not b;
    layer5_outputs(7965) <= not a;
    layer5_outputs(7966) <= 1'b1;
    layer5_outputs(7967) <= not a or b;
    layer5_outputs(7968) <= not (a and b);
    layer5_outputs(7969) <= not (a xor b);
    layer5_outputs(7970) <= not b;
    layer5_outputs(7971) <= not a or b;
    layer5_outputs(7972) <= not a;
    layer5_outputs(7973) <= not b;
    layer5_outputs(7974) <= not a or b;
    layer5_outputs(7975) <= not b;
    layer5_outputs(7976) <= not (a or b);
    layer5_outputs(7977) <= a or b;
    layer5_outputs(7978) <= not b or a;
    layer5_outputs(7979) <= not (a xor b);
    layer5_outputs(7980) <= a xor b;
    layer5_outputs(7981) <= b;
    layer5_outputs(7982) <= not b;
    layer5_outputs(7983) <= a or b;
    layer5_outputs(7984) <= a;
    layer5_outputs(7985) <= a and b;
    layer5_outputs(7986) <= not (a or b);
    layer5_outputs(7987) <= a and b;
    layer5_outputs(7988) <= b and not a;
    layer5_outputs(7989) <= not (a and b);
    layer5_outputs(7990) <= 1'b1;
    layer5_outputs(7991) <= a and not b;
    layer5_outputs(7992) <= not (a xor b);
    layer5_outputs(7993) <= b;
    layer5_outputs(7994) <= a xor b;
    layer5_outputs(7995) <= not (a xor b);
    layer5_outputs(7996) <= not (a or b);
    layer5_outputs(7997) <= not a;
    layer5_outputs(7998) <= a and not b;
    layer5_outputs(7999) <= not (a and b);
    layer5_outputs(8000) <= b and not a;
    layer5_outputs(8001) <= a or b;
    layer5_outputs(8002) <= not (a or b);
    layer5_outputs(8003) <= not a or b;
    layer5_outputs(8004) <= a xor b;
    layer5_outputs(8005) <= a;
    layer5_outputs(8006) <= not a;
    layer5_outputs(8007) <= a and not b;
    layer5_outputs(8008) <= b and not a;
    layer5_outputs(8009) <= 1'b0;
    layer5_outputs(8010) <= not (a and b);
    layer5_outputs(8011) <= 1'b1;
    layer5_outputs(8012) <= not (a xor b);
    layer5_outputs(8013) <= not (a xor b);
    layer5_outputs(8014) <= not (a and b);
    layer5_outputs(8015) <= a or b;
    layer5_outputs(8016) <= a;
    layer5_outputs(8017) <= not (a and b);
    layer5_outputs(8018) <= a;
    layer5_outputs(8019) <= a or b;
    layer5_outputs(8020) <= not (a xor b);
    layer5_outputs(8021) <= b and not a;
    layer5_outputs(8022) <= a;
    layer5_outputs(8023) <= not b;
    layer5_outputs(8024) <= not a or b;
    layer5_outputs(8025) <= not b;
    layer5_outputs(8026) <= b and not a;
    layer5_outputs(8027) <= not (a and b);
    layer5_outputs(8028) <= not b;
    layer5_outputs(8029) <= a and not b;
    layer5_outputs(8030) <= a and b;
    layer5_outputs(8031) <= a xor b;
    layer5_outputs(8032) <= a and b;
    layer5_outputs(8033) <= not a;
    layer5_outputs(8034) <= 1'b0;
    layer5_outputs(8035) <= not (a xor b);
    layer5_outputs(8036) <= a;
    layer5_outputs(8037) <= not (a and b);
    layer5_outputs(8038) <= not a or b;
    layer5_outputs(8039) <= not (a xor b);
    layer5_outputs(8040) <= a or b;
    layer5_outputs(8041) <= b;
    layer5_outputs(8042) <= 1'b0;
    layer5_outputs(8043) <= b;
    layer5_outputs(8044) <= not b;
    layer5_outputs(8045) <= not a;
    layer5_outputs(8046) <= a;
    layer5_outputs(8047) <= not b;
    layer5_outputs(8048) <= not a;
    layer5_outputs(8049) <= not a;
    layer5_outputs(8050) <= a xor b;
    layer5_outputs(8051) <= a and not b;
    layer5_outputs(8052) <= not (a or b);
    layer5_outputs(8053) <= 1'b0;
    layer5_outputs(8054) <= b and not a;
    layer5_outputs(8055) <= not a;
    layer5_outputs(8056) <= not (a xor b);
    layer5_outputs(8057) <= not b;
    layer5_outputs(8058) <= a or b;
    layer5_outputs(8059) <= not (a and b);
    layer5_outputs(8060) <= not a;
    layer5_outputs(8061) <= 1'b0;
    layer5_outputs(8062) <= a;
    layer5_outputs(8063) <= not (a and b);
    layer5_outputs(8064) <= b;
    layer5_outputs(8065) <= a and b;
    layer5_outputs(8066) <= not a;
    layer5_outputs(8067) <= not a or b;
    layer5_outputs(8068) <= b and not a;
    layer5_outputs(8069) <= a;
    layer5_outputs(8070) <= a xor b;
    layer5_outputs(8071) <= not b;
    layer5_outputs(8072) <= not (a and b);
    layer5_outputs(8073) <= a;
    layer5_outputs(8074) <= b;
    layer5_outputs(8075) <= a and b;
    layer5_outputs(8076) <= not a;
    layer5_outputs(8077) <= a xor b;
    layer5_outputs(8078) <= b;
    layer5_outputs(8079) <= a;
    layer5_outputs(8080) <= b and not a;
    layer5_outputs(8081) <= b;
    layer5_outputs(8082) <= a;
    layer5_outputs(8083) <= a and b;
    layer5_outputs(8084) <= not b or a;
    layer5_outputs(8085) <= not (a or b);
    layer5_outputs(8086) <= not a;
    layer5_outputs(8087) <= not (a xor b);
    layer5_outputs(8088) <= not a or b;
    layer5_outputs(8089) <= b;
    layer5_outputs(8090) <= a xor b;
    layer5_outputs(8091) <= a;
    layer5_outputs(8092) <= not a;
    layer5_outputs(8093) <= not (a xor b);
    layer5_outputs(8094) <= 1'b1;
    layer5_outputs(8095) <= b;
    layer5_outputs(8096) <= not (a and b);
    layer5_outputs(8097) <= not (a or b);
    layer5_outputs(8098) <= b;
    layer5_outputs(8099) <= not b;
    layer5_outputs(8100) <= not a or b;
    layer5_outputs(8101) <= not b or a;
    layer5_outputs(8102) <= a and not b;
    layer5_outputs(8103) <= a and not b;
    layer5_outputs(8104) <= b;
    layer5_outputs(8105) <= a or b;
    layer5_outputs(8106) <= 1'b1;
    layer5_outputs(8107) <= b and not a;
    layer5_outputs(8108) <= not a;
    layer5_outputs(8109) <= not a or b;
    layer5_outputs(8110) <= a;
    layer5_outputs(8111) <= a and b;
    layer5_outputs(8112) <= not a;
    layer5_outputs(8113) <= a or b;
    layer5_outputs(8114) <= a or b;
    layer5_outputs(8115) <= not (a or b);
    layer5_outputs(8116) <= not a;
    layer5_outputs(8117) <= 1'b0;
    layer5_outputs(8118) <= not (a or b);
    layer5_outputs(8119) <= a or b;
    layer5_outputs(8120) <= b;
    layer5_outputs(8121) <= a and not b;
    layer5_outputs(8122) <= a;
    layer5_outputs(8123) <= not a;
    layer5_outputs(8124) <= not (a or b);
    layer5_outputs(8125) <= a and not b;
    layer5_outputs(8126) <= not (a xor b);
    layer5_outputs(8127) <= b and not a;
    layer5_outputs(8128) <= not b or a;
    layer5_outputs(8129) <= not b;
    layer5_outputs(8130) <= not a or b;
    layer5_outputs(8131) <= a xor b;
    layer5_outputs(8132) <= 1'b1;
    layer5_outputs(8133) <= a and not b;
    layer5_outputs(8134) <= a and not b;
    layer5_outputs(8135) <= 1'b0;
    layer5_outputs(8136) <= not b;
    layer5_outputs(8137) <= not a or b;
    layer5_outputs(8138) <= not (a or b);
    layer5_outputs(8139) <= not (a or b);
    layer5_outputs(8140) <= not (a xor b);
    layer5_outputs(8141) <= 1'b1;
    layer5_outputs(8142) <= a and not b;
    layer5_outputs(8143) <= b;
    layer5_outputs(8144) <= not a;
    layer5_outputs(8145) <= not a;
    layer5_outputs(8146) <= b;
    layer5_outputs(8147) <= b and not a;
    layer5_outputs(8148) <= b and not a;
    layer5_outputs(8149) <= a xor b;
    layer5_outputs(8150) <= b;
    layer5_outputs(8151) <= not (a xor b);
    layer5_outputs(8152) <= not a or b;
    layer5_outputs(8153) <= not a or b;
    layer5_outputs(8154) <= a and not b;
    layer5_outputs(8155) <= not a or b;
    layer5_outputs(8156) <= not a;
    layer5_outputs(8157) <= not b or a;
    layer5_outputs(8158) <= a and not b;
    layer5_outputs(8159) <= a and b;
    layer5_outputs(8160) <= a;
    layer5_outputs(8161) <= a and not b;
    layer5_outputs(8162) <= not b;
    layer5_outputs(8163) <= not (a or b);
    layer5_outputs(8164) <= a or b;
    layer5_outputs(8165) <= not (a xor b);
    layer5_outputs(8166) <= not a;
    layer5_outputs(8167) <= a;
    layer5_outputs(8168) <= b;
    layer5_outputs(8169) <= a and not b;
    layer5_outputs(8170) <= a or b;
    layer5_outputs(8171) <= 1'b1;
    layer5_outputs(8172) <= 1'b0;
    layer5_outputs(8173) <= not b;
    layer5_outputs(8174) <= a xor b;
    layer5_outputs(8175) <= not b or a;
    layer5_outputs(8176) <= a and b;
    layer5_outputs(8177) <= b;
    layer5_outputs(8178) <= a and not b;
    layer5_outputs(8179) <= not b;
    layer5_outputs(8180) <= not b;
    layer5_outputs(8181) <= not a or b;
    layer5_outputs(8182) <= a;
    layer5_outputs(8183) <= not (a or b);
    layer5_outputs(8184) <= not (a and b);
    layer5_outputs(8185) <= a and not b;
    layer5_outputs(8186) <= not b;
    layer5_outputs(8187) <= b;
    layer5_outputs(8188) <= not a or b;
    layer5_outputs(8189) <= b and not a;
    layer5_outputs(8190) <= b and not a;
    layer5_outputs(8191) <= not b or a;
    layer5_outputs(8192) <= a;
    layer5_outputs(8193) <= not a;
    layer5_outputs(8194) <= not (a and b);
    layer5_outputs(8195) <= a;
    layer5_outputs(8196) <= not b;
    layer5_outputs(8197) <= not (a or b);
    layer5_outputs(8198) <= a;
    layer5_outputs(8199) <= not a;
    layer5_outputs(8200) <= a or b;
    layer5_outputs(8201) <= not b;
    layer5_outputs(8202) <= a or b;
    layer5_outputs(8203) <= not (a and b);
    layer5_outputs(8204) <= b;
    layer5_outputs(8205) <= not (a or b);
    layer5_outputs(8206) <= b;
    layer5_outputs(8207) <= a;
    layer5_outputs(8208) <= a;
    layer5_outputs(8209) <= a or b;
    layer5_outputs(8210) <= 1'b1;
    layer5_outputs(8211) <= not (a or b);
    layer5_outputs(8212) <= not b;
    layer5_outputs(8213) <= a;
    layer5_outputs(8214) <= b and not a;
    layer5_outputs(8215) <= not a;
    layer5_outputs(8216) <= not (a or b);
    layer5_outputs(8217) <= not a;
    layer5_outputs(8218) <= a;
    layer5_outputs(8219) <= a;
    layer5_outputs(8220) <= b;
    layer5_outputs(8221) <= a and not b;
    layer5_outputs(8222) <= 1'b1;
    layer5_outputs(8223) <= b;
    layer5_outputs(8224) <= not b;
    layer5_outputs(8225) <= 1'b0;
    layer5_outputs(8226) <= not (a xor b);
    layer5_outputs(8227) <= a;
    layer5_outputs(8228) <= a;
    layer5_outputs(8229) <= not a or b;
    layer5_outputs(8230) <= a or b;
    layer5_outputs(8231) <= not (a or b);
    layer5_outputs(8232) <= b;
    layer5_outputs(8233) <= b;
    layer5_outputs(8234) <= not b;
    layer5_outputs(8235) <= not (a and b);
    layer5_outputs(8236) <= not (a or b);
    layer5_outputs(8237) <= not (a or b);
    layer5_outputs(8238) <= not a;
    layer5_outputs(8239) <= a;
    layer5_outputs(8240) <= a or b;
    layer5_outputs(8241) <= a and not b;
    layer5_outputs(8242) <= not a or b;
    layer5_outputs(8243) <= b;
    layer5_outputs(8244) <= not a;
    layer5_outputs(8245) <= not (a or b);
    layer5_outputs(8246) <= b;
    layer5_outputs(8247) <= not b or a;
    layer5_outputs(8248) <= a and not b;
    layer5_outputs(8249) <= 1'b1;
    layer5_outputs(8250) <= a and not b;
    layer5_outputs(8251) <= b;
    layer5_outputs(8252) <= a or b;
    layer5_outputs(8253) <= b and not a;
    layer5_outputs(8254) <= a;
    layer5_outputs(8255) <= not (a or b);
    layer5_outputs(8256) <= not (a and b);
    layer5_outputs(8257) <= a and b;
    layer5_outputs(8258) <= not b or a;
    layer5_outputs(8259) <= a and b;
    layer5_outputs(8260) <= not b;
    layer5_outputs(8261) <= b;
    layer5_outputs(8262) <= a and not b;
    layer5_outputs(8263) <= not b or a;
    layer5_outputs(8264) <= not b;
    layer5_outputs(8265) <= not (a and b);
    layer5_outputs(8266) <= a and b;
    layer5_outputs(8267) <= a or b;
    layer5_outputs(8268) <= not (a and b);
    layer5_outputs(8269) <= not a;
    layer5_outputs(8270) <= b;
    layer5_outputs(8271) <= b;
    layer5_outputs(8272) <= b and not a;
    layer5_outputs(8273) <= not b;
    layer5_outputs(8274) <= a and not b;
    layer5_outputs(8275) <= not b;
    layer5_outputs(8276) <= not a;
    layer5_outputs(8277) <= not (a or b);
    layer5_outputs(8278) <= a xor b;
    layer5_outputs(8279) <= b;
    layer5_outputs(8280) <= not a;
    layer5_outputs(8281) <= a or b;
    layer5_outputs(8282) <= a and b;
    layer5_outputs(8283) <= not a;
    layer5_outputs(8284) <= b;
    layer5_outputs(8285) <= not b;
    layer5_outputs(8286) <= not b or a;
    layer5_outputs(8287) <= b;
    layer5_outputs(8288) <= b and not a;
    layer5_outputs(8289) <= not a;
    layer5_outputs(8290) <= a;
    layer5_outputs(8291) <= b;
    layer5_outputs(8292) <= a;
    layer5_outputs(8293) <= not (a or b);
    layer5_outputs(8294) <= not a;
    layer5_outputs(8295) <= a;
    layer5_outputs(8296) <= not a;
    layer5_outputs(8297) <= a xor b;
    layer5_outputs(8298) <= not b or a;
    layer5_outputs(8299) <= 1'b1;
    layer5_outputs(8300) <= not a;
    layer5_outputs(8301) <= a and b;
    layer5_outputs(8302) <= a;
    layer5_outputs(8303) <= a or b;
    layer5_outputs(8304) <= not a or b;
    layer5_outputs(8305) <= not (a or b);
    layer5_outputs(8306) <= not (a and b);
    layer5_outputs(8307) <= not a or b;
    layer5_outputs(8308) <= a or b;
    layer5_outputs(8309) <= a;
    layer5_outputs(8310) <= a or b;
    layer5_outputs(8311) <= not a;
    layer5_outputs(8312) <= a and b;
    layer5_outputs(8313) <= a xor b;
    layer5_outputs(8314) <= not a or b;
    layer5_outputs(8315) <= a and not b;
    layer5_outputs(8316) <= b and not a;
    layer5_outputs(8317) <= a and not b;
    layer5_outputs(8318) <= b and not a;
    layer5_outputs(8319) <= b;
    layer5_outputs(8320) <= a;
    layer5_outputs(8321) <= a xor b;
    layer5_outputs(8322) <= not b or a;
    layer5_outputs(8323) <= not a;
    layer5_outputs(8324) <= a xor b;
    layer5_outputs(8325) <= a and b;
    layer5_outputs(8326) <= not a;
    layer5_outputs(8327) <= not a;
    layer5_outputs(8328) <= b and not a;
    layer5_outputs(8329) <= a and not b;
    layer5_outputs(8330) <= not b;
    layer5_outputs(8331) <= 1'b0;
    layer5_outputs(8332) <= b;
    layer5_outputs(8333) <= not (a xor b);
    layer5_outputs(8334) <= a and not b;
    layer5_outputs(8335) <= 1'b0;
    layer5_outputs(8336) <= not b;
    layer5_outputs(8337) <= b;
    layer5_outputs(8338) <= not a;
    layer5_outputs(8339) <= not b;
    layer5_outputs(8340) <= not b;
    layer5_outputs(8341) <= not b;
    layer5_outputs(8342) <= not a or b;
    layer5_outputs(8343) <= a and b;
    layer5_outputs(8344) <= 1'b0;
    layer5_outputs(8345) <= a;
    layer5_outputs(8346) <= not b or a;
    layer5_outputs(8347) <= a and b;
    layer5_outputs(8348) <= not b or a;
    layer5_outputs(8349) <= 1'b1;
    layer5_outputs(8350) <= not a or b;
    layer5_outputs(8351) <= not b;
    layer5_outputs(8352) <= b;
    layer5_outputs(8353) <= not b;
    layer5_outputs(8354) <= a or b;
    layer5_outputs(8355) <= not a;
    layer5_outputs(8356) <= a and b;
    layer5_outputs(8357) <= a;
    layer5_outputs(8358) <= not (a and b);
    layer5_outputs(8359) <= not b;
    layer5_outputs(8360) <= a or b;
    layer5_outputs(8361) <= not (a xor b);
    layer5_outputs(8362) <= a;
    layer5_outputs(8363) <= not a;
    layer5_outputs(8364) <= not b;
    layer5_outputs(8365) <= not (a or b);
    layer5_outputs(8366) <= b and not a;
    layer5_outputs(8367) <= a or b;
    layer5_outputs(8368) <= not (a xor b);
    layer5_outputs(8369) <= a and b;
    layer5_outputs(8370) <= not b or a;
    layer5_outputs(8371) <= 1'b1;
    layer5_outputs(8372) <= a;
    layer5_outputs(8373) <= a and b;
    layer5_outputs(8374) <= not (a xor b);
    layer5_outputs(8375) <= a and not b;
    layer5_outputs(8376) <= 1'b0;
    layer5_outputs(8377) <= a xor b;
    layer5_outputs(8378) <= not a;
    layer5_outputs(8379) <= not b;
    layer5_outputs(8380) <= a;
    layer5_outputs(8381) <= b and not a;
    layer5_outputs(8382) <= not b;
    layer5_outputs(8383) <= a xor b;
    layer5_outputs(8384) <= not (a xor b);
    layer5_outputs(8385) <= b;
    layer5_outputs(8386) <= a;
    layer5_outputs(8387) <= a and not b;
    layer5_outputs(8388) <= a;
    layer5_outputs(8389) <= not b;
    layer5_outputs(8390) <= b and not a;
    layer5_outputs(8391) <= not (a or b);
    layer5_outputs(8392) <= a;
    layer5_outputs(8393) <= b;
    layer5_outputs(8394) <= 1'b0;
    layer5_outputs(8395) <= not a;
    layer5_outputs(8396) <= 1'b1;
    layer5_outputs(8397) <= a or b;
    layer5_outputs(8398) <= not (a and b);
    layer5_outputs(8399) <= 1'b1;
    layer5_outputs(8400) <= a xor b;
    layer5_outputs(8401) <= a and not b;
    layer5_outputs(8402) <= not a or b;
    layer5_outputs(8403) <= not (a or b);
    layer5_outputs(8404) <= b and not a;
    layer5_outputs(8405) <= not (a or b);
    layer5_outputs(8406) <= a and not b;
    layer5_outputs(8407) <= b;
    layer5_outputs(8408) <= a and not b;
    layer5_outputs(8409) <= not b or a;
    layer5_outputs(8410) <= not a;
    layer5_outputs(8411) <= a;
    layer5_outputs(8412) <= not a;
    layer5_outputs(8413) <= a xor b;
    layer5_outputs(8414) <= not a;
    layer5_outputs(8415) <= a and b;
    layer5_outputs(8416) <= b and not a;
    layer5_outputs(8417) <= not (a and b);
    layer5_outputs(8418) <= not b;
    layer5_outputs(8419) <= a;
    layer5_outputs(8420) <= b and not a;
    layer5_outputs(8421) <= 1'b0;
    layer5_outputs(8422) <= b;
    layer5_outputs(8423) <= not a or b;
    layer5_outputs(8424) <= 1'b0;
    layer5_outputs(8425) <= not a;
    layer5_outputs(8426) <= a and b;
    layer5_outputs(8427) <= not (a and b);
    layer5_outputs(8428) <= not b or a;
    layer5_outputs(8429) <= not b or a;
    layer5_outputs(8430) <= a;
    layer5_outputs(8431) <= not (a xor b);
    layer5_outputs(8432) <= not (a xor b);
    layer5_outputs(8433) <= not a or b;
    layer5_outputs(8434) <= not (a and b);
    layer5_outputs(8435) <= b and not a;
    layer5_outputs(8436) <= not b;
    layer5_outputs(8437) <= not a or b;
    layer5_outputs(8438) <= not b or a;
    layer5_outputs(8439) <= b and not a;
    layer5_outputs(8440) <= not (a and b);
    layer5_outputs(8441) <= a or b;
    layer5_outputs(8442) <= not (a and b);
    layer5_outputs(8443) <= a;
    layer5_outputs(8444) <= not a;
    layer5_outputs(8445) <= a;
    layer5_outputs(8446) <= a and not b;
    layer5_outputs(8447) <= b and not a;
    layer5_outputs(8448) <= 1'b0;
    layer5_outputs(8449) <= b and not a;
    layer5_outputs(8450) <= 1'b1;
    layer5_outputs(8451) <= a and not b;
    layer5_outputs(8452) <= a and b;
    layer5_outputs(8453) <= not a;
    layer5_outputs(8454) <= not (a and b);
    layer5_outputs(8455) <= a or b;
    layer5_outputs(8456) <= not b or a;
    layer5_outputs(8457) <= not (a or b);
    layer5_outputs(8458) <= a;
    layer5_outputs(8459) <= not b or a;
    layer5_outputs(8460) <= a;
    layer5_outputs(8461) <= a;
    layer5_outputs(8462) <= not b;
    layer5_outputs(8463) <= 1'b0;
    layer5_outputs(8464) <= not (a and b);
    layer5_outputs(8465) <= not b or a;
    layer5_outputs(8466) <= a and b;
    layer5_outputs(8467) <= b and not a;
    layer5_outputs(8468) <= a or b;
    layer5_outputs(8469) <= not b or a;
    layer5_outputs(8470) <= not a;
    layer5_outputs(8471) <= a or b;
    layer5_outputs(8472) <= not b;
    layer5_outputs(8473) <= a;
    layer5_outputs(8474) <= not b or a;
    layer5_outputs(8475) <= 1'b0;
    layer5_outputs(8476) <= a and b;
    layer5_outputs(8477) <= a or b;
    layer5_outputs(8478) <= a;
    layer5_outputs(8479) <= not (a and b);
    layer5_outputs(8480) <= not (a or b);
    layer5_outputs(8481) <= b;
    layer5_outputs(8482) <= 1'b1;
    layer5_outputs(8483) <= 1'b0;
    layer5_outputs(8484) <= a or b;
    layer5_outputs(8485) <= not b or a;
    layer5_outputs(8486) <= not (a or b);
    layer5_outputs(8487) <= not (a and b);
    layer5_outputs(8488) <= a or b;
    layer5_outputs(8489) <= a and not b;
    layer5_outputs(8490) <= not b or a;
    layer5_outputs(8491) <= a and b;
    layer5_outputs(8492) <= not (a or b);
    layer5_outputs(8493) <= a;
    layer5_outputs(8494) <= a and not b;
    layer5_outputs(8495) <= not (a and b);
    layer5_outputs(8496) <= a xor b;
    layer5_outputs(8497) <= 1'b0;
    layer5_outputs(8498) <= not (a and b);
    layer5_outputs(8499) <= not a or b;
    layer5_outputs(8500) <= b;
    layer5_outputs(8501) <= 1'b0;
    layer5_outputs(8502) <= not (a or b);
    layer5_outputs(8503) <= not (a and b);
    layer5_outputs(8504) <= not b or a;
    layer5_outputs(8505) <= not (a xor b);
    layer5_outputs(8506) <= not b or a;
    layer5_outputs(8507) <= a xor b;
    layer5_outputs(8508) <= 1'b1;
    layer5_outputs(8509) <= not a or b;
    layer5_outputs(8510) <= a and b;
    layer5_outputs(8511) <= not a or b;
    layer5_outputs(8512) <= not (a or b);
    layer5_outputs(8513) <= b and not a;
    layer5_outputs(8514) <= not b;
    layer5_outputs(8515) <= a;
    layer5_outputs(8516) <= b;
    layer5_outputs(8517) <= not (a and b);
    layer5_outputs(8518) <= a;
    layer5_outputs(8519) <= not (a xor b);
    layer5_outputs(8520) <= a;
    layer5_outputs(8521) <= not b or a;
    layer5_outputs(8522) <= a and b;
    layer5_outputs(8523) <= b;
    layer5_outputs(8524) <= a and not b;
    layer5_outputs(8525) <= not a or b;
    layer5_outputs(8526) <= not (a or b);
    layer5_outputs(8527) <= not a;
    layer5_outputs(8528) <= a xor b;
    layer5_outputs(8529) <= b and not a;
    layer5_outputs(8530) <= not a;
    layer5_outputs(8531) <= a xor b;
    layer5_outputs(8532) <= b;
    layer5_outputs(8533) <= b;
    layer5_outputs(8534) <= a;
    layer5_outputs(8535) <= not b;
    layer5_outputs(8536) <= not (a and b);
    layer5_outputs(8537) <= a and not b;
    layer5_outputs(8538) <= a;
    layer5_outputs(8539) <= not b;
    layer5_outputs(8540) <= a;
    layer5_outputs(8541) <= not a or b;
    layer5_outputs(8542) <= b;
    layer5_outputs(8543) <= a and not b;
    layer5_outputs(8544) <= not b;
    layer5_outputs(8545) <= a;
    layer5_outputs(8546) <= 1'b0;
    layer5_outputs(8547) <= not b or a;
    layer5_outputs(8548) <= not b or a;
    layer5_outputs(8549) <= not a;
    layer5_outputs(8550) <= not (a xor b);
    layer5_outputs(8551) <= a or b;
    layer5_outputs(8552) <= a and not b;
    layer5_outputs(8553) <= 1'b1;
    layer5_outputs(8554) <= b;
    layer5_outputs(8555) <= not a;
    layer5_outputs(8556) <= not (a and b);
    layer5_outputs(8557) <= b and not a;
    layer5_outputs(8558) <= b;
    layer5_outputs(8559) <= not b or a;
    layer5_outputs(8560) <= a;
    layer5_outputs(8561) <= a or b;
    layer5_outputs(8562) <= not (a and b);
    layer5_outputs(8563) <= not b or a;
    layer5_outputs(8564) <= not b or a;
    layer5_outputs(8565) <= not (a and b);
    layer5_outputs(8566) <= not b or a;
    layer5_outputs(8567) <= not b;
    layer5_outputs(8568) <= not a or b;
    layer5_outputs(8569) <= not b or a;
    layer5_outputs(8570) <= a;
    layer5_outputs(8571) <= not b;
    layer5_outputs(8572) <= 1'b1;
    layer5_outputs(8573) <= a;
    layer5_outputs(8574) <= not a;
    layer5_outputs(8575) <= 1'b1;
    layer5_outputs(8576) <= b and not a;
    layer5_outputs(8577) <= 1'b0;
    layer5_outputs(8578) <= not b;
    layer5_outputs(8579) <= not b or a;
    layer5_outputs(8580) <= not a or b;
    layer5_outputs(8581) <= a and not b;
    layer5_outputs(8582) <= a or b;
    layer5_outputs(8583) <= not (a or b);
    layer5_outputs(8584) <= a;
    layer5_outputs(8585) <= a and b;
    layer5_outputs(8586) <= not a;
    layer5_outputs(8587) <= not a;
    layer5_outputs(8588) <= not b;
    layer5_outputs(8589) <= a and b;
    layer5_outputs(8590) <= b and not a;
    layer5_outputs(8591) <= a;
    layer5_outputs(8592) <= b and not a;
    layer5_outputs(8593) <= not a;
    layer5_outputs(8594) <= not (a and b);
    layer5_outputs(8595) <= 1'b1;
    layer5_outputs(8596) <= not b or a;
    layer5_outputs(8597) <= not a;
    layer5_outputs(8598) <= a and not b;
    layer5_outputs(8599) <= b;
    layer5_outputs(8600) <= not (a and b);
    layer5_outputs(8601) <= a and b;
    layer5_outputs(8602) <= not b or a;
    layer5_outputs(8603) <= a and not b;
    layer5_outputs(8604) <= not (a xor b);
    layer5_outputs(8605) <= a and not b;
    layer5_outputs(8606) <= not b;
    layer5_outputs(8607) <= not b;
    layer5_outputs(8608) <= not b;
    layer5_outputs(8609) <= b and not a;
    layer5_outputs(8610) <= a and not b;
    layer5_outputs(8611) <= not a or b;
    layer5_outputs(8612) <= not b or a;
    layer5_outputs(8613) <= a xor b;
    layer5_outputs(8614) <= b;
    layer5_outputs(8615) <= not b or a;
    layer5_outputs(8616) <= not b;
    layer5_outputs(8617) <= a;
    layer5_outputs(8618) <= b and not a;
    layer5_outputs(8619) <= not (a or b);
    layer5_outputs(8620) <= a xor b;
    layer5_outputs(8621) <= a;
    layer5_outputs(8622) <= not b;
    layer5_outputs(8623) <= b;
    layer5_outputs(8624) <= not b or a;
    layer5_outputs(8625) <= not b;
    layer5_outputs(8626) <= 1'b0;
    layer5_outputs(8627) <= not (a or b);
    layer5_outputs(8628) <= b;
    layer5_outputs(8629) <= not a;
    layer5_outputs(8630) <= not b;
    layer5_outputs(8631) <= not b or a;
    layer5_outputs(8632) <= a or b;
    layer5_outputs(8633) <= 1'b0;
    layer5_outputs(8634) <= 1'b0;
    layer5_outputs(8635) <= 1'b1;
    layer5_outputs(8636) <= b and not a;
    layer5_outputs(8637) <= a and not b;
    layer5_outputs(8638) <= not b;
    layer5_outputs(8639) <= not a;
    layer5_outputs(8640) <= not b or a;
    layer5_outputs(8641) <= not b;
    layer5_outputs(8642) <= not b or a;
    layer5_outputs(8643) <= b;
    layer5_outputs(8644) <= not b;
    layer5_outputs(8645) <= not a;
    layer5_outputs(8646) <= not (a or b);
    layer5_outputs(8647) <= b;
    layer5_outputs(8648) <= a;
    layer5_outputs(8649) <= not b;
    layer5_outputs(8650) <= a;
    layer5_outputs(8651) <= b;
    layer5_outputs(8652) <= not (a and b);
    layer5_outputs(8653) <= a;
    layer5_outputs(8654) <= a;
    layer5_outputs(8655) <= b;
    layer5_outputs(8656) <= not a or b;
    layer5_outputs(8657) <= b and not a;
    layer5_outputs(8658) <= a or b;
    layer5_outputs(8659) <= not b;
    layer5_outputs(8660) <= not a or b;
    layer5_outputs(8661) <= a;
    layer5_outputs(8662) <= a or b;
    layer5_outputs(8663) <= not b;
    layer5_outputs(8664) <= not (a xor b);
    layer5_outputs(8665) <= a xor b;
    layer5_outputs(8666) <= not a or b;
    layer5_outputs(8667) <= a and not b;
    layer5_outputs(8668) <= a and b;
    layer5_outputs(8669) <= a;
    layer5_outputs(8670) <= a and b;
    layer5_outputs(8671) <= a or b;
    layer5_outputs(8672) <= not a;
    layer5_outputs(8673) <= b;
    layer5_outputs(8674) <= a;
    layer5_outputs(8675) <= not a;
    layer5_outputs(8676) <= not b;
    layer5_outputs(8677) <= a;
    layer5_outputs(8678) <= not a;
    layer5_outputs(8679) <= 1'b1;
    layer5_outputs(8680) <= not a;
    layer5_outputs(8681) <= not a;
    layer5_outputs(8682) <= 1'b1;
    layer5_outputs(8683) <= not (a and b);
    layer5_outputs(8684) <= 1'b1;
    layer5_outputs(8685) <= a xor b;
    layer5_outputs(8686) <= a or b;
    layer5_outputs(8687) <= a;
    layer5_outputs(8688) <= b;
    layer5_outputs(8689) <= 1'b0;
    layer5_outputs(8690) <= b;
    layer5_outputs(8691) <= not a or b;
    layer5_outputs(8692) <= not b or a;
    layer5_outputs(8693) <= not (a or b);
    layer5_outputs(8694) <= a and not b;
    layer5_outputs(8695) <= 1'b0;
    layer5_outputs(8696) <= not (a or b);
    layer5_outputs(8697) <= not (a xor b);
    layer5_outputs(8698) <= not a or b;
    layer5_outputs(8699) <= 1'b1;
    layer5_outputs(8700) <= not (a or b);
    layer5_outputs(8701) <= b;
    layer5_outputs(8702) <= not a;
    layer5_outputs(8703) <= not b or a;
    layer5_outputs(8704) <= a xor b;
    layer5_outputs(8705) <= 1'b0;
    layer5_outputs(8706) <= 1'b1;
    layer5_outputs(8707) <= a and not b;
    layer5_outputs(8708) <= a and not b;
    layer5_outputs(8709) <= a;
    layer5_outputs(8710) <= not (a and b);
    layer5_outputs(8711) <= not b;
    layer5_outputs(8712) <= a and not b;
    layer5_outputs(8713) <= a;
    layer5_outputs(8714) <= not (a and b);
    layer5_outputs(8715) <= a;
    layer5_outputs(8716) <= a xor b;
    layer5_outputs(8717) <= a xor b;
    layer5_outputs(8718) <= not b or a;
    layer5_outputs(8719) <= not a or b;
    layer5_outputs(8720) <= not b;
    layer5_outputs(8721) <= not b or a;
    layer5_outputs(8722) <= not b or a;
    layer5_outputs(8723) <= b;
    layer5_outputs(8724) <= b;
    layer5_outputs(8725) <= b and not a;
    layer5_outputs(8726) <= b;
    layer5_outputs(8727) <= not b;
    layer5_outputs(8728) <= not (a and b);
    layer5_outputs(8729) <= b and not a;
    layer5_outputs(8730) <= a xor b;
    layer5_outputs(8731) <= a xor b;
    layer5_outputs(8732) <= not (a xor b);
    layer5_outputs(8733) <= b;
    layer5_outputs(8734) <= a or b;
    layer5_outputs(8735) <= not b;
    layer5_outputs(8736) <= not (a or b);
    layer5_outputs(8737) <= a and b;
    layer5_outputs(8738) <= a;
    layer5_outputs(8739) <= not (a and b);
    layer5_outputs(8740) <= a and not b;
    layer5_outputs(8741) <= a and b;
    layer5_outputs(8742) <= not b;
    layer5_outputs(8743) <= a and not b;
    layer5_outputs(8744) <= 1'b0;
    layer5_outputs(8745) <= not b or a;
    layer5_outputs(8746) <= not b or a;
    layer5_outputs(8747) <= b;
    layer5_outputs(8748) <= not (a and b);
    layer5_outputs(8749) <= a and not b;
    layer5_outputs(8750) <= a or b;
    layer5_outputs(8751) <= a or b;
    layer5_outputs(8752) <= not a or b;
    layer5_outputs(8753) <= 1'b0;
    layer5_outputs(8754) <= not a;
    layer5_outputs(8755) <= a xor b;
    layer5_outputs(8756) <= b;
    layer5_outputs(8757) <= 1'b0;
    layer5_outputs(8758) <= a xor b;
    layer5_outputs(8759) <= a;
    layer5_outputs(8760) <= a xor b;
    layer5_outputs(8761) <= 1'b0;
    layer5_outputs(8762) <= b and not a;
    layer5_outputs(8763) <= 1'b1;
    layer5_outputs(8764) <= not b;
    layer5_outputs(8765) <= b;
    layer5_outputs(8766) <= a or b;
    layer5_outputs(8767) <= a and b;
    layer5_outputs(8768) <= not (a xor b);
    layer5_outputs(8769) <= 1'b0;
    layer5_outputs(8770) <= a and not b;
    layer5_outputs(8771) <= not b;
    layer5_outputs(8772) <= a and b;
    layer5_outputs(8773) <= a xor b;
    layer5_outputs(8774) <= b;
    layer5_outputs(8775) <= not (a and b);
    layer5_outputs(8776) <= 1'b1;
    layer5_outputs(8777) <= a;
    layer5_outputs(8778) <= a;
    layer5_outputs(8779) <= b;
    layer5_outputs(8780) <= not b;
    layer5_outputs(8781) <= not a;
    layer5_outputs(8782) <= a and not b;
    layer5_outputs(8783) <= not a;
    layer5_outputs(8784) <= 1'b1;
    layer5_outputs(8785) <= not (a and b);
    layer5_outputs(8786) <= a or b;
    layer5_outputs(8787) <= not b;
    layer5_outputs(8788) <= a;
    layer5_outputs(8789) <= not b or a;
    layer5_outputs(8790) <= 1'b1;
    layer5_outputs(8791) <= not a or b;
    layer5_outputs(8792) <= not a;
    layer5_outputs(8793) <= a;
    layer5_outputs(8794) <= a and not b;
    layer5_outputs(8795) <= not a or b;
    layer5_outputs(8796) <= b and not a;
    layer5_outputs(8797) <= not a;
    layer5_outputs(8798) <= a and b;
    layer5_outputs(8799) <= 1'b0;
    layer5_outputs(8800) <= not b;
    layer5_outputs(8801) <= not (a and b);
    layer5_outputs(8802) <= not b;
    layer5_outputs(8803) <= a and b;
    layer5_outputs(8804) <= not b or a;
    layer5_outputs(8805) <= 1'b1;
    layer5_outputs(8806) <= a and b;
    layer5_outputs(8807) <= a xor b;
    layer5_outputs(8808) <= not a or b;
    layer5_outputs(8809) <= not b;
    layer5_outputs(8810) <= 1'b1;
    layer5_outputs(8811) <= b;
    layer5_outputs(8812) <= b;
    layer5_outputs(8813) <= not (a and b);
    layer5_outputs(8814) <= not (a xor b);
    layer5_outputs(8815) <= b;
    layer5_outputs(8816) <= b;
    layer5_outputs(8817) <= not b or a;
    layer5_outputs(8818) <= b;
    layer5_outputs(8819) <= a;
    layer5_outputs(8820) <= not (a and b);
    layer5_outputs(8821) <= b and not a;
    layer5_outputs(8822) <= b;
    layer5_outputs(8823) <= not (a xor b);
    layer5_outputs(8824) <= not b;
    layer5_outputs(8825) <= b;
    layer5_outputs(8826) <= not b;
    layer5_outputs(8827) <= a;
    layer5_outputs(8828) <= a and not b;
    layer5_outputs(8829) <= a;
    layer5_outputs(8830) <= not (a xor b);
    layer5_outputs(8831) <= not a;
    layer5_outputs(8832) <= not b or a;
    layer5_outputs(8833) <= a xor b;
    layer5_outputs(8834) <= b and not a;
    layer5_outputs(8835) <= not b or a;
    layer5_outputs(8836) <= b and not a;
    layer5_outputs(8837) <= a;
    layer5_outputs(8838) <= b;
    layer5_outputs(8839) <= not (a or b);
    layer5_outputs(8840) <= a and b;
    layer5_outputs(8841) <= 1'b0;
    layer5_outputs(8842) <= a and b;
    layer5_outputs(8843) <= a or b;
    layer5_outputs(8844) <= not b or a;
    layer5_outputs(8845) <= a and not b;
    layer5_outputs(8846) <= a or b;
    layer5_outputs(8847) <= a xor b;
    layer5_outputs(8848) <= not b;
    layer5_outputs(8849) <= not b;
    layer5_outputs(8850) <= a xor b;
    layer5_outputs(8851) <= b;
    layer5_outputs(8852) <= not a;
    layer5_outputs(8853) <= a xor b;
    layer5_outputs(8854) <= not a;
    layer5_outputs(8855) <= not b;
    layer5_outputs(8856) <= not (a and b);
    layer5_outputs(8857) <= not a;
    layer5_outputs(8858) <= not (a or b);
    layer5_outputs(8859) <= a and b;
    layer5_outputs(8860) <= not a or b;
    layer5_outputs(8861) <= b and not a;
    layer5_outputs(8862) <= a and b;
    layer5_outputs(8863) <= not b or a;
    layer5_outputs(8864) <= not a or b;
    layer5_outputs(8865) <= a;
    layer5_outputs(8866) <= a;
    layer5_outputs(8867) <= b and not a;
    layer5_outputs(8868) <= not a or b;
    layer5_outputs(8869) <= a xor b;
    layer5_outputs(8870) <= not b or a;
    layer5_outputs(8871) <= not a;
    layer5_outputs(8872) <= b and not a;
    layer5_outputs(8873) <= not b;
    layer5_outputs(8874) <= not (a or b);
    layer5_outputs(8875) <= b;
    layer5_outputs(8876) <= a;
    layer5_outputs(8877) <= a and not b;
    layer5_outputs(8878) <= not b or a;
    layer5_outputs(8879) <= a or b;
    layer5_outputs(8880) <= a or b;
    layer5_outputs(8881) <= b;
    layer5_outputs(8882) <= 1'b1;
    layer5_outputs(8883) <= a xor b;
    layer5_outputs(8884) <= b;
    layer5_outputs(8885) <= not (a xor b);
    layer5_outputs(8886) <= not a;
    layer5_outputs(8887) <= a and b;
    layer5_outputs(8888) <= b and not a;
    layer5_outputs(8889) <= not (a xor b);
    layer5_outputs(8890) <= b and not a;
    layer5_outputs(8891) <= not a;
    layer5_outputs(8892) <= 1'b1;
    layer5_outputs(8893) <= not b or a;
    layer5_outputs(8894) <= not b or a;
    layer5_outputs(8895) <= 1'b1;
    layer5_outputs(8896) <= not (a xor b);
    layer5_outputs(8897) <= not (a xor b);
    layer5_outputs(8898) <= not b;
    layer5_outputs(8899) <= a xor b;
    layer5_outputs(8900) <= not a or b;
    layer5_outputs(8901) <= a and b;
    layer5_outputs(8902) <= a xor b;
    layer5_outputs(8903) <= not b or a;
    layer5_outputs(8904) <= not (a or b);
    layer5_outputs(8905) <= a and b;
    layer5_outputs(8906) <= not (a xor b);
    layer5_outputs(8907) <= a xor b;
    layer5_outputs(8908) <= a;
    layer5_outputs(8909) <= not b or a;
    layer5_outputs(8910) <= a;
    layer5_outputs(8911) <= not b or a;
    layer5_outputs(8912) <= a or b;
    layer5_outputs(8913) <= not (a xor b);
    layer5_outputs(8914) <= not b;
    layer5_outputs(8915) <= a xor b;
    layer5_outputs(8916) <= not a;
    layer5_outputs(8917) <= not b;
    layer5_outputs(8918) <= a xor b;
    layer5_outputs(8919) <= a or b;
    layer5_outputs(8920) <= a and not b;
    layer5_outputs(8921) <= 1'b1;
    layer5_outputs(8922) <= not a;
    layer5_outputs(8923) <= not b or a;
    layer5_outputs(8924) <= a;
    layer5_outputs(8925) <= not a or b;
    layer5_outputs(8926) <= a and not b;
    layer5_outputs(8927) <= not (a xor b);
    layer5_outputs(8928) <= b;
    layer5_outputs(8929) <= a and b;
    layer5_outputs(8930) <= a;
    layer5_outputs(8931) <= a;
    layer5_outputs(8932) <= not b;
    layer5_outputs(8933) <= a;
    layer5_outputs(8934) <= 1'b1;
    layer5_outputs(8935) <= a and not b;
    layer5_outputs(8936) <= 1'b1;
    layer5_outputs(8937) <= 1'b0;
    layer5_outputs(8938) <= a xor b;
    layer5_outputs(8939) <= b;
    layer5_outputs(8940) <= a and not b;
    layer5_outputs(8941) <= 1'b0;
    layer5_outputs(8942) <= not b;
    layer5_outputs(8943) <= 1'b1;
    layer5_outputs(8944) <= 1'b0;
    layer5_outputs(8945) <= not (a and b);
    layer5_outputs(8946) <= a xor b;
    layer5_outputs(8947) <= not b or a;
    layer5_outputs(8948) <= a;
    layer5_outputs(8949) <= a and not b;
    layer5_outputs(8950) <= not b or a;
    layer5_outputs(8951) <= 1'b0;
    layer5_outputs(8952) <= b and not a;
    layer5_outputs(8953) <= not a or b;
    layer5_outputs(8954) <= not b or a;
    layer5_outputs(8955) <= b;
    layer5_outputs(8956) <= b and not a;
    layer5_outputs(8957) <= not a;
    layer5_outputs(8958) <= not b;
    layer5_outputs(8959) <= a and b;
    layer5_outputs(8960) <= a;
    layer5_outputs(8961) <= not a or b;
    layer5_outputs(8962) <= not a or b;
    layer5_outputs(8963) <= not b or a;
    layer5_outputs(8964) <= b and not a;
    layer5_outputs(8965) <= not a;
    layer5_outputs(8966) <= b and not a;
    layer5_outputs(8967) <= not (a xor b);
    layer5_outputs(8968) <= not b;
    layer5_outputs(8969) <= b and not a;
    layer5_outputs(8970) <= b;
    layer5_outputs(8971) <= not b;
    layer5_outputs(8972) <= a and not b;
    layer5_outputs(8973) <= b and not a;
    layer5_outputs(8974) <= not (a xor b);
    layer5_outputs(8975) <= b;
    layer5_outputs(8976) <= b;
    layer5_outputs(8977) <= not b or a;
    layer5_outputs(8978) <= not b;
    layer5_outputs(8979) <= not b;
    layer5_outputs(8980) <= not a;
    layer5_outputs(8981) <= b;
    layer5_outputs(8982) <= a or b;
    layer5_outputs(8983) <= a;
    layer5_outputs(8984) <= not b or a;
    layer5_outputs(8985) <= b;
    layer5_outputs(8986) <= a xor b;
    layer5_outputs(8987) <= a;
    layer5_outputs(8988) <= b;
    layer5_outputs(8989) <= 1'b1;
    layer5_outputs(8990) <= not a;
    layer5_outputs(8991) <= a or b;
    layer5_outputs(8992) <= 1'b1;
    layer5_outputs(8993) <= not a;
    layer5_outputs(8994) <= not b;
    layer5_outputs(8995) <= 1'b1;
    layer5_outputs(8996) <= a and not b;
    layer5_outputs(8997) <= not b or a;
    layer5_outputs(8998) <= a and b;
    layer5_outputs(8999) <= not a;
    layer5_outputs(9000) <= 1'b0;
    layer5_outputs(9001) <= a or b;
    layer5_outputs(9002) <= a;
    layer5_outputs(9003) <= a and not b;
    layer5_outputs(9004) <= 1'b0;
    layer5_outputs(9005) <= 1'b0;
    layer5_outputs(9006) <= not a;
    layer5_outputs(9007) <= a;
    layer5_outputs(9008) <= b;
    layer5_outputs(9009) <= a or b;
    layer5_outputs(9010) <= not a;
    layer5_outputs(9011) <= a or b;
    layer5_outputs(9012) <= a and b;
    layer5_outputs(9013) <= not (a xor b);
    layer5_outputs(9014) <= not (a or b);
    layer5_outputs(9015) <= not b;
    layer5_outputs(9016) <= not a;
    layer5_outputs(9017) <= a and not b;
    layer5_outputs(9018) <= not b;
    layer5_outputs(9019) <= a or b;
    layer5_outputs(9020) <= not (a xor b);
    layer5_outputs(9021) <= not (a and b);
    layer5_outputs(9022) <= b;
    layer5_outputs(9023) <= not a or b;
    layer5_outputs(9024) <= not a or b;
    layer5_outputs(9025) <= a;
    layer5_outputs(9026) <= not a or b;
    layer5_outputs(9027) <= not (a and b);
    layer5_outputs(9028) <= not (a and b);
    layer5_outputs(9029) <= b;
    layer5_outputs(9030) <= not b or a;
    layer5_outputs(9031) <= not a;
    layer5_outputs(9032) <= a and b;
    layer5_outputs(9033) <= a;
    layer5_outputs(9034) <= a;
    layer5_outputs(9035) <= a and not b;
    layer5_outputs(9036) <= a;
    layer5_outputs(9037) <= a and b;
    layer5_outputs(9038) <= a and b;
    layer5_outputs(9039) <= not a;
    layer5_outputs(9040) <= a;
    layer5_outputs(9041) <= not a;
    layer5_outputs(9042) <= a;
    layer5_outputs(9043) <= a and not b;
    layer5_outputs(9044) <= a;
    layer5_outputs(9045) <= b;
    layer5_outputs(9046) <= a and b;
    layer5_outputs(9047) <= not (a and b);
    layer5_outputs(9048) <= a or b;
    layer5_outputs(9049) <= not b or a;
    layer5_outputs(9050) <= not (a xor b);
    layer5_outputs(9051) <= a;
    layer5_outputs(9052) <= 1'b0;
    layer5_outputs(9053) <= not b;
    layer5_outputs(9054) <= not b or a;
    layer5_outputs(9055) <= 1'b1;
    layer5_outputs(9056) <= 1'b0;
    layer5_outputs(9057) <= not a;
    layer5_outputs(9058) <= not b;
    layer5_outputs(9059) <= a and not b;
    layer5_outputs(9060) <= not a or b;
    layer5_outputs(9061) <= a or b;
    layer5_outputs(9062) <= a or b;
    layer5_outputs(9063) <= not (a or b);
    layer5_outputs(9064) <= a or b;
    layer5_outputs(9065) <= b;
    layer5_outputs(9066) <= b and not a;
    layer5_outputs(9067) <= not b;
    layer5_outputs(9068) <= 1'b1;
    layer5_outputs(9069) <= a and b;
    layer5_outputs(9070) <= not b;
    layer5_outputs(9071) <= not a;
    layer5_outputs(9072) <= not b;
    layer5_outputs(9073) <= not b or a;
    layer5_outputs(9074) <= not a or b;
    layer5_outputs(9075) <= a xor b;
    layer5_outputs(9076) <= a;
    layer5_outputs(9077) <= a and b;
    layer5_outputs(9078) <= not a;
    layer5_outputs(9079) <= 1'b1;
    layer5_outputs(9080) <= 1'b0;
    layer5_outputs(9081) <= not a;
    layer5_outputs(9082) <= b;
    layer5_outputs(9083) <= not b or a;
    layer5_outputs(9084) <= 1'b0;
    layer5_outputs(9085) <= 1'b1;
    layer5_outputs(9086) <= a;
    layer5_outputs(9087) <= not (a or b);
    layer5_outputs(9088) <= not (a or b);
    layer5_outputs(9089) <= not a or b;
    layer5_outputs(9090) <= not a;
    layer5_outputs(9091) <= not (a and b);
    layer5_outputs(9092) <= a xor b;
    layer5_outputs(9093) <= not b;
    layer5_outputs(9094) <= not b;
    layer5_outputs(9095) <= not b;
    layer5_outputs(9096) <= not (a or b);
    layer5_outputs(9097) <= b and not a;
    layer5_outputs(9098) <= not (a or b);
    layer5_outputs(9099) <= b;
    layer5_outputs(9100) <= not (a and b);
    layer5_outputs(9101) <= not b;
    layer5_outputs(9102) <= a and b;
    layer5_outputs(9103) <= not (a or b);
    layer5_outputs(9104) <= not b;
    layer5_outputs(9105) <= a and b;
    layer5_outputs(9106) <= b and not a;
    layer5_outputs(9107) <= a and not b;
    layer5_outputs(9108) <= a and b;
    layer5_outputs(9109) <= b;
    layer5_outputs(9110) <= not b or a;
    layer5_outputs(9111) <= not (a or b);
    layer5_outputs(9112) <= not a or b;
    layer5_outputs(9113) <= not (a xor b);
    layer5_outputs(9114) <= a;
    layer5_outputs(9115) <= not b or a;
    layer5_outputs(9116) <= not (a or b);
    layer5_outputs(9117) <= not a;
    layer5_outputs(9118) <= b;
    layer5_outputs(9119) <= a;
    layer5_outputs(9120) <= not b;
    layer5_outputs(9121) <= a and b;
    layer5_outputs(9122) <= not b or a;
    layer5_outputs(9123) <= 1'b0;
    layer5_outputs(9124) <= not (a and b);
    layer5_outputs(9125) <= a;
    layer5_outputs(9126) <= 1'b1;
    layer5_outputs(9127) <= a;
    layer5_outputs(9128) <= not a;
    layer5_outputs(9129) <= a xor b;
    layer5_outputs(9130) <= not a;
    layer5_outputs(9131) <= not (a xor b);
    layer5_outputs(9132) <= not b or a;
    layer5_outputs(9133) <= a;
    layer5_outputs(9134) <= a and b;
    layer5_outputs(9135) <= b;
    layer5_outputs(9136) <= not (a or b);
    layer5_outputs(9137) <= not (a xor b);
    layer5_outputs(9138) <= a xor b;
    layer5_outputs(9139) <= b;
    layer5_outputs(9140) <= not (a and b);
    layer5_outputs(9141) <= b and not a;
    layer5_outputs(9142) <= a;
    layer5_outputs(9143) <= a and not b;
    layer5_outputs(9144) <= not a or b;
    layer5_outputs(9145) <= a;
    layer5_outputs(9146) <= a and not b;
    layer5_outputs(9147) <= not (a xor b);
    layer5_outputs(9148) <= b and not a;
    layer5_outputs(9149) <= b;
    layer5_outputs(9150) <= a;
    layer5_outputs(9151) <= a;
    layer5_outputs(9152) <= a or b;
    layer5_outputs(9153) <= not a;
    layer5_outputs(9154) <= b;
    layer5_outputs(9155) <= b and not a;
    layer5_outputs(9156) <= not a or b;
    layer5_outputs(9157) <= not a;
    layer5_outputs(9158) <= not a;
    layer5_outputs(9159) <= a or b;
    layer5_outputs(9160) <= b and not a;
    layer5_outputs(9161) <= a and b;
    layer5_outputs(9162) <= not (a and b);
    layer5_outputs(9163) <= b;
    layer5_outputs(9164) <= not b or a;
    layer5_outputs(9165) <= 1'b0;
    layer5_outputs(9166) <= not a;
    layer5_outputs(9167) <= not a;
    layer5_outputs(9168) <= not b;
    layer5_outputs(9169) <= not (a xor b);
    layer5_outputs(9170) <= a xor b;
    layer5_outputs(9171) <= a;
    layer5_outputs(9172) <= not a;
    layer5_outputs(9173) <= a;
    layer5_outputs(9174) <= a xor b;
    layer5_outputs(9175) <= 1'b0;
    layer5_outputs(9176) <= 1'b1;
    layer5_outputs(9177) <= a and not b;
    layer5_outputs(9178) <= a;
    layer5_outputs(9179) <= a or b;
    layer5_outputs(9180) <= not (a xor b);
    layer5_outputs(9181) <= not b;
    layer5_outputs(9182) <= 1'b0;
    layer5_outputs(9183) <= not b;
    layer5_outputs(9184) <= b;
    layer5_outputs(9185) <= not a;
    layer5_outputs(9186) <= not (a or b);
    layer5_outputs(9187) <= b and not a;
    layer5_outputs(9188) <= not b;
    layer5_outputs(9189) <= a xor b;
    layer5_outputs(9190) <= not b;
    layer5_outputs(9191) <= b and not a;
    layer5_outputs(9192) <= not a or b;
    layer5_outputs(9193) <= 1'b1;
    layer5_outputs(9194) <= not (a or b);
    layer5_outputs(9195) <= b;
    layer5_outputs(9196) <= not b or a;
    layer5_outputs(9197) <= a and b;
    layer5_outputs(9198) <= not (a xor b);
    layer5_outputs(9199) <= b;
    layer5_outputs(9200) <= 1'b1;
    layer5_outputs(9201) <= b and not a;
    layer5_outputs(9202) <= 1'b1;
    layer5_outputs(9203) <= not (a and b);
    layer5_outputs(9204) <= not a or b;
    layer5_outputs(9205) <= 1'b1;
    layer5_outputs(9206) <= b;
    layer5_outputs(9207) <= not b;
    layer5_outputs(9208) <= a and not b;
    layer5_outputs(9209) <= a or b;
    layer5_outputs(9210) <= not (a xor b);
    layer5_outputs(9211) <= not b or a;
    layer5_outputs(9212) <= a and b;
    layer5_outputs(9213) <= not a or b;
    layer5_outputs(9214) <= not b;
    layer5_outputs(9215) <= not a;
    layer5_outputs(9216) <= a;
    layer5_outputs(9217) <= a and not b;
    layer5_outputs(9218) <= not a;
    layer5_outputs(9219) <= a;
    layer5_outputs(9220) <= not b;
    layer5_outputs(9221) <= not b or a;
    layer5_outputs(9222) <= not b;
    layer5_outputs(9223) <= not (a and b);
    layer5_outputs(9224) <= not a;
    layer5_outputs(9225) <= not b or a;
    layer5_outputs(9226) <= a;
    layer5_outputs(9227) <= not (a xor b);
    layer5_outputs(9228) <= not b;
    layer5_outputs(9229) <= a or b;
    layer5_outputs(9230) <= b and not a;
    layer5_outputs(9231) <= not a or b;
    layer5_outputs(9232) <= not b;
    layer5_outputs(9233) <= not (a xor b);
    layer5_outputs(9234) <= not (a and b);
    layer5_outputs(9235) <= 1'b1;
    layer5_outputs(9236) <= not a;
    layer5_outputs(9237) <= b;
    layer5_outputs(9238) <= not a;
    layer5_outputs(9239) <= b;
    layer5_outputs(9240) <= not a or b;
    layer5_outputs(9241) <= 1'b1;
    layer5_outputs(9242) <= a and b;
    layer5_outputs(9243) <= not (a xor b);
    layer5_outputs(9244) <= not a;
    layer5_outputs(9245) <= b;
    layer5_outputs(9246) <= a xor b;
    layer5_outputs(9247) <= a and not b;
    layer5_outputs(9248) <= not b;
    layer5_outputs(9249) <= not a or b;
    layer5_outputs(9250) <= not a;
    layer5_outputs(9251) <= not a or b;
    layer5_outputs(9252) <= a xor b;
    layer5_outputs(9253) <= not (a xor b);
    layer5_outputs(9254) <= not b or a;
    layer5_outputs(9255) <= b;
    layer5_outputs(9256) <= not a;
    layer5_outputs(9257) <= not (a and b);
    layer5_outputs(9258) <= a and not b;
    layer5_outputs(9259) <= not (a and b);
    layer5_outputs(9260) <= a xor b;
    layer5_outputs(9261) <= a and b;
    layer5_outputs(9262) <= a and not b;
    layer5_outputs(9263) <= a xor b;
    layer5_outputs(9264) <= b;
    layer5_outputs(9265) <= a;
    layer5_outputs(9266) <= a;
    layer5_outputs(9267) <= a;
    layer5_outputs(9268) <= not (a and b);
    layer5_outputs(9269) <= not (a and b);
    layer5_outputs(9270) <= not (a or b);
    layer5_outputs(9271) <= a and not b;
    layer5_outputs(9272) <= a;
    layer5_outputs(9273) <= not a;
    layer5_outputs(9274) <= not (a xor b);
    layer5_outputs(9275) <= 1'b0;
    layer5_outputs(9276) <= not a or b;
    layer5_outputs(9277) <= not a;
    layer5_outputs(9278) <= a xor b;
    layer5_outputs(9279) <= not (a xor b);
    layer5_outputs(9280) <= 1'b0;
    layer5_outputs(9281) <= a or b;
    layer5_outputs(9282) <= 1'b1;
    layer5_outputs(9283) <= a and not b;
    layer5_outputs(9284) <= 1'b0;
    layer5_outputs(9285) <= not (a xor b);
    layer5_outputs(9286) <= a and not b;
    layer5_outputs(9287) <= b;
    layer5_outputs(9288) <= not (a or b);
    layer5_outputs(9289) <= 1'b0;
    layer5_outputs(9290) <= a and b;
    layer5_outputs(9291) <= not a;
    layer5_outputs(9292) <= not a;
    layer5_outputs(9293) <= not (a and b);
    layer5_outputs(9294) <= not a;
    layer5_outputs(9295) <= not b or a;
    layer5_outputs(9296) <= b;
    layer5_outputs(9297) <= a and b;
    layer5_outputs(9298) <= a and not b;
    layer5_outputs(9299) <= a xor b;
    layer5_outputs(9300) <= a;
    layer5_outputs(9301) <= 1'b0;
    layer5_outputs(9302) <= not (a and b);
    layer5_outputs(9303) <= not a or b;
    layer5_outputs(9304) <= not (a xor b);
    layer5_outputs(9305) <= a;
    layer5_outputs(9306) <= 1'b0;
    layer5_outputs(9307) <= b;
    layer5_outputs(9308) <= b;
    layer5_outputs(9309) <= not b;
    layer5_outputs(9310) <= not a or b;
    layer5_outputs(9311) <= b;
    layer5_outputs(9312) <= b and not a;
    layer5_outputs(9313) <= b;
    layer5_outputs(9314) <= not b;
    layer5_outputs(9315) <= a and not b;
    layer5_outputs(9316) <= a and b;
    layer5_outputs(9317) <= a xor b;
    layer5_outputs(9318) <= a or b;
    layer5_outputs(9319) <= not b or a;
    layer5_outputs(9320) <= b and not a;
    layer5_outputs(9321) <= b and not a;
    layer5_outputs(9322) <= not (a xor b);
    layer5_outputs(9323) <= not a;
    layer5_outputs(9324) <= not (a and b);
    layer5_outputs(9325) <= a or b;
    layer5_outputs(9326) <= not (a xor b);
    layer5_outputs(9327) <= a;
    layer5_outputs(9328) <= b and not a;
    layer5_outputs(9329) <= a;
    layer5_outputs(9330) <= b;
    layer5_outputs(9331) <= a and b;
    layer5_outputs(9332) <= not (a and b);
    layer5_outputs(9333) <= not b;
    layer5_outputs(9334) <= b and not a;
    layer5_outputs(9335) <= a;
    layer5_outputs(9336) <= a or b;
    layer5_outputs(9337) <= not b or a;
    layer5_outputs(9338) <= not (a and b);
    layer5_outputs(9339) <= not (a or b);
    layer5_outputs(9340) <= not a or b;
    layer5_outputs(9341) <= not (a and b);
    layer5_outputs(9342) <= not b or a;
    layer5_outputs(9343) <= a and not b;
    layer5_outputs(9344) <= not b or a;
    layer5_outputs(9345) <= b;
    layer5_outputs(9346) <= not a;
    layer5_outputs(9347) <= not a or b;
    layer5_outputs(9348) <= not (a and b);
    layer5_outputs(9349) <= not (a and b);
    layer5_outputs(9350) <= not a;
    layer5_outputs(9351) <= not b;
    layer5_outputs(9352) <= not a;
    layer5_outputs(9353) <= a xor b;
    layer5_outputs(9354) <= a and b;
    layer5_outputs(9355) <= not (a xor b);
    layer5_outputs(9356) <= a or b;
    layer5_outputs(9357) <= a;
    layer5_outputs(9358) <= a or b;
    layer5_outputs(9359) <= not a or b;
    layer5_outputs(9360) <= not a;
    layer5_outputs(9361) <= not a;
    layer5_outputs(9362) <= not a or b;
    layer5_outputs(9363) <= not (a and b);
    layer5_outputs(9364) <= not (a and b);
    layer5_outputs(9365) <= not b or a;
    layer5_outputs(9366) <= b;
    layer5_outputs(9367) <= not a;
    layer5_outputs(9368) <= a or b;
    layer5_outputs(9369) <= not (a or b);
    layer5_outputs(9370) <= 1'b0;
    layer5_outputs(9371) <= a;
    layer5_outputs(9372) <= b and not a;
    layer5_outputs(9373) <= a;
    layer5_outputs(9374) <= not a;
    layer5_outputs(9375) <= not (a and b);
    layer5_outputs(9376) <= a xor b;
    layer5_outputs(9377) <= not (a xor b);
    layer5_outputs(9378) <= a or b;
    layer5_outputs(9379) <= a;
    layer5_outputs(9380) <= not b or a;
    layer5_outputs(9381) <= a;
    layer5_outputs(9382) <= a;
    layer5_outputs(9383) <= b;
    layer5_outputs(9384) <= not a;
    layer5_outputs(9385) <= not a or b;
    layer5_outputs(9386) <= not (a xor b);
    layer5_outputs(9387) <= not b or a;
    layer5_outputs(9388) <= a or b;
    layer5_outputs(9389) <= a;
    layer5_outputs(9390) <= a and not b;
    layer5_outputs(9391) <= a and not b;
    layer5_outputs(9392) <= 1'b0;
    layer5_outputs(9393) <= b and not a;
    layer5_outputs(9394) <= 1'b0;
    layer5_outputs(9395) <= a;
    layer5_outputs(9396) <= a and b;
    layer5_outputs(9397) <= a xor b;
    layer5_outputs(9398) <= not a;
    layer5_outputs(9399) <= b and not a;
    layer5_outputs(9400) <= not b;
    layer5_outputs(9401) <= not b;
    layer5_outputs(9402) <= not a;
    layer5_outputs(9403) <= a;
    layer5_outputs(9404) <= a and not b;
    layer5_outputs(9405) <= 1'b0;
    layer5_outputs(9406) <= not a;
    layer5_outputs(9407) <= not (a and b);
    layer5_outputs(9408) <= not b;
    layer5_outputs(9409) <= not (a or b);
    layer5_outputs(9410) <= not b;
    layer5_outputs(9411) <= a or b;
    layer5_outputs(9412) <= a and not b;
    layer5_outputs(9413) <= a and not b;
    layer5_outputs(9414) <= not a;
    layer5_outputs(9415) <= a;
    layer5_outputs(9416) <= not a;
    layer5_outputs(9417) <= a;
    layer5_outputs(9418) <= b and not a;
    layer5_outputs(9419) <= a and not b;
    layer5_outputs(9420) <= a xor b;
    layer5_outputs(9421) <= a and b;
    layer5_outputs(9422) <= a xor b;
    layer5_outputs(9423) <= b;
    layer5_outputs(9424) <= not a;
    layer5_outputs(9425) <= not b;
    layer5_outputs(9426) <= 1'b0;
    layer5_outputs(9427) <= not b;
    layer5_outputs(9428) <= b;
    layer5_outputs(9429) <= not a or b;
    layer5_outputs(9430) <= not b;
    layer5_outputs(9431) <= a;
    layer5_outputs(9432) <= not b;
    layer5_outputs(9433) <= 1'b0;
    layer5_outputs(9434) <= b;
    layer5_outputs(9435) <= a xor b;
    layer5_outputs(9436) <= a;
    layer5_outputs(9437) <= b;
    layer5_outputs(9438) <= b and not a;
    layer5_outputs(9439) <= a;
    layer5_outputs(9440) <= a and b;
    layer5_outputs(9441) <= a;
    layer5_outputs(9442) <= a;
    layer5_outputs(9443) <= not a or b;
    layer5_outputs(9444) <= a;
    layer5_outputs(9445) <= not b or a;
    layer5_outputs(9446) <= a;
    layer5_outputs(9447) <= 1'b1;
    layer5_outputs(9448) <= not (a or b);
    layer5_outputs(9449) <= not a;
    layer5_outputs(9450) <= a and b;
    layer5_outputs(9451) <= a or b;
    layer5_outputs(9452) <= not b;
    layer5_outputs(9453) <= not a or b;
    layer5_outputs(9454) <= a xor b;
    layer5_outputs(9455) <= not b;
    layer5_outputs(9456) <= a;
    layer5_outputs(9457) <= 1'b1;
    layer5_outputs(9458) <= not a;
    layer5_outputs(9459) <= not b;
    layer5_outputs(9460) <= not b;
    layer5_outputs(9461) <= b;
    layer5_outputs(9462) <= b;
    layer5_outputs(9463) <= not (a and b);
    layer5_outputs(9464) <= a and b;
    layer5_outputs(9465) <= not a or b;
    layer5_outputs(9466) <= b;
    layer5_outputs(9467) <= a or b;
    layer5_outputs(9468) <= not a or b;
    layer5_outputs(9469) <= b;
    layer5_outputs(9470) <= a and b;
    layer5_outputs(9471) <= not a or b;
    layer5_outputs(9472) <= a xor b;
    layer5_outputs(9473) <= not (a or b);
    layer5_outputs(9474) <= a and not b;
    layer5_outputs(9475) <= a and not b;
    layer5_outputs(9476) <= not a or b;
    layer5_outputs(9477) <= not b;
    layer5_outputs(9478) <= 1'b0;
    layer5_outputs(9479) <= a;
    layer5_outputs(9480) <= b;
    layer5_outputs(9481) <= not b;
    layer5_outputs(9482) <= a and not b;
    layer5_outputs(9483) <= a;
    layer5_outputs(9484) <= not b;
    layer5_outputs(9485) <= not b;
    layer5_outputs(9486) <= a;
    layer5_outputs(9487) <= a;
    layer5_outputs(9488) <= not b or a;
    layer5_outputs(9489) <= a and b;
    layer5_outputs(9490) <= b and not a;
    layer5_outputs(9491) <= b;
    layer5_outputs(9492) <= not a;
    layer5_outputs(9493) <= a or b;
    layer5_outputs(9494) <= a or b;
    layer5_outputs(9495) <= not a;
    layer5_outputs(9496) <= not (a and b);
    layer5_outputs(9497) <= b;
    layer5_outputs(9498) <= b and not a;
    layer5_outputs(9499) <= b;
    layer5_outputs(9500) <= 1'b0;
    layer5_outputs(9501) <= not (a and b);
    layer5_outputs(9502) <= not (a or b);
    layer5_outputs(9503) <= b;
    layer5_outputs(9504) <= not a;
    layer5_outputs(9505) <= not a;
    layer5_outputs(9506) <= b;
    layer5_outputs(9507) <= 1'b0;
    layer5_outputs(9508) <= not b;
    layer5_outputs(9509) <= not (a and b);
    layer5_outputs(9510) <= not a or b;
    layer5_outputs(9511) <= not (a or b);
    layer5_outputs(9512) <= b and not a;
    layer5_outputs(9513) <= not b;
    layer5_outputs(9514) <= not a;
    layer5_outputs(9515) <= not b;
    layer5_outputs(9516) <= not b or a;
    layer5_outputs(9517) <= not b;
    layer5_outputs(9518) <= not b or a;
    layer5_outputs(9519) <= a xor b;
    layer5_outputs(9520) <= a and not b;
    layer5_outputs(9521) <= not (a or b);
    layer5_outputs(9522) <= b;
    layer5_outputs(9523) <= 1'b0;
    layer5_outputs(9524) <= not (a xor b);
    layer5_outputs(9525) <= 1'b0;
    layer5_outputs(9526) <= not a or b;
    layer5_outputs(9527) <= not a;
    layer5_outputs(9528) <= not b or a;
    layer5_outputs(9529) <= 1'b1;
    layer5_outputs(9530) <= a;
    layer5_outputs(9531) <= not (a and b);
    layer5_outputs(9532) <= not b;
    layer5_outputs(9533) <= b;
    layer5_outputs(9534) <= a;
    layer5_outputs(9535) <= not (a xor b);
    layer5_outputs(9536) <= a;
    layer5_outputs(9537) <= a or b;
    layer5_outputs(9538) <= not (a xor b);
    layer5_outputs(9539) <= a or b;
    layer5_outputs(9540) <= a;
    layer5_outputs(9541) <= not a;
    layer5_outputs(9542) <= a;
    layer5_outputs(9543) <= b and not a;
    layer5_outputs(9544) <= 1'b0;
    layer5_outputs(9545) <= not b or a;
    layer5_outputs(9546) <= not a or b;
    layer5_outputs(9547) <= a and not b;
    layer5_outputs(9548) <= a;
    layer5_outputs(9549) <= not (a and b);
    layer5_outputs(9550) <= not (a xor b);
    layer5_outputs(9551) <= not b;
    layer5_outputs(9552) <= not a or b;
    layer5_outputs(9553) <= not (a and b);
    layer5_outputs(9554) <= not a;
    layer5_outputs(9555) <= not a;
    layer5_outputs(9556) <= not b;
    layer5_outputs(9557) <= 1'b0;
    layer5_outputs(9558) <= a and b;
    layer5_outputs(9559) <= 1'b1;
    layer5_outputs(9560) <= not (a and b);
    layer5_outputs(9561) <= a and not b;
    layer5_outputs(9562) <= not a;
    layer5_outputs(9563) <= a;
    layer5_outputs(9564) <= 1'b1;
    layer5_outputs(9565) <= not (a xor b);
    layer5_outputs(9566) <= 1'b1;
    layer5_outputs(9567) <= not a;
    layer5_outputs(9568) <= not a or b;
    layer5_outputs(9569) <= not a or b;
    layer5_outputs(9570) <= not b;
    layer5_outputs(9571) <= not a;
    layer5_outputs(9572) <= a and b;
    layer5_outputs(9573) <= not a or b;
    layer5_outputs(9574) <= not a or b;
    layer5_outputs(9575) <= not b;
    layer5_outputs(9576) <= not (a xor b);
    layer5_outputs(9577) <= not a;
    layer5_outputs(9578) <= a xor b;
    layer5_outputs(9579) <= a and b;
    layer5_outputs(9580) <= b;
    layer5_outputs(9581) <= not a;
    layer5_outputs(9582) <= not b or a;
    layer5_outputs(9583) <= not (a or b);
    layer5_outputs(9584) <= not b;
    layer5_outputs(9585) <= a;
    layer5_outputs(9586) <= not a or b;
    layer5_outputs(9587) <= not b or a;
    layer5_outputs(9588) <= a or b;
    layer5_outputs(9589) <= not a;
    layer5_outputs(9590) <= a;
    layer5_outputs(9591) <= a and b;
    layer5_outputs(9592) <= a;
    layer5_outputs(9593) <= not (a and b);
    layer5_outputs(9594) <= a or b;
    layer5_outputs(9595) <= a xor b;
    layer5_outputs(9596) <= a or b;
    layer5_outputs(9597) <= b;
    layer5_outputs(9598) <= not (a xor b);
    layer5_outputs(9599) <= not a;
    layer5_outputs(9600) <= not (a and b);
    layer5_outputs(9601) <= not a;
    layer5_outputs(9602) <= a or b;
    layer5_outputs(9603) <= not b;
    layer5_outputs(9604) <= b;
    layer5_outputs(9605) <= not (a and b);
    layer5_outputs(9606) <= a or b;
    layer5_outputs(9607) <= not b or a;
    layer5_outputs(9608) <= a and not b;
    layer5_outputs(9609) <= not a;
    layer5_outputs(9610) <= not b;
    layer5_outputs(9611) <= not a or b;
    layer5_outputs(9612) <= a and not b;
    layer5_outputs(9613) <= not (a or b);
    layer5_outputs(9614) <= b;
    layer5_outputs(9615) <= a and b;
    layer5_outputs(9616) <= not (a or b);
    layer5_outputs(9617) <= a and b;
    layer5_outputs(9618) <= b;
    layer5_outputs(9619) <= b and not a;
    layer5_outputs(9620) <= a;
    layer5_outputs(9621) <= not a;
    layer5_outputs(9622) <= a xor b;
    layer5_outputs(9623) <= not b;
    layer5_outputs(9624) <= b;
    layer5_outputs(9625) <= not b or a;
    layer5_outputs(9626) <= not a or b;
    layer5_outputs(9627) <= a;
    layer5_outputs(9628) <= not b or a;
    layer5_outputs(9629) <= not a or b;
    layer5_outputs(9630) <= a xor b;
    layer5_outputs(9631) <= not a or b;
    layer5_outputs(9632) <= not a;
    layer5_outputs(9633) <= 1'b0;
    layer5_outputs(9634) <= not a;
    layer5_outputs(9635) <= a or b;
    layer5_outputs(9636) <= b;
    layer5_outputs(9637) <= not a or b;
    layer5_outputs(9638) <= not b or a;
    layer5_outputs(9639) <= not b;
    layer5_outputs(9640) <= b and not a;
    layer5_outputs(9641) <= not (a or b);
    layer5_outputs(9642) <= not b;
    layer5_outputs(9643) <= 1'b1;
    layer5_outputs(9644) <= not (a and b);
    layer5_outputs(9645) <= a and not b;
    layer5_outputs(9646) <= a;
    layer5_outputs(9647) <= not a;
    layer5_outputs(9648) <= a and b;
    layer5_outputs(9649) <= not (a xor b);
    layer5_outputs(9650) <= not a;
    layer5_outputs(9651) <= not (a or b);
    layer5_outputs(9652) <= not a;
    layer5_outputs(9653) <= a and b;
    layer5_outputs(9654) <= a;
    layer5_outputs(9655) <= not a;
    layer5_outputs(9656) <= a and not b;
    layer5_outputs(9657) <= not b;
    layer5_outputs(9658) <= not b;
    layer5_outputs(9659) <= not a;
    layer5_outputs(9660) <= not a or b;
    layer5_outputs(9661) <= b and not a;
    layer5_outputs(9662) <= 1'b0;
    layer5_outputs(9663) <= b and not a;
    layer5_outputs(9664) <= b;
    layer5_outputs(9665) <= not b;
    layer5_outputs(9666) <= a and not b;
    layer5_outputs(9667) <= not b or a;
    layer5_outputs(9668) <= a and b;
    layer5_outputs(9669) <= a;
    layer5_outputs(9670) <= a xor b;
    layer5_outputs(9671) <= b and not a;
    layer5_outputs(9672) <= a and b;
    layer5_outputs(9673) <= a and b;
    layer5_outputs(9674) <= a;
    layer5_outputs(9675) <= not b;
    layer5_outputs(9676) <= not (a or b);
    layer5_outputs(9677) <= a and not b;
    layer5_outputs(9678) <= not (a and b);
    layer5_outputs(9679) <= not b;
    layer5_outputs(9680) <= a and not b;
    layer5_outputs(9681) <= a or b;
    layer5_outputs(9682) <= a and not b;
    layer5_outputs(9683) <= 1'b1;
    layer5_outputs(9684) <= a and b;
    layer5_outputs(9685) <= not b;
    layer5_outputs(9686) <= b;
    layer5_outputs(9687) <= not a or b;
    layer5_outputs(9688) <= a;
    layer5_outputs(9689) <= 1'b1;
    layer5_outputs(9690) <= a or b;
    layer5_outputs(9691) <= not a or b;
    layer5_outputs(9692) <= not (a or b);
    layer5_outputs(9693) <= not (a or b);
    layer5_outputs(9694) <= a;
    layer5_outputs(9695) <= a and not b;
    layer5_outputs(9696) <= a;
    layer5_outputs(9697) <= a or b;
    layer5_outputs(9698) <= not a;
    layer5_outputs(9699) <= not b;
    layer5_outputs(9700) <= a;
    layer5_outputs(9701) <= a and b;
    layer5_outputs(9702) <= not (a xor b);
    layer5_outputs(9703) <= not a;
    layer5_outputs(9704) <= 1'b0;
    layer5_outputs(9705) <= a and b;
    layer5_outputs(9706) <= b;
    layer5_outputs(9707) <= not (a or b);
    layer5_outputs(9708) <= 1'b0;
    layer5_outputs(9709) <= not a or b;
    layer5_outputs(9710) <= a and not b;
    layer5_outputs(9711) <= a and b;
    layer5_outputs(9712) <= not b;
    layer5_outputs(9713) <= 1'b0;
    layer5_outputs(9714) <= not (a and b);
    layer5_outputs(9715) <= b and not a;
    layer5_outputs(9716) <= a;
    layer5_outputs(9717) <= a;
    layer5_outputs(9718) <= not b or a;
    layer5_outputs(9719) <= not b;
    layer5_outputs(9720) <= a and b;
    layer5_outputs(9721) <= a and b;
    layer5_outputs(9722) <= not (a and b);
    layer5_outputs(9723) <= not a;
    layer5_outputs(9724) <= not b;
    layer5_outputs(9725) <= not (a or b);
    layer5_outputs(9726) <= 1'b1;
    layer5_outputs(9727) <= b;
    layer5_outputs(9728) <= a;
    layer5_outputs(9729) <= a and b;
    layer5_outputs(9730) <= b;
    layer5_outputs(9731) <= not b or a;
    layer5_outputs(9732) <= not a;
    layer5_outputs(9733) <= not b;
    layer5_outputs(9734) <= not (a and b);
    layer5_outputs(9735) <= not a;
    layer5_outputs(9736) <= a or b;
    layer5_outputs(9737) <= a;
    layer5_outputs(9738) <= not b;
    layer5_outputs(9739) <= a xor b;
    layer5_outputs(9740) <= 1'b1;
    layer5_outputs(9741) <= a and not b;
    layer5_outputs(9742) <= a;
    layer5_outputs(9743) <= not b;
    layer5_outputs(9744) <= b;
    layer5_outputs(9745) <= a and not b;
    layer5_outputs(9746) <= not b;
    layer5_outputs(9747) <= a;
    layer5_outputs(9748) <= b;
    layer5_outputs(9749) <= not (a or b);
    layer5_outputs(9750) <= a and b;
    layer5_outputs(9751) <= not a or b;
    layer5_outputs(9752) <= not a;
    layer5_outputs(9753) <= 1'b1;
    layer5_outputs(9754) <= not b;
    layer5_outputs(9755) <= b and not a;
    layer5_outputs(9756) <= not b or a;
    layer5_outputs(9757) <= not b;
    layer5_outputs(9758) <= b;
    layer5_outputs(9759) <= not a;
    layer5_outputs(9760) <= a xor b;
    layer5_outputs(9761) <= not b;
    layer5_outputs(9762) <= a;
    layer5_outputs(9763) <= a and not b;
    layer5_outputs(9764) <= a xor b;
    layer5_outputs(9765) <= a;
    layer5_outputs(9766) <= not b or a;
    layer5_outputs(9767) <= a and b;
    layer5_outputs(9768) <= b;
    layer5_outputs(9769) <= a;
    layer5_outputs(9770) <= b;
    layer5_outputs(9771) <= a xor b;
    layer5_outputs(9772) <= not b;
    layer5_outputs(9773) <= not (a and b);
    layer5_outputs(9774) <= not b;
    layer5_outputs(9775) <= b and not a;
    layer5_outputs(9776) <= not b;
    layer5_outputs(9777) <= b;
    layer5_outputs(9778) <= not b;
    layer5_outputs(9779) <= not b;
    layer5_outputs(9780) <= not a;
    layer5_outputs(9781) <= 1'b0;
    layer5_outputs(9782) <= a and not b;
    layer5_outputs(9783) <= 1'b1;
    layer5_outputs(9784) <= not b;
    layer5_outputs(9785) <= not a;
    layer5_outputs(9786) <= a and b;
    layer5_outputs(9787) <= not a;
    layer5_outputs(9788) <= not b or a;
    layer5_outputs(9789) <= not a;
    layer5_outputs(9790) <= b;
    layer5_outputs(9791) <= a and b;
    layer5_outputs(9792) <= a;
    layer5_outputs(9793) <= not b;
    layer5_outputs(9794) <= 1'b0;
    layer5_outputs(9795) <= not b;
    layer5_outputs(9796) <= 1'b0;
    layer5_outputs(9797) <= not a;
    layer5_outputs(9798) <= not a;
    layer5_outputs(9799) <= 1'b1;
    layer5_outputs(9800) <= not a or b;
    layer5_outputs(9801) <= a;
    layer5_outputs(9802) <= 1'b0;
    layer5_outputs(9803) <= a and not b;
    layer5_outputs(9804) <= a and not b;
    layer5_outputs(9805) <= b;
    layer5_outputs(9806) <= not (a or b);
    layer5_outputs(9807) <= b;
    layer5_outputs(9808) <= not (a or b);
    layer5_outputs(9809) <= not (a xor b);
    layer5_outputs(9810) <= not (a or b);
    layer5_outputs(9811) <= b and not a;
    layer5_outputs(9812) <= not b;
    layer5_outputs(9813) <= b and not a;
    layer5_outputs(9814) <= 1'b0;
    layer5_outputs(9815) <= a;
    layer5_outputs(9816) <= a and not b;
    layer5_outputs(9817) <= b and not a;
    layer5_outputs(9818) <= not (a or b);
    layer5_outputs(9819) <= b;
    layer5_outputs(9820) <= not (a xor b);
    layer5_outputs(9821) <= b;
    layer5_outputs(9822) <= b and not a;
    layer5_outputs(9823) <= a or b;
    layer5_outputs(9824) <= a;
    layer5_outputs(9825) <= a and b;
    layer5_outputs(9826) <= a;
    layer5_outputs(9827) <= not a;
    layer5_outputs(9828) <= not a;
    layer5_outputs(9829) <= a and b;
    layer5_outputs(9830) <= not a or b;
    layer5_outputs(9831) <= not b;
    layer5_outputs(9832) <= b and not a;
    layer5_outputs(9833) <= not b or a;
    layer5_outputs(9834) <= 1'b1;
    layer5_outputs(9835) <= a or b;
    layer5_outputs(9836) <= not a;
    layer5_outputs(9837) <= b and not a;
    layer5_outputs(9838) <= a and not b;
    layer5_outputs(9839) <= b;
    layer5_outputs(9840) <= not b;
    layer5_outputs(9841) <= a or b;
    layer5_outputs(9842) <= a;
    layer5_outputs(9843) <= not a or b;
    layer5_outputs(9844) <= 1'b0;
    layer5_outputs(9845) <= b;
    layer5_outputs(9846) <= not b or a;
    layer5_outputs(9847) <= a or b;
    layer5_outputs(9848) <= 1'b0;
    layer5_outputs(9849) <= a;
    layer5_outputs(9850) <= b;
    layer5_outputs(9851) <= not b or a;
    layer5_outputs(9852) <= 1'b1;
    layer5_outputs(9853) <= b and not a;
    layer5_outputs(9854) <= a;
    layer5_outputs(9855) <= not a;
    layer5_outputs(9856) <= not (a or b);
    layer5_outputs(9857) <= b;
    layer5_outputs(9858) <= not a or b;
    layer5_outputs(9859) <= b;
    layer5_outputs(9860) <= a and not b;
    layer5_outputs(9861) <= a xor b;
    layer5_outputs(9862) <= not a or b;
    layer5_outputs(9863) <= not a;
    layer5_outputs(9864) <= not (a or b);
    layer5_outputs(9865) <= 1'b1;
    layer5_outputs(9866) <= a xor b;
    layer5_outputs(9867) <= 1'b1;
    layer5_outputs(9868) <= a and b;
    layer5_outputs(9869) <= not a or b;
    layer5_outputs(9870) <= not (a and b);
    layer5_outputs(9871) <= a and not b;
    layer5_outputs(9872) <= a or b;
    layer5_outputs(9873) <= a or b;
    layer5_outputs(9874) <= 1'b1;
    layer5_outputs(9875) <= not (a or b);
    layer5_outputs(9876) <= a and not b;
    layer5_outputs(9877) <= b;
    layer5_outputs(9878) <= not a or b;
    layer5_outputs(9879) <= not (a or b);
    layer5_outputs(9880) <= not a;
    layer5_outputs(9881) <= not a or b;
    layer5_outputs(9882) <= a;
    layer5_outputs(9883) <= not a or b;
    layer5_outputs(9884) <= not b;
    layer5_outputs(9885) <= not (a xor b);
    layer5_outputs(9886) <= a and not b;
    layer5_outputs(9887) <= a;
    layer5_outputs(9888) <= 1'b0;
    layer5_outputs(9889) <= a;
    layer5_outputs(9890) <= not b;
    layer5_outputs(9891) <= not a or b;
    layer5_outputs(9892) <= a xor b;
    layer5_outputs(9893) <= not (a or b);
    layer5_outputs(9894) <= 1'b0;
    layer5_outputs(9895) <= not a;
    layer5_outputs(9896) <= 1'b1;
    layer5_outputs(9897) <= not (a and b);
    layer5_outputs(9898) <= a;
    layer5_outputs(9899) <= b;
    layer5_outputs(9900) <= b and not a;
    layer5_outputs(9901) <= a and b;
    layer5_outputs(9902) <= 1'b0;
    layer5_outputs(9903) <= 1'b0;
    layer5_outputs(9904) <= not (a or b);
    layer5_outputs(9905) <= a and not b;
    layer5_outputs(9906) <= not b or a;
    layer5_outputs(9907) <= a and b;
    layer5_outputs(9908) <= b and not a;
    layer5_outputs(9909) <= 1'b1;
    layer5_outputs(9910) <= b;
    layer5_outputs(9911) <= not a or b;
    layer5_outputs(9912) <= b;
    layer5_outputs(9913) <= 1'b0;
    layer5_outputs(9914) <= a;
    layer5_outputs(9915) <= a and b;
    layer5_outputs(9916) <= not (a and b);
    layer5_outputs(9917) <= 1'b1;
    layer5_outputs(9918) <= b and not a;
    layer5_outputs(9919) <= not b;
    layer5_outputs(9920) <= not a or b;
    layer5_outputs(9921) <= b and not a;
    layer5_outputs(9922) <= a or b;
    layer5_outputs(9923) <= a;
    layer5_outputs(9924) <= 1'b1;
    layer5_outputs(9925) <= a and b;
    layer5_outputs(9926) <= not a;
    layer5_outputs(9927) <= 1'b1;
    layer5_outputs(9928) <= a;
    layer5_outputs(9929) <= a or b;
    layer5_outputs(9930) <= b and not a;
    layer5_outputs(9931) <= not (a or b);
    layer5_outputs(9932) <= not b;
    layer5_outputs(9933) <= a or b;
    layer5_outputs(9934) <= not b or a;
    layer5_outputs(9935) <= not a;
    layer5_outputs(9936) <= not a or b;
    layer5_outputs(9937) <= not (a and b);
    layer5_outputs(9938) <= b and not a;
    layer5_outputs(9939) <= b;
    layer5_outputs(9940) <= not (a or b);
    layer5_outputs(9941) <= b;
    layer5_outputs(9942) <= a or b;
    layer5_outputs(9943) <= not b;
    layer5_outputs(9944) <= a;
    layer5_outputs(9945) <= b;
    layer5_outputs(9946) <= not (a or b);
    layer5_outputs(9947) <= b and not a;
    layer5_outputs(9948) <= not (a xor b);
    layer5_outputs(9949) <= 1'b0;
    layer5_outputs(9950) <= 1'b1;
    layer5_outputs(9951) <= a;
    layer5_outputs(9952) <= not b or a;
    layer5_outputs(9953) <= a;
    layer5_outputs(9954) <= a and not b;
    layer5_outputs(9955) <= not (a xor b);
    layer5_outputs(9956) <= not a or b;
    layer5_outputs(9957) <= 1'b1;
    layer5_outputs(9958) <= not b;
    layer5_outputs(9959) <= a or b;
    layer5_outputs(9960) <= not (a or b);
    layer5_outputs(9961) <= not (a and b);
    layer5_outputs(9962) <= not a;
    layer5_outputs(9963) <= not b;
    layer5_outputs(9964) <= b and not a;
    layer5_outputs(9965) <= not (a and b);
    layer5_outputs(9966) <= not b;
    layer5_outputs(9967) <= a or b;
    layer5_outputs(9968) <= a;
    layer5_outputs(9969) <= not a;
    layer5_outputs(9970) <= a;
    layer5_outputs(9971) <= b;
    layer5_outputs(9972) <= not (a and b);
    layer5_outputs(9973) <= a;
    layer5_outputs(9974) <= a or b;
    layer5_outputs(9975) <= not b;
    layer5_outputs(9976) <= a and not b;
    layer5_outputs(9977) <= a;
    layer5_outputs(9978) <= not a;
    layer5_outputs(9979) <= b and not a;
    layer5_outputs(9980) <= not b;
    layer5_outputs(9981) <= 1'b0;
    layer5_outputs(9982) <= not b;
    layer5_outputs(9983) <= not b;
    layer5_outputs(9984) <= not a;
    layer5_outputs(9985) <= not a;
    layer5_outputs(9986) <= not b or a;
    layer5_outputs(9987) <= not b;
    layer5_outputs(9988) <= not a;
    layer5_outputs(9989) <= 1'b0;
    layer5_outputs(9990) <= a xor b;
    layer5_outputs(9991) <= not b or a;
    layer5_outputs(9992) <= not b or a;
    layer5_outputs(9993) <= a or b;
    layer5_outputs(9994) <= b;
    layer5_outputs(9995) <= not b or a;
    layer5_outputs(9996) <= 1'b1;
    layer5_outputs(9997) <= not b or a;
    layer5_outputs(9998) <= b;
    layer5_outputs(9999) <= not b;
    layer5_outputs(10000) <= a xor b;
    layer5_outputs(10001) <= a or b;
    layer5_outputs(10002) <= a;
    layer5_outputs(10003) <= not b;
    layer5_outputs(10004) <= not b;
    layer5_outputs(10005) <= b and not a;
    layer5_outputs(10006) <= a xor b;
    layer5_outputs(10007) <= not a or b;
    layer5_outputs(10008) <= b;
    layer5_outputs(10009) <= a;
    layer5_outputs(10010) <= not (a xor b);
    layer5_outputs(10011) <= a and not b;
    layer5_outputs(10012) <= b and not a;
    layer5_outputs(10013) <= a;
    layer5_outputs(10014) <= a;
    layer5_outputs(10015) <= a;
    layer5_outputs(10016) <= not b;
    layer5_outputs(10017) <= a or b;
    layer5_outputs(10018) <= a or b;
    layer5_outputs(10019) <= not b;
    layer5_outputs(10020) <= not b;
    layer5_outputs(10021) <= not (a or b);
    layer5_outputs(10022) <= b;
    layer5_outputs(10023) <= not (a or b);
    layer5_outputs(10024) <= not (a and b);
    layer5_outputs(10025) <= b and not a;
    layer5_outputs(10026) <= b and not a;
    layer5_outputs(10027) <= not b or a;
    layer5_outputs(10028) <= a and not b;
    layer5_outputs(10029) <= a and not b;
    layer5_outputs(10030) <= b;
    layer5_outputs(10031) <= not (a xor b);
    layer5_outputs(10032) <= not b or a;
    layer5_outputs(10033) <= not (a xor b);
    layer5_outputs(10034) <= not a;
    layer5_outputs(10035) <= not (a or b);
    layer5_outputs(10036) <= not b;
    layer5_outputs(10037) <= not (a and b);
    layer5_outputs(10038) <= not b or a;
    layer5_outputs(10039) <= not a;
    layer5_outputs(10040) <= 1'b0;
    layer5_outputs(10041) <= a xor b;
    layer5_outputs(10042) <= not b;
    layer5_outputs(10043) <= not b or a;
    layer5_outputs(10044) <= not b or a;
    layer5_outputs(10045) <= a and not b;
    layer5_outputs(10046) <= not (a xor b);
    layer5_outputs(10047) <= a;
    layer5_outputs(10048) <= a xor b;
    layer5_outputs(10049) <= a and not b;
    layer5_outputs(10050) <= a or b;
    layer5_outputs(10051) <= b;
    layer5_outputs(10052) <= b and not a;
    layer5_outputs(10053) <= a;
    layer5_outputs(10054) <= not b;
    layer5_outputs(10055) <= a xor b;
    layer5_outputs(10056) <= b;
    layer5_outputs(10057) <= a xor b;
    layer5_outputs(10058) <= a and b;
    layer5_outputs(10059) <= a xor b;
    layer5_outputs(10060) <= not b or a;
    layer5_outputs(10061) <= not a;
    layer5_outputs(10062) <= not b or a;
    layer5_outputs(10063) <= a xor b;
    layer5_outputs(10064) <= not (a xor b);
    layer5_outputs(10065) <= not a or b;
    layer5_outputs(10066) <= not (a xor b);
    layer5_outputs(10067) <= b and not a;
    layer5_outputs(10068) <= b;
    layer5_outputs(10069) <= b;
    layer5_outputs(10070) <= a or b;
    layer5_outputs(10071) <= a and b;
    layer5_outputs(10072) <= not b;
    layer5_outputs(10073) <= a;
    layer5_outputs(10074) <= a;
    layer5_outputs(10075) <= not a or b;
    layer5_outputs(10076) <= a or b;
    layer5_outputs(10077) <= 1'b0;
    layer5_outputs(10078) <= not (a or b);
    layer5_outputs(10079) <= not (a or b);
    layer5_outputs(10080) <= a or b;
    layer5_outputs(10081) <= b;
    layer5_outputs(10082) <= not a;
    layer5_outputs(10083) <= not a or b;
    layer5_outputs(10084) <= a or b;
    layer5_outputs(10085) <= b and not a;
    layer5_outputs(10086) <= a or b;
    layer5_outputs(10087) <= a;
    layer5_outputs(10088) <= not (a xor b);
    layer5_outputs(10089) <= b and not a;
    layer5_outputs(10090) <= not a;
    layer5_outputs(10091) <= not (a and b);
    layer5_outputs(10092) <= b;
    layer5_outputs(10093) <= not a;
    layer5_outputs(10094) <= not (a xor b);
    layer5_outputs(10095) <= not (a and b);
    layer5_outputs(10096) <= not (a and b);
    layer5_outputs(10097) <= a and b;
    layer5_outputs(10098) <= a;
    layer5_outputs(10099) <= a and b;
    layer5_outputs(10100) <= not a or b;
    layer5_outputs(10101) <= b;
    layer5_outputs(10102) <= not b;
    layer5_outputs(10103) <= not (a xor b);
    layer5_outputs(10104) <= not (a and b);
    layer5_outputs(10105) <= b;
    layer5_outputs(10106) <= not b;
    layer5_outputs(10107) <= b and not a;
    layer5_outputs(10108) <= a or b;
    layer5_outputs(10109) <= not b or a;
    layer5_outputs(10110) <= not a or b;
    layer5_outputs(10111) <= b;
    layer5_outputs(10112) <= not b or a;
    layer5_outputs(10113) <= not (a or b);
    layer5_outputs(10114) <= 1'b0;
    layer5_outputs(10115) <= b;
    layer5_outputs(10116) <= not b;
    layer5_outputs(10117) <= not a or b;
    layer5_outputs(10118) <= 1'b0;
    layer5_outputs(10119) <= not (a or b);
    layer5_outputs(10120) <= not b or a;
    layer5_outputs(10121) <= a and b;
    layer5_outputs(10122) <= a;
    layer5_outputs(10123) <= not (a xor b);
    layer5_outputs(10124) <= not a;
    layer5_outputs(10125) <= b;
    layer5_outputs(10126) <= b;
    layer5_outputs(10127) <= a or b;
    layer5_outputs(10128) <= not (a and b);
    layer5_outputs(10129) <= not a;
    layer5_outputs(10130) <= not (a or b);
    layer5_outputs(10131) <= not b or a;
    layer5_outputs(10132) <= a or b;
    layer5_outputs(10133) <= not b;
    layer5_outputs(10134) <= not (a or b);
    layer5_outputs(10135) <= not (a xor b);
    layer5_outputs(10136) <= not (a and b);
    layer5_outputs(10137) <= a xor b;
    layer5_outputs(10138) <= b and not a;
    layer5_outputs(10139) <= not b;
    layer5_outputs(10140) <= a;
    layer5_outputs(10141) <= not a;
    layer5_outputs(10142) <= not a or b;
    layer5_outputs(10143) <= b and not a;
    layer5_outputs(10144) <= b;
    layer5_outputs(10145) <= a or b;
    layer5_outputs(10146) <= not a;
    layer5_outputs(10147) <= not a;
    layer5_outputs(10148) <= not b or a;
    layer5_outputs(10149) <= not a;
    layer5_outputs(10150) <= a and not b;
    layer5_outputs(10151) <= a and b;
    layer5_outputs(10152) <= not b;
    layer5_outputs(10153) <= a or b;
    layer5_outputs(10154) <= not (a xor b);
    layer5_outputs(10155) <= a;
    layer5_outputs(10156) <= not b or a;
    layer5_outputs(10157) <= a;
    layer5_outputs(10158) <= not b or a;
    layer5_outputs(10159) <= b;
    layer5_outputs(10160) <= a and not b;
    layer5_outputs(10161) <= b;
    layer5_outputs(10162) <= a;
    layer5_outputs(10163) <= not b;
    layer5_outputs(10164) <= b;
    layer5_outputs(10165) <= not b;
    layer5_outputs(10166) <= not b;
    layer5_outputs(10167) <= a or b;
    layer5_outputs(10168) <= a or b;
    layer5_outputs(10169) <= 1'b1;
    layer5_outputs(10170) <= a and not b;
    layer5_outputs(10171) <= not a;
    layer5_outputs(10172) <= not a;
    layer5_outputs(10173) <= not b;
    layer5_outputs(10174) <= not a or b;
    layer5_outputs(10175) <= a and b;
    layer5_outputs(10176) <= not (a xor b);
    layer5_outputs(10177) <= not (a and b);
    layer5_outputs(10178) <= a and b;
    layer5_outputs(10179) <= 1'b0;
    layer5_outputs(10180) <= not a;
    layer5_outputs(10181) <= not b or a;
    layer5_outputs(10182) <= not (a and b);
    layer5_outputs(10183) <= b;
    layer5_outputs(10184) <= a;
    layer5_outputs(10185) <= a;
    layer5_outputs(10186) <= not (a and b);
    layer5_outputs(10187) <= not b;
    layer5_outputs(10188) <= b;
    layer5_outputs(10189) <= a and b;
    layer5_outputs(10190) <= b;
    layer5_outputs(10191) <= not b or a;
    layer5_outputs(10192) <= a or b;
    layer5_outputs(10193) <= 1'b0;
    layer5_outputs(10194) <= 1'b1;
    layer5_outputs(10195) <= not (a xor b);
    layer5_outputs(10196) <= a;
    layer5_outputs(10197) <= a or b;
    layer5_outputs(10198) <= b;
    layer5_outputs(10199) <= not a;
    layer5_outputs(10200) <= a or b;
    layer5_outputs(10201) <= not b or a;
    layer5_outputs(10202) <= not b or a;
    layer5_outputs(10203) <= not b or a;
    layer5_outputs(10204) <= 1'b1;
    layer5_outputs(10205) <= b;
    layer5_outputs(10206) <= not (a or b);
    layer5_outputs(10207) <= b and not a;
    layer5_outputs(10208) <= a and b;
    layer5_outputs(10209) <= a;
    layer5_outputs(10210) <= not a;
    layer5_outputs(10211) <= b and not a;
    layer5_outputs(10212) <= a;
    layer5_outputs(10213) <= not b or a;
    layer5_outputs(10214) <= not a or b;
    layer5_outputs(10215) <= not b;
    layer5_outputs(10216) <= not a or b;
    layer5_outputs(10217) <= not b;
    layer5_outputs(10218) <= a;
    layer5_outputs(10219) <= a or b;
    layer5_outputs(10220) <= b;
    layer5_outputs(10221) <= a;
    layer5_outputs(10222) <= not a or b;
    layer5_outputs(10223) <= a or b;
    layer5_outputs(10224) <= 1'b1;
    layer5_outputs(10225) <= not b;
    layer5_outputs(10226) <= not b;
    layer5_outputs(10227) <= a;
    layer5_outputs(10228) <= not (a xor b);
    layer5_outputs(10229) <= not a or b;
    layer5_outputs(10230) <= not b;
    layer5_outputs(10231) <= not (a and b);
    layer5_outputs(10232) <= b and not a;
    layer5_outputs(10233) <= not a;
    layer5_outputs(10234) <= not (a or b);
    layer5_outputs(10235) <= b and not a;
    layer5_outputs(10236) <= not (a and b);
    layer5_outputs(10237) <= not (a and b);
    layer5_outputs(10238) <= not b;
    layer5_outputs(10239) <= a xor b;
    layer6_outputs(0) <= not (a or b);
    layer6_outputs(1) <= not (a xor b);
    layer6_outputs(2) <= b;
    layer6_outputs(3) <= a and not b;
    layer6_outputs(4) <= a;
    layer6_outputs(5) <= not (a and b);
    layer6_outputs(6) <= a and b;
    layer6_outputs(7) <= 1'b1;
    layer6_outputs(8) <= a xor b;
    layer6_outputs(9) <= a or b;
    layer6_outputs(10) <= not (a or b);
    layer6_outputs(11) <= b;
    layer6_outputs(12) <= not b;
    layer6_outputs(13) <= not (a or b);
    layer6_outputs(14) <= 1'b1;
    layer6_outputs(15) <= not (a xor b);
    layer6_outputs(16) <= a;
    layer6_outputs(17) <= b;
    layer6_outputs(18) <= not a;
    layer6_outputs(19) <= not (a or b);
    layer6_outputs(20) <= not b;
    layer6_outputs(21) <= not b;
    layer6_outputs(22) <= not b;
    layer6_outputs(23) <= a or b;
    layer6_outputs(24) <= not b;
    layer6_outputs(25) <= not b or a;
    layer6_outputs(26) <= not a;
    layer6_outputs(27) <= not (a and b);
    layer6_outputs(28) <= not b or a;
    layer6_outputs(29) <= a;
    layer6_outputs(30) <= b and not a;
    layer6_outputs(31) <= not a;
    layer6_outputs(32) <= a;
    layer6_outputs(33) <= not (a xor b);
    layer6_outputs(34) <= a;
    layer6_outputs(35) <= not b;
    layer6_outputs(36) <= not (a and b);
    layer6_outputs(37) <= not a or b;
    layer6_outputs(38) <= a and b;
    layer6_outputs(39) <= a and b;
    layer6_outputs(40) <= a and b;
    layer6_outputs(41) <= b and not a;
    layer6_outputs(42) <= not b;
    layer6_outputs(43) <= not b;
    layer6_outputs(44) <= a and b;
    layer6_outputs(45) <= not a;
    layer6_outputs(46) <= not b or a;
    layer6_outputs(47) <= b and not a;
    layer6_outputs(48) <= not b;
    layer6_outputs(49) <= not b or a;
    layer6_outputs(50) <= a or b;
    layer6_outputs(51) <= a and b;
    layer6_outputs(52) <= a and b;
    layer6_outputs(53) <= b and not a;
    layer6_outputs(54) <= a or b;
    layer6_outputs(55) <= a xor b;
    layer6_outputs(56) <= b and not a;
    layer6_outputs(57) <= b;
    layer6_outputs(58) <= not (a xor b);
    layer6_outputs(59) <= b;
    layer6_outputs(60) <= b and not a;
    layer6_outputs(61) <= not (a xor b);
    layer6_outputs(62) <= b;
    layer6_outputs(63) <= b;
    layer6_outputs(64) <= not a or b;
    layer6_outputs(65) <= not b or a;
    layer6_outputs(66) <= a and b;
    layer6_outputs(67) <= not (a or b);
    layer6_outputs(68) <= a or b;
    layer6_outputs(69) <= not (a xor b);
    layer6_outputs(70) <= not (a or b);
    layer6_outputs(71) <= a xor b;
    layer6_outputs(72) <= not a;
    layer6_outputs(73) <= not (a and b);
    layer6_outputs(74) <= b and not a;
    layer6_outputs(75) <= not (a or b);
    layer6_outputs(76) <= not a or b;
    layer6_outputs(77) <= b;
    layer6_outputs(78) <= not b;
    layer6_outputs(79) <= not a;
    layer6_outputs(80) <= not b or a;
    layer6_outputs(81) <= not a;
    layer6_outputs(82) <= a xor b;
    layer6_outputs(83) <= b;
    layer6_outputs(84) <= not a;
    layer6_outputs(85) <= not a;
    layer6_outputs(86) <= not a or b;
    layer6_outputs(87) <= not (a or b);
    layer6_outputs(88) <= not (a and b);
    layer6_outputs(89) <= not a or b;
    layer6_outputs(90) <= not (a or b);
    layer6_outputs(91) <= not (a or b);
    layer6_outputs(92) <= not (a and b);
    layer6_outputs(93) <= not (a and b);
    layer6_outputs(94) <= a or b;
    layer6_outputs(95) <= 1'b0;
    layer6_outputs(96) <= not (a and b);
    layer6_outputs(97) <= a xor b;
    layer6_outputs(98) <= not (a or b);
    layer6_outputs(99) <= a xor b;
    layer6_outputs(100) <= b and not a;
    layer6_outputs(101) <= a;
    layer6_outputs(102) <= a xor b;
    layer6_outputs(103) <= b;
    layer6_outputs(104) <= a and not b;
    layer6_outputs(105) <= b;
    layer6_outputs(106) <= not (a and b);
    layer6_outputs(107) <= not (a and b);
    layer6_outputs(108) <= not b;
    layer6_outputs(109) <= a and not b;
    layer6_outputs(110) <= a;
    layer6_outputs(111) <= not a or b;
    layer6_outputs(112) <= not b;
    layer6_outputs(113) <= a and b;
    layer6_outputs(114) <= not (a and b);
    layer6_outputs(115) <= a and b;
    layer6_outputs(116) <= b;
    layer6_outputs(117) <= a;
    layer6_outputs(118) <= a or b;
    layer6_outputs(119) <= not (a xor b);
    layer6_outputs(120) <= b;
    layer6_outputs(121) <= a or b;
    layer6_outputs(122) <= a and not b;
    layer6_outputs(123) <= a xor b;
    layer6_outputs(124) <= not (a xor b);
    layer6_outputs(125) <= b;
    layer6_outputs(126) <= a xor b;
    layer6_outputs(127) <= not b;
    layer6_outputs(128) <= a;
    layer6_outputs(129) <= 1'b0;
    layer6_outputs(130) <= not (a or b);
    layer6_outputs(131) <= not a;
    layer6_outputs(132) <= not a;
    layer6_outputs(133) <= not a;
    layer6_outputs(134) <= 1'b0;
    layer6_outputs(135) <= a and b;
    layer6_outputs(136) <= a and not b;
    layer6_outputs(137) <= not b;
    layer6_outputs(138) <= not a;
    layer6_outputs(139) <= not b or a;
    layer6_outputs(140) <= b;
    layer6_outputs(141) <= a;
    layer6_outputs(142) <= b;
    layer6_outputs(143) <= not (a and b);
    layer6_outputs(144) <= a or b;
    layer6_outputs(145) <= a or b;
    layer6_outputs(146) <= b;
    layer6_outputs(147) <= not b;
    layer6_outputs(148) <= a;
    layer6_outputs(149) <= b;
    layer6_outputs(150) <= b and not a;
    layer6_outputs(151) <= not a;
    layer6_outputs(152) <= b;
    layer6_outputs(153) <= a;
    layer6_outputs(154) <= a xor b;
    layer6_outputs(155) <= 1'b1;
    layer6_outputs(156) <= not a;
    layer6_outputs(157) <= not b or a;
    layer6_outputs(158) <= not a or b;
    layer6_outputs(159) <= a or b;
    layer6_outputs(160) <= a and not b;
    layer6_outputs(161) <= not (a or b);
    layer6_outputs(162) <= a or b;
    layer6_outputs(163) <= a and not b;
    layer6_outputs(164) <= a xor b;
    layer6_outputs(165) <= not b or a;
    layer6_outputs(166) <= b;
    layer6_outputs(167) <= a;
    layer6_outputs(168) <= not (a or b);
    layer6_outputs(169) <= not (a and b);
    layer6_outputs(170) <= not b or a;
    layer6_outputs(171) <= b;
    layer6_outputs(172) <= b;
    layer6_outputs(173) <= not b or a;
    layer6_outputs(174) <= a or b;
    layer6_outputs(175) <= a or b;
    layer6_outputs(176) <= b;
    layer6_outputs(177) <= b;
    layer6_outputs(178) <= not (a or b);
    layer6_outputs(179) <= not a or b;
    layer6_outputs(180) <= b and not a;
    layer6_outputs(181) <= not b;
    layer6_outputs(182) <= not a;
    layer6_outputs(183) <= not b or a;
    layer6_outputs(184) <= not a;
    layer6_outputs(185) <= b and not a;
    layer6_outputs(186) <= not (a xor b);
    layer6_outputs(187) <= b;
    layer6_outputs(188) <= not a or b;
    layer6_outputs(189) <= b;
    layer6_outputs(190) <= 1'b1;
    layer6_outputs(191) <= a or b;
    layer6_outputs(192) <= a;
    layer6_outputs(193) <= not b or a;
    layer6_outputs(194) <= not (a xor b);
    layer6_outputs(195) <= not (a xor b);
    layer6_outputs(196) <= not b or a;
    layer6_outputs(197) <= not (a and b);
    layer6_outputs(198) <= b;
    layer6_outputs(199) <= not b or a;
    layer6_outputs(200) <= a and b;
    layer6_outputs(201) <= a;
    layer6_outputs(202) <= a;
    layer6_outputs(203) <= not (a or b);
    layer6_outputs(204) <= not b or a;
    layer6_outputs(205) <= not (a and b);
    layer6_outputs(206) <= a and b;
    layer6_outputs(207) <= a and b;
    layer6_outputs(208) <= not b;
    layer6_outputs(209) <= b;
    layer6_outputs(210) <= not a or b;
    layer6_outputs(211) <= b and not a;
    layer6_outputs(212) <= not b or a;
    layer6_outputs(213) <= a xor b;
    layer6_outputs(214) <= 1'b0;
    layer6_outputs(215) <= not (a xor b);
    layer6_outputs(216) <= not (a or b);
    layer6_outputs(217) <= a and not b;
    layer6_outputs(218) <= not a;
    layer6_outputs(219) <= a;
    layer6_outputs(220) <= not b;
    layer6_outputs(221) <= a or b;
    layer6_outputs(222) <= b;
    layer6_outputs(223) <= b;
    layer6_outputs(224) <= not b or a;
    layer6_outputs(225) <= not a;
    layer6_outputs(226) <= 1'b1;
    layer6_outputs(227) <= not a;
    layer6_outputs(228) <= b and not a;
    layer6_outputs(229) <= b;
    layer6_outputs(230) <= not b;
    layer6_outputs(231) <= not a;
    layer6_outputs(232) <= not b;
    layer6_outputs(233) <= b;
    layer6_outputs(234) <= b;
    layer6_outputs(235) <= not b;
    layer6_outputs(236) <= a;
    layer6_outputs(237) <= b;
    layer6_outputs(238) <= not b;
    layer6_outputs(239) <= b;
    layer6_outputs(240) <= not b or a;
    layer6_outputs(241) <= not b;
    layer6_outputs(242) <= a and not b;
    layer6_outputs(243) <= b and not a;
    layer6_outputs(244) <= a;
    layer6_outputs(245) <= not a;
    layer6_outputs(246) <= a and b;
    layer6_outputs(247) <= b;
    layer6_outputs(248) <= not (a or b);
    layer6_outputs(249) <= not b;
    layer6_outputs(250) <= not (a and b);
    layer6_outputs(251) <= not a;
    layer6_outputs(252) <= b;
    layer6_outputs(253) <= a or b;
    layer6_outputs(254) <= a xor b;
    layer6_outputs(255) <= b and not a;
    layer6_outputs(256) <= not b or a;
    layer6_outputs(257) <= not b;
    layer6_outputs(258) <= a and b;
    layer6_outputs(259) <= not a;
    layer6_outputs(260) <= a;
    layer6_outputs(261) <= a and not b;
    layer6_outputs(262) <= not b;
    layer6_outputs(263) <= not b;
    layer6_outputs(264) <= not a;
    layer6_outputs(265) <= not (a xor b);
    layer6_outputs(266) <= not (a xor b);
    layer6_outputs(267) <= not b;
    layer6_outputs(268) <= not (a or b);
    layer6_outputs(269) <= b;
    layer6_outputs(270) <= b and not a;
    layer6_outputs(271) <= b;
    layer6_outputs(272) <= a xor b;
    layer6_outputs(273) <= not b;
    layer6_outputs(274) <= not b;
    layer6_outputs(275) <= not a or b;
    layer6_outputs(276) <= not a;
    layer6_outputs(277) <= 1'b0;
    layer6_outputs(278) <= not b or a;
    layer6_outputs(279) <= not (a or b);
    layer6_outputs(280) <= not b;
    layer6_outputs(281) <= a or b;
    layer6_outputs(282) <= b and not a;
    layer6_outputs(283) <= not (a or b);
    layer6_outputs(284) <= b;
    layer6_outputs(285) <= a and b;
    layer6_outputs(286) <= not b;
    layer6_outputs(287) <= not (a xor b);
    layer6_outputs(288) <= 1'b1;
    layer6_outputs(289) <= b;
    layer6_outputs(290) <= not b;
    layer6_outputs(291) <= a;
    layer6_outputs(292) <= not a or b;
    layer6_outputs(293) <= not (a and b);
    layer6_outputs(294) <= not (a or b);
    layer6_outputs(295) <= not b;
    layer6_outputs(296) <= a and not b;
    layer6_outputs(297) <= 1'b1;
    layer6_outputs(298) <= a and not b;
    layer6_outputs(299) <= b;
    layer6_outputs(300) <= 1'b1;
    layer6_outputs(301) <= not b;
    layer6_outputs(302) <= not (a and b);
    layer6_outputs(303) <= not (a or b);
    layer6_outputs(304) <= not b or a;
    layer6_outputs(305) <= b;
    layer6_outputs(306) <= not (a and b);
    layer6_outputs(307) <= a and not b;
    layer6_outputs(308) <= a or b;
    layer6_outputs(309) <= a;
    layer6_outputs(310) <= not a;
    layer6_outputs(311) <= b;
    layer6_outputs(312) <= not a or b;
    layer6_outputs(313) <= a xor b;
    layer6_outputs(314) <= a;
    layer6_outputs(315) <= 1'b0;
    layer6_outputs(316) <= not a;
    layer6_outputs(317) <= not (a xor b);
    layer6_outputs(318) <= not b or a;
    layer6_outputs(319) <= not b;
    layer6_outputs(320) <= a xor b;
    layer6_outputs(321) <= not (a and b);
    layer6_outputs(322) <= b;
    layer6_outputs(323) <= not a;
    layer6_outputs(324) <= not b;
    layer6_outputs(325) <= not a;
    layer6_outputs(326) <= not a;
    layer6_outputs(327) <= a xor b;
    layer6_outputs(328) <= not a or b;
    layer6_outputs(329) <= not b or a;
    layer6_outputs(330) <= a xor b;
    layer6_outputs(331) <= not a;
    layer6_outputs(332) <= not (a or b);
    layer6_outputs(333) <= not (a xor b);
    layer6_outputs(334) <= not a or b;
    layer6_outputs(335) <= not a or b;
    layer6_outputs(336) <= a;
    layer6_outputs(337) <= 1'b1;
    layer6_outputs(338) <= b and not a;
    layer6_outputs(339) <= b;
    layer6_outputs(340) <= b and not a;
    layer6_outputs(341) <= a xor b;
    layer6_outputs(342) <= b;
    layer6_outputs(343) <= a or b;
    layer6_outputs(344) <= not (a or b);
    layer6_outputs(345) <= not b;
    layer6_outputs(346) <= not (a xor b);
    layer6_outputs(347) <= not b;
    layer6_outputs(348) <= not b;
    layer6_outputs(349) <= not b or a;
    layer6_outputs(350) <= a and b;
    layer6_outputs(351) <= not b;
    layer6_outputs(352) <= b;
    layer6_outputs(353) <= not (a or b);
    layer6_outputs(354) <= a;
    layer6_outputs(355) <= a xor b;
    layer6_outputs(356) <= b;
    layer6_outputs(357) <= a;
    layer6_outputs(358) <= a;
    layer6_outputs(359) <= not a;
    layer6_outputs(360) <= not (a xor b);
    layer6_outputs(361) <= not b;
    layer6_outputs(362) <= a xor b;
    layer6_outputs(363) <= a;
    layer6_outputs(364) <= not a;
    layer6_outputs(365) <= not a or b;
    layer6_outputs(366) <= a and b;
    layer6_outputs(367) <= not a;
    layer6_outputs(368) <= not (a or b);
    layer6_outputs(369) <= a xor b;
    layer6_outputs(370) <= a;
    layer6_outputs(371) <= a;
    layer6_outputs(372) <= a or b;
    layer6_outputs(373) <= b and not a;
    layer6_outputs(374) <= a;
    layer6_outputs(375) <= not a;
    layer6_outputs(376) <= not (a and b);
    layer6_outputs(377) <= not b;
    layer6_outputs(378) <= not a;
    layer6_outputs(379) <= a and not b;
    layer6_outputs(380) <= not (a xor b);
    layer6_outputs(381) <= b and not a;
    layer6_outputs(382) <= not a or b;
    layer6_outputs(383) <= a;
    layer6_outputs(384) <= b;
    layer6_outputs(385) <= a or b;
    layer6_outputs(386) <= not b;
    layer6_outputs(387) <= a;
    layer6_outputs(388) <= b;
    layer6_outputs(389) <= not a or b;
    layer6_outputs(390) <= a;
    layer6_outputs(391) <= not b;
    layer6_outputs(392) <= a and b;
    layer6_outputs(393) <= not b or a;
    layer6_outputs(394) <= not b or a;
    layer6_outputs(395) <= a or b;
    layer6_outputs(396) <= not a;
    layer6_outputs(397) <= not a;
    layer6_outputs(398) <= not (a xor b);
    layer6_outputs(399) <= b and not a;
    layer6_outputs(400) <= not a;
    layer6_outputs(401) <= a;
    layer6_outputs(402) <= b;
    layer6_outputs(403) <= not (a and b);
    layer6_outputs(404) <= b;
    layer6_outputs(405) <= not a or b;
    layer6_outputs(406) <= not (a or b);
    layer6_outputs(407) <= a;
    layer6_outputs(408) <= not a;
    layer6_outputs(409) <= a or b;
    layer6_outputs(410) <= a and not b;
    layer6_outputs(411) <= not (a or b);
    layer6_outputs(412) <= a or b;
    layer6_outputs(413) <= a and b;
    layer6_outputs(414) <= not a;
    layer6_outputs(415) <= not b or a;
    layer6_outputs(416) <= b;
    layer6_outputs(417) <= 1'b1;
    layer6_outputs(418) <= a;
    layer6_outputs(419) <= not b or a;
    layer6_outputs(420) <= 1'b0;
    layer6_outputs(421) <= b;
    layer6_outputs(422) <= not b;
    layer6_outputs(423) <= not b;
    layer6_outputs(424) <= b and not a;
    layer6_outputs(425) <= a xor b;
    layer6_outputs(426) <= not a or b;
    layer6_outputs(427) <= not (a xor b);
    layer6_outputs(428) <= a;
    layer6_outputs(429) <= b;
    layer6_outputs(430) <= a;
    layer6_outputs(431) <= not a or b;
    layer6_outputs(432) <= not (a and b);
    layer6_outputs(433) <= not b;
    layer6_outputs(434) <= b;
    layer6_outputs(435) <= not (a and b);
    layer6_outputs(436) <= not b;
    layer6_outputs(437) <= 1'b1;
    layer6_outputs(438) <= not b;
    layer6_outputs(439) <= a and b;
    layer6_outputs(440) <= 1'b1;
    layer6_outputs(441) <= not (a or b);
    layer6_outputs(442) <= a xor b;
    layer6_outputs(443) <= a and b;
    layer6_outputs(444) <= a;
    layer6_outputs(445) <= b and not a;
    layer6_outputs(446) <= a and b;
    layer6_outputs(447) <= not a;
    layer6_outputs(448) <= not a;
    layer6_outputs(449) <= not b or a;
    layer6_outputs(450) <= not a;
    layer6_outputs(451) <= not a;
    layer6_outputs(452) <= b and not a;
    layer6_outputs(453) <= a and b;
    layer6_outputs(454) <= not a;
    layer6_outputs(455) <= 1'b1;
    layer6_outputs(456) <= 1'b1;
    layer6_outputs(457) <= not b or a;
    layer6_outputs(458) <= a and b;
    layer6_outputs(459) <= not (a and b);
    layer6_outputs(460) <= not a or b;
    layer6_outputs(461) <= not a;
    layer6_outputs(462) <= a;
    layer6_outputs(463) <= b;
    layer6_outputs(464) <= b;
    layer6_outputs(465) <= not a;
    layer6_outputs(466) <= not (a or b);
    layer6_outputs(467) <= not a;
    layer6_outputs(468) <= a;
    layer6_outputs(469) <= b and not a;
    layer6_outputs(470) <= not a;
    layer6_outputs(471) <= b and not a;
    layer6_outputs(472) <= b and not a;
    layer6_outputs(473) <= not (a or b);
    layer6_outputs(474) <= not (a xor b);
    layer6_outputs(475) <= not (a xor b);
    layer6_outputs(476) <= b;
    layer6_outputs(477) <= b;
    layer6_outputs(478) <= not b;
    layer6_outputs(479) <= not (a or b);
    layer6_outputs(480) <= a and b;
    layer6_outputs(481) <= a and b;
    layer6_outputs(482) <= a;
    layer6_outputs(483) <= not a;
    layer6_outputs(484) <= b;
    layer6_outputs(485) <= not (a or b);
    layer6_outputs(486) <= a and b;
    layer6_outputs(487) <= not b or a;
    layer6_outputs(488) <= not b;
    layer6_outputs(489) <= a;
    layer6_outputs(490) <= not b;
    layer6_outputs(491) <= b and not a;
    layer6_outputs(492) <= not b;
    layer6_outputs(493) <= a and b;
    layer6_outputs(494) <= a;
    layer6_outputs(495) <= a or b;
    layer6_outputs(496) <= not a;
    layer6_outputs(497) <= b and not a;
    layer6_outputs(498) <= a and b;
    layer6_outputs(499) <= a;
    layer6_outputs(500) <= b;
    layer6_outputs(501) <= b;
    layer6_outputs(502) <= not (a and b);
    layer6_outputs(503) <= b;
    layer6_outputs(504) <= not a or b;
    layer6_outputs(505) <= b;
    layer6_outputs(506) <= not b or a;
    layer6_outputs(507) <= not a or b;
    layer6_outputs(508) <= not (a xor b);
    layer6_outputs(509) <= not (a or b);
    layer6_outputs(510) <= not b or a;
    layer6_outputs(511) <= a or b;
    layer6_outputs(512) <= not (a xor b);
    layer6_outputs(513) <= b;
    layer6_outputs(514) <= a and b;
    layer6_outputs(515) <= not b or a;
    layer6_outputs(516) <= 1'b0;
    layer6_outputs(517) <= not a or b;
    layer6_outputs(518) <= not (a or b);
    layer6_outputs(519) <= not a;
    layer6_outputs(520) <= not (a and b);
    layer6_outputs(521) <= a;
    layer6_outputs(522) <= 1'b1;
    layer6_outputs(523) <= b;
    layer6_outputs(524) <= b;
    layer6_outputs(525) <= not (a or b);
    layer6_outputs(526) <= b;
    layer6_outputs(527) <= not b or a;
    layer6_outputs(528) <= not a;
    layer6_outputs(529) <= a;
    layer6_outputs(530) <= not b;
    layer6_outputs(531) <= not a or b;
    layer6_outputs(532) <= not b;
    layer6_outputs(533) <= a;
    layer6_outputs(534) <= a or b;
    layer6_outputs(535) <= 1'b0;
    layer6_outputs(536) <= b;
    layer6_outputs(537) <= a xor b;
    layer6_outputs(538) <= a or b;
    layer6_outputs(539) <= not (a or b);
    layer6_outputs(540) <= a xor b;
    layer6_outputs(541) <= a xor b;
    layer6_outputs(542) <= not a or b;
    layer6_outputs(543) <= not (a xor b);
    layer6_outputs(544) <= b and not a;
    layer6_outputs(545) <= not a;
    layer6_outputs(546) <= not b or a;
    layer6_outputs(547) <= not a;
    layer6_outputs(548) <= a xor b;
    layer6_outputs(549) <= a xor b;
    layer6_outputs(550) <= b;
    layer6_outputs(551) <= not b or a;
    layer6_outputs(552) <= not (a or b);
    layer6_outputs(553) <= not a or b;
    layer6_outputs(554) <= not a or b;
    layer6_outputs(555) <= a xor b;
    layer6_outputs(556) <= a xor b;
    layer6_outputs(557) <= not b or a;
    layer6_outputs(558) <= a or b;
    layer6_outputs(559) <= not (a xor b);
    layer6_outputs(560) <= not (a or b);
    layer6_outputs(561) <= not b;
    layer6_outputs(562) <= not a;
    layer6_outputs(563) <= a xor b;
    layer6_outputs(564) <= b and not a;
    layer6_outputs(565) <= 1'b1;
    layer6_outputs(566) <= not b;
    layer6_outputs(567) <= not b;
    layer6_outputs(568) <= not b;
    layer6_outputs(569) <= not a or b;
    layer6_outputs(570) <= a or b;
    layer6_outputs(571) <= a and b;
    layer6_outputs(572) <= not a or b;
    layer6_outputs(573) <= not b or a;
    layer6_outputs(574) <= b;
    layer6_outputs(575) <= not a;
    layer6_outputs(576) <= a and b;
    layer6_outputs(577) <= b and not a;
    layer6_outputs(578) <= not (a and b);
    layer6_outputs(579) <= not a;
    layer6_outputs(580) <= not b;
    layer6_outputs(581) <= b;
    layer6_outputs(582) <= not b;
    layer6_outputs(583) <= b;
    layer6_outputs(584) <= 1'b1;
    layer6_outputs(585) <= a or b;
    layer6_outputs(586) <= not (a xor b);
    layer6_outputs(587) <= a;
    layer6_outputs(588) <= not (a xor b);
    layer6_outputs(589) <= not a or b;
    layer6_outputs(590) <= b;
    layer6_outputs(591) <= a and b;
    layer6_outputs(592) <= a or b;
    layer6_outputs(593) <= a and b;
    layer6_outputs(594) <= a;
    layer6_outputs(595) <= not b or a;
    layer6_outputs(596) <= not (a xor b);
    layer6_outputs(597) <= a;
    layer6_outputs(598) <= not b;
    layer6_outputs(599) <= 1'b1;
    layer6_outputs(600) <= not b;
    layer6_outputs(601) <= not b or a;
    layer6_outputs(602) <= 1'b0;
    layer6_outputs(603) <= not b;
    layer6_outputs(604) <= not b;
    layer6_outputs(605) <= b and not a;
    layer6_outputs(606) <= a xor b;
    layer6_outputs(607) <= a;
    layer6_outputs(608) <= 1'b0;
    layer6_outputs(609) <= a or b;
    layer6_outputs(610) <= not (a xor b);
    layer6_outputs(611) <= b and not a;
    layer6_outputs(612) <= a and b;
    layer6_outputs(613) <= not a;
    layer6_outputs(614) <= b and not a;
    layer6_outputs(615) <= not a;
    layer6_outputs(616) <= b and not a;
    layer6_outputs(617) <= a;
    layer6_outputs(618) <= a or b;
    layer6_outputs(619) <= not (a or b);
    layer6_outputs(620) <= not (a or b);
    layer6_outputs(621) <= a xor b;
    layer6_outputs(622) <= a or b;
    layer6_outputs(623) <= not (a and b);
    layer6_outputs(624) <= not (a or b);
    layer6_outputs(625) <= b and not a;
    layer6_outputs(626) <= not (a or b);
    layer6_outputs(627) <= not (a or b);
    layer6_outputs(628) <= b;
    layer6_outputs(629) <= not (a xor b);
    layer6_outputs(630) <= a xor b;
    layer6_outputs(631) <= not (a and b);
    layer6_outputs(632) <= a and not b;
    layer6_outputs(633) <= a;
    layer6_outputs(634) <= not b;
    layer6_outputs(635) <= not a;
    layer6_outputs(636) <= not a or b;
    layer6_outputs(637) <= not (a xor b);
    layer6_outputs(638) <= not b or a;
    layer6_outputs(639) <= b;
    layer6_outputs(640) <= not (a and b);
    layer6_outputs(641) <= a;
    layer6_outputs(642) <= not a;
    layer6_outputs(643) <= b;
    layer6_outputs(644) <= not b;
    layer6_outputs(645) <= not b;
    layer6_outputs(646) <= not (a xor b);
    layer6_outputs(647) <= a and not b;
    layer6_outputs(648) <= not a;
    layer6_outputs(649) <= not (a or b);
    layer6_outputs(650) <= not a;
    layer6_outputs(651) <= b;
    layer6_outputs(652) <= a and not b;
    layer6_outputs(653) <= not b or a;
    layer6_outputs(654) <= b;
    layer6_outputs(655) <= not b or a;
    layer6_outputs(656) <= not (a or b);
    layer6_outputs(657) <= not b;
    layer6_outputs(658) <= a and not b;
    layer6_outputs(659) <= not a;
    layer6_outputs(660) <= b and not a;
    layer6_outputs(661) <= b;
    layer6_outputs(662) <= a and not b;
    layer6_outputs(663) <= not a;
    layer6_outputs(664) <= 1'b1;
    layer6_outputs(665) <= not (a xor b);
    layer6_outputs(666) <= not (a or b);
    layer6_outputs(667) <= a;
    layer6_outputs(668) <= not b;
    layer6_outputs(669) <= a or b;
    layer6_outputs(670) <= not b;
    layer6_outputs(671) <= not (a or b);
    layer6_outputs(672) <= not a;
    layer6_outputs(673) <= b and not a;
    layer6_outputs(674) <= not (a and b);
    layer6_outputs(675) <= not a or b;
    layer6_outputs(676) <= a;
    layer6_outputs(677) <= b;
    layer6_outputs(678) <= not b;
    layer6_outputs(679) <= not b;
    layer6_outputs(680) <= not b or a;
    layer6_outputs(681) <= a;
    layer6_outputs(682) <= a or b;
    layer6_outputs(683) <= not (a xor b);
    layer6_outputs(684) <= not b;
    layer6_outputs(685) <= not b;
    layer6_outputs(686) <= not a;
    layer6_outputs(687) <= a and not b;
    layer6_outputs(688) <= 1'b1;
    layer6_outputs(689) <= b;
    layer6_outputs(690) <= a or b;
    layer6_outputs(691) <= not b or a;
    layer6_outputs(692) <= a;
    layer6_outputs(693) <= a;
    layer6_outputs(694) <= not (a or b);
    layer6_outputs(695) <= not a;
    layer6_outputs(696) <= not a or b;
    layer6_outputs(697) <= not a or b;
    layer6_outputs(698) <= b;
    layer6_outputs(699) <= a;
    layer6_outputs(700) <= not b;
    layer6_outputs(701) <= not (a or b);
    layer6_outputs(702) <= not b;
    layer6_outputs(703) <= a;
    layer6_outputs(704) <= a or b;
    layer6_outputs(705) <= not a;
    layer6_outputs(706) <= a or b;
    layer6_outputs(707) <= a;
    layer6_outputs(708) <= b;
    layer6_outputs(709) <= not a or b;
    layer6_outputs(710) <= not b;
    layer6_outputs(711) <= not b;
    layer6_outputs(712) <= a or b;
    layer6_outputs(713) <= a and not b;
    layer6_outputs(714) <= not a;
    layer6_outputs(715) <= not a;
    layer6_outputs(716) <= b;
    layer6_outputs(717) <= not b;
    layer6_outputs(718) <= a and not b;
    layer6_outputs(719) <= not b;
    layer6_outputs(720) <= not b or a;
    layer6_outputs(721) <= a xor b;
    layer6_outputs(722) <= not a;
    layer6_outputs(723) <= a or b;
    layer6_outputs(724) <= not b;
    layer6_outputs(725) <= not a;
    layer6_outputs(726) <= not b;
    layer6_outputs(727) <= not b;
    layer6_outputs(728) <= a;
    layer6_outputs(729) <= not (a xor b);
    layer6_outputs(730) <= not b or a;
    layer6_outputs(731) <= not (a or b);
    layer6_outputs(732) <= b and not a;
    layer6_outputs(733) <= not a;
    layer6_outputs(734) <= not b or a;
    layer6_outputs(735) <= not (a xor b);
    layer6_outputs(736) <= not (a and b);
    layer6_outputs(737) <= a;
    layer6_outputs(738) <= not (a xor b);
    layer6_outputs(739) <= not (a xor b);
    layer6_outputs(740) <= b;
    layer6_outputs(741) <= a and b;
    layer6_outputs(742) <= b;
    layer6_outputs(743) <= not (a xor b);
    layer6_outputs(744) <= not a;
    layer6_outputs(745) <= a or b;
    layer6_outputs(746) <= not b;
    layer6_outputs(747) <= not b or a;
    layer6_outputs(748) <= b;
    layer6_outputs(749) <= a and b;
    layer6_outputs(750) <= 1'b0;
    layer6_outputs(751) <= a;
    layer6_outputs(752) <= not (a and b);
    layer6_outputs(753) <= 1'b1;
    layer6_outputs(754) <= not b or a;
    layer6_outputs(755) <= a;
    layer6_outputs(756) <= not a or b;
    layer6_outputs(757) <= a;
    layer6_outputs(758) <= not (a and b);
    layer6_outputs(759) <= 1'b1;
    layer6_outputs(760) <= a;
    layer6_outputs(761) <= not (a or b);
    layer6_outputs(762) <= a;
    layer6_outputs(763) <= a xor b;
    layer6_outputs(764) <= not (a or b);
    layer6_outputs(765) <= not b or a;
    layer6_outputs(766) <= not a;
    layer6_outputs(767) <= not (a xor b);
    layer6_outputs(768) <= not a or b;
    layer6_outputs(769) <= b;
    layer6_outputs(770) <= b and not a;
    layer6_outputs(771) <= not b;
    layer6_outputs(772) <= not a;
    layer6_outputs(773) <= not b;
    layer6_outputs(774) <= not a;
    layer6_outputs(775) <= not b;
    layer6_outputs(776) <= not b;
    layer6_outputs(777) <= b and not a;
    layer6_outputs(778) <= b and not a;
    layer6_outputs(779) <= 1'b1;
    layer6_outputs(780) <= b;
    layer6_outputs(781) <= not (a and b);
    layer6_outputs(782) <= not (a xor b);
    layer6_outputs(783) <= not a;
    layer6_outputs(784) <= b;
    layer6_outputs(785) <= not a or b;
    layer6_outputs(786) <= not (a xor b);
    layer6_outputs(787) <= 1'b0;
    layer6_outputs(788) <= b;
    layer6_outputs(789) <= a;
    layer6_outputs(790) <= not b;
    layer6_outputs(791) <= b and not a;
    layer6_outputs(792) <= not a;
    layer6_outputs(793) <= a xor b;
    layer6_outputs(794) <= b;
    layer6_outputs(795) <= 1'b1;
    layer6_outputs(796) <= a or b;
    layer6_outputs(797) <= a or b;
    layer6_outputs(798) <= a xor b;
    layer6_outputs(799) <= not b;
    layer6_outputs(800) <= not (a or b);
    layer6_outputs(801) <= a and not b;
    layer6_outputs(802) <= a and not b;
    layer6_outputs(803) <= not a;
    layer6_outputs(804) <= not b;
    layer6_outputs(805) <= not (a xor b);
    layer6_outputs(806) <= not a or b;
    layer6_outputs(807) <= b;
    layer6_outputs(808) <= not (a and b);
    layer6_outputs(809) <= a and not b;
    layer6_outputs(810) <= b;
    layer6_outputs(811) <= not a;
    layer6_outputs(812) <= not b;
    layer6_outputs(813) <= not a or b;
    layer6_outputs(814) <= not a;
    layer6_outputs(815) <= 1'b1;
    layer6_outputs(816) <= not (a xor b);
    layer6_outputs(817) <= not b;
    layer6_outputs(818) <= a xor b;
    layer6_outputs(819) <= a xor b;
    layer6_outputs(820) <= 1'b0;
    layer6_outputs(821) <= 1'b0;
    layer6_outputs(822) <= a and b;
    layer6_outputs(823) <= not b;
    layer6_outputs(824) <= b;
    layer6_outputs(825) <= not b or a;
    layer6_outputs(826) <= b;
    layer6_outputs(827) <= a and b;
    layer6_outputs(828) <= b and not a;
    layer6_outputs(829) <= not b or a;
    layer6_outputs(830) <= a and b;
    layer6_outputs(831) <= a and not b;
    layer6_outputs(832) <= a;
    layer6_outputs(833) <= a or b;
    layer6_outputs(834) <= a;
    layer6_outputs(835) <= a and b;
    layer6_outputs(836) <= a xor b;
    layer6_outputs(837) <= a;
    layer6_outputs(838) <= a and b;
    layer6_outputs(839) <= not (a and b);
    layer6_outputs(840) <= a or b;
    layer6_outputs(841) <= a and b;
    layer6_outputs(842) <= a;
    layer6_outputs(843) <= a;
    layer6_outputs(844) <= a or b;
    layer6_outputs(845) <= a and not b;
    layer6_outputs(846) <= not a or b;
    layer6_outputs(847) <= a or b;
    layer6_outputs(848) <= a xor b;
    layer6_outputs(849) <= b;
    layer6_outputs(850) <= b;
    layer6_outputs(851) <= b and not a;
    layer6_outputs(852) <= a xor b;
    layer6_outputs(853) <= not a;
    layer6_outputs(854) <= not (a and b);
    layer6_outputs(855) <= b;
    layer6_outputs(856) <= not (a xor b);
    layer6_outputs(857) <= not b;
    layer6_outputs(858) <= b and not a;
    layer6_outputs(859) <= not b;
    layer6_outputs(860) <= not (a and b);
    layer6_outputs(861) <= a xor b;
    layer6_outputs(862) <= not b or a;
    layer6_outputs(863) <= a;
    layer6_outputs(864) <= not b;
    layer6_outputs(865) <= not b;
    layer6_outputs(866) <= not b or a;
    layer6_outputs(867) <= not (a or b);
    layer6_outputs(868) <= a and not b;
    layer6_outputs(869) <= not a or b;
    layer6_outputs(870) <= not (a xor b);
    layer6_outputs(871) <= b;
    layer6_outputs(872) <= a xor b;
    layer6_outputs(873) <= a;
    layer6_outputs(874) <= a;
    layer6_outputs(875) <= not a;
    layer6_outputs(876) <= a or b;
    layer6_outputs(877) <= not (a xor b);
    layer6_outputs(878) <= not a;
    layer6_outputs(879) <= b and not a;
    layer6_outputs(880) <= not b or a;
    layer6_outputs(881) <= a xor b;
    layer6_outputs(882) <= a and not b;
    layer6_outputs(883) <= a and not b;
    layer6_outputs(884) <= a;
    layer6_outputs(885) <= not a;
    layer6_outputs(886) <= a and not b;
    layer6_outputs(887) <= a;
    layer6_outputs(888) <= b;
    layer6_outputs(889) <= not (a and b);
    layer6_outputs(890) <= not (a or b);
    layer6_outputs(891) <= not (a and b);
    layer6_outputs(892) <= not b;
    layer6_outputs(893) <= not (a and b);
    layer6_outputs(894) <= a;
    layer6_outputs(895) <= a;
    layer6_outputs(896) <= a and not b;
    layer6_outputs(897) <= not b;
    layer6_outputs(898) <= b;
    layer6_outputs(899) <= not a;
    layer6_outputs(900) <= a;
    layer6_outputs(901) <= not a;
    layer6_outputs(902) <= b and not a;
    layer6_outputs(903) <= not b;
    layer6_outputs(904) <= b;
    layer6_outputs(905) <= not b;
    layer6_outputs(906) <= a;
    layer6_outputs(907) <= not a or b;
    layer6_outputs(908) <= not (a and b);
    layer6_outputs(909) <= 1'b0;
    layer6_outputs(910) <= a;
    layer6_outputs(911) <= a or b;
    layer6_outputs(912) <= a and b;
    layer6_outputs(913) <= not a;
    layer6_outputs(914) <= a or b;
    layer6_outputs(915) <= a and b;
    layer6_outputs(916) <= a or b;
    layer6_outputs(917) <= a or b;
    layer6_outputs(918) <= not (a or b);
    layer6_outputs(919) <= not b or a;
    layer6_outputs(920) <= not (a xor b);
    layer6_outputs(921) <= a and not b;
    layer6_outputs(922) <= not b or a;
    layer6_outputs(923) <= b and not a;
    layer6_outputs(924) <= a;
    layer6_outputs(925) <= b;
    layer6_outputs(926) <= not b or a;
    layer6_outputs(927) <= not b or a;
    layer6_outputs(928) <= not (a and b);
    layer6_outputs(929) <= a xor b;
    layer6_outputs(930) <= not b;
    layer6_outputs(931) <= a;
    layer6_outputs(932) <= not (a xor b);
    layer6_outputs(933) <= b and not a;
    layer6_outputs(934) <= not (a xor b);
    layer6_outputs(935) <= a;
    layer6_outputs(936) <= b and not a;
    layer6_outputs(937) <= a;
    layer6_outputs(938) <= not b or a;
    layer6_outputs(939) <= not a;
    layer6_outputs(940) <= not (a and b);
    layer6_outputs(941) <= not a or b;
    layer6_outputs(942) <= a xor b;
    layer6_outputs(943) <= not (a xor b);
    layer6_outputs(944) <= a or b;
    layer6_outputs(945) <= not b;
    layer6_outputs(946) <= a and b;
    layer6_outputs(947) <= a or b;
    layer6_outputs(948) <= not b;
    layer6_outputs(949) <= not (a xor b);
    layer6_outputs(950) <= not a or b;
    layer6_outputs(951) <= b;
    layer6_outputs(952) <= b;
    layer6_outputs(953) <= not (a and b);
    layer6_outputs(954) <= not (a or b);
    layer6_outputs(955) <= a;
    layer6_outputs(956) <= a or b;
    layer6_outputs(957) <= not a;
    layer6_outputs(958) <= not (a and b);
    layer6_outputs(959) <= not b;
    layer6_outputs(960) <= a;
    layer6_outputs(961) <= not b or a;
    layer6_outputs(962) <= a;
    layer6_outputs(963) <= b;
    layer6_outputs(964) <= a xor b;
    layer6_outputs(965) <= a and b;
    layer6_outputs(966) <= not (a or b);
    layer6_outputs(967) <= not (a or b);
    layer6_outputs(968) <= not (a xor b);
    layer6_outputs(969) <= a and b;
    layer6_outputs(970) <= not a or b;
    layer6_outputs(971) <= not (a or b);
    layer6_outputs(972) <= not a;
    layer6_outputs(973) <= not a;
    layer6_outputs(974) <= not (a and b);
    layer6_outputs(975) <= b;
    layer6_outputs(976) <= not b;
    layer6_outputs(977) <= b and not a;
    layer6_outputs(978) <= b and not a;
    layer6_outputs(979) <= a xor b;
    layer6_outputs(980) <= not (a and b);
    layer6_outputs(981) <= a and b;
    layer6_outputs(982) <= a xor b;
    layer6_outputs(983) <= not b;
    layer6_outputs(984) <= b and not a;
    layer6_outputs(985) <= not b or a;
    layer6_outputs(986) <= not b;
    layer6_outputs(987) <= not b or a;
    layer6_outputs(988) <= not b;
    layer6_outputs(989) <= b and not a;
    layer6_outputs(990) <= not b;
    layer6_outputs(991) <= a;
    layer6_outputs(992) <= a and not b;
    layer6_outputs(993) <= a xor b;
    layer6_outputs(994) <= a and b;
    layer6_outputs(995) <= b and not a;
    layer6_outputs(996) <= b;
    layer6_outputs(997) <= not b;
    layer6_outputs(998) <= not b;
    layer6_outputs(999) <= not (a or b);
    layer6_outputs(1000) <= not (a xor b);
    layer6_outputs(1001) <= a or b;
    layer6_outputs(1002) <= not a;
    layer6_outputs(1003) <= not a;
    layer6_outputs(1004) <= not (a xor b);
    layer6_outputs(1005) <= a or b;
    layer6_outputs(1006) <= not b or a;
    layer6_outputs(1007) <= b;
    layer6_outputs(1008) <= not (a xor b);
    layer6_outputs(1009) <= a xor b;
    layer6_outputs(1010) <= a;
    layer6_outputs(1011) <= not a;
    layer6_outputs(1012) <= 1'b1;
    layer6_outputs(1013) <= b and not a;
    layer6_outputs(1014) <= a;
    layer6_outputs(1015) <= a;
    layer6_outputs(1016) <= a and b;
    layer6_outputs(1017) <= not b or a;
    layer6_outputs(1018) <= b;
    layer6_outputs(1019) <= not a;
    layer6_outputs(1020) <= a or b;
    layer6_outputs(1021) <= not b;
    layer6_outputs(1022) <= not (a and b);
    layer6_outputs(1023) <= not a;
    layer6_outputs(1024) <= not b or a;
    layer6_outputs(1025) <= b;
    layer6_outputs(1026) <= b;
    layer6_outputs(1027) <= a;
    layer6_outputs(1028) <= not a;
    layer6_outputs(1029) <= a and b;
    layer6_outputs(1030) <= a and not b;
    layer6_outputs(1031) <= a or b;
    layer6_outputs(1032) <= not (a xor b);
    layer6_outputs(1033) <= not (a or b);
    layer6_outputs(1034) <= a and b;
    layer6_outputs(1035) <= a;
    layer6_outputs(1036) <= a or b;
    layer6_outputs(1037) <= a and not b;
    layer6_outputs(1038) <= a;
    layer6_outputs(1039) <= not a;
    layer6_outputs(1040) <= not a;
    layer6_outputs(1041) <= a and not b;
    layer6_outputs(1042) <= a and b;
    layer6_outputs(1043) <= not (a xor b);
    layer6_outputs(1044) <= b and not a;
    layer6_outputs(1045) <= b;
    layer6_outputs(1046) <= not b;
    layer6_outputs(1047) <= b and not a;
    layer6_outputs(1048) <= a;
    layer6_outputs(1049) <= not a;
    layer6_outputs(1050) <= not b or a;
    layer6_outputs(1051) <= not b or a;
    layer6_outputs(1052) <= not a or b;
    layer6_outputs(1053) <= 1'b1;
    layer6_outputs(1054) <= not b or a;
    layer6_outputs(1055) <= a and b;
    layer6_outputs(1056) <= not a;
    layer6_outputs(1057) <= not (a and b);
    layer6_outputs(1058) <= not (a and b);
    layer6_outputs(1059) <= a xor b;
    layer6_outputs(1060) <= not a;
    layer6_outputs(1061) <= not a or b;
    layer6_outputs(1062) <= a or b;
    layer6_outputs(1063) <= a and b;
    layer6_outputs(1064) <= 1'b1;
    layer6_outputs(1065) <= b;
    layer6_outputs(1066) <= a xor b;
    layer6_outputs(1067) <= not a;
    layer6_outputs(1068) <= not a;
    layer6_outputs(1069) <= a or b;
    layer6_outputs(1070) <= b;
    layer6_outputs(1071) <= not (a and b);
    layer6_outputs(1072) <= b;
    layer6_outputs(1073) <= b;
    layer6_outputs(1074) <= not (a xor b);
    layer6_outputs(1075) <= not b;
    layer6_outputs(1076) <= not b;
    layer6_outputs(1077) <= 1'b1;
    layer6_outputs(1078) <= a xor b;
    layer6_outputs(1079) <= not a;
    layer6_outputs(1080) <= b and not a;
    layer6_outputs(1081) <= not a;
    layer6_outputs(1082) <= a;
    layer6_outputs(1083) <= not b;
    layer6_outputs(1084) <= a or b;
    layer6_outputs(1085) <= not a or b;
    layer6_outputs(1086) <= not b;
    layer6_outputs(1087) <= not a;
    layer6_outputs(1088) <= not a or b;
    layer6_outputs(1089) <= not b;
    layer6_outputs(1090) <= a or b;
    layer6_outputs(1091) <= a;
    layer6_outputs(1092) <= a and b;
    layer6_outputs(1093) <= not b;
    layer6_outputs(1094) <= not a;
    layer6_outputs(1095) <= not b;
    layer6_outputs(1096) <= b;
    layer6_outputs(1097) <= b;
    layer6_outputs(1098) <= not b;
    layer6_outputs(1099) <= not b;
    layer6_outputs(1100) <= a;
    layer6_outputs(1101) <= 1'b1;
    layer6_outputs(1102) <= a xor b;
    layer6_outputs(1103) <= not b;
    layer6_outputs(1104) <= b and not a;
    layer6_outputs(1105) <= a and not b;
    layer6_outputs(1106) <= not (a and b);
    layer6_outputs(1107) <= a and not b;
    layer6_outputs(1108) <= 1'b1;
    layer6_outputs(1109) <= not a;
    layer6_outputs(1110) <= not a;
    layer6_outputs(1111) <= not b or a;
    layer6_outputs(1112) <= b;
    layer6_outputs(1113) <= not (a or b);
    layer6_outputs(1114) <= not b;
    layer6_outputs(1115) <= b;
    layer6_outputs(1116) <= not (a or b);
    layer6_outputs(1117) <= a;
    layer6_outputs(1118) <= a xor b;
    layer6_outputs(1119) <= a;
    layer6_outputs(1120) <= not (a or b);
    layer6_outputs(1121) <= not a;
    layer6_outputs(1122) <= not a;
    layer6_outputs(1123) <= not a or b;
    layer6_outputs(1124) <= not b;
    layer6_outputs(1125) <= not (a xor b);
    layer6_outputs(1126) <= a;
    layer6_outputs(1127) <= not b;
    layer6_outputs(1128) <= b;
    layer6_outputs(1129) <= not a;
    layer6_outputs(1130) <= a;
    layer6_outputs(1131) <= not a;
    layer6_outputs(1132) <= a;
    layer6_outputs(1133) <= a and b;
    layer6_outputs(1134) <= 1'b1;
    layer6_outputs(1135) <= not b or a;
    layer6_outputs(1136) <= not b;
    layer6_outputs(1137) <= not a or b;
    layer6_outputs(1138) <= not (a or b);
    layer6_outputs(1139) <= not a;
    layer6_outputs(1140) <= not (a or b);
    layer6_outputs(1141) <= not a;
    layer6_outputs(1142) <= a and b;
    layer6_outputs(1143) <= b and not a;
    layer6_outputs(1144) <= not a;
    layer6_outputs(1145) <= not b;
    layer6_outputs(1146) <= b and not a;
    layer6_outputs(1147) <= not (a or b);
    layer6_outputs(1148) <= b;
    layer6_outputs(1149) <= b;
    layer6_outputs(1150) <= not b;
    layer6_outputs(1151) <= not (a or b);
    layer6_outputs(1152) <= not (a or b);
    layer6_outputs(1153) <= not a;
    layer6_outputs(1154) <= a;
    layer6_outputs(1155) <= a and not b;
    layer6_outputs(1156) <= not (a or b);
    layer6_outputs(1157) <= not a or b;
    layer6_outputs(1158) <= a or b;
    layer6_outputs(1159) <= not a;
    layer6_outputs(1160) <= b and not a;
    layer6_outputs(1161) <= not a or b;
    layer6_outputs(1162) <= not a;
    layer6_outputs(1163) <= a or b;
    layer6_outputs(1164) <= a xor b;
    layer6_outputs(1165) <= a or b;
    layer6_outputs(1166) <= a and b;
    layer6_outputs(1167) <= a and b;
    layer6_outputs(1168) <= a xor b;
    layer6_outputs(1169) <= a xor b;
    layer6_outputs(1170) <= not (a or b);
    layer6_outputs(1171) <= not (a and b);
    layer6_outputs(1172) <= not a;
    layer6_outputs(1173) <= not a;
    layer6_outputs(1174) <= a and b;
    layer6_outputs(1175) <= b and not a;
    layer6_outputs(1176) <= not a;
    layer6_outputs(1177) <= b;
    layer6_outputs(1178) <= 1'b0;
    layer6_outputs(1179) <= not b;
    layer6_outputs(1180) <= a xor b;
    layer6_outputs(1181) <= not b;
    layer6_outputs(1182) <= not a;
    layer6_outputs(1183) <= a xor b;
    layer6_outputs(1184) <= not (a or b);
    layer6_outputs(1185) <= not a;
    layer6_outputs(1186) <= not a;
    layer6_outputs(1187) <= not a;
    layer6_outputs(1188) <= a xor b;
    layer6_outputs(1189) <= b and not a;
    layer6_outputs(1190) <= not (a or b);
    layer6_outputs(1191) <= not b;
    layer6_outputs(1192) <= b;
    layer6_outputs(1193) <= b;
    layer6_outputs(1194) <= a or b;
    layer6_outputs(1195) <= b and not a;
    layer6_outputs(1196) <= not (a or b);
    layer6_outputs(1197) <= not b or a;
    layer6_outputs(1198) <= a or b;
    layer6_outputs(1199) <= b;
    layer6_outputs(1200) <= a or b;
    layer6_outputs(1201) <= a xor b;
    layer6_outputs(1202) <= a or b;
    layer6_outputs(1203) <= b;
    layer6_outputs(1204) <= not b;
    layer6_outputs(1205) <= b;
    layer6_outputs(1206) <= a;
    layer6_outputs(1207) <= not b;
    layer6_outputs(1208) <= not (a or b);
    layer6_outputs(1209) <= a;
    layer6_outputs(1210) <= a;
    layer6_outputs(1211) <= not a;
    layer6_outputs(1212) <= a and b;
    layer6_outputs(1213) <= b and not a;
    layer6_outputs(1214) <= 1'b0;
    layer6_outputs(1215) <= b;
    layer6_outputs(1216) <= not (a or b);
    layer6_outputs(1217) <= not (a or b);
    layer6_outputs(1218) <= not a or b;
    layer6_outputs(1219) <= a and not b;
    layer6_outputs(1220) <= not a;
    layer6_outputs(1221) <= a;
    layer6_outputs(1222) <= a and b;
    layer6_outputs(1223) <= not a;
    layer6_outputs(1224) <= b and not a;
    layer6_outputs(1225) <= a and b;
    layer6_outputs(1226) <= not (a and b);
    layer6_outputs(1227) <= b;
    layer6_outputs(1228) <= a or b;
    layer6_outputs(1229) <= not (a and b);
    layer6_outputs(1230) <= not a;
    layer6_outputs(1231) <= a;
    layer6_outputs(1232) <= a;
    layer6_outputs(1233) <= not b or a;
    layer6_outputs(1234) <= not a;
    layer6_outputs(1235) <= b;
    layer6_outputs(1236) <= a and b;
    layer6_outputs(1237) <= a or b;
    layer6_outputs(1238) <= not a;
    layer6_outputs(1239) <= a or b;
    layer6_outputs(1240) <= not b or a;
    layer6_outputs(1241) <= a and b;
    layer6_outputs(1242) <= not a or b;
    layer6_outputs(1243) <= not (a or b);
    layer6_outputs(1244) <= not a;
    layer6_outputs(1245) <= a and b;
    layer6_outputs(1246) <= not a;
    layer6_outputs(1247) <= not b;
    layer6_outputs(1248) <= not a or b;
    layer6_outputs(1249) <= a or b;
    layer6_outputs(1250) <= a and b;
    layer6_outputs(1251) <= not a;
    layer6_outputs(1252) <= b and not a;
    layer6_outputs(1253) <= not b;
    layer6_outputs(1254) <= not (a and b);
    layer6_outputs(1255) <= not a;
    layer6_outputs(1256) <= not (a or b);
    layer6_outputs(1257) <= a xor b;
    layer6_outputs(1258) <= not (a and b);
    layer6_outputs(1259) <= not b or a;
    layer6_outputs(1260) <= not a;
    layer6_outputs(1261) <= not b;
    layer6_outputs(1262) <= not (a xor b);
    layer6_outputs(1263) <= b;
    layer6_outputs(1264) <= a or b;
    layer6_outputs(1265) <= a;
    layer6_outputs(1266) <= b and not a;
    layer6_outputs(1267) <= not (a and b);
    layer6_outputs(1268) <= not b;
    layer6_outputs(1269) <= a and not b;
    layer6_outputs(1270) <= a;
    layer6_outputs(1271) <= not a;
    layer6_outputs(1272) <= a;
    layer6_outputs(1273) <= not a;
    layer6_outputs(1274) <= a xor b;
    layer6_outputs(1275) <= b;
    layer6_outputs(1276) <= not (a xor b);
    layer6_outputs(1277) <= not a;
    layer6_outputs(1278) <= a or b;
    layer6_outputs(1279) <= a xor b;
    layer6_outputs(1280) <= not b;
    layer6_outputs(1281) <= b;
    layer6_outputs(1282) <= a;
    layer6_outputs(1283) <= a;
    layer6_outputs(1284) <= b;
    layer6_outputs(1285) <= a;
    layer6_outputs(1286) <= b;
    layer6_outputs(1287) <= b and not a;
    layer6_outputs(1288) <= a;
    layer6_outputs(1289) <= not a;
    layer6_outputs(1290) <= not b;
    layer6_outputs(1291) <= not a or b;
    layer6_outputs(1292) <= a;
    layer6_outputs(1293) <= a and b;
    layer6_outputs(1294) <= 1'b1;
    layer6_outputs(1295) <= not b;
    layer6_outputs(1296) <= a;
    layer6_outputs(1297) <= a and b;
    layer6_outputs(1298) <= not b or a;
    layer6_outputs(1299) <= not b;
    layer6_outputs(1300) <= not a;
    layer6_outputs(1301) <= not (a or b);
    layer6_outputs(1302) <= not b or a;
    layer6_outputs(1303) <= not (a and b);
    layer6_outputs(1304) <= b and not a;
    layer6_outputs(1305) <= not b or a;
    layer6_outputs(1306) <= not b;
    layer6_outputs(1307) <= not a or b;
    layer6_outputs(1308) <= b;
    layer6_outputs(1309) <= a and not b;
    layer6_outputs(1310) <= a;
    layer6_outputs(1311) <= not a or b;
    layer6_outputs(1312) <= a xor b;
    layer6_outputs(1313) <= a and not b;
    layer6_outputs(1314) <= not b;
    layer6_outputs(1315) <= a;
    layer6_outputs(1316) <= not a or b;
    layer6_outputs(1317) <= not a;
    layer6_outputs(1318) <= not (a xor b);
    layer6_outputs(1319) <= not (a or b);
    layer6_outputs(1320) <= not a;
    layer6_outputs(1321) <= a and b;
    layer6_outputs(1322) <= not (a or b);
    layer6_outputs(1323) <= not (a and b);
    layer6_outputs(1324) <= not a or b;
    layer6_outputs(1325) <= not a or b;
    layer6_outputs(1326) <= not a;
    layer6_outputs(1327) <= not b;
    layer6_outputs(1328) <= not a or b;
    layer6_outputs(1329) <= b;
    layer6_outputs(1330) <= not b;
    layer6_outputs(1331) <= b and not a;
    layer6_outputs(1332) <= not a;
    layer6_outputs(1333) <= not a or b;
    layer6_outputs(1334) <= not a or b;
    layer6_outputs(1335) <= not b;
    layer6_outputs(1336) <= b and not a;
    layer6_outputs(1337) <= a and b;
    layer6_outputs(1338) <= a and not b;
    layer6_outputs(1339) <= not a or b;
    layer6_outputs(1340) <= a or b;
    layer6_outputs(1341) <= not b;
    layer6_outputs(1342) <= a and b;
    layer6_outputs(1343) <= a;
    layer6_outputs(1344) <= not (a or b);
    layer6_outputs(1345) <= not b;
    layer6_outputs(1346) <= a and b;
    layer6_outputs(1347) <= not a;
    layer6_outputs(1348) <= not b;
    layer6_outputs(1349) <= not (a or b);
    layer6_outputs(1350) <= 1'b1;
    layer6_outputs(1351) <= b and not a;
    layer6_outputs(1352) <= a and not b;
    layer6_outputs(1353) <= not a;
    layer6_outputs(1354) <= not a or b;
    layer6_outputs(1355) <= a xor b;
    layer6_outputs(1356) <= a and not b;
    layer6_outputs(1357) <= a;
    layer6_outputs(1358) <= not b;
    layer6_outputs(1359) <= not (a or b);
    layer6_outputs(1360) <= not b or a;
    layer6_outputs(1361) <= 1'b1;
    layer6_outputs(1362) <= a;
    layer6_outputs(1363) <= not b or a;
    layer6_outputs(1364) <= not b;
    layer6_outputs(1365) <= a and b;
    layer6_outputs(1366) <= b;
    layer6_outputs(1367) <= not a;
    layer6_outputs(1368) <= b;
    layer6_outputs(1369) <= not b;
    layer6_outputs(1370) <= not (a xor b);
    layer6_outputs(1371) <= b and not a;
    layer6_outputs(1372) <= not (a xor b);
    layer6_outputs(1373) <= a and not b;
    layer6_outputs(1374) <= not a or b;
    layer6_outputs(1375) <= not (a xor b);
    layer6_outputs(1376) <= not b;
    layer6_outputs(1377) <= a;
    layer6_outputs(1378) <= a and b;
    layer6_outputs(1379) <= not (a or b);
    layer6_outputs(1380) <= not b or a;
    layer6_outputs(1381) <= not a;
    layer6_outputs(1382) <= a xor b;
    layer6_outputs(1383) <= not (a xor b);
    layer6_outputs(1384) <= b;
    layer6_outputs(1385) <= a and not b;
    layer6_outputs(1386) <= not b or a;
    layer6_outputs(1387) <= a and not b;
    layer6_outputs(1388) <= not b;
    layer6_outputs(1389) <= a and not b;
    layer6_outputs(1390) <= not (a or b);
    layer6_outputs(1391) <= not (a xor b);
    layer6_outputs(1392) <= 1'b1;
    layer6_outputs(1393) <= not b or a;
    layer6_outputs(1394) <= 1'b1;
    layer6_outputs(1395) <= b;
    layer6_outputs(1396) <= b and not a;
    layer6_outputs(1397) <= a and b;
    layer6_outputs(1398) <= a and b;
    layer6_outputs(1399) <= b and not a;
    layer6_outputs(1400) <= b and not a;
    layer6_outputs(1401) <= a or b;
    layer6_outputs(1402) <= not a or b;
    layer6_outputs(1403) <= not a;
    layer6_outputs(1404) <= a and b;
    layer6_outputs(1405) <= not b;
    layer6_outputs(1406) <= 1'b0;
    layer6_outputs(1407) <= b and not a;
    layer6_outputs(1408) <= not (a or b);
    layer6_outputs(1409) <= not (a or b);
    layer6_outputs(1410) <= not (a xor b);
    layer6_outputs(1411) <= a;
    layer6_outputs(1412) <= not (a xor b);
    layer6_outputs(1413) <= 1'b0;
    layer6_outputs(1414) <= a;
    layer6_outputs(1415) <= not a or b;
    layer6_outputs(1416) <= a and not b;
    layer6_outputs(1417) <= not b;
    layer6_outputs(1418) <= not a;
    layer6_outputs(1419) <= not a;
    layer6_outputs(1420) <= not (a xor b);
    layer6_outputs(1421) <= not (a xor b);
    layer6_outputs(1422) <= a xor b;
    layer6_outputs(1423) <= not (a and b);
    layer6_outputs(1424) <= a xor b;
    layer6_outputs(1425) <= not a;
    layer6_outputs(1426) <= not a;
    layer6_outputs(1427) <= not (a xor b);
    layer6_outputs(1428) <= not a or b;
    layer6_outputs(1429) <= not (a or b);
    layer6_outputs(1430) <= not (a xor b);
    layer6_outputs(1431) <= not (a or b);
    layer6_outputs(1432) <= not a;
    layer6_outputs(1433) <= b;
    layer6_outputs(1434) <= a;
    layer6_outputs(1435) <= not b;
    layer6_outputs(1436) <= a or b;
    layer6_outputs(1437) <= a and b;
    layer6_outputs(1438) <= a or b;
    layer6_outputs(1439) <= a or b;
    layer6_outputs(1440) <= not a;
    layer6_outputs(1441) <= b;
    layer6_outputs(1442) <= a and not b;
    layer6_outputs(1443) <= not a;
    layer6_outputs(1444) <= a or b;
    layer6_outputs(1445) <= not b;
    layer6_outputs(1446) <= a or b;
    layer6_outputs(1447) <= a and not b;
    layer6_outputs(1448) <= a xor b;
    layer6_outputs(1449) <= a;
    layer6_outputs(1450) <= not a;
    layer6_outputs(1451) <= not (a or b);
    layer6_outputs(1452) <= not b or a;
    layer6_outputs(1453) <= not (a and b);
    layer6_outputs(1454) <= not (a or b);
    layer6_outputs(1455) <= b;
    layer6_outputs(1456) <= not b;
    layer6_outputs(1457) <= b and not a;
    layer6_outputs(1458) <= b;
    layer6_outputs(1459) <= not (a xor b);
    layer6_outputs(1460) <= not b or a;
    layer6_outputs(1461) <= not a;
    layer6_outputs(1462) <= not (a and b);
    layer6_outputs(1463) <= not a;
    layer6_outputs(1464) <= a xor b;
    layer6_outputs(1465) <= b and not a;
    layer6_outputs(1466) <= b;
    layer6_outputs(1467) <= a;
    layer6_outputs(1468) <= b;
    layer6_outputs(1469) <= not b;
    layer6_outputs(1470) <= a;
    layer6_outputs(1471) <= not (a and b);
    layer6_outputs(1472) <= a;
    layer6_outputs(1473) <= 1'b0;
    layer6_outputs(1474) <= not b;
    layer6_outputs(1475) <= a or b;
    layer6_outputs(1476) <= b;
    layer6_outputs(1477) <= not b or a;
    layer6_outputs(1478) <= b;
    layer6_outputs(1479) <= a or b;
    layer6_outputs(1480) <= a or b;
    layer6_outputs(1481) <= not b or a;
    layer6_outputs(1482) <= b and not a;
    layer6_outputs(1483) <= not (a or b);
    layer6_outputs(1484) <= a and not b;
    layer6_outputs(1485) <= not (a and b);
    layer6_outputs(1486) <= a and not b;
    layer6_outputs(1487) <= not a;
    layer6_outputs(1488) <= a and b;
    layer6_outputs(1489) <= b;
    layer6_outputs(1490) <= b;
    layer6_outputs(1491) <= not (a xor b);
    layer6_outputs(1492) <= 1'b1;
    layer6_outputs(1493) <= b;
    layer6_outputs(1494) <= a and not b;
    layer6_outputs(1495) <= not a;
    layer6_outputs(1496) <= a xor b;
    layer6_outputs(1497) <= a xor b;
    layer6_outputs(1498) <= a or b;
    layer6_outputs(1499) <= not b or a;
    layer6_outputs(1500) <= a or b;
    layer6_outputs(1501) <= a;
    layer6_outputs(1502) <= not b or a;
    layer6_outputs(1503) <= a;
    layer6_outputs(1504) <= not b;
    layer6_outputs(1505) <= not b;
    layer6_outputs(1506) <= not (a and b);
    layer6_outputs(1507) <= a or b;
    layer6_outputs(1508) <= b and not a;
    layer6_outputs(1509) <= not (a or b);
    layer6_outputs(1510) <= not b;
    layer6_outputs(1511) <= not (a or b);
    layer6_outputs(1512) <= not b;
    layer6_outputs(1513) <= 1'b0;
    layer6_outputs(1514) <= b and not a;
    layer6_outputs(1515) <= a and not b;
    layer6_outputs(1516) <= not (a xor b);
    layer6_outputs(1517) <= not b;
    layer6_outputs(1518) <= b;
    layer6_outputs(1519) <= not a or b;
    layer6_outputs(1520) <= b;
    layer6_outputs(1521) <= not (a or b);
    layer6_outputs(1522) <= not (a and b);
    layer6_outputs(1523) <= a xor b;
    layer6_outputs(1524) <= b;
    layer6_outputs(1525) <= b;
    layer6_outputs(1526) <= a or b;
    layer6_outputs(1527) <= b;
    layer6_outputs(1528) <= a or b;
    layer6_outputs(1529) <= b and not a;
    layer6_outputs(1530) <= not a;
    layer6_outputs(1531) <= not a;
    layer6_outputs(1532) <= not (a or b);
    layer6_outputs(1533) <= b and not a;
    layer6_outputs(1534) <= a or b;
    layer6_outputs(1535) <= not b;
    layer6_outputs(1536) <= a;
    layer6_outputs(1537) <= a or b;
    layer6_outputs(1538) <= a xor b;
    layer6_outputs(1539) <= a;
    layer6_outputs(1540) <= not b or a;
    layer6_outputs(1541) <= not b;
    layer6_outputs(1542) <= not a or b;
    layer6_outputs(1543) <= not (a and b);
    layer6_outputs(1544) <= b;
    layer6_outputs(1545) <= not b;
    layer6_outputs(1546) <= b;
    layer6_outputs(1547) <= not (a xor b);
    layer6_outputs(1548) <= not a or b;
    layer6_outputs(1549) <= not b or a;
    layer6_outputs(1550) <= a and b;
    layer6_outputs(1551) <= not (a or b);
    layer6_outputs(1552) <= not b;
    layer6_outputs(1553) <= not a or b;
    layer6_outputs(1554) <= not b;
    layer6_outputs(1555) <= not (a or b);
    layer6_outputs(1556) <= b;
    layer6_outputs(1557) <= b;
    layer6_outputs(1558) <= not b;
    layer6_outputs(1559) <= not a;
    layer6_outputs(1560) <= b;
    layer6_outputs(1561) <= a;
    layer6_outputs(1562) <= not (a xor b);
    layer6_outputs(1563) <= not (a xor b);
    layer6_outputs(1564) <= a;
    layer6_outputs(1565) <= not a or b;
    layer6_outputs(1566) <= not (a xor b);
    layer6_outputs(1567) <= not (a and b);
    layer6_outputs(1568) <= a or b;
    layer6_outputs(1569) <= not (a and b);
    layer6_outputs(1570) <= not a;
    layer6_outputs(1571) <= a and not b;
    layer6_outputs(1572) <= a or b;
    layer6_outputs(1573) <= not b or a;
    layer6_outputs(1574) <= not (a and b);
    layer6_outputs(1575) <= not b;
    layer6_outputs(1576) <= a xor b;
    layer6_outputs(1577) <= not a or b;
    layer6_outputs(1578) <= b and not a;
    layer6_outputs(1579) <= 1'b1;
    layer6_outputs(1580) <= not a;
    layer6_outputs(1581) <= not a;
    layer6_outputs(1582) <= a and not b;
    layer6_outputs(1583) <= a;
    layer6_outputs(1584) <= not a or b;
    layer6_outputs(1585) <= not (a or b);
    layer6_outputs(1586) <= 1'b1;
    layer6_outputs(1587) <= a;
    layer6_outputs(1588) <= not b;
    layer6_outputs(1589) <= not a;
    layer6_outputs(1590) <= not (a or b);
    layer6_outputs(1591) <= a;
    layer6_outputs(1592) <= not b or a;
    layer6_outputs(1593) <= not (a or b);
    layer6_outputs(1594) <= a;
    layer6_outputs(1595) <= not (a or b);
    layer6_outputs(1596) <= a or b;
    layer6_outputs(1597) <= not (a and b);
    layer6_outputs(1598) <= a and not b;
    layer6_outputs(1599) <= not b or a;
    layer6_outputs(1600) <= a;
    layer6_outputs(1601) <= not b;
    layer6_outputs(1602) <= a;
    layer6_outputs(1603) <= a;
    layer6_outputs(1604) <= not a;
    layer6_outputs(1605) <= a or b;
    layer6_outputs(1606) <= not b or a;
    layer6_outputs(1607) <= a xor b;
    layer6_outputs(1608) <= a and not b;
    layer6_outputs(1609) <= a or b;
    layer6_outputs(1610) <= a;
    layer6_outputs(1611) <= a and b;
    layer6_outputs(1612) <= not a;
    layer6_outputs(1613) <= not b;
    layer6_outputs(1614) <= not (a xor b);
    layer6_outputs(1615) <= b and not a;
    layer6_outputs(1616) <= not b;
    layer6_outputs(1617) <= a and not b;
    layer6_outputs(1618) <= not a;
    layer6_outputs(1619) <= not b;
    layer6_outputs(1620) <= b and not a;
    layer6_outputs(1621) <= not a;
    layer6_outputs(1622) <= 1'b0;
    layer6_outputs(1623) <= not (a or b);
    layer6_outputs(1624) <= not b;
    layer6_outputs(1625) <= not b;
    layer6_outputs(1626) <= a and not b;
    layer6_outputs(1627) <= not (a or b);
    layer6_outputs(1628) <= a;
    layer6_outputs(1629) <= 1'b1;
    layer6_outputs(1630) <= not (a and b);
    layer6_outputs(1631) <= 1'b1;
    layer6_outputs(1632) <= not a or b;
    layer6_outputs(1633) <= not (a xor b);
    layer6_outputs(1634) <= b;
    layer6_outputs(1635) <= not a;
    layer6_outputs(1636) <= a;
    layer6_outputs(1637) <= not a;
    layer6_outputs(1638) <= not b;
    layer6_outputs(1639) <= a xor b;
    layer6_outputs(1640) <= not (a xor b);
    layer6_outputs(1641) <= not (a and b);
    layer6_outputs(1642) <= not a or b;
    layer6_outputs(1643) <= not a or b;
    layer6_outputs(1644) <= a xor b;
    layer6_outputs(1645) <= not (a or b);
    layer6_outputs(1646) <= not (a xor b);
    layer6_outputs(1647) <= not a or b;
    layer6_outputs(1648) <= not b;
    layer6_outputs(1649) <= not b or a;
    layer6_outputs(1650) <= not a;
    layer6_outputs(1651) <= not a;
    layer6_outputs(1652) <= not a;
    layer6_outputs(1653) <= not b or a;
    layer6_outputs(1654) <= b and not a;
    layer6_outputs(1655) <= a or b;
    layer6_outputs(1656) <= not (a and b);
    layer6_outputs(1657) <= b and not a;
    layer6_outputs(1658) <= not a or b;
    layer6_outputs(1659) <= not b;
    layer6_outputs(1660) <= 1'b0;
    layer6_outputs(1661) <= not (a and b);
    layer6_outputs(1662) <= a xor b;
    layer6_outputs(1663) <= not b or a;
    layer6_outputs(1664) <= a xor b;
    layer6_outputs(1665) <= not (a or b);
    layer6_outputs(1666) <= a xor b;
    layer6_outputs(1667) <= not a or b;
    layer6_outputs(1668) <= not (a and b);
    layer6_outputs(1669) <= not a or b;
    layer6_outputs(1670) <= not a;
    layer6_outputs(1671) <= b;
    layer6_outputs(1672) <= a;
    layer6_outputs(1673) <= not b;
    layer6_outputs(1674) <= not b;
    layer6_outputs(1675) <= not (a xor b);
    layer6_outputs(1676) <= a;
    layer6_outputs(1677) <= not a;
    layer6_outputs(1678) <= a;
    layer6_outputs(1679) <= a and b;
    layer6_outputs(1680) <= not a;
    layer6_outputs(1681) <= not a;
    layer6_outputs(1682) <= not (a or b);
    layer6_outputs(1683) <= not b or a;
    layer6_outputs(1684) <= not a or b;
    layer6_outputs(1685) <= b and not a;
    layer6_outputs(1686) <= a;
    layer6_outputs(1687) <= b;
    layer6_outputs(1688) <= a and not b;
    layer6_outputs(1689) <= a;
    layer6_outputs(1690) <= not b;
    layer6_outputs(1691) <= b and not a;
    layer6_outputs(1692) <= a and b;
    layer6_outputs(1693) <= not (a and b);
    layer6_outputs(1694) <= not (a and b);
    layer6_outputs(1695) <= a and not b;
    layer6_outputs(1696) <= a or b;
    layer6_outputs(1697) <= a and b;
    layer6_outputs(1698) <= not (a and b);
    layer6_outputs(1699) <= not b or a;
    layer6_outputs(1700) <= not b or a;
    layer6_outputs(1701) <= not a;
    layer6_outputs(1702) <= a;
    layer6_outputs(1703) <= a and not b;
    layer6_outputs(1704) <= b;
    layer6_outputs(1705) <= a;
    layer6_outputs(1706) <= b and not a;
    layer6_outputs(1707) <= not (a or b);
    layer6_outputs(1708) <= a;
    layer6_outputs(1709) <= a xor b;
    layer6_outputs(1710) <= not a or b;
    layer6_outputs(1711) <= a or b;
    layer6_outputs(1712) <= a xor b;
    layer6_outputs(1713) <= 1'b0;
    layer6_outputs(1714) <= b;
    layer6_outputs(1715) <= not a;
    layer6_outputs(1716) <= not (a or b);
    layer6_outputs(1717) <= not (a and b);
    layer6_outputs(1718) <= not b;
    layer6_outputs(1719) <= b and not a;
    layer6_outputs(1720) <= a or b;
    layer6_outputs(1721) <= b;
    layer6_outputs(1722) <= not a;
    layer6_outputs(1723) <= not b or a;
    layer6_outputs(1724) <= not (a xor b);
    layer6_outputs(1725) <= a xor b;
    layer6_outputs(1726) <= b;
    layer6_outputs(1727) <= not a;
    layer6_outputs(1728) <= a and b;
    layer6_outputs(1729) <= a or b;
    layer6_outputs(1730) <= b and not a;
    layer6_outputs(1731) <= b;
    layer6_outputs(1732) <= b and not a;
    layer6_outputs(1733) <= not b;
    layer6_outputs(1734) <= b and not a;
    layer6_outputs(1735) <= 1'b0;
    layer6_outputs(1736) <= not b or a;
    layer6_outputs(1737) <= not b or a;
    layer6_outputs(1738) <= a and b;
    layer6_outputs(1739) <= not (a and b);
    layer6_outputs(1740) <= not a or b;
    layer6_outputs(1741) <= not b;
    layer6_outputs(1742) <= not b;
    layer6_outputs(1743) <= b;
    layer6_outputs(1744) <= a;
    layer6_outputs(1745) <= not a;
    layer6_outputs(1746) <= b;
    layer6_outputs(1747) <= not b or a;
    layer6_outputs(1748) <= not a;
    layer6_outputs(1749) <= not (a and b);
    layer6_outputs(1750) <= not a;
    layer6_outputs(1751) <= not (a or b);
    layer6_outputs(1752) <= not b or a;
    layer6_outputs(1753) <= not (a and b);
    layer6_outputs(1754) <= 1'b1;
    layer6_outputs(1755) <= not (a or b);
    layer6_outputs(1756) <= a or b;
    layer6_outputs(1757) <= b;
    layer6_outputs(1758) <= b;
    layer6_outputs(1759) <= not b;
    layer6_outputs(1760) <= a or b;
    layer6_outputs(1761) <= a and b;
    layer6_outputs(1762) <= not b or a;
    layer6_outputs(1763) <= a and not b;
    layer6_outputs(1764) <= not a;
    layer6_outputs(1765) <= not a;
    layer6_outputs(1766) <= a xor b;
    layer6_outputs(1767) <= a or b;
    layer6_outputs(1768) <= a and not b;
    layer6_outputs(1769) <= a and not b;
    layer6_outputs(1770) <= not a;
    layer6_outputs(1771) <= a and b;
    layer6_outputs(1772) <= a;
    layer6_outputs(1773) <= not a;
    layer6_outputs(1774) <= a;
    layer6_outputs(1775) <= not a or b;
    layer6_outputs(1776) <= not a;
    layer6_outputs(1777) <= b;
    layer6_outputs(1778) <= b;
    layer6_outputs(1779) <= b;
    layer6_outputs(1780) <= not a;
    layer6_outputs(1781) <= b and not a;
    layer6_outputs(1782) <= a;
    layer6_outputs(1783) <= not b or a;
    layer6_outputs(1784) <= not b;
    layer6_outputs(1785) <= a;
    layer6_outputs(1786) <= not a or b;
    layer6_outputs(1787) <= not b;
    layer6_outputs(1788) <= b;
    layer6_outputs(1789) <= a and b;
    layer6_outputs(1790) <= not a or b;
    layer6_outputs(1791) <= a and not b;
    layer6_outputs(1792) <= not a or b;
    layer6_outputs(1793) <= not b;
    layer6_outputs(1794) <= b;
    layer6_outputs(1795) <= a xor b;
    layer6_outputs(1796) <= a and b;
    layer6_outputs(1797) <= a;
    layer6_outputs(1798) <= a;
    layer6_outputs(1799) <= not (a and b);
    layer6_outputs(1800) <= 1'b1;
    layer6_outputs(1801) <= 1'b0;
    layer6_outputs(1802) <= b;
    layer6_outputs(1803) <= 1'b0;
    layer6_outputs(1804) <= a;
    layer6_outputs(1805) <= not b;
    layer6_outputs(1806) <= not b;
    layer6_outputs(1807) <= not (a and b);
    layer6_outputs(1808) <= not (a xor b);
    layer6_outputs(1809) <= b and not a;
    layer6_outputs(1810) <= not a;
    layer6_outputs(1811) <= a;
    layer6_outputs(1812) <= a;
    layer6_outputs(1813) <= not (a or b);
    layer6_outputs(1814) <= a;
    layer6_outputs(1815) <= b and not a;
    layer6_outputs(1816) <= a and b;
    layer6_outputs(1817) <= not (a and b);
    layer6_outputs(1818) <= not b or a;
    layer6_outputs(1819) <= not b or a;
    layer6_outputs(1820) <= b;
    layer6_outputs(1821) <= not (a xor b);
    layer6_outputs(1822) <= not a or b;
    layer6_outputs(1823) <= not b;
    layer6_outputs(1824) <= 1'b1;
    layer6_outputs(1825) <= not a;
    layer6_outputs(1826) <= a and b;
    layer6_outputs(1827) <= not b or a;
    layer6_outputs(1828) <= not (a or b);
    layer6_outputs(1829) <= not (a or b);
    layer6_outputs(1830) <= not b;
    layer6_outputs(1831) <= not b;
    layer6_outputs(1832) <= not (a and b);
    layer6_outputs(1833) <= not b;
    layer6_outputs(1834) <= 1'b0;
    layer6_outputs(1835) <= a;
    layer6_outputs(1836) <= not a;
    layer6_outputs(1837) <= a and not b;
    layer6_outputs(1838) <= a;
    layer6_outputs(1839) <= not a or b;
    layer6_outputs(1840) <= not a;
    layer6_outputs(1841) <= b and not a;
    layer6_outputs(1842) <= a;
    layer6_outputs(1843) <= not b;
    layer6_outputs(1844) <= not (a xor b);
    layer6_outputs(1845) <= a xor b;
    layer6_outputs(1846) <= 1'b1;
    layer6_outputs(1847) <= not (a xor b);
    layer6_outputs(1848) <= not b or a;
    layer6_outputs(1849) <= b and not a;
    layer6_outputs(1850) <= not a;
    layer6_outputs(1851) <= a xor b;
    layer6_outputs(1852) <= a;
    layer6_outputs(1853) <= not (a xor b);
    layer6_outputs(1854) <= b and not a;
    layer6_outputs(1855) <= b;
    layer6_outputs(1856) <= not b;
    layer6_outputs(1857) <= 1'b0;
    layer6_outputs(1858) <= a;
    layer6_outputs(1859) <= a;
    layer6_outputs(1860) <= not b;
    layer6_outputs(1861) <= b and not a;
    layer6_outputs(1862) <= a and b;
    layer6_outputs(1863) <= b and not a;
    layer6_outputs(1864) <= not b or a;
    layer6_outputs(1865) <= b;
    layer6_outputs(1866) <= not b or a;
    layer6_outputs(1867) <= not (a or b);
    layer6_outputs(1868) <= not b;
    layer6_outputs(1869) <= not a or b;
    layer6_outputs(1870) <= a xor b;
    layer6_outputs(1871) <= a and not b;
    layer6_outputs(1872) <= not a;
    layer6_outputs(1873) <= not a;
    layer6_outputs(1874) <= a;
    layer6_outputs(1875) <= b;
    layer6_outputs(1876) <= a or b;
    layer6_outputs(1877) <= 1'b0;
    layer6_outputs(1878) <= not (a or b);
    layer6_outputs(1879) <= not (a or b);
    layer6_outputs(1880) <= 1'b0;
    layer6_outputs(1881) <= not (a xor b);
    layer6_outputs(1882) <= b;
    layer6_outputs(1883) <= 1'b0;
    layer6_outputs(1884) <= not b or a;
    layer6_outputs(1885) <= a;
    layer6_outputs(1886) <= not a or b;
    layer6_outputs(1887) <= a and not b;
    layer6_outputs(1888) <= b;
    layer6_outputs(1889) <= not b;
    layer6_outputs(1890) <= not b;
    layer6_outputs(1891) <= not a;
    layer6_outputs(1892) <= not (a xor b);
    layer6_outputs(1893) <= a and not b;
    layer6_outputs(1894) <= a and b;
    layer6_outputs(1895) <= not b;
    layer6_outputs(1896) <= not b or a;
    layer6_outputs(1897) <= a;
    layer6_outputs(1898) <= 1'b1;
    layer6_outputs(1899) <= a;
    layer6_outputs(1900) <= a xor b;
    layer6_outputs(1901) <= not a;
    layer6_outputs(1902) <= a;
    layer6_outputs(1903) <= 1'b0;
    layer6_outputs(1904) <= b;
    layer6_outputs(1905) <= a or b;
    layer6_outputs(1906) <= not (a or b);
    layer6_outputs(1907) <= not a;
    layer6_outputs(1908) <= a;
    layer6_outputs(1909) <= a xor b;
    layer6_outputs(1910) <= not (a or b);
    layer6_outputs(1911) <= a or b;
    layer6_outputs(1912) <= a;
    layer6_outputs(1913) <= not b;
    layer6_outputs(1914) <= not b;
    layer6_outputs(1915) <= not b;
    layer6_outputs(1916) <= not (a or b);
    layer6_outputs(1917) <= not a;
    layer6_outputs(1918) <= not (a or b);
    layer6_outputs(1919) <= a xor b;
    layer6_outputs(1920) <= not a;
    layer6_outputs(1921) <= a;
    layer6_outputs(1922) <= not (a xor b);
    layer6_outputs(1923) <= 1'b1;
    layer6_outputs(1924) <= a;
    layer6_outputs(1925) <= a;
    layer6_outputs(1926) <= b and not a;
    layer6_outputs(1927) <= not b;
    layer6_outputs(1928) <= a or b;
    layer6_outputs(1929) <= a xor b;
    layer6_outputs(1930) <= a and b;
    layer6_outputs(1931) <= not (a xor b);
    layer6_outputs(1932) <= a;
    layer6_outputs(1933) <= not b or a;
    layer6_outputs(1934) <= b;
    layer6_outputs(1935) <= a;
    layer6_outputs(1936) <= not (a or b);
    layer6_outputs(1937) <= not a or b;
    layer6_outputs(1938) <= not a or b;
    layer6_outputs(1939) <= not b or a;
    layer6_outputs(1940) <= not b;
    layer6_outputs(1941) <= a;
    layer6_outputs(1942) <= not b;
    layer6_outputs(1943) <= a and not b;
    layer6_outputs(1944) <= not b;
    layer6_outputs(1945) <= a;
    layer6_outputs(1946) <= not b or a;
    layer6_outputs(1947) <= a and not b;
    layer6_outputs(1948) <= not b or a;
    layer6_outputs(1949) <= not a;
    layer6_outputs(1950) <= not b or a;
    layer6_outputs(1951) <= 1'b0;
    layer6_outputs(1952) <= not b;
    layer6_outputs(1953) <= 1'b0;
    layer6_outputs(1954) <= a xor b;
    layer6_outputs(1955) <= not b;
    layer6_outputs(1956) <= not a;
    layer6_outputs(1957) <= not b;
    layer6_outputs(1958) <= b;
    layer6_outputs(1959) <= a;
    layer6_outputs(1960) <= not (a and b);
    layer6_outputs(1961) <= b;
    layer6_outputs(1962) <= not b;
    layer6_outputs(1963) <= a;
    layer6_outputs(1964) <= not a;
    layer6_outputs(1965) <= not b;
    layer6_outputs(1966) <= a and b;
    layer6_outputs(1967) <= not (a xor b);
    layer6_outputs(1968) <= a and b;
    layer6_outputs(1969) <= a;
    layer6_outputs(1970) <= not (a and b);
    layer6_outputs(1971) <= not (a and b);
    layer6_outputs(1972) <= a and not b;
    layer6_outputs(1973) <= a;
    layer6_outputs(1974) <= a and not b;
    layer6_outputs(1975) <= a or b;
    layer6_outputs(1976) <= not (a and b);
    layer6_outputs(1977) <= a or b;
    layer6_outputs(1978) <= not b;
    layer6_outputs(1979) <= not (a xor b);
    layer6_outputs(1980) <= not (a or b);
    layer6_outputs(1981) <= a;
    layer6_outputs(1982) <= a;
    layer6_outputs(1983) <= a;
    layer6_outputs(1984) <= a and not b;
    layer6_outputs(1985) <= not b or a;
    layer6_outputs(1986) <= a xor b;
    layer6_outputs(1987) <= b;
    layer6_outputs(1988) <= not b;
    layer6_outputs(1989) <= not b;
    layer6_outputs(1990) <= not a;
    layer6_outputs(1991) <= not a;
    layer6_outputs(1992) <= a or b;
    layer6_outputs(1993) <= not (a or b);
    layer6_outputs(1994) <= not b;
    layer6_outputs(1995) <= not (a or b);
    layer6_outputs(1996) <= not b;
    layer6_outputs(1997) <= b;
    layer6_outputs(1998) <= not a;
    layer6_outputs(1999) <= a;
    layer6_outputs(2000) <= b;
    layer6_outputs(2001) <= b and not a;
    layer6_outputs(2002) <= a;
    layer6_outputs(2003) <= not a;
    layer6_outputs(2004) <= a or b;
    layer6_outputs(2005) <= b;
    layer6_outputs(2006) <= not b;
    layer6_outputs(2007) <= not b;
    layer6_outputs(2008) <= b;
    layer6_outputs(2009) <= not b or a;
    layer6_outputs(2010) <= a and not b;
    layer6_outputs(2011) <= b;
    layer6_outputs(2012) <= a xor b;
    layer6_outputs(2013) <= a and not b;
    layer6_outputs(2014) <= not a;
    layer6_outputs(2015) <= 1'b0;
    layer6_outputs(2016) <= 1'b0;
    layer6_outputs(2017) <= not a;
    layer6_outputs(2018) <= a xor b;
    layer6_outputs(2019) <= a;
    layer6_outputs(2020) <= a or b;
    layer6_outputs(2021) <= not (a xor b);
    layer6_outputs(2022) <= not (a xor b);
    layer6_outputs(2023) <= a;
    layer6_outputs(2024) <= b and not a;
    layer6_outputs(2025) <= b;
    layer6_outputs(2026) <= 1'b1;
    layer6_outputs(2027) <= 1'b0;
    layer6_outputs(2028) <= not b;
    layer6_outputs(2029) <= not b or a;
    layer6_outputs(2030) <= not b or a;
    layer6_outputs(2031) <= not a;
    layer6_outputs(2032) <= b;
    layer6_outputs(2033) <= b;
    layer6_outputs(2034) <= not a or b;
    layer6_outputs(2035) <= b and not a;
    layer6_outputs(2036) <= 1'b1;
    layer6_outputs(2037) <= a;
    layer6_outputs(2038) <= b;
    layer6_outputs(2039) <= not b or a;
    layer6_outputs(2040) <= b and not a;
    layer6_outputs(2041) <= a and not b;
    layer6_outputs(2042) <= 1'b0;
    layer6_outputs(2043) <= not (a or b);
    layer6_outputs(2044) <= b and not a;
    layer6_outputs(2045) <= not a or b;
    layer6_outputs(2046) <= a and not b;
    layer6_outputs(2047) <= not (a xor b);
    layer6_outputs(2048) <= 1'b0;
    layer6_outputs(2049) <= a xor b;
    layer6_outputs(2050) <= a xor b;
    layer6_outputs(2051) <= a and not b;
    layer6_outputs(2052) <= b and not a;
    layer6_outputs(2053) <= a and not b;
    layer6_outputs(2054) <= not (a or b);
    layer6_outputs(2055) <= not (a xor b);
    layer6_outputs(2056) <= b and not a;
    layer6_outputs(2057) <= a and not b;
    layer6_outputs(2058) <= not b or a;
    layer6_outputs(2059) <= b and not a;
    layer6_outputs(2060) <= b;
    layer6_outputs(2061) <= not a;
    layer6_outputs(2062) <= a;
    layer6_outputs(2063) <= a xor b;
    layer6_outputs(2064) <= not b;
    layer6_outputs(2065) <= a and b;
    layer6_outputs(2066) <= a;
    layer6_outputs(2067) <= b and not a;
    layer6_outputs(2068) <= b;
    layer6_outputs(2069) <= a xor b;
    layer6_outputs(2070) <= b and not a;
    layer6_outputs(2071) <= not (a and b);
    layer6_outputs(2072) <= a and b;
    layer6_outputs(2073) <= a;
    layer6_outputs(2074) <= not b;
    layer6_outputs(2075) <= not b;
    layer6_outputs(2076) <= not b;
    layer6_outputs(2077) <= not a;
    layer6_outputs(2078) <= not b;
    layer6_outputs(2079) <= not (a xor b);
    layer6_outputs(2080) <= a or b;
    layer6_outputs(2081) <= not b;
    layer6_outputs(2082) <= not (a and b);
    layer6_outputs(2083) <= b and not a;
    layer6_outputs(2084) <= b;
    layer6_outputs(2085) <= not b or a;
    layer6_outputs(2086) <= not a;
    layer6_outputs(2087) <= not b;
    layer6_outputs(2088) <= a xor b;
    layer6_outputs(2089) <= not (a and b);
    layer6_outputs(2090) <= b;
    layer6_outputs(2091) <= not b;
    layer6_outputs(2092) <= not a or b;
    layer6_outputs(2093) <= a and b;
    layer6_outputs(2094) <= a and not b;
    layer6_outputs(2095) <= not (a and b);
    layer6_outputs(2096) <= not a;
    layer6_outputs(2097) <= b and not a;
    layer6_outputs(2098) <= not a;
    layer6_outputs(2099) <= not b;
    layer6_outputs(2100) <= a;
    layer6_outputs(2101) <= not b;
    layer6_outputs(2102) <= not a;
    layer6_outputs(2103) <= 1'b1;
    layer6_outputs(2104) <= b and not a;
    layer6_outputs(2105) <= a xor b;
    layer6_outputs(2106) <= a;
    layer6_outputs(2107) <= not a;
    layer6_outputs(2108) <= a;
    layer6_outputs(2109) <= not a;
    layer6_outputs(2110) <= not (a and b);
    layer6_outputs(2111) <= a and not b;
    layer6_outputs(2112) <= not b;
    layer6_outputs(2113) <= not (a or b);
    layer6_outputs(2114) <= not a or b;
    layer6_outputs(2115) <= a and b;
    layer6_outputs(2116) <= not a or b;
    layer6_outputs(2117) <= not (a or b);
    layer6_outputs(2118) <= b;
    layer6_outputs(2119) <= b;
    layer6_outputs(2120) <= not (a or b);
    layer6_outputs(2121) <= a and b;
    layer6_outputs(2122) <= a or b;
    layer6_outputs(2123) <= a;
    layer6_outputs(2124) <= not (a and b);
    layer6_outputs(2125) <= a;
    layer6_outputs(2126) <= b and not a;
    layer6_outputs(2127) <= a;
    layer6_outputs(2128) <= 1'b0;
    layer6_outputs(2129) <= not a;
    layer6_outputs(2130) <= not a;
    layer6_outputs(2131) <= a and not b;
    layer6_outputs(2132) <= not (a xor b);
    layer6_outputs(2133) <= not (a or b);
    layer6_outputs(2134) <= a xor b;
    layer6_outputs(2135) <= not (a or b);
    layer6_outputs(2136) <= not a or b;
    layer6_outputs(2137) <= not a;
    layer6_outputs(2138) <= not b;
    layer6_outputs(2139) <= b;
    layer6_outputs(2140) <= not a or b;
    layer6_outputs(2141) <= 1'b0;
    layer6_outputs(2142) <= a or b;
    layer6_outputs(2143) <= a or b;
    layer6_outputs(2144) <= not b;
    layer6_outputs(2145) <= not a or b;
    layer6_outputs(2146) <= a or b;
    layer6_outputs(2147) <= b;
    layer6_outputs(2148) <= a;
    layer6_outputs(2149) <= not a;
    layer6_outputs(2150) <= b;
    layer6_outputs(2151) <= a and not b;
    layer6_outputs(2152) <= not a;
    layer6_outputs(2153) <= not a;
    layer6_outputs(2154) <= b;
    layer6_outputs(2155) <= not (a or b);
    layer6_outputs(2156) <= a;
    layer6_outputs(2157) <= b and not a;
    layer6_outputs(2158) <= b;
    layer6_outputs(2159) <= not b;
    layer6_outputs(2160) <= not a or b;
    layer6_outputs(2161) <= b;
    layer6_outputs(2162) <= not b;
    layer6_outputs(2163) <= a or b;
    layer6_outputs(2164) <= not a;
    layer6_outputs(2165) <= not b;
    layer6_outputs(2166) <= a;
    layer6_outputs(2167) <= a and b;
    layer6_outputs(2168) <= 1'b0;
    layer6_outputs(2169) <= a and b;
    layer6_outputs(2170) <= not (a or b);
    layer6_outputs(2171) <= a;
    layer6_outputs(2172) <= not a;
    layer6_outputs(2173) <= a;
    layer6_outputs(2174) <= b and not a;
    layer6_outputs(2175) <= a or b;
    layer6_outputs(2176) <= not b or a;
    layer6_outputs(2177) <= not a;
    layer6_outputs(2178) <= a xor b;
    layer6_outputs(2179) <= not a or b;
    layer6_outputs(2180) <= not b;
    layer6_outputs(2181) <= not (a xor b);
    layer6_outputs(2182) <= not b;
    layer6_outputs(2183) <= not (a and b);
    layer6_outputs(2184) <= b and not a;
    layer6_outputs(2185) <= a xor b;
    layer6_outputs(2186) <= 1'b0;
    layer6_outputs(2187) <= not a;
    layer6_outputs(2188) <= b;
    layer6_outputs(2189) <= not a;
    layer6_outputs(2190) <= b;
    layer6_outputs(2191) <= not b or a;
    layer6_outputs(2192) <= not (a and b);
    layer6_outputs(2193) <= b and not a;
    layer6_outputs(2194) <= not (a xor b);
    layer6_outputs(2195) <= not (a or b);
    layer6_outputs(2196) <= not (a or b);
    layer6_outputs(2197) <= a and b;
    layer6_outputs(2198) <= not b or a;
    layer6_outputs(2199) <= not a;
    layer6_outputs(2200) <= b;
    layer6_outputs(2201) <= a and not b;
    layer6_outputs(2202) <= b and not a;
    layer6_outputs(2203) <= b;
    layer6_outputs(2204) <= not a or b;
    layer6_outputs(2205) <= a xor b;
    layer6_outputs(2206) <= a;
    layer6_outputs(2207) <= a xor b;
    layer6_outputs(2208) <= not b or a;
    layer6_outputs(2209) <= not (a xor b);
    layer6_outputs(2210) <= not (a xor b);
    layer6_outputs(2211) <= a or b;
    layer6_outputs(2212) <= not a;
    layer6_outputs(2213) <= a xor b;
    layer6_outputs(2214) <= a xor b;
    layer6_outputs(2215) <= 1'b1;
    layer6_outputs(2216) <= b;
    layer6_outputs(2217) <= not b;
    layer6_outputs(2218) <= 1'b1;
    layer6_outputs(2219) <= not b or a;
    layer6_outputs(2220) <= a xor b;
    layer6_outputs(2221) <= not b or a;
    layer6_outputs(2222) <= a and b;
    layer6_outputs(2223) <= a and not b;
    layer6_outputs(2224) <= a;
    layer6_outputs(2225) <= not (a or b);
    layer6_outputs(2226) <= not a;
    layer6_outputs(2227) <= a;
    layer6_outputs(2228) <= a;
    layer6_outputs(2229) <= not (a and b);
    layer6_outputs(2230) <= 1'b1;
    layer6_outputs(2231) <= a;
    layer6_outputs(2232) <= a xor b;
    layer6_outputs(2233) <= not a;
    layer6_outputs(2234) <= a;
    layer6_outputs(2235) <= not b;
    layer6_outputs(2236) <= a;
    layer6_outputs(2237) <= a;
    layer6_outputs(2238) <= not a or b;
    layer6_outputs(2239) <= not b or a;
    layer6_outputs(2240) <= 1'b1;
    layer6_outputs(2241) <= b;
    layer6_outputs(2242) <= not b;
    layer6_outputs(2243) <= b;
    layer6_outputs(2244) <= not b;
    layer6_outputs(2245) <= not b;
    layer6_outputs(2246) <= not (a xor b);
    layer6_outputs(2247) <= not (a and b);
    layer6_outputs(2248) <= a or b;
    layer6_outputs(2249) <= b;
    layer6_outputs(2250) <= b;
    layer6_outputs(2251) <= not (a xor b);
    layer6_outputs(2252) <= a xor b;
    layer6_outputs(2253) <= a or b;
    layer6_outputs(2254) <= not (a and b);
    layer6_outputs(2255) <= not (a or b);
    layer6_outputs(2256) <= a and b;
    layer6_outputs(2257) <= a and b;
    layer6_outputs(2258) <= not a;
    layer6_outputs(2259) <= a;
    layer6_outputs(2260) <= not a or b;
    layer6_outputs(2261) <= not a or b;
    layer6_outputs(2262) <= not (a xor b);
    layer6_outputs(2263) <= not a or b;
    layer6_outputs(2264) <= a or b;
    layer6_outputs(2265) <= not (a xor b);
    layer6_outputs(2266) <= b;
    layer6_outputs(2267) <= not (a or b);
    layer6_outputs(2268) <= not (a and b);
    layer6_outputs(2269) <= not b or a;
    layer6_outputs(2270) <= a;
    layer6_outputs(2271) <= not b;
    layer6_outputs(2272) <= not b or a;
    layer6_outputs(2273) <= a;
    layer6_outputs(2274) <= not (a xor b);
    layer6_outputs(2275) <= not (a and b);
    layer6_outputs(2276) <= a and not b;
    layer6_outputs(2277) <= b and not a;
    layer6_outputs(2278) <= b;
    layer6_outputs(2279) <= a;
    layer6_outputs(2280) <= not a;
    layer6_outputs(2281) <= b and not a;
    layer6_outputs(2282) <= a and not b;
    layer6_outputs(2283) <= a or b;
    layer6_outputs(2284) <= a;
    layer6_outputs(2285) <= a and b;
    layer6_outputs(2286) <= not (a xor b);
    layer6_outputs(2287) <= a;
    layer6_outputs(2288) <= not a;
    layer6_outputs(2289) <= a or b;
    layer6_outputs(2290) <= not (a or b);
    layer6_outputs(2291) <= not b;
    layer6_outputs(2292) <= not a or b;
    layer6_outputs(2293) <= b;
    layer6_outputs(2294) <= a xor b;
    layer6_outputs(2295) <= not (a and b);
    layer6_outputs(2296) <= 1'b1;
    layer6_outputs(2297) <= a xor b;
    layer6_outputs(2298) <= not b;
    layer6_outputs(2299) <= not b;
    layer6_outputs(2300) <= not a;
    layer6_outputs(2301) <= not (a xor b);
    layer6_outputs(2302) <= not b or a;
    layer6_outputs(2303) <= a or b;
    layer6_outputs(2304) <= not b;
    layer6_outputs(2305) <= not a;
    layer6_outputs(2306) <= not a;
    layer6_outputs(2307) <= a;
    layer6_outputs(2308) <= a and not b;
    layer6_outputs(2309) <= b;
    layer6_outputs(2310) <= a xor b;
    layer6_outputs(2311) <= a and b;
    layer6_outputs(2312) <= not b;
    layer6_outputs(2313) <= a or b;
    layer6_outputs(2314) <= 1'b0;
    layer6_outputs(2315) <= b and not a;
    layer6_outputs(2316) <= not b;
    layer6_outputs(2317) <= a;
    layer6_outputs(2318) <= b;
    layer6_outputs(2319) <= a or b;
    layer6_outputs(2320) <= not a;
    layer6_outputs(2321) <= a and not b;
    layer6_outputs(2322) <= a;
    layer6_outputs(2323) <= a or b;
    layer6_outputs(2324) <= a or b;
    layer6_outputs(2325) <= 1'b0;
    layer6_outputs(2326) <= a;
    layer6_outputs(2327) <= a;
    layer6_outputs(2328) <= not a;
    layer6_outputs(2329) <= b and not a;
    layer6_outputs(2330) <= a or b;
    layer6_outputs(2331) <= a or b;
    layer6_outputs(2332) <= a xor b;
    layer6_outputs(2333) <= not b;
    layer6_outputs(2334) <= not a;
    layer6_outputs(2335) <= a or b;
    layer6_outputs(2336) <= not (a or b);
    layer6_outputs(2337) <= not (a and b);
    layer6_outputs(2338) <= a;
    layer6_outputs(2339) <= a or b;
    layer6_outputs(2340) <= a or b;
    layer6_outputs(2341) <= not a or b;
    layer6_outputs(2342) <= a xor b;
    layer6_outputs(2343) <= not a or b;
    layer6_outputs(2344) <= not a or b;
    layer6_outputs(2345) <= not b or a;
    layer6_outputs(2346) <= not b;
    layer6_outputs(2347) <= not b;
    layer6_outputs(2348) <= not b;
    layer6_outputs(2349) <= not b;
    layer6_outputs(2350) <= 1'b1;
    layer6_outputs(2351) <= not (a xor b);
    layer6_outputs(2352) <= a;
    layer6_outputs(2353) <= not b;
    layer6_outputs(2354) <= not a;
    layer6_outputs(2355) <= not a or b;
    layer6_outputs(2356) <= a;
    layer6_outputs(2357) <= b and not a;
    layer6_outputs(2358) <= not (a xor b);
    layer6_outputs(2359) <= a;
    layer6_outputs(2360) <= 1'b0;
    layer6_outputs(2361) <= a;
    layer6_outputs(2362) <= b;
    layer6_outputs(2363) <= not (a xor b);
    layer6_outputs(2364) <= not a or b;
    layer6_outputs(2365) <= a;
    layer6_outputs(2366) <= not a;
    layer6_outputs(2367) <= b;
    layer6_outputs(2368) <= 1'b0;
    layer6_outputs(2369) <= b and not a;
    layer6_outputs(2370) <= b;
    layer6_outputs(2371) <= not a;
    layer6_outputs(2372) <= not b or a;
    layer6_outputs(2373) <= a;
    layer6_outputs(2374) <= a;
    layer6_outputs(2375) <= not (a and b);
    layer6_outputs(2376) <= b;
    layer6_outputs(2377) <= not a;
    layer6_outputs(2378) <= not a;
    layer6_outputs(2379) <= a and b;
    layer6_outputs(2380) <= not b;
    layer6_outputs(2381) <= not b or a;
    layer6_outputs(2382) <= b;
    layer6_outputs(2383) <= not b;
    layer6_outputs(2384) <= b;
    layer6_outputs(2385) <= not a or b;
    layer6_outputs(2386) <= not a;
    layer6_outputs(2387) <= not a;
    layer6_outputs(2388) <= not a or b;
    layer6_outputs(2389) <= not b;
    layer6_outputs(2390) <= a;
    layer6_outputs(2391) <= b and not a;
    layer6_outputs(2392) <= not a or b;
    layer6_outputs(2393) <= b;
    layer6_outputs(2394) <= a;
    layer6_outputs(2395) <= 1'b0;
    layer6_outputs(2396) <= b;
    layer6_outputs(2397) <= not a;
    layer6_outputs(2398) <= not b;
    layer6_outputs(2399) <= b;
    layer6_outputs(2400) <= not b;
    layer6_outputs(2401) <= a;
    layer6_outputs(2402) <= a;
    layer6_outputs(2403) <= not b;
    layer6_outputs(2404) <= a xor b;
    layer6_outputs(2405) <= 1'b1;
    layer6_outputs(2406) <= not a or b;
    layer6_outputs(2407) <= 1'b1;
    layer6_outputs(2408) <= not b or a;
    layer6_outputs(2409) <= not (a and b);
    layer6_outputs(2410) <= b;
    layer6_outputs(2411) <= not b or a;
    layer6_outputs(2412) <= b;
    layer6_outputs(2413) <= not a or b;
    layer6_outputs(2414) <= not (a and b);
    layer6_outputs(2415) <= not (a xor b);
    layer6_outputs(2416) <= b;
    layer6_outputs(2417) <= not a;
    layer6_outputs(2418) <= a or b;
    layer6_outputs(2419) <= not b or a;
    layer6_outputs(2420) <= a;
    layer6_outputs(2421) <= not a;
    layer6_outputs(2422) <= not b or a;
    layer6_outputs(2423) <= not a;
    layer6_outputs(2424) <= not (a xor b);
    layer6_outputs(2425) <= a xor b;
    layer6_outputs(2426) <= not a or b;
    layer6_outputs(2427) <= a;
    layer6_outputs(2428) <= not b;
    layer6_outputs(2429) <= not b;
    layer6_outputs(2430) <= not a or b;
    layer6_outputs(2431) <= not a or b;
    layer6_outputs(2432) <= a;
    layer6_outputs(2433) <= a;
    layer6_outputs(2434) <= b;
    layer6_outputs(2435) <= not (a xor b);
    layer6_outputs(2436) <= a;
    layer6_outputs(2437) <= a and not b;
    layer6_outputs(2438) <= not (a and b);
    layer6_outputs(2439) <= a;
    layer6_outputs(2440) <= not (a or b);
    layer6_outputs(2441) <= a and not b;
    layer6_outputs(2442) <= a;
    layer6_outputs(2443) <= a and not b;
    layer6_outputs(2444) <= b and not a;
    layer6_outputs(2445) <= a xor b;
    layer6_outputs(2446) <= a;
    layer6_outputs(2447) <= not (a xor b);
    layer6_outputs(2448) <= b and not a;
    layer6_outputs(2449) <= a or b;
    layer6_outputs(2450) <= b;
    layer6_outputs(2451) <= not a or b;
    layer6_outputs(2452) <= not (a or b);
    layer6_outputs(2453) <= not (a and b);
    layer6_outputs(2454) <= not a or b;
    layer6_outputs(2455) <= not b;
    layer6_outputs(2456) <= not a;
    layer6_outputs(2457) <= b;
    layer6_outputs(2458) <= b;
    layer6_outputs(2459) <= a;
    layer6_outputs(2460) <= not (a xor b);
    layer6_outputs(2461) <= a;
    layer6_outputs(2462) <= a;
    layer6_outputs(2463) <= not a or b;
    layer6_outputs(2464) <= b;
    layer6_outputs(2465) <= b;
    layer6_outputs(2466) <= not (a or b);
    layer6_outputs(2467) <= b;
    layer6_outputs(2468) <= not (a xor b);
    layer6_outputs(2469) <= a xor b;
    layer6_outputs(2470) <= b;
    layer6_outputs(2471) <= not b;
    layer6_outputs(2472) <= a or b;
    layer6_outputs(2473) <= not (a and b);
    layer6_outputs(2474) <= not b;
    layer6_outputs(2475) <= not b;
    layer6_outputs(2476) <= a;
    layer6_outputs(2477) <= a and not b;
    layer6_outputs(2478) <= b and not a;
    layer6_outputs(2479) <= b and not a;
    layer6_outputs(2480) <= not a;
    layer6_outputs(2481) <= not a or b;
    layer6_outputs(2482) <= a and not b;
    layer6_outputs(2483) <= not (a and b);
    layer6_outputs(2484) <= b and not a;
    layer6_outputs(2485) <= b and not a;
    layer6_outputs(2486) <= a xor b;
    layer6_outputs(2487) <= not b;
    layer6_outputs(2488) <= not (a and b);
    layer6_outputs(2489) <= not a;
    layer6_outputs(2490) <= a and not b;
    layer6_outputs(2491) <= not b;
    layer6_outputs(2492) <= a xor b;
    layer6_outputs(2493) <= b;
    layer6_outputs(2494) <= a and b;
    layer6_outputs(2495) <= b and not a;
    layer6_outputs(2496) <= not (a xor b);
    layer6_outputs(2497) <= not (a and b);
    layer6_outputs(2498) <= not a;
    layer6_outputs(2499) <= a and not b;
    layer6_outputs(2500) <= b;
    layer6_outputs(2501) <= not b;
    layer6_outputs(2502) <= not a;
    layer6_outputs(2503) <= not a or b;
    layer6_outputs(2504) <= not (a xor b);
    layer6_outputs(2505) <= 1'b1;
    layer6_outputs(2506) <= a xor b;
    layer6_outputs(2507) <= a and b;
    layer6_outputs(2508) <= a xor b;
    layer6_outputs(2509) <= a xor b;
    layer6_outputs(2510) <= not a;
    layer6_outputs(2511) <= not a;
    layer6_outputs(2512) <= not b;
    layer6_outputs(2513) <= not b or a;
    layer6_outputs(2514) <= a xor b;
    layer6_outputs(2515) <= a or b;
    layer6_outputs(2516) <= b;
    layer6_outputs(2517) <= not b;
    layer6_outputs(2518) <= a or b;
    layer6_outputs(2519) <= not a;
    layer6_outputs(2520) <= a or b;
    layer6_outputs(2521) <= not a;
    layer6_outputs(2522) <= not a;
    layer6_outputs(2523) <= a and b;
    layer6_outputs(2524) <= not b;
    layer6_outputs(2525) <= not a or b;
    layer6_outputs(2526) <= a or b;
    layer6_outputs(2527) <= a xor b;
    layer6_outputs(2528) <= not (a xor b);
    layer6_outputs(2529) <= a;
    layer6_outputs(2530) <= not (a or b);
    layer6_outputs(2531) <= b and not a;
    layer6_outputs(2532) <= not (a and b);
    layer6_outputs(2533) <= a;
    layer6_outputs(2534) <= b and not a;
    layer6_outputs(2535) <= not b or a;
    layer6_outputs(2536) <= 1'b1;
    layer6_outputs(2537) <= not (a or b);
    layer6_outputs(2538) <= a;
    layer6_outputs(2539) <= a and not b;
    layer6_outputs(2540) <= not (a xor b);
    layer6_outputs(2541) <= b and not a;
    layer6_outputs(2542) <= not b;
    layer6_outputs(2543) <= not (a and b);
    layer6_outputs(2544) <= a xor b;
    layer6_outputs(2545) <= not b or a;
    layer6_outputs(2546) <= b;
    layer6_outputs(2547) <= not (a or b);
    layer6_outputs(2548) <= not b;
    layer6_outputs(2549) <= not a or b;
    layer6_outputs(2550) <= a;
    layer6_outputs(2551) <= a xor b;
    layer6_outputs(2552) <= not b;
    layer6_outputs(2553) <= a xor b;
    layer6_outputs(2554) <= not a or b;
    layer6_outputs(2555) <= not (a and b);
    layer6_outputs(2556) <= not (a or b);
    layer6_outputs(2557) <= not a;
    layer6_outputs(2558) <= a or b;
    layer6_outputs(2559) <= a;
    layer6_outputs(2560) <= not b;
    layer6_outputs(2561) <= not (a and b);
    layer6_outputs(2562) <= not b;
    layer6_outputs(2563) <= not a;
    layer6_outputs(2564) <= not a;
    layer6_outputs(2565) <= not a;
    layer6_outputs(2566) <= a;
    layer6_outputs(2567) <= a xor b;
    layer6_outputs(2568) <= a xor b;
    layer6_outputs(2569) <= not b;
    layer6_outputs(2570) <= not (a and b);
    layer6_outputs(2571) <= not b;
    layer6_outputs(2572) <= a;
    layer6_outputs(2573) <= a;
    layer6_outputs(2574) <= not b;
    layer6_outputs(2575) <= a;
    layer6_outputs(2576) <= not b;
    layer6_outputs(2577) <= a and b;
    layer6_outputs(2578) <= not b or a;
    layer6_outputs(2579) <= not a;
    layer6_outputs(2580) <= not (a xor b);
    layer6_outputs(2581) <= not (a xor b);
    layer6_outputs(2582) <= b;
    layer6_outputs(2583) <= a or b;
    layer6_outputs(2584) <= not (a xor b);
    layer6_outputs(2585) <= not (a or b);
    layer6_outputs(2586) <= a;
    layer6_outputs(2587) <= not a;
    layer6_outputs(2588) <= not (a and b);
    layer6_outputs(2589) <= not a;
    layer6_outputs(2590) <= not (a and b);
    layer6_outputs(2591) <= b and not a;
    layer6_outputs(2592) <= not a or b;
    layer6_outputs(2593) <= not (a and b);
    layer6_outputs(2594) <= not b;
    layer6_outputs(2595) <= not a;
    layer6_outputs(2596) <= not (a xor b);
    layer6_outputs(2597) <= a xor b;
    layer6_outputs(2598) <= b;
    layer6_outputs(2599) <= not (a and b);
    layer6_outputs(2600) <= not (a and b);
    layer6_outputs(2601) <= not a or b;
    layer6_outputs(2602) <= not b;
    layer6_outputs(2603) <= a and b;
    layer6_outputs(2604) <= a and b;
    layer6_outputs(2605) <= not (a or b);
    layer6_outputs(2606) <= not a;
    layer6_outputs(2607) <= not b or a;
    layer6_outputs(2608) <= a;
    layer6_outputs(2609) <= not (a and b);
    layer6_outputs(2610) <= a;
    layer6_outputs(2611) <= a and not b;
    layer6_outputs(2612) <= a;
    layer6_outputs(2613) <= not b;
    layer6_outputs(2614) <= a;
    layer6_outputs(2615) <= not b;
    layer6_outputs(2616) <= a and b;
    layer6_outputs(2617) <= a xor b;
    layer6_outputs(2618) <= not a;
    layer6_outputs(2619) <= not (a or b);
    layer6_outputs(2620) <= a and not b;
    layer6_outputs(2621) <= a and b;
    layer6_outputs(2622) <= a and b;
    layer6_outputs(2623) <= a or b;
    layer6_outputs(2624) <= not b or a;
    layer6_outputs(2625) <= not a;
    layer6_outputs(2626) <= 1'b0;
    layer6_outputs(2627) <= b;
    layer6_outputs(2628) <= a and b;
    layer6_outputs(2629) <= a;
    layer6_outputs(2630) <= b;
    layer6_outputs(2631) <= not b;
    layer6_outputs(2632) <= not b or a;
    layer6_outputs(2633) <= not a;
    layer6_outputs(2634) <= b;
    layer6_outputs(2635) <= b and not a;
    layer6_outputs(2636) <= a xor b;
    layer6_outputs(2637) <= a and b;
    layer6_outputs(2638) <= not (a xor b);
    layer6_outputs(2639) <= a;
    layer6_outputs(2640) <= not b;
    layer6_outputs(2641) <= not (a and b);
    layer6_outputs(2642) <= not (a and b);
    layer6_outputs(2643) <= b;
    layer6_outputs(2644) <= a and not b;
    layer6_outputs(2645) <= a and not b;
    layer6_outputs(2646) <= b;
    layer6_outputs(2647) <= a;
    layer6_outputs(2648) <= a and not b;
    layer6_outputs(2649) <= not a or b;
    layer6_outputs(2650) <= a;
    layer6_outputs(2651) <= a or b;
    layer6_outputs(2652) <= a;
    layer6_outputs(2653) <= a;
    layer6_outputs(2654) <= not (a and b);
    layer6_outputs(2655) <= a and not b;
    layer6_outputs(2656) <= not (a or b);
    layer6_outputs(2657) <= not (a xor b);
    layer6_outputs(2658) <= b;
    layer6_outputs(2659) <= b;
    layer6_outputs(2660) <= 1'b0;
    layer6_outputs(2661) <= not (a and b);
    layer6_outputs(2662) <= not (a and b);
    layer6_outputs(2663) <= b;
    layer6_outputs(2664) <= not a;
    layer6_outputs(2665) <= a or b;
    layer6_outputs(2666) <= a and b;
    layer6_outputs(2667) <= not b;
    layer6_outputs(2668) <= not b;
    layer6_outputs(2669) <= not b;
    layer6_outputs(2670) <= a and b;
    layer6_outputs(2671) <= b;
    layer6_outputs(2672) <= not a;
    layer6_outputs(2673) <= a;
    layer6_outputs(2674) <= b and not a;
    layer6_outputs(2675) <= not (a or b);
    layer6_outputs(2676) <= not b;
    layer6_outputs(2677) <= not a or b;
    layer6_outputs(2678) <= a or b;
    layer6_outputs(2679) <= not b or a;
    layer6_outputs(2680) <= not (a xor b);
    layer6_outputs(2681) <= not b;
    layer6_outputs(2682) <= not a or b;
    layer6_outputs(2683) <= not (a xor b);
    layer6_outputs(2684) <= b;
    layer6_outputs(2685) <= b;
    layer6_outputs(2686) <= a and b;
    layer6_outputs(2687) <= a and b;
    layer6_outputs(2688) <= not b or a;
    layer6_outputs(2689) <= not b or a;
    layer6_outputs(2690) <= b and not a;
    layer6_outputs(2691) <= not b;
    layer6_outputs(2692) <= b;
    layer6_outputs(2693) <= a;
    layer6_outputs(2694) <= a and not b;
    layer6_outputs(2695) <= a;
    layer6_outputs(2696) <= a and b;
    layer6_outputs(2697) <= not b;
    layer6_outputs(2698) <= a and not b;
    layer6_outputs(2699) <= a xor b;
    layer6_outputs(2700) <= not b;
    layer6_outputs(2701) <= b;
    layer6_outputs(2702) <= a;
    layer6_outputs(2703) <= a;
    layer6_outputs(2704) <= not b or a;
    layer6_outputs(2705) <= a;
    layer6_outputs(2706) <= not (a and b);
    layer6_outputs(2707) <= not b;
    layer6_outputs(2708) <= not a or b;
    layer6_outputs(2709) <= a and b;
    layer6_outputs(2710) <= not b or a;
    layer6_outputs(2711) <= a or b;
    layer6_outputs(2712) <= a or b;
    layer6_outputs(2713) <= not a;
    layer6_outputs(2714) <= a and not b;
    layer6_outputs(2715) <= not (a or b);
    layer6_outputs(2716) <= b;
    layer6_outputs(2717) <= not (a or b);
    layer6_outputs(2718) <= a and b;
    layer6_outputs(2719) <= b;
    layer6_outputs(2720) <= a;
    layer6_outputs(2721) <= 1'b1;
    layer6_outputs(2722) <= not (a or b);
    layer6_outputs(2723) <= b;
    layer6_outputs(2724) <= a;
    layer6_outputs(2725) <= 1'b1;
    layer6_outputs(2726) <= not b;
    layer6_outputs(2727) <= not (a xor b);
    layer6_outputs(2728) <= not a;
    layer6_outputs(2729) <= a;
    layer6_outputs(2730) <= b;
    layer6_outputs(2731) <= not b;
    layer6_outputs(2732) <= not (a and b);
    layer6_outputs(2733) <= not (a xor b);
    layer6_outputs(2734) <= 1'b1;
    layer6_outputs(2735) <= not (a and b);
    layer6_outputs(2736) <= a;
    layer6_outputs(2737) <= b and not a;
    layer6_outputs(2738) <= a xor b;
    layer6_outputs(2739) <= a;
    layer6_outputs(2740) <= b;
    layer6_outputs(2741) <= not (a xor b);
    layer6_outputs(2742) <= not b or a;
    layer6_outputs(2743) <= a xor b;
    layer6_outputs(2744) <= not (a xor b);
    layer6_outputs(2745) <= not (a and b);
    layer6_outputs(2746) <= 1'b0;
    layer6_outputs(2747) <= not a;
    layer6_outputs(2748) <= b;
    layer6_outputs(2749) <= a or b;
    layer6_outputs(2750) <= a and not b;
    layer6_outputs(2751) <= not a;
    layer6_outputs(2752) <= a;
    layer6_outputs(2753) <= not (a and b);
    layer6_outputs(2754) <= not a or b;
    layer6_outputs(2755) <= a;
    layer6_outputs(2756) <= not b;
    layer6_outputs(2757) <= a or b;
    layer6_outputs(2758) <= not b;
    layer6_outputs(2759) <= b and not a;
    layer6_outputs(2760) <= not a;
    layer6_outputs(2761) <= a and b;
    layer6_outputs(2762) <= a and b;
    layer6_outputs(2763) <= not (a and b);
    layer6_outputs(2764) <= b;
    layer6_outputs(2765) <= not a;
    layer6_outputs(2766) <= not (a or b);
    layer6_outputs(2767) <= b;
    layer6_outputs(2768) <= b and not a;
    layer6_outputs(2769) <= a or b;
    layer6_outputs(2770) <= a and b;
    layer6_outputs(2771) <= not (a xor b);
    layer6_outputs(2772) <= not (a and b);
    layer6_outputs(2773) <= b;
    layer6_outputs(2774) <= not b;
    layer6_outputs(2775) <= not b;
    layer6_outputs(2776) <= not a;
    layer6_outputs(2777) <= not a;
    layer6_outputs(2778) <= a or b;
    layer6_outputs(2779) <= not a;
    layer6_outputs(2780) <= a or b;
    layer6_outputs(2781) <= a xor b;
    layer6_outputs(2782) <= a;
    layer6_outputs(2783) <= not a;
    layer6_outputs(2784) <= b;
    layer6_outputs(2785) <= a and not b;
    layer6_outputs(2786) <= not (a xor b);
    layer6_outputs(2787) <= not b;
    layer6_outputs(2788) <= not b;
    layer6_outputs(2789) <= not b;
    layer6_outputs(2790) <= b;
    layer6_outputs(2791) <= b;
    layer6_outputs(2792) <= a and b;
    layer6_outputs(2793) <= not b or a;
    layer6_outputs(2794) <= a;
    layer6_outputs(2795) <= a and b;
    layer6_outputs(2796) <= not b;
    layer6_outputs(2797) <= a;
    layer6_outputs(2798) <= a xor b;
    layer6_outputs(2799) <= not b;
    layer6_outputs(2800) <= not (a xor b);
    layer6_outputs(2801) <= 1'b0;
    layer6_outputs(2802) <= a xor b;
    layer6_outputs(2803) <= not b or a;
    layer6_outputs(2804) <= a;
    layer6_outputs(2805) <= not a or b;
    layer6_outputs(2806) <= a;
    layer6_outputs(2807) <= not a or b;
    layer6_outputs(2808) <= not b;
    layer6_outputs(2809) <= not a;
    layer6_outputs(2810) <= not a;
    layer6_outputs(2811) <= not a;
    layer6_outputs(2812) <= not a;
    layer6_outputs(2813) <= 1'b1;
    layer6_outputs(2814) <= a and b;
    layer6_outputs(2815) <= 1'b0;
    layer6_outputs(2816) <= not a or b;
    layer6_outputs(2817) <= not a;
    layer6_outputs(2818) <= b;
    layer6_outputs(2819) <= b;
    layer6_outputs(2820) <= a and not b;
    layer6_outputs(2821) <= not a;
    layer6_outputs(2822) <= not (a or b);
    layer6_outputs(2823) <= a and b;
    layer6_outputs(2824) <= not b;
    layer6_outputs(2825) <= not a;
    layer6_outputs(2826) <= not b;
    layer6_outputs(2827) <= a and b;
    layer6_outputs(2828) <= b and not a;
    layer6_outputs(2829) <= a;
    layer6_outputs(2830) <= a or b;
    layer6_outputs(2831) <= a;
    layer6_outputs(2832) <= not b;
    layer6_outputs(2833) <= a and b;
    layer6_outputs(2834) <= a and b;
    layer6_outputs(2835) <= a and not b;
    layer6_outputs(2836) <= not b;
    layer6_outputs(2837) <= b;
    layer6_outputs(2838) <= not b or a;
    layer6_outputs(2839) <= not a or b;
    layer6_outputs(2840) <= a and not b;
    layer6_outputs(2841) <= not b or a;
    layer6_outputs(2842) <= not (a xor b);
    layer6_outputs(2843) <= 1'b0;
    layer6_outputs(2844) <= not b;
    layer6_outputs(2845) <= a and not b;
    layer6_outputs(2846) <= b and not a;
    layer6_outputs(2847) <= 1'b1;
    layer6_outputs(2848) <= b;
    layer6_outputs(2849) <= a;
    layer6_outputs(2850) <= not b;
    layer6_outputs(2851) <= b;
    layer6_outputs(2852) <= a and not b;
    layer6_outputs(2853) <= a;
    layer6_outputs(2854) <= not a or b;
    layer6_outputs(2855) <= b;
    layer6_outputs(2856) <= b;
    layer6_outputs(2857) <= not (a or b);
    layer6_outputs(2858) <= b;
    layer6_outputs(2859) <= b;
    layer6_outputs(2860) <= not (a or b);
    layer6_outputs(2861) <= b and not a;
    layer6_outputs(2862) <= b;
    layer6_outputs(2863) <= not b or a;
    layer6_outputs(2864) <= not a;
    layer6_outputs(2865) <= not b or a;
    layer6_outputs(2866) <= b and not a;
    layer6_outputs(2867) <= a or b;
    layer6_outputs(2868) <= a and b;
    layer6_outputs(2869) <= not a;
    layer6_outputs(2870) <= not a;
    layer6_outputs(2871) <= not b;
    layer6_outputs(2872) <= a;
    layer6_outputs(2873) <= not b or a;
    layer6_outputs(2874) <= a and not b;
    layer6_outputs(2875) <= 1'b1;
    layer6_outputs(2876) <= not a;
    layer6_outputs(2877) <= b and not a;
    layer6_outputs(2878) <= a;
    layer6_outputs(2879) <= b;
    layer6_outputs(2880) <= not a or b;
    layer6_outputs(2881) <= not a;
    layer6_outputs(2882) <= a xor b;
    layer6_outputs(2883) <= not a;
    layer6_outputs(2884) <= a or b;
    layer6_outputs(2885) <= not (a xor b);
    layer6_outputs(2886) <= 1'b0;
    layer6_outputs(2887) <= not (a or b);
    layer6_outputs(2888) <= 1'b0;
    layer6_outputs(2889) <= b;
    layer6_outputs(2890) <= not (a xor b);
    layer6_outputs(2891) <= a xor b;
    layer6_outputs(2892) <= not (a and b);
    layer6_outputs(2893) <= b;
    layer6_outputs(2894) <= a and not b;
    layer6_outputs(2895) <= b;
    layer6_outputs(2896) <= not (a xor b);
    layer6_outputs(2897) <= a;
    layer6_outputs(2898) <= a;
    layer6_outputs(2899) <= b;
    layer6_outputs(2900) <= b and not a;
    layer6_outputs(2901) <= b;
    layer6_outputs(2902) <= not a;
    layer6_outputs(2903) <= a;
    layer6_outputs(2904) <= not (a or b);
    layer6_outputs(2905) <= a or b;
    layer6_outputs(2906) <= a and b;
    layer6_outputs(2907) <= not a or b;
    layer6_outputs(2908) <= not b or a;
    layer6_outputs(2909) <= not a or b;
    layer6_outputs(2910) <= not (a and b);
    layer6_outputs(2911) <= not (a and b);
    layer6_outputs(2912) <= not (a or b);
    layer6_outputs(2913) <= 1'b0;
    layer6_outputs(2914) <= a and b;
    layer6_outputs(2915) <= not a;
    layer6_outputs(2916) <= not (a and b);
    layer6_outputs(2917) <= b;
    layer6_outputs(2918) <= not a;
    layer6_outputs(2919) <= not b or a;
    layer6_outputs(2920) <= not (a and b);
    layer6_outputs(2921) <= not (a or b);
    layer6_outputs(2922) <= not (a xor b);
    layer6_outputs(2923) <= a and b;
    layer6_outputs(2924) <= a;
    layer6_outputs(2925) <= a xor b;
    layer6_outputs(2926) <= not b;
    layer6_outputs(2927) <= b and not a;
    layer6_outputs(2928) <= a;
    layer6_outputs(2929) <= b;
    layer6_outputs(2930) <= not a or b;
    layer6_outputs(2931) <= 1'b0;
    layer6_outputs(2932) <= b;
    layer6_outputs(2933) <= not a;
    layer6_outputs(2934) <= a xor b;
    layer6_outputs(2935) <= b;
    layer6_outputs(2936) <= not (a xor b);
    layer6_outputs(2937) <= b and not a;
    layer6_outputs(2938) <= b and not a;
    layer6_outputs(2939) <= a xor b;
    layer6_outputs(2940) <= not b;
    layer6_outputs(2941) <= a xor b;
    layer6_outputs(2942) <= a;
    layer6_outputs(2943) <= a;
    layer6_outputs(2944) <= 1'b1;
    layer6_outputs(2945) <= a;
    layer6_outputs(2946) <= not (a and b);
    layer6_outputs(2947) <= not (a xor b);
    layer6_outputs(2948) <= not a;
    layer6_outputs(2949) <= a or b;
    layer6_outputs(2950) <= a and not b;
    layer6_outputs(2951) <= a and b;
    layer6_outputs(2952) <= a xor b;
    layer6_outputs(2953) <= a;
    layer6_outputs(2954) <= a or b;
    layer6_outputs(2955) <= a or b;
    layer6_outputs(2956) <= not (a or b);
    layer6_outputs(2957) <= b and not a;
    layer6_outputs(2958) <= not (a and b);
    layer6_outputs(2959) <= b and not a;
    layer6_outputs(2960) <= not b;
    layer6_outputs(2961) <= not (a xor b);
    layer6_outputs(2962) <= not b;
    layer6_outputs(2963) <= not (a xor b);
    layer6_outputs(2964) <= not a or b;
    layer6_outputs(2965) <= not (a and b);
    layer6_outputs(2966) <= a and b;
    layer6_outputs(2967) <= not (a and b);
    layer6_outputs(2968) <= a or b;
    layer6_outputs(2969) <= not (a or b);
    layer6_outputs(2970) <= a xor b;
    layer6_outputs(2971) <= not a;
    layer6_outputs(2972) <= 1'b0;
    layer6_outputs(2973) <= not b;
    layer6_outputs(2974) <= not b;
    layer6_outputs(2975) <= 1'b0;
    layer6_outputs(2976) <= not (a and b);
    layer6_outputs(2977) <= not b;
    layer6_outputs(2978) <= a and b;
    layer6_outputs(2979) <= a xor b;
    layer6_outputs(2980) <= b and not a;
    layer6_outputs(2981) <= a and b;
    layer6_outputs(2982) <= not b;
    layer6_outputs(2983) <= 1'b0;
    layer6_outputs(2984) <= not a or b;
    layer6_outputs(2985) <= not a or b;
    layer6_outputs(2986) <= not b or a;
    layer6_outputs(2987) <= a and not b;
    layer6_outputs(2988) <= b and not a;
    layer6_outputs(2989) <= a and not b;
    layer6_outputs(2990) <= not b;
    layer6_outputs(2991) <= b and not a;
    layer6_outputs(2992) <= a xor b;
    layer6_outputs(2993) <= not (a xor b);
    layer6_outputs(2994) <= a xor b;
    layer6_outputs(2995) <= not (a or b);
    layer6_outputs(2996) <= not a;
    layer6_outputs(2997) <= not a;
    layer6_outputs(2998) <= a xor b;
    layer6_outputs(2999) <= a;
    layer6_outputs(3000) <= not (a and b);
    layer6_outputs(3001) <= not b;
    layer6_outputs(3002) <= not a;
    layer6_outputs(3003) <= not b;
    layer6_outputs(3004) <= b and not a;
    layer6_outputs(3005) <= a xor b;
    layer6_outputs(3006) <= not a or b;
    layer6_outputs(3007) <= not b;
    layer6_outputs(3008) <= a and not b;
    layer6_outputs(3009) <= not a;
    layer6_outputs(3010) <= a and b;
    layer6_outputs(3011) <= a or b;
    layer6_outputs(3012) <= a;
    layer6_outputs(3013) <= not a;
    layer6_outputs(3014) <= not a or b;
    layer6_outputs(3015) <= not (a and b);
    layer6_outputs(3016) <= not b or a;
    layer6_outputs(3017) <= 1'b0;
    layer6_outputs(3018) <= not (a xor b);
    layer6_outputs(3019) <= not (a or b);
    layer6_outputs(3020) <= b;
    layer6_outputs(3021) <= not a;
    layer6_outputs(3022) <= not (a xor b);
    layer6_outputs(3023) <= not a;
    layer6_outputs(3024) <= a xor b;
    layer6_outputs(3025) <= b and not a;
    layer6_outputs(3026) <= a and b;
    layer6_outputs(3027) <= not (a and b);
    layer6_outputs(3028) <= a and b;
    layer6_outputs(3029) <= b;
    layer6_outputs(3030) <= b;
    layer6_outputs(3031) <= a xor b;
    layer6_outputs(3032) <= not a or b;
    layer6_outputs(3033) <= a xor b;
    layer6_outputs(3034) <= not (a or b);
    layer6_outputs(3035) <= a;
    layer6_outputs(3036) <= a xor b;
    layer6_outputs(3037) <= 1'b1;
    layer6_outputs(3038) <= a and not b;
    layer6_outputs(3039) <= a and not b;
    layer6_outputs(3040) <= not (a and b);
    layer6_outputs(3041) <= not b or a;
    layer6_outputs(3042) <= not b;
    layer6_outputs(3043) <= a;
    layer6_outputs(3044) <= not a or b;
    layer6_outputs(3045) <= b and not a;
    layer6_outputs(3046) <= b;
    layer6_outputs(3047) <= a and not b;
    layer6_outputs(3048) <= not b;
    layer6_outputs(3049) <= not a;
    layer6_outputs(3050) <= not a;
    layer6_outputs(3051) <= not (a xor b);
    layer6_outputs(3052) <= a and not b;
    layer6_outputs(3053) <= not a;
    layer6_outputs(3054) <= a;
    layer6_outputs(3055) <= not a;
    layer6_outputs(3056) <= not a;
    layer6_outputs(3057) <= b and not a;
    layer6_outputs(3058) <= 1'b1;
    layer6_outputs(3059) <= a or b;
    layer6_outputs(3060) <= b and not a;
    layer6_outputs(3061) <= a xor b;
    layer6_outputs(3062) <= b and not a;
    layer6_outputs(3063) <= not (a or b);
    layer6_outputs(3064) <= not (a or b);
    layer6_outputs(3065) <= not (a and b);
    layer6_outputs(3066) <= 1'b1;
    layer6_outputs(3067) <= a and b;
    layer6_outputs(3068) <= 1'b1;
    layer6_outputs(3069) <= 1'b1;
    layer6_outputs(3070) <= a and not b;
    layer6_outputs(3071) <= not a;
    layer6_outputs(3072) <= a or b;
    layer6_outputs(3073) <= not a or b;
    layer6_outputs(3074) <= not a;
    layer6_outputs(3075) <= b;
    layer6_outputs(3076) <= a or b;
    layer6_outputs(3077) <= not b;
    layer6_outputs(3078) <= not a;
    layer6_outputs(3079) <= b and not a;
    layer6_outputs(3080) <= not a;
    layer6_outputs(3081) <= not (a and b);
    layer6_outputs(3082) <= not b;
    layer6_outputs(3083) <= a or b;
    layer6_outputs(3084) <= b;
    layer6_outputs(3085) <= a or b;
    layer6_outputs(3086) <= not a or b;
    layer6_outputs(3087) <= 1'b0;
    layer6_outputs(3088) <= not a;
    layer6_outputs(3089) <= a or b;
    layer6_outputs(3090) <= a and not b;
    layer6_outputs(3091) <= 1'b1;
    layer6_outputs(3092) <= a xor b;
    layer6_outputs(3093) <= b;
    layer6_outputs(3094) <= not (a or b);
    layer6_outputs(3095) <= b;
    layer6_outputs(3096) <= not (a and b);
    layer6_outputs(3097) <= b and not a;
    layer6_outputs(3098) <= not b;
    layer6_outputs(3099) <= b and not a;
    layer6_outputs(3100) <= not a;
    layer6_outputs(3101) <= b;
    layer6_outputs(3102) <= b;
    layer6_outputs(3103) <= a;
    layer6_outputs(3104) <= b and not a;
    layer6_outputs(3105) <= b;
    layer6_outputs(3106) <= not a;
    layer6_outputs(3107) <= not b;
    layer6_outputs(3108) <= 1'b1;
    layer6_outputs(3109) <= a and not b;
    layer6_outputs(3110) <= a xor b;
    layer6_outputs(3111) <= a and b;
    layer6_outputs(3112) <= a or b;
    layer6_outputs(3113) <= not (a and b);
    layer6_outputs(3114) <= not a or b;
    layer6_outputs(3115) <= b and not a;
    layer6_outputs(3116) <= a;
    layer6_outputs(3117) <= 1'b0;
    layer6_outputs(3118) <= a and b;
    layer6_outputs(3119) <= not (a xor b);
    layer6_outputs(3120) <= a or b;
    layer6_outputs(3121) <= a;
    layer6_outputs(3122) <= not a;
    layer6_outputs(3123) <= not (a and b);
    layer6_outputs(3124) <= not b;
    layer6_outputs(3125) <= b and not a;
    layer6_outputs(3126) <= not b;
    layer6_outputs(3127) <= not b or a;
    layer6_outputs(3128) <= a and b;
    layer6_outputs(3129) <= a xor b;
    layer6_outputs(3130) <= a and not b;
    layer6_outputs(3131) <= not b;
    layer6_outputs(3132) <= not (a or b);
    layer6_outputs(3133) <= not (a and b);
    layer6_outputs(3134) <= not b;
    layer6_outputs(3135) <= b;
    layer6_outputs(3136) <= not (a xor b);
    layer6_outputs(3137) <= b;
    layer6_outputs(3138) <= a;
    layer6_outputs(3139) <= a;
    layer6_outputs(3140) <= not a or b;
    layer6_outputs(3141) <= not a;
    layer6_outputs(3142) <= not (a and b);
    layer6_outputs(3143) <= a;
    layer6_outputs(3144) <= not (a xor b);
    layer6_outputs(3145) <= 1'b0;
    layer6_outputs(3146) <= not b;
    layer6_outputs(3147) <= not (a and b);
    layer6_outputs(3148) <= not b or a;
    layer6_outputs(3149) <= b and not a;
    layer6_outputs(3150) <= a or b;
    layer6_outputs(3151) <= not b;
    layer6_outputs(3152) <= not a or b;
    layer6_outputs(3153) <= a and b;
    layer6_outputs(3154) <= not b;
    layer6_outputs(3155) <= not (a xor b);
    layer6_outputs(3156) <= not (a or b);
    layer6_outputs(3157) <= 1'b0;
    layer6_outputs(3158) <= b and not a;
    layer6_outputs(3159) <= not a or b;
    layer6_outputs(3160) <= not (a and b);
    layer6_outputs(3161) <= a or b;
    layer6_outputs(3162) <= not a;
    layer6_outputs(3163) <= a xor b;
    layer6_outputs(3164) <= a and not b;
    layer6_outputs(3165) <= a and not b;
    layer6_outputs(3166) <= b and not a;
    layer6_outputs(3167) <= not (a xor b);
    layer6_outputs(3168) <= not (a or b);
    layer6_outputs(3169) <= not (a xor b);
    layer6_outputs(3170) <= not a;
    layer6_outputs(3171) <= b and not a;
    layer6_outputs(3172) <= not a or b;
    layer6_outputs(3173) <= not (a xor b);
    layer6_outputs(3174) <= a xor b;
    layer6_outputs(3175) <= 1'b0;
    layer6_outputs(3176) <= not (a xor b);
    layer6_outputs(3177) <= a and b;
    layer6_outputs(3178) <= b;
    layer6_outputs(3179) <= b;
    layer6_outputs(3180) <= not a;
    layer6_outputs(3181) <= a;
    layer6_outputs(3182) <= a and not b;
    layer6_outputs(3183) <= not (a xor b);
    layer6_outputs(3184) <= a xor b;
    layer6_outputs(3185) <= a;
    layer6_outputs(3186) <= a and b;
    layer6_outputs(3187) <= not b;
    layer6_outputs(3188) <= not (a xor b);
    layer6_outputs(3189) <= a and not b;
    layer6_outputs(3190) <= not (a xor b);
    layer6_outputs(3191) <= b and not a;
    layer6_outputs(3192) <= not a or b;
    layer6_outputs(3193) <= a and not b;
    layer6_outputs(3194) <= not a;
    layer6_outputs(3195) <= not a or b;
    layer6_outputs(3196) <= not b;
    layer6_outputs(3197) <= a;
    layer6_outputs(3198) <= a and b;
    layer6_outputs(3199) <= b and not a;
    layer6_outputs(3200) <= a;
    layer6_outputs(3201) <= 1'b1;
    layer6_outputs(3202) <= not (a or b);
    layer6_outputs(3203) <= a;
    layer6_outputs(3204) <= a xor b;
    layer6_outputs(3205) <= 1'b0;
    layer6_outputs(3206) <= a xor b;
    layer6_outputs(3207) <= b and not a;
    layer6_outputs(3208) <= a or b;
    layer6_outputs(3209) <= not b or a;
    layer6_outputs(3210) <= not a;
    layer6_outputs(3211) <= a and b;
    layer6_outputs(3212) <= b and not a;
    layer6_outputs(3213) <= a and not b;
    layer6_outputs(3214) <= not a;
    layer6_outputs(3215) <= a;
    layer6_outputs(3216) <= a;
    layer6_outputs(3217) <= not b or a;
    layer6_outputs(3218) <= a;
    layer6_outputs(3219) <= a or b;
    layer6_outputs(3220) <= a xor b;
    layer6_outputs(3221) <= a and b;
    layer6_outputs(3222) <= not b;
    layer6_outputs(3223) <= a;
    layer6_outputs(3224) <= not a or b;
    layer6_outputs(3225) <= a and b;
    layer6_outputs(3226) <= not a;
    layer6_outputs(3227) <= not b;
    layer6_outputs(3228) <= not a or b;
    layer6_outputs(3229) <= a and not b;
    layer6_outputs(3230) <= a xor b;
    layer6_outputs(3231) <= not a or b;
    layer6_outputs(3232) <= not a or b;
    layer6_outputs(3233) <= not (a and b);
    layer6_outputs(3234) <= not b;
    layer6_outputs(3235) <= not b;
    layer6_outputs(3236) <= not b;
    layer6_outputs(3237) <= not (a xor b);
    layer6_outputs(3238) <= b;
    layer6_outputs(3239) <= not b or a;
    layer6_outputs(3240) <= b and not a;
    layer6_outputs(3241) <= not b;
    layer6_outputs(3242) <= b and not a;
    layer6_outputs(3243) <= 1'b0;
    layer6_outputs(3244) <= not a or b;
    layer6_outputs(3245) <= not b;
    layer6_outputs(3246) <= not a;
    layer6_outputs(3247) <= b;
    layer6_outputs(3248) <= not b or a;
    layer6_outputs(3249) <= a;
    layer6_outputs(3250) <= not b or a;
    layer6_outputs(3251) <= not a or b;
    layer6_outputs(3252) <= a or b;
    layer6_outputs(3253) <= b and not a;
    layer6_outputs(3254) <= a;
    layer6_outputs(3255) <= not b;
    layer6_outputs(3256) <= not (a xor b);
    layer6_outputs(3257) <= a and not b;
    layer6_outputs(3258) <= not b or a;
    layer6_outputs(3259) <= not b;
    layer6_outputs(3260) <= not b or a;
    layer6_outputs(3261) <= not (a or b);
    layer6_outputs(3262) <= a and not b;
    layer6_outputs(3263) <= not (a or b);
    layer6_outputs(3264) <= b;
    layer6_outputs(3265) <= a xor b;
    layer6_outputs(3266) <= not b;
    layer6_outputs(3267) <= not b;
    layer6_outputs(3268) <= not a;
    layer6_outputs(3269) <= not b;
    layer6_outputs(3270) <= a;
    layer6_outputs(3271) <= 1'b1;
    layer6_outputs(3272) <= not b;
    layer6_outputs(3273) <= 1'b0;
    layer6_outputs(3274) <= not b;
    layer6_outputs(3275) <= a or b;
    layer6_outputs(3276) <= not a;
    layer6_outputs(3277) <= a and not b;
    layer6_outputs(3278) <= 1'b1;
    layer6_outputs(3279) <= b;
    layer6_outputs(3280) <= a xor b;
    layer6_outputs(3281) <= a or b;
    layer6_outputs(3282) <= b;
    layer6_outputs(3283) <= not a;
    layer6_outputs(3284) <= not a;
    layer6_outputs(3285) <= a and b;
    layer6_outputs(3286) <= not (a or b);
    layer6_outputs(3287) <= a;
    layer6_outputs(3288) <= not (a and b);
    layer6_outputs(3289) <= a and b;
    layer6_outputs(3290) <= not a or b;
    layer6_outputs(3291) <= not (a and b);
    layer6_outputs(3292) <= a or b;
    layer6_outputs(3293) <= 1'b1;
    layer6_outputs(3294) <= a and not b;
    layer6_outputs(3295) <= b and not a;
    layer6_outputs(3296) <= not a;
    layer6_outputs(3297) <= not (a or b);
    layer6_outputs(3298) <= a and not b;
    layer6_outputs(3299) <= not (a xor b);
    layer6_outputs(3300) <= not (a xor b);
    layer6_outputs(3301) <= a and b;
    layer6_outputs(3302) <= a;
    layer6_outputs(3303) <= b;
    layer6_outputs(3304) <= not b;
    layer6_outputs(3305) <= not a;
    layer6_outputs(3306) <= not (a or b);
    layer6_outputs(3307) <= not a or b;
    layer6_outputs(3308) <= not (a or b);
    layer6_outputs(3309) <= not b or a;
    layer6_outputs(3310) <= b and not a;
    layer6_outputs(3311) <= not b or a;
    layer6_outputs(3312) <= b;
    layer6_outputs(3313) <= not (a or b);
    layer6_outputs(3314) <= not a;
    layer6_outputs(3315) <= 1'b1;
    layer6_outputs(3316) <= b;
    layer6_outputs(3317) <= not (a xor b);
    layer6_outputs(3318) <= a xor b;
    layer6_outputs(3319) <= a;
    layer6_outputs(3320) <= a;
    layer6_outputs(3321) <= b;
    layer6_outputs(3322) <= a or b;
    layer6_outputs(3323) <= not (a and b);
    layer6_outputs(3324) <= 1'b0;
    layer6_outputs(3325) <= a xor b;
    layer6_outputs(3326) <= not (a or b);
    layer6_outputs(3327) <= b;
    layer6_outputs(3328) <= 1'b0;
    layer6_outputs(3329) <= not b;
    layer6_outputs(3330) <= not a;
    layer6_outputs(3331) <= a;
    layer6_outputs(3332) <= not b or a;
    layer6_outputs(3333) <= 1'b0;
    layer6_outputs(3334) <= b;
    layer6_outputs(3335) <= a and b;
    layer6_outputs(3336) <= not b;
    layer6_outputs(3337) <= not (a or b);
    layer6_outputs(3338) <= not a;
    layer6_outputs(3339) <= not b;
    layer6_outputs(3340) <= not b;
    layer6_outputs(3341) <= a or b;
    layer6_outputs(3342) <= 1'b0;
    layer6_outputs(3343) <= not b or a;
    layer6_outputs(3344) <= a and b;
    layer6_outputs(3345) <= a xor b;
    layer6_outputs(3346) <= not (a and b);
    layer6_outputs(3347) <= not (a or b);
    layer6_outputs(3348) <= not b;
    layer6_outputs(3349) <= b;
    layer6_outputs(3350) <= not (a xor b);
    layer6_outputs(3351) <= not b;
    layer6_outputs(3352) <= not b;
    layer6_outputs(3353) <= not a or b;
    layer6_outputs(3354) <= not b;
    layer6_outputs(3355) <= b;
    layer6_outputs(3356) <= b;
    layer6_outputs(3357) <= not b;
    layer6_outputs(3358) <= not b;
    layer6_outputs(3359) <= not (a and b);
    layer6_outputs(3360) <= a;
    layer6_outputs(3361) <= b and not a;
    layer6_outputs(3362) <= a;
    layer6_outputs(3363) <= not b;
    layer6_outputs(3364) <= not b or a;
    layer6_outputs(3365) <= a;
    layer6_outputs(3366) <= not a or b;
    layer6_outputs(3367) <= a or b;
    layer6_outputs(3368) <= a;
    layer6_outputs(3369) <= a;
    layer6_outputs(3370) <= b;
    layer6_outputs(3371) <= not (a or b);
    layer6_outputs(3372) <= not b or a;
    layer6_outputs(3373) <= a and b;
    layer6_outputs(3374) <= b;
    layer6_outputs(3375) <= not (a xor b);
    layer6_outputs(3376) <= a;
    layer6_outputs(3377) <= not a or b;
    layer6_outputs(3378) <= not b;
    layer6_outputs(3379) <= b;
    layer6_outputs(3380) <= not (a or b);
    layer6_outputs(3381) <= not b;
    layer6_outputs(3382) <= b and not a;
    layer6_outputs(3383) <= a;
    layer6_outputs(3384) <= b and not a;
    layer6_outputs(3385) <= not a;
    layer6_outputs(3386) <= b and not a;
    layer6_outputs(3387) <= 1'b0;
    layer6_outputs(3388) <= not (a or b);
    layer6_outputs(3389) <= a;
    layer6_outputs(3390) <= not (a or b);
    layer6_outputs(3391) <= 1'b0;
    layer6_outputs(3392) <= b;
    layer6_outputs(3393) <= not a or b;
    layer6_outputs(3394) <= not a;
    layer6_outputs(3395) <= not b;
    layer6_outputs(3396) <= b;
    layer6_outputs(3397) <= b;
    layer6_outputs(3398) <= b;
    layer6_outputs(3399) <= not b or a;
    layer6_outputs(3400) <= not (a xor b);
    layer6_outputs(3401) <= not a;
    layer6_outputs(3402) <= not (a and b);
    layer6_outputs(3403) <= 1'b0;
    layer6_outputs(3404) <= not a or b;
    layer6_outputs(3405) <= not a;
    layer6_outputs(3406) <= not a or b;
    layer6_outputs(3407) <= not (a and b);
    layer6_outputs(3408) <= 1'b0;
    layer6_outputs(3409) <= not a or b;
    layer6_outputs(3410) <= not b;
    layer6_outputs(3411) <= not b;
    layer6_outputs(3412) <= a;
    layer6_outputs(3413) <= 1'b0;
    layer6_outputs(3414) <= b and not a;
    layer6_outputs(3415) <= not a;
    layer6_outputs(3416) <= b and not a;
    layer6_outputs(3417) <= not (a xor b);
    layer6_outputs(3418) <= a or b;
    layer6_outputs(3419) <= b;
    layer6_outputs(3420) <= not a or b;
    layer6_outputs(3421) <= a or b;
    layer6_outputs(3422) <= not b;
    layer6_outputs(3423) <= not b or a;
    layer6_outputs(3424) <= a;
    layer6_outputs(3425) <= a xor b;
    layer6_outputs(3426) <= not a;
    layer6_outputs(3427) <= not b or a;
    layer6_outputs(3428) <= not b;
    layer6_outputs(3429) <= not a;
    layer6_outputs(3430) <= a xor b;
    layer6_outputs(3431) <= a or b;
    layer6_outputs(3432) <= not (a xor b);
    layer6_outputs(3433) <= not b;
    layer6_outputs(3434) <= not b;
    layer6_outputs(3435) <= a and b;
    layer6_outputs(3436) <= not b or a;
    layer6_outputs(3437) <= a and not b;
    layer6_outputs(3438) <= not a;
    layer6_outputs(3439) <= not b;
    layer6_outputs(3440) <= b and not a;
    layer6_outputs(3441) <= a and b;
    layer6_outputs(3442) <= not a;
    layer6_outputs(3443) <= a or b;
    layer6_outputs(3444) <= a xor b;
    layer6_outputs(3445) <= a;
    layer6_outputs(3446) <= not (a xor b);
    layer6_outputs(3447) <= a and not b;
    layer6_outputs(3448) <= a xor b;
    layer6_outputs(3449) <= not b;
    layer6_outputs(3450) <= not a;
    layer6_outputs(3451) <= a and not b;
    layer6_outputs(3452) <= not (a xor b);
    layer6_outputs(3453) <= a and b;
    layer6_outputs(3454) <= not b;
    layer6_outputs(3455) <= a;
    layer6_outputs(3456) <= b;
    layer6_outputs(3457) <= not a;
    layer6_outputs(3458) <= not b;
    layer6_outputs(3459) <= b and not a;
    layer6_outputs(3460) <= b and not a;
    layer6_outputs(3461) <= not (a or b);
    layer6_outputs(3462) <= b;
    layer6_outputs(3463) <= not b;
    layer6_outputs(3464) <= a or b;
    layer6_outputs(3465) <= not a;
    layer6_outputs(3466) <= not a;
    layer6_outputs(3467) <= not a;
    layer6_outputs(3468) <= a;
    layer6_outputs(3469) <= not b;
    layer6_outputs(3470) <= not (a or b);
    layer6_outputs(3471) <= not (a xor b);
    layer6_outputs(3472) <= not (a or b);
    layer6_outputs(3473) <= not (a xor b);
    layer6_outputs(3474) <= a xor b;
    layer6_outputs(3475) <= a xor b;
    layer6_outputs(3476) <= not (a and b);
    layer6_outputs(3477) <= not b;
    layer6_outputs(3478) <= a and not b;
    layer6_outputs(3479) <= not b;
    layer6_outputs(3480) <= b and not a;
    layer6_outputs(3481) <= a or b;
    layer6_outputs(3482) <= not (a xor b);
    layer6_outputs(3483) <= not (a xor b);
    layer6_outputs(3484) <= not (a or b);
    layer6_outputs(3485) <= a or b;
    layer6_outputs(3486) <= a or b;
    layer6_outputs(3487) <= a;
    layer6_outputs(3488) <= a;
    layer6_outputs(3489) <= a;
    layer6_outputs(3490) <= a and b;
    layer6_outputs(3491) <= a and b;
    layer6_outputs(3492) <= a or b;
    layer6_outputs(3493) <= not (a or b);
    layer6_outputs(3494) <= b;
    layer6_outputs(3495) <= not (a or b);
    layer6_outputs(3496) <= b;
    layer6_outputs(3497) <= b;
    layer6_outputs(3498) <= a xor b;
    layer6_outputs(3499) <= not a;
    layer6_outputs(3500) <= not b;
    layer6_outputs(3501) <= not (a and b);
    layer6_outputs(3502) <= a;
    layer6_outputs(3503) <= a and not b;
    layer6_outputs(3504) <= a and b;
    layer6_outputs(3505) <= not b;
    layer6_outputs(3506) <= a;
    layer6_outputs(3507) <= not (a xor b);
    layer6_outputs(3508) <= 1'b0;
    layer6_outputs(3509) <= a xor b;
    layer6_outputs(3510) <= b and not a;
    layer6_outputs(3511) <= a;
    layer6_outputs(3512) <= b;
    layer6_outputs(3513) <= b and not a;
    layer6_outputs(3514) <= a and not b;
    layer6_outputs(3515) <= a;
    layer6_outputs(3516) <= not (a or b);
    layer6_outputs(3517) <= not b or a;
    layer6_outputs(3518) <= a and not b;
    layer6_outputs(3519) <= a;
    layer6_outputs(3520) <= not b;
    layer6_outputs(3521) <= a xor b;
    layer6_outputs(3522) <= not b or a;
    layer6_outputs(3523) <= not (a xor b);
    layer6_outputs(3524) <= b;
    layer6_outputs(3525) <= not a;
    layer6_outputs(3526) <= not (a and b);
    layer6_outputs(3527) <= a and b;
    layer6_outputs(3528) <= a and not b;
    layer6_outputs(3529) <= a;
    layer6_outputs(3530) <= a xor b;
    layer6_outputs(3531) <= not b;
    layer6_outputs(3532) <= not (a or b);
    layer6_outputs(3533) <= not (a xor b);
    layer6_outputs(3534) <= not (a and b);
    layer6_outputs(3535) <= not (a and b);
    layer6_outputs(3536) <= b and not a;
    layer6_outputs(3537) <= not a;
    layer6_outputs(3538) <= 1'b0;
    layer6_outputs(3539) <= not b or a;
    layer6_outputs(3540) <= not a or b;
    layer6_outputs(3541) <= b;
    layer6_outputs(3542) <= b;
    layer6_outputs(3543) <= not a;
    layer6_outputs(3544) <= not a;
    layer6_outputs(3545) <= not b;
    layer6_outputs(3546) <= not a;
    layer6_outputs(3547) <= not a;
    layer6_outputs(3548) <= not b;
    layer6_outputs(3549) <= not b;
    layer6_outputs(3550) <= a or b;
    layer6_outputs(3551) <= 1'b0;
    layer6_outputs(3552) <= a;
    layer6_outputs(3553) <= not (a and b);
    layer6_outputs(3554) <= 1'b0;
    layer6_outputs(3555) <= not a;
    layer6_outputs(3556) <= b;
    layer6_outputs(3557) <= b;
    layer6_outputs(3558) <= b and not a;
    layer6_outputs(3559) <= not b or a;
    layer6_outputs(3560) <= a;
    layer6_outputs(3561) <= a and not b;
    layer6_outputs(3562) <= a and not b;
    layer6_outputs(3563) <= not a or b;
    layer6_outputs(3564) <= a;
    layer6_outputs(3565) <= a;
    layer6_outputs(3566) <= b;
    layer6_outputs(3567) <= not (a or b);
    layer6_outputs(3568) <= b and not a;
    layer6_outputs(3569) <= not a;
    layer6_outputs(3570) <= a and b;
    layer6_outputs(3571) <= not (a or b);
    layer6_outputs(3572) <= b and not a;
    layer6_outputs(3573) <= b;
    layer6_outputs(3574) <= not b;
    layer6_outputs(3575) <= not (a and b);
    layer6_outputs(3576) <= a or b;
    layer6_outputs(3577) <= not b or a;
    layer6_outputs(3578) <= a;
    layer6_outputs(3579) <= not b or a;
    layer6_outputs(3580) <= not (a xor b);
    layer6_outputs(3581) <= b;
    layer6_outputs(3582) <= not b;
    layer6_outputs(3583) <= a and not b;
    layer6_outputs(3584) <= b and not a;
    layer6_outputs(3585) <= not (a or b);
    layer6_outputs(3586) <= not b or a;
    layer6_outputs(3587) <= a and not b;
    layer6_outputs(3588) <= a;
    layer6_outputs(3589) <= b and not a;
    layer6_outputs(3590) <= b and not a;
    layer6_outputs(3591) <= b;
    layer6_outputs(3592) <= not a;
    layer6_outputs(3593) <= not (a and b);
    layer6_outputs(3594) <= not a;
    layer6_outputs(3595) <= a xor b;
    layer6_outputs(3596) <= not (a or b);
    layer6_outputs(3597) <= not (a or b);
    layer6_outputs(3598) <= not a;
    layer6_outputs(3599) <= not a or b;
    layer6_outputs(3600) <= a or b;
    layer6_outputs(3601) <= b;
    layer6_outputs(3602) <= not b;
    layer6_outputs(3603) <= a or b;
    layer6_outputs(3604) <= 1'b1;
    layer6_outputs(3605) <= not a;
    layer6_outputs(3606) <= not b;
    layer6_outputs(3607) <= a or b;
    layer6_outputs(3608) <= b and not a;
    layer6_outputs(3609) <= not (a and b);
    layer6_outputs(3610) <= b;
    layer6_outputs(3611) <= 1'b1;
    layer6_outputs(3612) <= not a;
    layer6_outputs(3613) <= b;
    layer6_outputs(3614) <= not a or b;
    layer6_outputs(3615) <= not a;
    layer6_outputs(3616) <= a xor b;
    layer6_outputs(3617) <= b and not a;
    layer6_outputs(3618) <= a or b;
    layer6_outputs(3619) <= a;
    layer6_outputs(3620) <= a;
    layer6_outputs(3621) <= not b;
    layer6_outputs(3622) <= b;
    layer6_outputs(3623) <= not b or a;
    layer6_outputs(3624) <= not a;
    layer6_outputs(3625) <= a or b;
    layer6_outputs(3626) <= a;
    layer6_outputs(3627) <= not (a xor b);
    layer6_outputs(3628) <= not a;
    layer6_outputs(3629) <= b and not a;
    layer6_outputs(3630) <= a;
    layer6_outputs(3631) <= not (a or b);
    layer6_outputs(3632) <= not (a xor b);
    layer6_outputs(3633) <= not (a xor b);
    layer6_outputs(3634) <= not b;
    layer6_outputs(3635) <= not a;
    layer6_outputs(3636) <= a or b;
    layer6_outputs(3637) <= not a;
    layer6_outputs(3638) <= not b;
    layer6_outputs(3639) <= not a;
    layer6_outputs(3640) <= b;
    layer6_outputs(3641) <= not (a or b);
    layer6_outputs(3642) <= not b or a;
    layer6_outputs(3643) <= 1'b1;
    layer6_outputs(3644) <= not b;
    layer6_outputs(3645) <= not (a xor b);
    layer6_outputs(3646) <= not b;
    layer6_outputs(3647) <= a xor b;
    layer6_outputs(3648) <= not (a xor b);
    layer6_outputs(3649) <= b;
    layer6_outputs(3650) <= a;
    layer6_outputs(3651) <= b;
    layer6_outputs(3652) <= a and b;
    layer6_outputs(3653) <= not b;
    layer6_outputs(3654) <= not a;
    layer6_outputs(3655) <= a or b;
    layer6_outputs(3656) <= b;
    layer6_outputs(3657) <= not b or a;
    layer6_outputs(3658) <= a and b;
    layer6_outputs(3659) <= not (a and b);
    layer6_outputs(3660) <= a and not b;
    layer6_outputs(3661) <= not (a xor b);
    layer6_outputs(3662) <= not a or b;
    layer6_outputs(3663) <= a and not b;
    layer6_outputs(3664) <= not a;
    layer6_outputs(3665) <= a and b;
    layer6_outputs(3666) <= a and b;
    layer6_outputs(3667) <= b;
    layer6_outputs(3668) <= a xor b;
    layer6_outputs(3669) <= not a;
    layer6_outputs(3670) <= a and b;
    layer6_outputs(3671) <= b;
    layer6_outputs(3672) <= 1'b0;
    layer6_outputs(3673) <= a;
    layer6_outputs(3674) <= b;
    layer6_outputs(3675) <= not (a or b);
    layer6_outputs(3676) <= not (a or b);
    layer6_outputs(3677) <= a and b;
    layer6_outputs(3678) <= not b or a;
    layer6_outputs(3679) <= not b or a;
    layer6_outputs(3680) <= b and not a;
    layer6_outputs(3681) <= not b;
    layer6_outputs(3682) <= not b;
    layer6_outputs(3683) <= a;
    layer6_outputs(3684) <= a;
    layer6_outputs(3685) <= not a;
    layer6_outputs(3686) <= not (a xor b);
    layer6_outputs(3687) <= b;
    layer6_outputs(3688) <= not b;
    layer6_outputs(3689) <= not b;
    layer6_outputs(3690) <= not (a or b);
    layer6_outputs(3691) <= a and not b;
    layer6_outputs(3692) <= not (a or b);
    layer6_outputs(3693) <= not a or b;
    layer6_outputs(3694) <= not b;
    layer6_outputs(3695) <= not b;
    layer6_outputs(3696) <= 1'b0;
    layer6_outputs(3697) <= a or b;
    layer6_outputs(3698) <= b;
    layer6_outputs(3699) <= a and b;
    layer6_outputs(3700) <= a and b;
    layer6_outputs(3701) <= not (a or b);
    layer6_outputs(3702) <= not (a and b);
    layer6_outputs(3703) <= not (a and b);
    layer6_outputs(3704) <= a and b;
    layer6_outputs(3705) <= a and b;
    layer6_outputs(3706) <= not (a or b);
    layer6_outputs(3707) <= not (a and b);
    layer6_outputs(3708) <= b;
    layer6_outputs(3709) <= not a or b;
    layer6_outputs(3710) <= not a;
    layer6_outputs(3711) <= not (a xor b);
    layer6_outputs(3712) <= not a;
    layer6_outputs(3713) <= not a;
    layer6_outputs(3714) <= not b;
    layer6_outputs(3715) <= not b;
    layer6_outputs(3716) <= a and not b;
    layer6_outputs(3717) <= a and b;
    layer6_outputs(3718) <= a or b;
    layer6_outputs(3719) <= b;
    layer6_outputs(3720) <= a;
    layer6_outputs(3721) <= b;
    layer6_outputs(3722) <= not a or b;
    layer6_outputs(3723) <= 1'b1;
    layer6_outputs(3724) <= not b or a;
    layer6_outputs(3725) <= not a;
    layer6_outputs(3726) <= not b or a;
    layer6_outputs(3727) <= a;
    layer6_outputs(3728) <= not (a xor b);
    layer6_outputs(3729) <= not b or a;
    layer6_outputs(3730) <= b and not a;
    layer6_outputs(3731) <= not b;
    layer6_outputs(3732) <= a and b;
    layer6_outputs(3733) <= 1'b0;
    layer6_outputs(3734) <= not b;
    layer6_outputs(3735) <= b;
    layer6_outputs(3736) <= not b;
    layer6_outputs(3737) <= a;
    layer6_outputs(3738) <= not b;
    layer6_outputs(3739) <= b and not a;
    layer6_outputs(3740) <= not a or b;
    layer6_outputs(3741) <= not b;
    layer6_outputs(3742) <= not b;
    layer6_outputs(3743) <= a and not b;
    layer6_outputs(3744) <= b and not a;
    layer6_outputs(3745) <= a and not b;
    layer6_outputs(3746) <= a or b;
    layer6_outputs(3747) <= not b;
    layer6_outputs(3748) <= a;
    layer6_outputs(3749) <= a or b;
    layer6_outputs(3750) <= b;
    layer6_outputs(3751) <= a or b;
    layer6_outputs(3752) <= a xor b;
    layer6_outputs(3753) <= a;
    layer6_outputs(3754) <= a;
    layer6_outputs(3755) <= not b;
    layer6_outputs(3756) <= not b;
    layer6_outputs(3757) <= not a or b;
    layer6_outputs(3758) <= not b or a;
    layer6_outputs(3759) <= b;
    layer6_outputs(3760) <= not (a xor b);
    layer6_outputs(3761) <= not b;
    layer6_outputs(3762) <= a or b;
    layer6_outputs(3763) <= a xor b;
    layer6_outputs(3764) <= a and b;
    layer6_outputs(3765) <= not (a or b);
    layer6_outputs(3766) <= not b;
    layer6_outputs(3767) <= b;
    layer6_outputs(3768) <= not (a and b);
    layer6_outputs(3769) <= not a or b;
    layer6_outputs(3770) <= not b;
    layer6_outputs(3771) <= b and not a;
    layer6_outputs(3772) <= a and b;
    layer6_outputs(3773) <= a;
    layer6_outputs(3774) <= a and not b;
    layer6_outputs(3775) <= a and not b;
    layer6_outputs(3776) <= not b;
    layer6_outputs(3777) <= a xor b;
    layer6_outputs(3778) <= not b;
    layer6_outputs(3779) <= not (a and b);
    layer6_outputs(3780) <= b;
    layer6_outputs(3781) <= b;
    layer6_outputs(3782) <= b;
    layer6_outputs(3783) <= b;
    layer6_outputs(3784) <= not b or a;
    layer6_outputs(3785) <= not b or a;
    layer6_outputs(3786) <= 1'b1;
    layer6_outputs(3787) <= a and not b;
    layer6_outputs(3788) <= not a or b;
    layer6_outputs(3789) <= b;
    layer6_outputs(3790) <= b and not a;
    layer6_outputs(3791) <= b;
    layer6_outputs(3792) <= 1'b1;
    layer6_outputs(3793) <= a or b;
    layer6_outputs(3794) <= a xor b;
    layer6_outputs(3795) <= not a;
    layer6_outputs(3796) <= a and not b;
    layer6_outputs(3797) <= not b or a;
    layer6_outputs(3798) <= not b or a;
    layer6_outputs(3799) <= not a;
    layer6_outputs(3800) <= a xor b;
    layer6_outputs(3801) <= b and not a;
    layer6_outputs(3802) <= 1'b0;
    layer6_outputs(3803) <= not b or a;
    layer6_outputs(3804) <= b;
    layer6_outputs(3805) <= not b or a;
    layer6_outputs(3806) <= not a or b;
    layer6_outputs(3807) <= a;
    layer6_outputs(3808) <= a or b;
    layer6_outputs(3809) <= b;
    layer6_outputs(3810) <= not (a or b);
    layer6_outputs(3811) <= not (a or b);
    layer6_outputs(3812) <= not a;
    layer6_outputs(3813) <= a and b;
    layer6_outputs(3814) <= b;
    layer6_outputs(3815) <= 1'b1;
    layer6_outputs(3816) <= b;
    layer6_outputs(3817) <= not a;
    layer6_outputs(3818) <= a;
    layer6_outputs(3819) <= a;
    layer6_outputs(3820) <= not a;
    layer6_outputs(3821) <= a;
    layer6_outputs(3822) <= a and not b;
    layer6_outputs(3823) <= not b;
    layer6_outputs(3824) <= a and b;
    layer6_outputs(3825) <= b;
    layer6_outputs(3826) <= a;
    layer6_outputs(3827) <= a and b;
    layer6_outputs(3828) <= not b or a;
    layer6_outputs(3829) <= not (a or b);
    layer6_outputs(3830) <= b;
    layer6_outputs(3831) <= a;
    layer6_outputs(3832) <= not b or a;
    layer6_outputs(3833) <= not a;
    layer6_outputs(3834) <= b and not a;
    layer6_outputs(3835) <= a and b;
    layer6_outputs(3836) <= a and not b;
    layer6_outputs(3837) <= not (a or b);
    layer6_outputs(3838) <= a;
    layer6_outputs(3839) <= b;
    layer6_outputs(3840) <= a;
    layer6_outputs(3841) <= a and not b;
    layer6_outputs(3842) <= not b;
    layer6_outputs(3843) <= not b;
    layer6_outputs(3844) <= a and b;
    layer6_outputs(3845) <= not a;
    layer6_outputs(3846) <= not a;
    layer6_outputs(3847) <= a and not b;
    layer6_outputs(3848) <= a or b;
    layer6_outputs(3849) <= b and not a;
    layer6_outputs(3850) <= a;
    layer6_outputs(3851) <= a xor b;
    layer6_outputs(3852) <= a and b;
    layer6_outputs(3853) <= not b;
    layer6_outputs(3854) <= a xor b;
    layer6_outputs(3855) <= a and not b;
    layer6_outputs(3856) <= b;
    layer6_outputs(3857) <= a and b;
    layer6_outputs(3858) <= not (a xor b);
    layer6_outputs(3859) <= not b or a;
    layer6_outputs(3860) <= not b or a;
    layer6_outputs(3861) <= not b or a;
    layer6_outputs(3862) <= not (a and b);
    layer6_outputs(3863) <= not a;
    layer6_outputs(3864) <= not (a and b);
    layer6_outputs(3865) <= 1'b0;
    layer6_outputs(3866) <= a and b;
    layer6_outputs(3867) <= not (a xor b);
    layer6_outputs(3868) <= not b or a;
    layer6_outputs(3869) <= a;
    layer6_outputs(3870) <= b;
    layer6_outputs(3871) <= not (a or b);
    layer6_outputs(3872) <= not b;
    layer6_outputs(3873) <= not a or b;
    layer6_outputs(3874) <= not a;
    layer6_outputs(3875) <= not b or a;
    layer6_outputs(3876) <= b;
    layer6_outputs(3877) <= b;
    layer6_outputs(3878) <= not (a xor b);
    layer6_outputs(3879) <= not a;
    layer6_outputs(3880) <= not (a and b);
    layer6_outputs(3881) <= not b;
    layer6_outputs(3882) <= a and b;
    layer6_outputs(3883) <= a;
    layer6_outputs(3884) <= not b or a;
    layer6_outputs(3885) <= not b or a;
    layer6_outputs(3886) <= not a or b;
    layer6_outputs(3887) <= not b;
    layer6_outputs(3888) <= 1'b1;
    layer6_outputs(3889) <= not b;
    layer6_outputs(3890) <= not (a and b);
    layer6_outputs(3891) <= not b;
    layer6_outputs(3892) <= not b or a;
    layer6_outputs(3893) <= not a or b;
    layer6_outputs(3894) <= a and not b;
    layer6_outputs(3895) <= a;
    layer6_outputs(3896) <= a;
    layer6_outputs(3897) <= not a;
    layer6_outputs(3898) <= 1'b1;
    layer6_outputs(3899) <= not a;
    layer6_outputs(3900) <= a and b;
    layer6_outputs(3901) <= not (a xor b);
    layer6_outputs(3902) <= not a;
    layer6_outputs(3903) <= b;
    layer6_outputs(3904) <= a or b;
    layer6_outputs(3905) <= a and b;
    layer6_outputs(3906) <= b;
    layer6_outputs(3907) <= a;
    layer6_outputs(3908) <= not b;
    layer6_outputs(3909) <= a or b;
    layer6_outputs(3910) <= not a;
    layer6_outputs(3911) <= not b;
    layer6_outputs(3912) <= not a or b;
    layer6_outputs(3913) <= not (a xor b);
    layer6_outputs(3914) <= 1'b0;
    layer6_outputs(3915) <= not a;
    layer6_outputs(3916) <= not a or b;
    layer6_outputs(3917) <= not a;
    layer6_outputs(3918) <= not (a and b);
    layer6_outputs(3919) <= b and not a;
    layer6_outputs(3920) <= b;
    layer6_outputs(3921) <= b;
    layer6_outputs(3922) <= a xor b;
    layer6_outputs(3923) <= not a or b;
    layer6_outputs(3924) <= a;
    layer6_outputs(3925) <= a or b;
    layer6_outputs(3926) <= 1'b0;
    layer6_outputs(3927) <= a or b;
    layer6_outputs(3928) <= not (a and b);
    layer6_outputs(3929) <= a;
    layer6_outputs(3930) <= not a or b;
    layer6_outputs(3931) <= not a or b;
    layer6_outputs(3932) <= not (a or b);
    layer6_outputs(3933) <= not (a or b);
    layer6_outputs(3934) <= b;
    layer6_outputs(3935) <= a and not b;
    layer6_outputs(3936) <= not b;
    layer6_outputs(3937) <= not (a and b);
    layer6_outputs(3938) <= a and b;
    layer6_outputs(3939) <= a and not b;
    layer6_outputs(3940) <= b;
    layer6_outputs(3941) <= not b;
    layer6_outputs(3942) <= b;
    layer6_outputs(3943) <= b and not a;
    layer6_outputs(3944) <= b and not a;
    layer6_outputs(3945) <= not b;
    layer6_outputs(3946) <= 1'b0;
    layer6_outputs(3947) <= b;
    layer6_outputs(3948) <= not (a xor b);
    layer6_outputs(3949) <= not a;
    layer6_outputs(3950) <= a and not b;
    layer6_outputs(3951) <= b;
    layer6_outputs(3952) <= a;
    layer6_outputs(3953) <= not (a or b);
    layer6_outputs(3954) <= b and not a;
    layer6_outputs(3955) <= a and not b;
    layer6_outputs(3956) <= not a or b;
    layer6_outputs(3957) <= a xor b;
    layer6_outputs(3958) <= not b;
    layer6_outputs(3959) <= b and not a;
    layer6_outputs(3960) <= not b or a;
    layer6_outputs(3961) <= b;
    layer6_outputs(3962) <= a;
    layer6_outputs(3963) <= not a;
    layer6_outputs(3964) <= a and not b;
    layer6_outputs(3965) <= not b;
    layer6_outputs(3966) <= a and not b;
    layer6_outputs(3967) <= a xor b;
    layer6_outputs(3968) <= b;
    layer6_outputs(3969) <= a xor b;
    layer6_outputs(3970) <= b;
    layer6_outputs(3971) <= not a or b;
    layer6_outputs(3972) <= b and not a;
    layer6_outputs(3973) <= a and b;
    layer6_outputs(3974) <= a or b;
    layer6_outputs(3975) <= not (a and b);
    layer6_outputs(3976) <= 1'b1;
    layer6_outputs(3977) <= not (a or b);
    layer6_outputs(3978) <= not (a xor b);
    layer6_outputs(3979) <= b and not a;
    layer6_outputs(3980) <= b;
    layer6_outputs(3981) <= not a;
    layer6_outputs(3982) <= a and b;
    layer6_outputs(3983) <= a;
    layer6_outputs(3984) <= not b or a;
    layer6_outputs(3985) <= a xor b;
    layer6_outputs(3986) <= b;
    layer6_outputs(3987) <= not (a or b);
    layer6_outputs(3988) <= not a;
    layer6_outputs(3989) <= a and not b;
    layer6_outputs(3990) <= not (a or b);
    layer6_outputs(3991) <= 1'b1;
    layer6_outputs(3992) <= not b;
    layer6_outputs(3993) <= a xor b;
    layer6_outputs(3994) <= not a or b;
    layer6_outputs(3995) <= not b;
    layer6_outputs(3996) <= not a;
    layer6_outputs(3997) <= not (a xor b);
    layer6_outputs(3998) <= not (a xor b);
    layer6_outputs(3999) <= not (a or b);
    layer6_outputs(4000) <= b and not a;
    layer6_outputs(4001) <= not a;
    layer6_outputs(4002) <= not a or b;
    layer6_outputs(4003) <= not a or b;
    layer6_outputs(4004) <= 1'b1;
    layer6_outputs(4005) <= not a;
    layer6_outputs(4006) <= b;
    layer6_outputs(4007) <= not b;
    layer6_outputs(4008) <= not (a and b);
    layer6_outputs(4009) <= a;
    layer6_outputs(4010) <= not a;
    layer6_outputs(4011) <= not (a xor b);
    layer6_outputs(4012) <= a;
    layer6_outputs(4013) <= b;
    layer6_outputs(4014) <= not a or b;
    layer6_outputs(4015) <= b and not a;
    layer6_outputs(4016) <= not a;
    layer6_outputs(4017) <= not b;
    layer6_outputs(4018) <= a or b;
    layer6_outputs(4019) <= a and b;
    layer6_outputs(4020) <= 1'b0;
    layer6_outputs(4021) <= not a;
    layer6_outputs(4022) <= a or b;
    layer6_outputs(4023) <= b and not a;
    layer6_outputs(4024) <= not (a and b);
    layer6_outputs(4025) <= 1'b0;
    layer6_outputs(4026) <= not (a xor b);
    layer6_outputs(4027) <= not (a xor b);
    layer6_outputs(4028) <= a and not b;
    layer6_outputs(4029) <= a;
    layer6_outputs(4030) <= a or b;
    layer6_outputs(4031) <= not (a xor b);
    layer6_outputs(4032) <= not a;
    layer6_outputs(4033) <= a and not b;
    layer6_outputs(4034) <= not b or a;
    layer6_outputs(4035) <= not b or a;
    layer6_outputs(4036) <= not a;
    layer6_outputs(4037) <= a;
    layer6_outputs(4038) <= a and b;
    layer6_outputs(4039) <= a;
    layer6_outputs(4040) <= not b or a;
    layer6_outputs(4041) <= b;
    layer6_outputs(4042) <= not a or b;
    layer6_outputs(4043) <= b and not a;
    layer6_outputs(4044) <= not a or b;
    layer6_outputs(4045) <= a and not b;
    layer6_outputs(4046) <= a xor b;
    layer6_outputs(4047) <= not (a or b);
    layer6_outputs(4048) <= b;
    layer6_outputs(4049) <= not b or a;
    layer6_outputs(4050) <= not a;
    layer6_outputs(4051) <= not b;
    layer6_outputs(4052) <= a and b;
    layer6_outputs(4053) <= not a or b;
    layer6_outputs(4054) <= a;
    layer6_outputs(4055) <= not b or a;
    layer6_outputs(4056) <= not (a and b);
    layer6_outputs(4057) <= not b;
    layer6_outputs(4058) <= a and b;
    layer6_outputs(4059) <= a and not b;
    layer6_outputs(4060) <= not a;
    layer6_outputs(4061) <= not (a and b);
    layer6_outputs(4062) <= not b;
    layer6_outputs(4063) <= b;
    layer6_outputs(4064) <= not a;
    layer6_outputs(4065) <= not a;
    layer6_outputs(4066) <= 1'b1;
    layer6_outputs(4067) <= not a;
    layer6_outputs(4068) <= not a or b;
    layer6_outputs(4069) <= a;
    layer6_outputs(4070) <= a xor b;
    layer6_outputs(4071) <= not a or b;
    layer6_outputs(4072) <= not a;
    layer6_outputs(4073) <= not a or b;
    layer6_outputs(4074) <= a;
    layer6_outputs(4075) <= a or b;
    layer6_outputs(4076) <= b;
    layer6_outputs(4077) <= not b or a;
    layer6_outputs(4078) <= not b;
    layer6_outputs(4079) <= a or b;
    layer6_outputs(4080) <= not b;
    layer6_outputs(4081) <= not a or b;
    layer6_outputs(4082) <= a or b;
    layer6_outputs(4083) <= a and not b;
    layer6_outputs(4084) <= b and not a;
    layer6_outputs(4085) <= not (a xor b);
    layer6_outputs(4086) <= not a;
    layer6_outputs(4087) <= not a;
    layer6_outputs(4088) <= a;
    layer6_outputs(4089) <= not b or a;
    layer6_outputs(4090) <= not a;
    layer6_outputs(4091) <= b;
    layer6_outputs(4092) <= not b or a;
    layer6_outputs(4093) <= 1'b0;
    layer6_outputs(4094) <= a;
    layer6_outputs(4095) <= not b;
    layer6_outputs(4096) <= not b;
    layer6_outputs(4097) <= a xor b;
    layer6_outputs(4098) <= a and not b;
    layer6_outputs(4099) <= a and b;
    layer6_outputs(4100) <= not a or b;
    layer6_outputs(4101) <= 1'b0;
    layer6_outputs(4102) <= not a;
    layer6_outputs(4103) <= b and not a;
    layer6_outputs(4104) <= not a or b;
    layer6_outputs(4105) <= a xor b;
    layer6_outputs(4106) <= a xor b;
    layer6_outputs(4107) <= not a or b;
    layer6_outputs(4108) <= not (a and b);
    layer6_outputs(4109) <= a xor b;
    layer6_outputs(4110) <= a;
    layer6_outputs(4111) <= not b;
    layer6_outputs(4112) <= a;
    layer6_outputs(4113) <= 1'b1;
    layer6_outputs(4114) <= not b;
    layer6_outputs(4115) <= 1'b1;
    layer6_outputs(4116) <= not (a xor b);
    layer6_outputs(4117) <= 1'b1;
    layer6_outputs(4118) <= not b;
    layer6_outputs(4119) <= not (a or b);
    layer6_outputs(4120) <= a;
    layer6_outputs(4121) <= a;
    layer6_outputs(4122) <= not a;
    layer6_outputs(4123) <= not (a or b);
    layer6_outputs(4124) <= not b or a;
    layer6_outputs(4125) <= a xor b;
    layer6_outputs(4126) <= not b;
    layer6_outputs(4127) <= not (a xor b);
    layer6_outputs(4128) <= b;
    layer6_outputs(4129) <= a xor b;
    layer6_outputs(4130) <= b;
    layer6_outputs(4131) <= not b;
    layer6_outputs(4132) <= 1'b1;
    layer6_outputs(4133) <= not a;
    layer6_outputs(4134) <= b;
    layer6_outputs(4135) <= a or b;
    layer6_outputs(4136) <= not b or a;
    layer6_outputs(4137) <= not a;
    layer6_outputs(4138) <= a;
    layer6_outputs(4139) <= 1'b1;
    layer6_outputs(4140) <= a;
    layer6_outputs(4141) <= not b;
    layer6_outputs(4142) <= not a or b;
    layer6_outputs(4143) <= not (a xor b);
    layer6_outputs(4144) <= b;
    layer6_outputs(4145) <= not a;
    layer6_outputs(4146) <= a xor b;
    layer6_outputs(4147) <= b;
    layer6_outputs(4148) <= a and not b;
    layer6_outputs(4149) <= not a or b;
    layer6_outputs(4150) <= b;
    layer6_outputs(4151) <= a and b;
    layer6_outputs(4152) <= a and not b;
    layer6_outputs(4153) <= not b;
    layer6_outputs(4154) <= b;
    layer6_outputs(4155) <= a xor b;
    layer6_outputs(4156) <= b and not a;
    layer6_outputs(4157) <= a or b;
    layer6_outputs(4158) <= b and not a;
    layer6_outputs(4159) <= 1'b0;
    layer6_outputs(4160) <= b and not a;
    layer6_outputs(4161) <= a;
    layer6_outputs(4162) <= not (a and b);
    layer6_outputs(4163) <= not a or b;
    layer6_outputs(4164) <= b and not a;
    layer6_outputs(4165) <= not a;
    layer6_outputs(4166) <= not (a xor b);
    layer6_outputs(4167) <= 1'b1;
    layer6_outputs(4168) <= a and b;
    layer6_outputs(4169) <= a and b;
    layer6_outputs(4170) <= a and not b;
    layer6_outputs(4171) <= a or b;
    layer6_outputs(4172) <= not (a xor b);
    layer6_outputs(4173) <= not a;
    layer6_outputs(4174) <= 1'b1;
    layer6_outputs(4175) <= a xor b;
    layer6_outputs(4176) <= a;
    layer6_outputs(4177) <= not a;
    layer6_outputs(4178) <= a xor b;
    layer6_outputs(4179) <= a and not b;
    layer6_outputs(4180) <= b;
    layer6_outputs(4181) <= a or b;
    layer6_outputs(4182) <= a and not b;
    layer6_outputs(4183) <= not b;
    layer6_outputs(4184) <= a;
    layer6_outputs(4185) <= b;
    layer6_outputs(4186) <= a and b;
    layer6_outputs(4187) <= not (a and b);
    layer6_outputs(4188) <= b;
    layer6_outputs(4189) <= not b;
    layer6_outputs(4190) <= a and not b;
    layer6_outputs(4191) <= b and not a;
    layer6_outputs(4192) <= a and not b;
    layer6_outputs(4193) <= a and b;
    layer6_outputs(4194) <= 1'b0;
    layer6_outputs(4195) <= a and not b;
    layer6_outputs(4196) <= not b;
    layer6_outputs(4197) <= not a;
    layer6_outputs(4198) <= a and b;
    layer6_outputs(4199) <= not a;
    layer6_outputs(4200) <= a xor b;
    layer6_outputs(4201) <= a and b;
    layer6_outputs(4202) <= not a or b;
    layer6_outputs(4203) <= b;
    layer6_outputs(4204) <= not a;
    layer6_outputs(4205) <= a and not b;
    layer6_outputs(4206) <= b;
    layer6_outputs(4207) <= not (a and b);
    layer6_outputs(4208) <= b;
    layer6_outputs(4209) <= a xor b;
    layer6_outputs(4210) <= not b or a;
    layer6_outputs(4211) <= not (a and b);
    layer6_outputs(4212) <= a and b;
    layer6_outputs(4213) <= b;
    layer6_outputs(4214) <= a or b;
    layer6_outputs(4215) <= a and b;
    layer6_outputs(4216) <= b;
    layer6_outputs(4217) <= a xor b;
    layer6_outputs(4218) <= a;
    layer6_outputs(4219) <= not b;
    layer6_outputs(4220) <= not a;
    layer6_outputs(4221) <= a;
    layer6_outputs(4222) <= a and b;
    layer6_outputs(4223) <= b;
    layer6_outputs(4224) <= not a;
    layer6_outputs(4225) <= not b;
    layer6_outputs(4226) <= b;
    layer6_outputs(4227) <= a;
    layer6_outputs(4228) <= not a or b;
    layer6_outputs(4229) <= a xor b;
    layer6_outputs(4230) <= not b;
    layer6_outputs(4231) <= a and not b;
    layer6_outputs(4232) <= not b;
    layer6_outputs(4233) <= not (a or b);
    layer6_outputs(4234) <= b;
    layer6_outputs(4235) <= a xor b;
    layer6_outputs(4236) <= b;
    layer6_outputs(4237) <= a;
    layer6_outputs(4238) <= a and not b;
    layer6_outputs(4239) <= b and not a;
    layer6_outputs(4240) <= b;
    layer6_outputs(4241) <= a xor b;
    layer6_outputs(4242) <= a and not b;
    layer6_outputs(4243) <= not b;
    layer6_outputs(4244) <= b;
    layer6_outputs(4245) <= a;
    layer6_outputs(4246) <= a xor b;
    layer6_outputs(4247) <= a;
    layer6_outputs(4248) <= not a;
    layer6_outputs(4249) <= not a;
    layer6_outputs(4250) <= not a;
    layer6_outputs(4251) <= a and b;
    layer6_outputs(4252) <= a;
    layer6_outputs(4253) <= a or b;
    layer6_outputs(4254) <= not a;
    layer6_outputs(4255) <= a;
    layer6_outputs(4256) <= a;
    layer6_outputs(4257) <= a;
    layer6_outputs(4258) <= not b;
    layer6_outputs(4259) <= a and not b;
    layer6_outputs(4260) <= 1'b1;
    layer6_outputs(4261) <= not a;
    layer6_outputs(4262) <= a and b;
    layer6_outputs(4263) <= 1'b1;
    layer6_outputs(4264) <= 1'b1;
    layer6_outputs(4265) <= a and not b;
    layer6_outputs(4266) <= a or b;
    layer6_outputs(4267) <= a;
    layer6_outputs(4268) <= a xor b;
    layer6_outputs(4269) <= not (a or b);
    layer6_outputs(4270) <= a and b;
    layer6_outputs(4271) <= not (a xor b);
    layer6_outputs(4272) <= 1'b0;
    layer6_outputs(4273) <= not a;
    layer6_outputs(4274) <= b and not a;
    layer6_outputs(4275) <= not a or b;
    layer6_outputs(4276) <= a and not b;
    layer6_outputs(4277) <= a xor b;
    layer6_outputs(4278) <= a and not b;
    layer6_outputs(4279) <= not b;
    layer6_outputs(4280) <= not (a and b);
    layer6_outputs(4281) <= not (a or b);
    layer6_outputs(4282) <= not a or b;
    layer6_outputs(4283) <= not b or a;
    layer6_outputs(4284) <= b and not a;
    layer6_outputs(4285) <= not b;
    layer6_outputs(4286) <= a or b;
    layer6_outputs(4287) <= not a;
    layer6_outputs(4288) <= 1'b0;
    layer6_outputs(4289) <= b;
    layer6_outputs(4290) <= not b or a;
    layer6_outputs(4291) <= not (a xor b);
    layer6_outputs(4292) <= not a or b;
    layer6_outputs(4293) <= not a;
    layer6_outputs(4294) <= not (a xor b);
    layer6_outputs(4295) <= not (a and b);
    layer6_outputs(4296) <= not (a and b);
    layer6_outputs(4297) <= a xor b;
    layer6_outputs(4298) <= a or b;
    layer6_outputs(4299) <= not b or a;
    layer6_outputs(4300) <= not (a or b);
    layer6_outputs(4301) <= a and not b;
    layer6_outputs(4302) <= b;
    layer6_outputs(4303) <= not b;
    layer6_outputs(4304) <= not a or b;
    layer6_outputs(4305) <= not a;
    layer6_outputs(4306) <= b and not a;
    layer6_outputs(4307) <= a and not b;
    layer6_outputs(4308) <= not a or b;
    layer6_outputs(4309) <= a or b;
    layer6_outputs(4310) <= b;
    layer6_outputs(4311) <= not (a xor b);
    layer6_outputs(4312) <= not a;
    layer6_outputs(4313) <= a or b;
    layer6_outputs(4314) <= a or b;
    layer6_outputs(4315) <= a and b;
    layer6_outputs(4316) <= not b;
    layer6_outputs(4317) <= a and not b;
    layer6_outputs(4318) <= not b or a;
    layer6_outputs(4319) <= b;
    layer6_outputs(4320) <= a and b;
    layer6_outputs(4321) <= b;
    layer6_outputs(4322) <= not a;
    layer6_outputs(4323) <= a and not b;
    layer6_outputs(4324) <= not a or b;
    layer6_outputs(4325) <= b;
    layer6_outputs(4326) <= not a or b;
    layer6_outputs(4327) <= b;
    layer6_outputs(4328) <= a;
    layer6_outputs(4329) <= not a or b;
    layer6_outputs(4330) <= not a or b;
    layer6_outputs(4331) <= a or b;
    layer6_outputs(4332) <= b;
    layer6_outputs(4333) <= not a;
    layer6_outputs(4334) <= 1'b0;
    layer6_outputs(4335) <= a;
    layer6_outputs(4336) <= not a;
    layer6_outputs(4337) <= not (a xor b);
    layer6_outputs(4338) <= a;
    layer6_outputs(4339) <= a;
    layer6_outputs(4340) <= not (a and b);
    layer6_outputs(4341) <= not a or b;
    layer6_outputs(4342) <= not (a or b);
    layer6_outputs(4343) <= not a;
    layer6_outputs(4344) <= not b;
    layer6_outputs(4345) <= b;
    layer6_outputs(4346) <= not a or b;
    layer6_outputs(4347) <= a;
    layer6_outputs(4348) <= not (a or b);
    layer6_outputs(4349) <= a xor b;
    layer6_outputs(4350) <= not a;
    layer6_outputs(4351) <= not a;
    layer6_outputs(4352) <= b;
    layer6_outputs(4353) <= not (a or b);
    layer6_outputs(4354) <= a and b;
    layer6_outputs(4355) <= b and not a;
    layer6_outputs(4356) <= b;
    layer6_outputs(4357) <= b and not a;
    layer6_outputs(4358) <= a;
    layer6_outputs(4359) <= b;
    layer6_outputs(4360) <= a and not b;
    layer6_outputs(4361) <= a xor b;
    layer6_outputs(4362) <= not (a and b);
    layer6_outputs(4363) <= not a or b;
    layer6_outputs(4364) <= b;
    layer6_outputs(4365) <= not (a or b);
    layer6_outputs(4366) <= not b;
    layer6_outputs(4367) <= b;
    layer6_outputs(4368) <= a and not b;
    layer6_outputs(4369) <= not b or a;
    layer6_outputs(4370) <= a and not b;
    layer6_outputs(4371) <= a;
    layer6_outputs(4372) <= a and not b;
    layer6_outputs(4373) <= not b or a;
    layer6_outputs(4374) <= a or b;
    layer6_outputs(4375) <= 1'b1;
    layer6_outputs(4376) <= not a;
    layer6_outputs(4377) <= not (a or b);
    layer6_outputs(4378) <= 1'b0;
    layer6_outputs(4379) <= not (a and b);
    layer6_outputs(4380) <= b;
    layer6_outputs(4381) <= not b or a;
    layer6_outputs(4382) <= b and not a;
    layer6_outputs(4383) <= not (a xor b);
    layer6_outputs(4384) <= not (a xor b);
    layer6_outputs(4385) <= a or b;
    layer6_outputs(4386) <= not (a and b);
    layer6_outputs(4387) <= a or b;
    layer6_outputs(4388) <= a;
    layer6_outputs(4389) <= not a or b;
    layer6_outputs(4390) <= b and not a;
    layer6_outputs(4391) <= not (a or b);
    layer6_outputs(4392) <= not b;
    layer6_outputs(4393) <= not (a or b);
    layer6_outputs(4394) <= a and not b;
    layer6_outputs(4395) <= not b;
    layer6_outputs(4396) <= a xor b;
    layer6_outputs(4397) <= not a;
    layer6_outputs(4398) <= a;
    layer6_outputs(4399) <= not a;
    layer6_outputs(4400) <= a xor b;
    layer6_outputs(4401) <= a and not b;
    layer6_outputs(4402) <= a or b;
    layer6_outputs(4403) <= not b or a;
    layer6_outputs(4404) <= not a;
    layer6_outputs(4405) <= a and not b;
    layer6_outputs(4406) <= a and b;
    layer6_outputs(4407) <= not b or a;
    layer6_outputs(4408) <= not (a and b);
    layer6_outputs(4409) <= not b;
    layer6_outputs(4410) <= b;
    layer6_outputs(4411) <= b;
    layer6_outputs(4412) <= not (a xor b);
    layer6_outputs(4413) <= a;
    layer6_outputs(4414) <= not (a and b);
    layer6_outputs(4415) <= a;
    layer6_outputs(4416) <= b;
    layer6_outputs(4417) <= a;
    layer6_outputs(4418) <= a or b;
    layer6_outputs(4419) <= not b or a;
    layer6_outputs(4420) <= not b or a;
    layer6_outputs(4421) <= not a;
    layer6_outputs(4422) <= not b;
    layer6_outputs(4423) <= b;
    layer6_outputs(4424) <= not (a or b);
    layer6_outputs(4425) <= a and not b;
    layer6_outputs(4426) <= not a or b;
    layer6_outputs(4427) <= a or b;
    layer6_outputs(4428) <= a;
    layer6_outputs(4429) <= a;
    layer6_outputs(4430) <= not a;
    layer6_outputs(4431) <= not b;
    layer6_outputs(4432) <= a and b;
    layer6_outputs(4433) <= not (a xor b);
    layer6_outputs(4434) <= not (a and b);
    layer6_outputs(4435) <= a;
    layer6_outputs(4436) <= 1'b0;
    layer6_outputs(4437) <= b;
    layer6_outputs(4438) <= a;
    layer6_outputs(4439) <= b and not a;
    layer6_outputs(4440) <= a;
    layer6_outputs(4441) <= a and b;
    layer6_outputs(4442) <= not (a or b);
    layer6_outputs(4443) <= a and b;
    layer6_outputs(4444) <= not b;
    layer6_outputs(4445) <= not a or b;
    layer6_outputs(4446) <= b;
    layer6_outputs(4447) <= a xor b;
    layer6_outputs(4448) <= b;
    layer6_outputs(4449) <= not (a or b);
    layer6_outputs(4450) <= not b;
    layer6_outputs(4451) <= 1'b1;
    layer6_outputs(4452) <= b and not a;
    layer6_outputs(4453) <= 1'b1;
    layer6_outputs(4454) <= a;
    layer6_outputs(4455) <= not b;
    layer6_outputs(4456) <= not a;
    layer6_outputs(4457) <= a xor b;
    layer6_outputs(4458) <= 1'b0;
    layer6_outputs(4459) <= a xor b;
    layer6_outputs(4460) <= a;
    layer6_outputs(4461) <= not b or a;
    layer6_outputs(4462) <= a and not b;
    layer6_outputs(4463) <= b;
    layer6_outputs(4464) <= not (a xor b);
    layer6_outputs(4465) <= b;
    layer6_outputs(4466) <= b;
    layer6_outputs(4467) <= not b or a;
    layer6_outputs(4468) <= not (a xor b);
    layer6_outputs(4469) <= a and not b;
    layer6_outputs(4470) <= a and b;
    layer6_outputs(4471) <= not b;
    layer6_outputs(4472) <= not b;
    layer6_outputs(4473) <= not b;
    layer6_outputs(4474) <= a;
    layer6_outputs(4475) <= not (a xor b);
    layer6_outputs(4476) <= not a;
    layer6_outputs(4477) <= not (a xor b);
    layer6_outputs(4478) <= b;
    layer6_outputs(4479) <= not b;
    layer6_outputs(4480) <= b and not a;
    layer6_outputs(4481) <= not b;
    layer6_outputs(4482) <= not (a or b);
    layer6_outputs(4483) <= a and b;
    layer6_outputs(4484) <= not a or b;
    layer6_outputs(4485) <= not b or a;
    layer6_outputs(4486) <= not (a and b);
    layer6_outputs(4487) <= not a;
    layer6_outputs(4488) <= a and not b;
    layer6_outputs(4489) <= not b;
    layer6_outputs(4490) <= not (a xor b);
    layer6_outputs(4491) <= not (a or b);
    layer6_outputs(4492) <= a;
    layer6_outputs(4493) <= a xor b;
    layer6_outputs(4494) <= not a;
    layer6_outputs(4495) <= a;
    layer6_outputs(4496) <= not a;
    layer6_outputs(4497) <= not (a xor b);
    layer6_outputs(4498) <= b and not a;
    layer6_outputs(4499) <= not (a or b);
    layer6_outputs(4500) <= 1'b1;
    layer6_outputs(4501) <= not b;
    layer6_outputs(4502) <= a;
    layer6_outputs(4503) <= 1'b1;
    layer6_outputs(4504) <= a and b;
    layer6_outputs(4505) <= 1'b1;
    layer6_outputs(4506) <= not a;
    layer6_outputs(4507) <= not a;
    layer6_outputs(4508) <= not (a xor b);
    layer6_outputs(4509) <= b;
    layer6_outputs(4510) <= a;
    layer6_outputs(4511) <= a and b;
    layer6_outputs(4512) <= a or b;
    layer6_outputs(4513) <= b and not a;
    layer6_outputs(4514) <= not a or b;
    layer6_outputs(4515) <= not (a and b);
    layer6_outputs(4516) <= b and not a;
    layer6_outputs(4517) <= a or b;
    layer6_outputs(4518) <= not a;
    layer6_outputs(4519) <= a and b;
    layer6_outputs(4520) <= a and not b;
    layer6_outputs(4521) <= a and b;
    layer6_outputs(4522) <= not a;
    layer6_outputs(4523) <= a xor b;
    layer6_outputs(4524) <= b and not a;
    layer6_outputs(4525) <= not (a and b);
    layer6_outputs(4526) <= not (a or b);
    layer6_outputs(4527) <= not a or b;
    layer6_outputs(4528) <= not (a and b);
    layer6_outputs(4529) <= not (a xor b);
    layer6_outputs(4530) <= b;
    layer6_outputs(4531) <= not a;
    layer6_outputs(4532) <= not a;
    layer6_outputs(4533) <= not a;
    layer6_outputs(4534) <= a xor b;
    layer6_outputs(4535) <= a and not b;
    layer6_outputs(4536) <= not b;
    layer6_outputs(4537) <= b;
    layer6_outputs(4538) <= not (a and b);
    layer6_outputs(4539) <= not (a and b);
    layer6_outputs(4540) <= a xor b;
    layer6_outputs(4541) <= not b;
    layer6_outputs(4542) <= a;
    layer6_outputs(4543) <= a;
    layer6_outputs(4544) <= a;
    layer6_outputs(4545) <= a or b;
    layer6_outputs(4546) <= not a or b;
    layer6_outputs(4547) <= b;
    layer6_outputs(4548) <= 1'b0;
    layer6_outputs(4549) <= a xor b;
    layer6_outputs(4550) <= a and not b;
    layer6_outputs(4551) <= not (a or b);
    layer6_outputs(4552) <= b and not a;
    layer6_outputs(4553) <= not a;
    layer6_outputs(4554) <= a and not b;
    layer6_outputs(4555) <= not b;
    layer6_outputs(4556) <= a;
    layer6_outputs(4557) <= a;
    layer6_outputs(4558) <= a;
    layer6_outputs(4559) <= not b;
    layer6_outputs(4560) <= a xor b;
    layer6_outputs(4561) <= not a;
    layer6_outputs(4562) <= not a;
    layer6_outputs(4563) <= not b;
    layer6_outputs(4564) <= b;
    layer6_outputs(4565) <= not b;
    layer6_outputs(4566) <= 1'b1;
    layer6_outputs(4567) <= not (a and b);
    layer6_outputs(4568) <= not b;
    layer6_outputs(4569) <= not a or b;
    layer6_outputs(4570) <= 1'b0;
    layer6_outputs(4571) <= not b or a;
    layer6_outputs(4572) <= b;
    layer6_outputs(4573) <= not b;
    layer6_outputs(4574) <= a;
    layer6_outputs(4575) <= a;
    layer6_outputs(4576) <= not (a xor b);
    layer6_outputs(4577) <= a and b;
    layer6_outputs(4578) <= not a;
    layer6_outputs(4579) <= not (a xor b);
    layer6_outputs(4580) <= b and not a;
    layer6_outputs(4581) <= a and not b;
    layer6_outputs(4582) <= not a;
    layer6_outputs(4583) <= not b;
    layer6_outputs(4584) <= not a or b;
    layer6_outputs(4585) <= b;
    layer6_outputs(4586) <= not b;
    layer6_outputs(4587) <= not (a and b);
    layer6_outputs(4588) <= not (a and b);
    layer6_outputs(4589) <= a or b;
    layer6_outputs(4590) <= a;
    layer6_outputs(4591) <= not b;
    layer6_outputs(4592) <= a or b;
    layer6_outputs(4593) <= a xor b;
    layer6_outputs(4594) <= b;
    layer6_outputs(4595) <= a and not b;
    layer6_outputs(4596) <= not a or b;
    layer6_outputs(4597) <= not (a and b);
    layer6_outputs(4598) <= a;
    layer6_outputs(4599) <= a and b;
    layer6_outputs(4600) <= b;
    layer6_outputs(4601) <= a or b;
    layer6_outputs(4602) <= a;
    layer6_outputs(4603) <= not (a and b);
    layer6_outputs(4604) <= b;
    layer6_outputs(4605) <= not a;
    layer6_outputs(4606) <= b;
    layer6_outputs(4607) <= not (a and b);
    layer6_outputs(4608) <= not (a xor b);
    layer6_outputs(4609) <= a or b;
    layer6_outputs(4610) <= not (a or b);
    layer6_outputs(4611) <= a or b;
    layer6_outputs(4612) <= not a or b;
    layer6_outputs(4613) <= not b or a;
    layer6_outputs(4614) <= not b or a;
    layer6_outputs(4615) <= a;
    layer6_outputs(4616) <= b and not a;
    layer6_outputs(4617) <= a or b;
    layer6_outputs(4618) <= not a or b;
    layer6_outputs(4619) <= not (a xor b);
    layer6_outputs(4620) <= not a or b;
    layer6_outputs(4621) <= a;
    layer6_outputs(4622) <= not (a or b);
    layer6_outputs(4623) <= not (a xor b);
    layer6_outputs(4624) <= not (a xor b);
    layer6_outputs(4625) <= not a;
    layer6_outputs(4626) <= b;
    layer6_outputs(4627) <= 1'b1;
    layer6_outputs(4628) <= not b or a;
    layer6_outputs(4629) <= 1'b1;
    layer6_outputs(4630) <= not b;
    layer6_outputs(4631) <= not b or a;
    layer6_outputs(4632) <= not a;
    layer6_outputs(4633) <= 1'b0;
    layer6_outputs(4634) <= a xor b;
    layer6_outputs(4635) <= b and not a;
    layer6_outputs(4636) <= not (a xor b);
    layer6_outputs(4637) <= b;
    layer6_outputs(4638) <= not b or a;
    layer6_outputs(4639) <= b and not a;
    layer6_outputs(4640) <= not a or b;
    layer6_outputs(4641) <= a;
    layer6_outputs(4642) <= not b;
    layer6_outputs(4643) <= a or b;
    layer6_outputs(4644) <= not a or b;
    layer6_outputs(4645) <= not b;
    layer6_outputs(4646) <= a and not b;
    layer6_outputs(4647) <= b and not a;
    layer6_outputs(4648) <= not (a or b);
    layer6_outputs(4649) <= not (a and b);
    layer6_outputs(4650) <= 1'b1;
    layer6_outputs(4651) <= not b or a;
    layer6_outputs(4652) <= a or b;
    layer6_outputs(4653) <= not a;
    layer6_outputs(4654) <= a and not b;
    layer6_outputs(4655) <= not b;
    layer6_outputs(4656) <= not (a and b);
    layer6_outputs(4657) <= a and b;
    layer6_outputs(4658) <= a;
    layer6_outputs(4659) <= a and not b;
    layer6_outputs(4660) <= not (a xor b);
    layer6_outputs(4661) <= a and not b;
    layer6_outputs(4662) <= not b;
    layer6_outputs(4663) <= not a;
    layer6_outputs(4664) <= not (a xor b);
    layer6_outputs(4665) <= not b or a;
    layer6_outputs(4666) <= not (a and b);
    layer6_outputs(4667) <= a;
    layer6_outputs(4668) <= not b;
    layer6_outputs(4669) <= a or b;
    layer6_outputs(4670) <= a;
    layer6_outputs(4671) <= not b or a;
    layer6_outputs(4672) <= b;
    layer6_outputs(4673) <= not (a or b);
    layer6_outputs(4674) <= a and not b;
    layer6_outputs(4675) <= b;
    layer6_outputs(4676) <= b;
    layer6_outputs(4677) <= b;
    layer6_outputs(4678) <= not b;
    layer6_outputs(4679) <= a xor b;
    layer6_outputs(4680) <= b and not a;
    layer6_outputs(4681) <= not (a or b);
    layer6_outputs(4682) <= not b;
    layer6_outputs(4683) <= not b;
    layer6_outputs(4684) <= a and not b;
    layer6_outputs(4685) <= a;
    layer6_outputs(4686) <= a and not b;
    layer6_outputs(4687) <= not a or b;
    layer6_outputs(4688) <= a and not b;
    layer6_outputs(4689) <= not a or b;
    layer6_outputs(4690) <= a and b;
    layer6_outputs(4691) <= a and not b;
    layer6_outputs(4692) <= not a;
    layer6_outputs(4693) <= a xor b;
    layer6_outputs(4694) <= a and b;
    layer6_outputs(4695) <= not (a and b);
    layer6_outputs(4696) <= a;
    layer6_outputs(4697) <= not a or b;
    layer6_outputs(4698) <= a;
    layer6_outputs(4699) <= b and not a;
    layer6_outputs(4700) <= not a or b;
    layer6_outputs(4701) <= not (a and b);
    layer6_outputs(4702) <= b and not a;
    layer6_outputs(4703) <= not b;
    layer6_outputs(4704) <= a and not b;
    layer6_outputs(4705) <= a;
    layer6_outputs(4706) <= 1'b0;
    layer6_outputs(4707) <= not (a and b);
    layer6_outputs(4708) <= a or b;
    layer6_outputs(4709) <= a;
    layer6_outputs(4710) <= a;
    layer6_outputs(4711) <= a;
    layer6_outputs(4712) <= b and not a;
    layer6_outputs(4713) <= not a or b;
    layer6_outputs(4714) <= b;
    layer6_outputs(4715) <= b;
    layer6_outputs(4716) <= not (a and b);
    layer6_outputs(4717) <= not a or b;
    layer6_outputs(4718) <= not (a and b);
    layer6_outputs(4719) <= not a;
    layer6_outputs(4720) <= a;
    layer6_outputs(4721) <= not b or a;
    layer6_outputs(4722) <= not b or a;
    layer6_outputs(4723) <= a and not b;
    layer6_outputs(4724) <= not (a or b);
    layer6_outputs(4725) <= a;
    layer6_outputs(4726) <= a or b;
    layer6_outputs(4727) <= not (a or b);
    layer6_outputs(4728) <= b;
    layer6_outputs(4729) <= a and not b;
    layer6_outputs(4730) <= a;
    layer6_outputs(4731) <= a xor b;
    layer6_outputs(4732) <= a;
    layer6_outputs(4733) <= not a;
    layer6_outputs(4734) <= a and not b;
    layer6_outputs(4735) <= not (a and b);
    layer6_outputs(4736) <= b;
    layer6_outputs(4737) <= a or b;
    layer6_outputs(4738) <= a xor b;
    layer6_outputs(4739) <= a and not b;
    layer6_outputs(4740) <= not (a or b);
    layer6_outputs(4741) <= not (a or b);
    layer6_outputs(4742) <= b and not a;
    layer6_outputs(4743) <= b;
    layer6_outputs(4744) <= 1'b0;
    layer6_outputs(4745) <= not b;
    layer6_outputs(4746) <= not (a and b);
    layer6_outputs(4747) <= b and not a;
    layer6_outputs(4748) <= not (a xor b);
    layer6_outputs(4749) <= a;
    layer6_outputs(4750) <= not (a and b);
    layer6_outputs(4751) <= a;
    layer6_outputs(4752) <= a;
    layer6_outputs(4753) <= a or b;
    layer6_outputs(4754) <= a or b;
    layer6_outputs(4755) <= not (a or b);
    layer6_outputs(4756) <= a xor b;
    layer6_outputs(4757) <= not (a xor b);
    layer6_outputs(4758) <= not b;
    layer6_outputs(4759) <= not a or b;
    layer6_outputs(4760) <= a and not b;
    layer6_outputs(4761) <= not b;
    layer6_outputs(4762) <= a or b;
    layer6_outputs(4763) <= not b or a;
    layer6_outputs(4764) <= a or b;
    layer6_outputs(4765) <= a;
    layer6_outputs(4766) <= not b;
    layer6_outputs(4767) <= not a;
    layer6_outputs(4768) <= b;
    layer6_outputs(4769) <= b;
    layer6_outputs(4770) <= not a;
    layer6_outputs(4771) <= not (a and b);
    layer6_outputs(4772) <= a and b;
    layer6_outputs(4773) <= a and b;
    layer6_outputs(4774) <= not a;
    layer6_outputs(4775) <= a xor b;
    layer6_outputs(4776) <= a;
    layer6_outputs(4777) <= not a;
    layer6_outputs(4778) <= not b or a;
    layer6_outputs(4779) <= 1'b0;
    layer6_outputs(4780) <= not b;
    layer6_outputs(4781) <= b;
    layer6_outputs(4782) <= b and not a;
    layer6_outputs(4783) <= not b;
    layer6_outputs(4784) <= a;
    layer6_outputs(4785) <= a and not b;
    layer6_outputs(4786) <= a;
    layer6_outputs(4787) <= not b;
    layer6_outputs(4788) <= b;
    layer6_outputs(4789) <= 1'b1;
    layer6_outputs(4790) <= b and not a;
    layer6_outputs(4791) <= a xor b;
    layer6_outputs(4792) <= 1'b0;
    layer6_outputs(4793) <= b and not a;
    layer6_outputs(4794) <= not a or b;
    layer6_outputs(4795) <= not b or a;
    layer6_outputs(4796) <= a;
    layer6_outputs(4797) <= not a or b;
    layer6_outputs(4798) <= a and b;
    layer6_outputs(4799) <= not b or a;
    layer6_outputs(4800) <= a and not b;
    layer6_outputs(4801) <= not b;
    layer6_outputs(4802) <= a;
    layer6_outputs(4803) <= not a;
    layer6_outputs(4804) <= not b;
    layer6_outputs(4805) <= a or b;
    layer6_outputs(4806) <= b and not a;
    layer6_outputs(4807) <= not a;
    layer6_outputs(4808) <= not a;
    layer6_outputs(4809) <= not a;
    layer6_outputs(4810) <= not a;
    layer6_outputs(4811) <= not (a and b);
    layer6_outputs(4812) <= not (a or b);
    layer6_outputs(4813) <= not b or a;
    layer6_outputs(4814) <= not b or a;
    layer6_outputs(4815) <= not b;
    layer6_outputs(4816) <= not b;
    layer6_outputs(4817) <= not b;
    layer6_outputs(4818) <= b;
    layer6_outputs(4819) <= not b or a;
    layer6_outputs(4820) <= not a;
    layer6_outputs(4821) <= not a or b;
    layer6_outputs(4822) <= not (a or b);
    layer6_outputs(4823) <= a;
    layer6_outputs(4824) <= not a or b;
    layer6_outputs(4825) <= a and not b;
    layer6_outputs(4826) <= not b;
    layer6_outputs(4827) <= not a or b;
    layer6_outputs(4828) <= b;
    layer6_outputs(4829) <= a;
    layer6_outputs(4830) <= not a or b;
    layer6_outputs(4831) <= 1'b0;
    layer6_outputs(4832) <= not a;
    layer6_outputs(4833) <= not b;
    layer6_outputs(4834) <= not a;
    layer6_outputs(4835) <= a;
    layer6_outputs(4836) <= a;
    layer6_outputs(4837) <= a and b;
    layer6_outputs(4838) <= b;
    layer6_outputs(4839) <= not (a xor b);
    layer6_outputs(4840) <= not a;
    layer6_outputs(4841) <= a and b;
    layer6_outputs(4842) <= not b or a;
    layer6_outputs(4843) <= not a or b;
    layer6_outputs(4844) <= b;
    layer6_outputs(4845) <= not (a xor b);
    layer6_outputs(4846) <= not b;
    layer6_outputs(4847) <= not a;
    layer6_outputs(4848) <= not b;
    layer6_outputs(4849) <= b and not a;
    layer6_outputs(4850) <= not a;
    layer6_outputs(4851) <= a or b;
    layer6_outputs(4852) <= 1'b0;
    layer6_outputs(4853) <= a xor b;
    layer6_outputs(4854) <= not (a xor b);
    layer6_outputs(4855) <= a and not b;
    layer6_outputs(4856) <= not a;
    layer6_outputs(4857) <= b;
    layer6_outputs(4858) <= not (a and b);
    layer6_outputs(4859) <= not b or a;
    layer6_outputs(4860) <= not a;
    layer6_outputs(4861) <= a and not b;
    layer6_outputs(4862) <= a and b;
    layer6_outputs(4863) <= a;
    layer6_outputs(4864) <= not b or a;
    layer6_outputs(4865) <= 1'b0;
    layer6_outputs(4866) <= a or b;
    layer6_outputs(4867) <= b;
    layer6_outputs(4868) <= a;
    layer6_outputs(4869) <= not b;
    layer6_outputs(4870) <= not a;
    layer6_outputs(4871) <= a and not b;
    layer6_outputs(4872) <= not (a or b);
    layer6_outputs(4873) <= b;
    layer6_outputs(4874) <= a;
    layer6_outputs(4875) <= not b;
    layer6_outputs(4876) <= a and b;
    layer6_outputs(4877) <= 1'b1;
    layer6_outputs(4878) <= a xor b;
    layer6_outputs(4879) <= not (a and b);
    layer6_outputs(4880) <= not b or a;
    layer6_outputs(4881) <= b and not a;
    layer6_outputs(4882) <= a;
    layer6_outputs(4883) <= a and not b;
    layer6_outputs(4884) <= not a or b;
    layer6_outputs(4885) <= not (a or b);
    layer6_outputs(4886) <= not (a or b);
    layer6_outputs(4887) <= b;
    layer6_outputs(4888) <= a;
    layer6_outputs(4889) <= a xor b;
    layer6_outputs(4890) <= b;
    layer6_outputs(4891) <= a and not b;
    layer6_outputs(4892) <= not (a xor b);
    layer6_outputs(4893) <= not b;
    layer6_outputs(4894) <= a xor b;
    layer6_outputs(4895) <= not (a or b);
    layer6_outputs(4896) <= a;
    layer6_outputs(4897) <= not (a xor b);
    layer6_outputs(4898) <= not b;
    layer6_outputs(4899) <= not (a and b);
    layer6_outputs(4900) <= not (a and b);
    layer6_outputs(4901) <= not a;
    layer6_outputs(4902) <= not a or b;
    layer6_outputs(4903) <= a or b;
    layer6_outputs(4904) <= not a;
    layer6_outputs(4905) <= not (a or b);
    layer6_outputs(4906) <= b;
    layer6_outputs(4907) <= a or b;
    layer6_outputs(4908) <= not (a and b);
    layer6_outputs(4909) <= not (a or b);
    layer6_outputs(4910) <= not b;
    layer6_outputs(4911) <= 1'b1;
    layer6_outputs(4912) <= b and not a;
    layer6_outputs(4913) <= b;
    layer6_outputs(4914) <= a;
    layer6_outputs(4915) <= not (a or b);
    layer6_outputs(4916) <= not b;
    layer6_outputs(4917) <= a and b;
    layer6_outputs(4918) <= not a;
    layer6_outputs(4919) <= b and not a;
    layer6_outputs(4920) <= a;
    layer6_outputs(4921) <= not a;
    layer6_outputs(4922) <= b and not a;
    layer6_outputs(4923) <= a or b;
    layer6_outputs(4924) <= b;
    layer6_outputs(4925) <= a or b;
    layer6_outputs(4926) <= b;
    layer6_outputs(4927) <= 1'b0;
    layer6_outputs(4928) <= not a;
    layer6_outputs(4929) <= not b;
    layer6_outputs(4930) <= not b;
    layer6_outputs(4931) <= not b;
    layer6_outputs(4932) <= a and not b;
    layer6_outputs(4933) <= 1'b1;
    layer6_outputs(4934) <= a xor b;
    layer6_outputs(4935) <= not a or b;
    layer6_outputs(4936) <= not b;
    layer6_outputs(4937) <= not (a or b);
    layer6_outputs(4938) <= b;
    layer6_outputs(4939) <= b;
    layer6_outputs(4940) <= not (a xor b);
    layer6_outputs(4941) <= not (a xor b);
    layer6_outputs(4942) <= b and not a;
    layer6_outputs(4943) <= not b;
    layer6_outputs(4944) <= a and not b;
    layer6_outputs(4945) <= not (a and b);
    layer6_outputs(4946) <= a;
    layer6_outputs(4947) <= a and not b;
    layer6_outputs(4948) <= a;
    layer6_outputs(4949) <= not (a and b);
    layer6_outputs(4950) <= a;
    layer6_outputs(4951) <= 1'b0;
    layer6_outputs(4952) <= a;
    layer6_outputs(4953) <= a xor b;
    layer6_outputs(4954) <= not a;
    layer6_outputs(4955) <= a or b;
    layer6_outputs(4956) <= b and not a;
    layer6_outputs(4957) <= b and not a;
    layer6_outputs(4958) <= not b;
    layer6_outputs(4959) <= b;
    layer6_outputs(4960) <= a and b;
    layer6_outputs(4961) <= not a or b;
    layer6_outputs(4962) <= not (a xor b);
    layer6_outputs(4963) <= 1'b0;
    layer6_outputs(4964) <= not a or b;
    layer6_outputs(4965) <= not b or a;
    layer6_outputs(4966) <= b;
    layer6_outputs(4967) <= b and not a;
    layer6_outputs(4968) <= a and not b;
    layer6_outputs(4969) <= not a or b;
    layer6_outputs(4970) <= not a;
    layer6_outputs(4971) <= a xor b;
    layer6_outputs(4972) <= a xor b;
    layer6_outputs(4973) <= a;
    layer6_outputs(4974) <= not b;
    layer6_outputs(4975) <= not (a or b);
    layer6_outputs(4976) <= a;
    layer6_outputs(4977) <= a or b;
    layer6_outputs(4978) <= not a;
    layer6_outputs(4979) <= a and not b;
    layer6_outputs(4980) <= not (a xor b);
    layer6_outputs(4981) <= not (a xor b);
    layer6_outputs(4982) <= not b;
    layer6_outputs(4983) <= b;
    layer6_outputs(4984) <= not (a or b);
    layer6_outputs(4985) <= a or b;
    layer6_outputs(4986) <= not a or b;
    layer6_outputs(4987) <= not b;
    layer6_outputs(4988) <= not b;
    layer6_outputs(4989) <= not (a or b);
    layer6_outputs(4990) <= a or b;
    layer6_outputs(4991) <= not a or b;
    layer6_outputs(4992) <= not b;
    layer6_outputs(4993) <= a xor b;
    layer6_outputs(4994) <= not a;
    layer6_outputs(4995) <= not b or a;
    layer6_outputs(4996) <= not (a xor b);
    layer6_outputs(4997) <= a and b;
    layer6_outputs(4998) <= a and b;
    layer6_outputs(4999) <= a;
    layer6_outputs(5000) <= a and not b;
    layer6_outputs(5001) <= a;
    layer6_outputs(5002) <= a;
    layer6_outputs(5003) <= not b or a;
    layer6_outputs(5004) <= not a or b;
    layer6_outputs(5005) <= a and b;
    layer6_outputs(5006) <= a;
    layer6_outputs(5007) <= not b or a;
    layer6_outputs(5008) <= not (a and b);
    layer6_outputs(5009) <= not (a and b);
    layer6_outputs(5010) <= b and not a;
    layer6_outputs(5011) <= not (a xor b);
    layer6_outputs(5012) <= a xor b;
    layer6_outputs(5013) <= b;
    layer6_outputs(5014) <= a;
    layer6_outputs(5015) <= a and not b;
    layer6_outputs(5016) <= not b or a;
    layer6_outputs(5017) <= not a;
    layer6_outputs(5018) <= not (a and b);
    layer6_outputs(5019) <= not (a xor b);
    layer6_outputs(5020) <= a;
    layer6_outputs(5021) <= not a;
    layer6_outputs(5022) <= not a;
    layer6_outputs(5023) <= b and not a;
    layer6_outputs(5024) <= a and b;
    layer6_outputs(5025) <= a or b;
    layer6_outputs(5026) <= not (a and b);
    layer6_outputs(5027) <= a and not b;
    layer6_outputs(5028) <= not b or a;
    layer6_outputs(5029) <= b and not a;
    layer6_outputs(5030) <= not (a xor b);
    layer6_outputs(5031) <= not a;
    layer6_outputs(5032) <= not (a and b);
    layer6_outputs(5033) <= not (a and b);
    layer6_outputs(5034) <= not (a and b);
    layer6_outputs(5035) <= not a or b;
    layer6_outputs(5036) <= a and not b;
    layer6_outputs(5037) <= a or b;
    layer6_outputs(5038) <= a xor b;
    layer6_outputs(5039) <= a xor b;
    layer6_outputs(5040) <= not a;
    layer6_outputs(5041) <= a;
    layer6_outputs(5042) <= not a or b;
    layer6_outputs(5043) <= a and not b;
    layer6_outputs(5044) <= not b;
    layer6_outputs(5045) <= not a or b;
    layer6_outputs(5046) <= b;
    layer6_outputs(5047) <= b;
    layer6_outputs(5048) <= not b;
    layer6_outputs(5049) <= a;
    layer6_outputs(5050) <= not b or a;
    layer6_outputs(5051) <= not (a or b);
    layer6_outputs(5052) <= 1'b0;
    layer6_outputs(5053) <= b and not a;
    layer6_outputs(5054) <= not b;
    layer6_outputs(5055) <= a or b;
    layer6_outputs(5056) <= not b;
    layer6_outputs(5057) <= not (a and b);
    layer6_outputs(5058) <= b and not a;
    layer6_outputs(5059) <= not a;
    layer6_outputs(5060) <= 1'b0;
    layer6_outputs(5061) <= not a;
    layer6_outputs(5062) <= not a or b;
    layer6_outputs(5063) <= not a or b;
    layer6_outputs(5064) <= a xor b;
    layer6_outputs(5065) <= a and b;
    layer6_outputs(5066) <= not (a or b);
    layer6_outputs(5067) <= not (a xor b);
    layer6_outputs(5068) <= a and b;
    layer6_outputs(5069) <= a xor b;
    layer6_outputs(5070) <= a;
    layer6_outputs(5071) <= not b;
    layer6_outputs(5072) <= b and not a;
    layer6_outputs(5073) <= not b;
    layer6_outputs(5074) <= a or b;
    layer6_outputs(5075) <= not a or b;
    layer6_outputs(5076) <= not b or a;
    layer6_outputs(5077) <= b;
    layer6_outputs(5078) <= not b;
    layer6_outputs(5079) <= not (a xor b);
    layer6_outputs(5080) <= not a;
    layer6_outputs(5081) <= not a or b;
    layer6_outputs(5082) <= not b;
    layer6_outputs(5083) <= a xor b;
    layer6_outputs(5084) <= not a or b;
    layer6_outputs(5085) <= a;
    layer6_outputs(5086) <= not (a xor b);
    layer6_outputs(5087) <= 1'b0;
    layer6_outputs(5088) <= not b or a;
    layer6_outputs(5089) <= not a or b;
    layer6_outputs(5090) <= not (a xor b);
    layer6_outputs(5091) <= not (a xor b);
    layer6_outputs(5092) <= not (a and b);
    layer6_outputs(5093) <= not a;
    layer6_outputs(5094) <= not a;
    layer6_outputs(5095) <= b and not a;
    layer6_outputs(5096) <= a and not b;
    layer6_outputs(5097) <= not b;
    layer6_outputs(5098) <= not (a or b);
    layer6_outputs(5099) <= not b;
    layer6_outputs(5100) <= not b;
    layer6_outputs(5101) <= b;
    layer6_outputs(5102) <= 1'b1;
    layer6_outputs(5103) <= a;
    layer6_outputs(5104) <= b;
    layer6_outputs(5105) <= a and b;
    layer6_outputs(5106) <= not a or b;
    layer6_outputs(5107) <= not (a and b);
    layer6_outputs(5108) <= b;
    layer6_outputs(5109) <= not b;
    layer6_outputs(5110) <= a;
    layer6_outputs(5111) <= a;
    layer6_outputs(5112) <= not (a xor b);
    layer6_outputs(5113) <= not b or a;
    layer6_outputs(5114) <= not (a or b);
    layer6_outputs(5115) <= a xor b;
    layer6_outputs(5116) <= a and b;
    layer6_outputs(5117) <= not a;
    layer6_outputs(5118) <= a xor b;
    layer6_outputs(5119) <= b and not a;
    layer6_outputs(5120) <= a;
    layer6_outputs(5121) <= a;
    layer6_outputs(5122) <= not (a and b);
    layer6_outputs(5123) <= not (a xor b);
    layer6_outputs(5124) <= a xor b;
    layer6_outputs(5125) <= not b;
    layer6_outputs(5126) <= not b or a;
    layer6_outputs(5127) <= not a;
    layer6_outputs(5128) <= a or b;
    layer6_outputs(5129) <= a;
    layer6_outputs(5130) <= not a or b;
    layer6_outputs(5131) <= a and not b;
    layer6_outputs(5132) <= a and not b;
    layer6_outputs(5133) <= not (a xor b);
    layer6_outputs(5134) <= b;
    layer6_outputs(5135) <= a;
    layer6_outputs(5136) <= not b;
    layer6_outputs(5137) <= b and not a;
    layer6_outputs(5138) <= not (a or b);
    layer6_outputs(5139) <= b and not a;
    layer6_outputs(5140) <= not b or a;
    layer6_outputs(5141) <= not a;
    layer6_outputs(5142) <= not (a or b);
    layer6_outputs(5143) <= b;
    layer6_outputs(5144) <= not (a and b);
    layer6_outputs(5145) <= a or b;
    layer6_outputs(5146) <= not b;
    layer6_outputs(5147) <= b;
    layer6_outputs(5148) <= not a or b;
    layer6_outputs(5149) <= a xor b;
    layer6_outputs(5150) <= a xor b;
    layer6_outputs(5151) <= 1'b0;
    layer6_outputs(5152) <= a xor b;
    layer6_outputs(5153) <= not b;
    layer6_outputs(5154) <= not b;
    layer6_outputs(5155) <= 1'b1;
    layer6_outputs(5156) <= a or b;
    layer6_outputs(5157) <= b;
    layer6_outputs(5158) <= a and not b;
    layer6_outputs(5159) <= b and not a;
    layer6_outputs(5160) <= a;
    layer6_outputs(5161) <= 1'b0;
    layer6_outputs(5162) <= not b;
    layer6_outputs(5163) <= not a;
    layer6_outputs(5164) <= a;
    layer6_outputs(5165) <= a xor b;
    layer6_outputs(5166) <= not a;
    layer6_outputs(5167) <= not b;
    layer6_outputs(5168) <= not a;
    layer6_outputs(5169) <= not (a or b);
    layer6_outputs(5170) <= b;
    layer6_outputs(5171) <= not (a xor b);
    layer6_outputs(5172) <= a or b;
    layer6_outputs(5173) <= not b;
    layer6_outputs(5174) <= not a;
    layer6_outputs(5175) <= a xor b;
    layer6_outputs(5176) <= not b or a;
    layer6_outputs(5177) <= not (a xor b);
    layer6_outputs(5178) <= 1'b1;
    layer6_outputs(5179) <= a and not b;
    layer6_outputs(5180) <= b;
    layer6_outputs(5181) <= a;
    layer6_outputs(5182) <= 1'b1;
    layer6_outputs(5183) <= b and not a;
    layer6_outputs(5184) <= not b;
    layer6_outputs(5185) <= not (a or b);
    layer6_outputs(5186) <= not b;
    layer6_outputs(5187) <= a;
    layer6_outputs(5188) <= a;
    layer6_outputs(5189) <= not a;
    layer6_outputs(5190) <= b and not a;
    layer6_outputs(5191) <= a;
    layer6_outputs(5192) <= 1'b1;
    layer6_outputs(5193) <= a and not b;
    layer6_outputs(5194) <= not b;
    layer6_outputs(5195) <= not b or a;
    layer6_outputs(5196) <= a;
    layer6_outputs(5197) <= b and not a;
    layer6_outputs(5198) <= not (a and b);
    layer6_outputs(5199) <= a and not b;
    layer6_outputs(5200) <= a and not b;
    layer6_outputs(5201) <= not a;
    layer6_outputs(5202) <= a;
    layer6_outputs(5203) <= a;
    layer6_outputs(5204) <= not (a xor b);
    layer6_outputs(5205) <= not (a or b);
    layer6_outputs(5206) <= a and not b;
    layer6_outputs(5207) <= b and not a;
    layer6_outputs(5208) <= not (a xor b);
    layer6_outputs(5209) <= a or b;
    layer6_outputs(5210) <= b;
    layer6_outputs(5211) <= not b;
    layer6_outputs(5212) <= a xor b;
    layer6_outputs(5213) <= b;
    layer6_outputs(5214) <= not (a and b);
    layer6_outputs(5215) <= not b or a;
    layer6_outputs(5216) <= a or b;
    layer6_outputs(5217) <= b and not a;
    layer6_outputs(5218) <= not a or b;
    layer6_outputs(5219) <= not (a or b);
    layer6_outputs(5220) <= not (a xor b);
    layer6_outputs(5221) <= a;
    layer6_outputs(5222) <= not a;
    layer6_outputs(5223) <= not a;
    layer6_outputs(5224) <= not b or a;
    layer6_outputs(5225) <= a or b;
    layer6_outputs(5226) <= not a;
    layer6_outputs(5227) <= a and b;
    layer6_outputs(5228) <= a xor b;
    layer6_outputs(5229) <= not (a and b);
    layer6_outputs(5230) <= not b or a;
    layer6_outputs(5231) <= not b;
    layer6_outputs(5232) <= b and not a;
    layer6_outputs(5233) <= not a or b;
    layer6_outputs(5234) <= not a or b;
    layer6_outputs(5235) <= a or b;
    layer6_outputs(5236) <= not (a xor b);
    layer6_outputs(5237) <= not b;
    layer6_outputs(5238) <= a and b;
    layer6_outputs(5239) <= a;
    layer6_outputs(5240) <= not (a or b);
    layer6_outputs(5241) <= not a or b;
    layer6_outputs(5242) <= a and b;
    layer6_outputs(5243) <= not b or a;
    layer6_outputs(5244) <= b;
    layer6_outputs(5245) <= not (a or b);
    layer6_outputs(5246) <= a;
    layer6_outputs(5247) <= b;
    layer6_outputs(5248) <= not b;
    layer6_outputs(5249) <= a;
    layer6_outputs(5250) <= a and b;
    layer6_outputs(5251) <= b;
    layer6_outputs(5252) <= 1'b0;
    layer6_outputs(5253) <= not b;
    layer6_outputs(5254) <= not b;
    layer6_outputs(5255) <= a;
    layer6_outputs(5256) <= 1'b0;
    layer6_outputs(5257) <= not a or b;
    layer6_outputs(5258) <= a;
    layer6_outputs(5259) <= not (a xor b);
    layer6_outputs(5260) <= a or b;
    layer6_outputs(5261) <= not b or a;
    layer6_outputs(5262) <= b;
    layer6_outputs(5263) <= not (a or b);
    layer6_outputs(5264) <= a;
    layer6_outputs(5265) <= not a or b;
    layer6_outputs(5266) <= a and not b;
    layer6_outputs(5267) <= not a;
    layer6_outputs(5268) <= not a;
    layer6_outputs(5269) <= b;
    layer6_outputs(5270) <= not b;
    layer6_outputs(5271) <= a and not b;
    layer6_outputs(5272) <= not b;
    layer6_outputs(5273) <= not a or b;
    layer6_outputs(5274) <= a or b;
    layer6_outputs(5275) <= not a or b;
    layer6_outputs(5276) <= not (a xor b);
    layer6_outputs(5277) <= a;
    layer6_outputs(5278) <= not (a or b);
    layer6_outputs(5279) <= b and not a;
    layer6_outputs(5280) <= not (a xor b);
    layer6_outputs(5281) <= a and b;
    layer6_outputs(5282) <= not (a or b);
    layer6_outputs(5283) <= b and not a;
    layer6_outputs(5284) <= a and b;
    layer6_outputs(5285) <= a;
    layer6_outputs(5286) <= not (a or b);
    layer6_outputs(5287) <= not a or b;
    layer6_outputs(5288) <= a and b;
    layer6_outputs(5289) <= not a;
    layer6_outputs(5290) <= a;
    layer6_outputs(5291) <= b;
    layer6_outputs(5292) <= not (a xor b);
    layer6_outputs(5293) <= not (a xor b);
    layer6_outputs(5294) <= not b or a;
    layer6_outputs(5295) <= a xor b;
    layer6_outputs(5296) <= a and b;
    layer6_outputs(5297) <= b;
    layer6_outputs(5298) <= a or b;
    layer6_outputs(5299) <= not (a or b);
    layer6_outputs(5300) <= a;
    layer6_outputs(5301) <= not a;
    layer6_outputs(5302) <= not b;
    layer6_outputs(5303) <= b;
    layer6_outputs(5304) <= b;
    layer6_outputs(5305) <= b and not a;
    layer6_outputs(5306) <= not a;
    layer6_outputs(5307) <= not (a and b);
    layer6_outputs(5308) <= not a;
    layer6_outputs(5309) <= a;
    layer6_outputs(5310) <= b;
    layer6_outputs(5311) <= not b;
    layer6_outputs(5312) <= not b;
    layer6_outputs(5313) <= not (a xor b);
    layer6_outputs(5314) <= not b or a;
    layer6_outputs(5315) <= not b;
    layer6_outputs(5316) <= a or b;
    layer6_outputs(5317) <= not (a and b);
    layer6_outputs(5318) <= a xor b;
    layer6_outputs(5319) <= a;
    layer6_outputs(5320) <= a and not b;
    layer6_outputs(5321) <= b;
    layer6_outputs(5322) <= 1'b0;
    layer6_outputs(5323) <= not a;
    layer6_outputs(5324) <= not a;
    layer6_outputs(5325) <= b;
    layer6_outputs(5326) <= b and not a;
    layer6_outputs(5327) <= a;
    layer6_outputs(5328) <= a and not b;
    layer6_outputs(5329) <= a;
    layer6_outputs(5330) <= b and not a;
    layer6_outputs(5331) <= a;
    layer6_outputs(5332) <= not a;
    layer6_outputs(5333) <= not a or b;
    layer6_outputs(5334) <= 1'b1;
    layer6_outputs(5335) <= a or b;
    layer6_outputs(5336) <= a or b;
    layer6_outputs(5337) <= not b or a;
    layer6_outputs(5338) <= a;
    layer6_outputs(5339) <= b;
    layer6_outputs(5340) <= not (a or b);
    layer6_outputs(5341) <= not a;
    layer6_outputs(5342) <= 1'b0;
    layer6_outputs(5343) <= not b;
    layer6_outputs(5344) <= not b;
    layer6_outputs(5345) <= not b or a;
    layer6_outputs(5346) <= a;
    layer6_outputs(5347) <= b;
    layer6_outputs(5348) <= not a;
    layer6_outputs(5349) <= a or b;
    layer6_outputs(5350) <= not b;
    layer6_outputs(5351) <= not a;
    layer6_outputs(5352) <= not b or a;
    layer6_outputs(5353) <= 1'b0;
    layer6_outputs(5354) <= a xor b;
    layer6_outputs(5355) <= not a;
    layer6_outputs(5356) <= not (a xor b);
    layer6_outputs(5357) <= a and b;
    layer6_outputs(5358) <= not b;
    layer6_outputs(5359) <= not b or a;
    layer6_outputs(5360) <= b;
    layer6_outputs(5361) <= not b;
    layer6_outputs(5362) <= not (a xor b);
    layer6_outputs(5363) <= not (a and b);
    layer6_outputs(5364) <= not a;
    layer6_outputs(5365) <= b and not a;
    layer6_outputs(5366) <= not (a xor b);
    layer6_outputs(5367) <= 1'b0;
    layer6_outputs(5368) <= not (a or b);
    layer6_outputs(5369) <= not a;
    layer6_outputs(5370) <= not a;
    layer6_outputs(5371) <= not (a xor b);
    layer6_outputs(5372) <= not a or b;
    layer6_outputs(5373) <= b;
    layer6_outputs(5374) <= not b;
    layer6_outputs(5375) <= a or b;
    layer6_outputs(5376) <= a;
    layer6_outputs(5377) <= not b;
    layer6_outputs(5378) <= not b or a;
    layer6_outputs(5379) <= not (a xor b);
    layer6_outputs(5380) <= not b;
    layer6_outputs(5381) <= not b or a;
    layer6_outputs(5382) <= not a;
    layer6_outputs(5383) <= a;
    layer6_outputs(5384) <= a xor b;
    layer6_outputs(5385) <= b;
    layer6_outputs(5386) <= not b;
    layer6_outputs(5387) <= b and not a;
    layer6_outputs(5388) <= not b;
    layer6_outputs(5389) <= not a or b;
    layer6_outputs(5390) <= 1'b0;
    layer6_outputs(5391) <= not b or a;
    layer6_outputs(5392) <= not b;
    layer6_outputs(5393) <= not (a xor b);
    layer6_outputs(5394) <= a xor b;
    layer6_outputs(5395) <= not b;
    layer6_outputs(5396) <= not a;
    layer6_outputs(5397) <= a xor b;
    layer6_outputs(5398) <= a;
    layer6_outputs(5399) <= a xor b;
    layer6_outputs(5400) <= a or b;
    layer6_outputs(5401) <= not b or a;
    layer6_outputs(5402) <= not a or b;
    layer6_outputs(5403) <= a;
    layer6_outputs(5404) <= not (a or b);
    layer6_outputs(5405) <= not b or a;
    layer6_outputs(5406) <= a;
    layer6_outputs(5407) <= b;
    layer6_outputs(5408) <= a and not b;
    layer6_outputs(5409) <= a xor b;
    layer6_outputs(5410) <= not a;
    layer6_outputs(5411) <= a;
    layer6_outputs(5412) <= not b;
    layer6_outputs(5413) <= a or b;
    layer6_outputs(5414) <= a;
    layer6_outputs(5415) <= b and not a;
    layer6_outputs(5416) <= a or b;
    layer6_outputs(5417) <= a;
    layer6_outputs(5418) <= 1'b0;
    layer6_outputs(5419) <= not a;
    layer6_outputs(5420) <= b;
    layer6_outputs(5421) <= not (a xor b);
    layer6_outputs(5422) <= not a;
    layer6_outputs(5423) <= a or b;
    layer6_outputs(5424) <= not a or b;
    layer6_outputs(5425) <= a and not b;
    layer6_outputs(5426) <= a or b;
    layer6_outputs(5427) <= not b;
    layer6_outputs(5428) <= a and b;
    layer6_outputs(5429) <= b;
    layer6_outputs(5430) <= a xor b;
    layer6_outputs(5431) <= b;
    layer6_outputs(5432) <= not (a or b);
    layer6_outputs(5433) <= not (a and b);
    layer6_outputs(5434) <= not b or a;
    layer6_outputs(5435) <= b;
    layer6_outputs(5436) <= a;
    layer6_outputs(5437) <= a xor b;
    layer6_outputs(5438) <= not a;
    layer6_outputs(5439) <= not (a xor b);
    layer6_outputs(5440) <= not b;
    layer6_outputs(5441) <= a or b;
    layer6_outputs(5442) <= not (a or b);
    layer6_outputs(5443) <= not a or b;
    layer6_outputs(5444) <= b;
    layer6_outputs(5445) <= a;
    layer6_outputs(5446) <= a and b;
    layer6_outputs(5447) <= not (a and b);
    layer6_outputs(5448) <= a and b;
    layer6_outputs(5449) <= b;
    layer6_outputs(5450) <= not a;
    layer6_outputs(5451) <= a xor b;
    layer6_outputs(5452) <= not (a xor b);
    layer6_outputs(5453) <= not b or a;
    layer6_outputs(5454) <= b;
    layer6_outputs(5455) <= b;
    layer6_outputs(5456) <= a;
    layer6_outputs(5457) <= a;
    layer6_outputs(5458) <= not a or b;
    layer6_outputs(5459) <= a or b;
    layer6_outputs(5460) <= not a;
    layer6_outputs(5461) <= b;
    layer6_outputs(5462) <= a and not b;
    layer6_outputs(5463) <= not b or a;
    layer6_outputs(5464) <= a and not b;
    layer6_outputs(5465) <= a xor b;
    layer6_outputs(5466) <= not a or b;
    layer6_outputs(5467) <= a and not b;
    layer6_outputs(5468) <= not (a and b);
    layer6_outputs(5469) <= not b;
    layer6_outputs(5470) <= b and not a;
    layer6_outputs(5471) <= not a;
    layer6_outputs(5472) <= not (a and b);
    layer6_outputs(5473) <= not b or a;
    layer6_outputs(5474) <= a or b;
    layer6_outputs(5475) <= not (a or b);
    layer6_outputs(5476) <= not b;
    layer6_outputs(5477) <= not a;
    layer6_outputs(5478) <= not (a or b);
    layer6_outputs(5479) <= not b;
    layer6_outputs(5480) <= a;
    layer6_outputs(5481) <= not a or b;
    layer6_outputs(5482) <= 1'b1;
    layer6_outputs(5483) <= b and not a;
    layer6_outputs(5484) <= not (a or b);
    layer6_outputs(5485) <= not (a xor b);
    layer6_outputs(5486) <= 1'b1;
    layer6_outputs(5487) <= not (a and b);
    layer6_outputs(5488) <= a;
    layer6_outputs(5489) <= 1'b0;
    layer6_outputs(5490) <= a;
    layer6_outputs(5491) <= not (a and b);
    layer6_outputs(5492) <= a;
    layer6_outputs(5493) <= a or b;
    layer6_outputs(5494) <= a xor b;
    layer6_outputs(5495) <= not b;
    layer6_outputs(5496) <= a xor b;
    layer6_outputs(5497) <= a;
    layer6_outputs(5498) <= b;
    layer6_outputs(5499) <= not (a or b);
    layer6_outputs(5500) <= not b;
    layer6_outputs(5501) <= b;
    layer6_outputs(5502) <= not a;
    layer6_outputs(5503) <= a and b;
    layer6_outputs(5504) <= b and not a;
    layer6_outputs(5505) <= not b or a;
    layer6_outputs(5506) <= not a;
    layer6_outputs(5507) <= a;
    layer6_outputs(5508) <= not b;
    layer6_outputs(5509) <= 1'b1;
    layer6_outputs(5510) <= not (a or b);
    layer6_outputs(5511) <= not a or b;
    layer6_outputs(5512) <= b;
    layer6_outputs(5513) <= not (a and b);
    layer6_outputs(5514) <= a xor b;
    layer6_outputs(5515) <= not (a and b);
    layer6_outputs(5516) <= a or b;
    layer6_outputs(5517) <= a;
    layer6_outputs(5518) <= not b;
    layer6_outputs(5519) <= a;
    layer6_outputs(5520) <= a;
    layer6_outputs(5521) <= not b;
    layer6_outputs(5522) <= a and b;
    layer6_outputs(5523) <= a;
    layer6_outputs(5524) <= not (a and b);
    layer6_outputs(5525) <= not a;
    layer6_outputs(5526) <= not a;
    layer6_outputs(5527) <= a;
    layer6_outputs(5528) <= a and not b;
    layer6_outputs(5529) <= a and not b;
    layer6_outputs(5530) <= not a;
    layer6_outputs(5531) <= a xor b;
    layer6_outputs(5532) <= a;
    layer6_outputs(5533) <= not b;
    layer6_outputs(5534) <= a xor b;
    layer6_outputs(5535) <= not a;
    layer6_outputs(5536) <= a and b;
    layer6_outputs(5537) <= a or b;
    layer6_outputs(5538) <= a and not b;
    layer6_outputs(5539) <= a xor b;
    layer6_outputs(5540) <= a;
    layer6_outputs(5541) <= not (a and b);
    layer6_outputs(5542) <= b;
    layer6_outputs(5543) <= b and not a;
    layer6_outputs(5544) <= a;
    layer6_outputs(5545) <= not b;
    layer6_outputs(5546) <= not (a and b);
    layer6_outputs(5547) <= a and b;
    layer6_outputs(5548) <= not (a and b);
    layer6_outputs(5549) <= b;
    layer6_outputs(5550) <= not a or b;
    layer6_outputs(5551) <= b and not a;
    layer6_outputs(5552) <= b;
    layer6_outputs(5553) <= not (a or b);
    layer6_outputs(5554) <= a;
    layer6_outputs(5555) <= a or b;
    layer6_outputs(5556) <= not (a or b);
    layer6_outputs(5557) <= a and not b;
    layer6_outputs(5558) <= not a;
    layer6_outputs(5559) <= not (a and b);
    layer6_outputs(5560) <= not b;
    layer6_outputs(5561) <= a or b;
    layer6_outputs(5562) <= not (a or b);
    layer6_outputs(5563) <= 1'b1;
    layer6_outputs(5564) <= a and not b;
    layer6_outputs(5565) <= a and b;
    layer6_outputs(5566) <= a and b;
    layer6_outputs(5567) <= b;
    layer6_outputs(5568) <= not (a xor b);
    layer6_outputs(5569) <= not (a and b);
    layer6_outputs(5570) <= not (a and b);
    layer6_outputs(5571) <= not b;
    layer6_outputs(5572) <= a or b;
    layer6_outputs(5573) <= not (a or b);
    layer6_outputs(5574) <= a;
    layer6_outputs(5575) <= not (a or b);
    layer6_outputs(5576) <= not (a xor b);
    layer6_outputs(5577) <= a;
    layer6_outputs(5578) <= a;
    layer6_outputs(5579) <= not (a or b);
    layer6_outputs(5580) <= not b;
    layer6_outputs(5581) <= a and b;
    layer6_outputs(5582) <= not b or a;
    layer6_outputs(5583) <= b;
    layer6_outputs(5584) <= not b;
    layer6_outputs(5585) <= a;
    layer6_outputs(5586) <= 1'b1;
    layer6_outputs(5587) <= b;
    layer6_outputs(5588) <= a;
    layer6_outputs(5589) <= a and not b;
    layer6_outputs(5590) <= 1'b1;
    layer6_outputs(5591) <= a or b;
    layer6_outputs(5592) <= a and not b;
    layer6_outputs(5593) <= not a;
    layer6_outputs(5594) <= b and not a;
    layer6_outputs(5595) <= a xor b;
    layer6_outputs(5596) <= not (a and b);
    layer6_outputs(5597) <= a or b;
    layer6_outputs(5598) <= not a or b;
    layer6_outputs(5599) <= not (a or b);
    layer6_outputs(5600) <= a;
    layer6_outputs(5601) <= b;
    layer6_outputs(5602) <= a;
    layer6_outputs(5603) <= a;
    layer6_outputs(5604) <= not b;
    layer6_outputs(5605) <= a and not b;
    layer6_outputs(5606) <= b;
    layer6_outputs(5607) <= a and not b;
    layer6_outputs(5608) <= not a or b;
    layer6_outputs(5609) <= b;
    layer6_outputs(5610) <= not b;
    layer6_outputs(5611) <= not (a xor b);
    layer6_outputs(5612) <= 1'b1;
    layer6_outputs(5613) <= not a or b;
    layer6_outputs(5614) <= not b;
    layer6_outputs(5615) <= not a or b;
    layer6_outputs(5616) <= not b;
    layer6_outputs(5617) <= not a or b;
    layer6_outputs(5618) <= not (a and b);
    layer6_outputs(5619) <= not a;
    layer6_outputs(5620) <= a and not b;
    layer6_outputs(5621) <= a and not b;
    layer6_outputs(5622) <= 1'b0;
    layer6_outputs(5623) <= not a;
    layer6_outputs(5624) <= a;
    layer6_outputs(5625) <= not (a or b);
    layer6_outputs(5626) <= b;
    layer6_outputs(5627) <= not b;
    layer6_outputs(5628) <= not b;
    layer6_outputs(5629) <= not b;
    layer6_outputs(5630) <= a or b;
    layer6_outputs(5631) <= b;
    layer6_outputs(5632) <= a xor b;
    layer6_outputs(5633) <= not a;
    layer6_outputs(5634) <= b;
    layer6_outputs(5635) <= a and not b;
    layer6_outputs(5636) <= b and not a;
    layer6_outputs(5637) <= not (a and b);
    layer6_outputs(5638) <= b;
    layer6_outputs(5639) <= not (a or b);
    layer6_outputs(5640) <= not (a and b);
    layer6_outputs(5641) <= a;
    layer6_outputs(5642) <= a;
    layer6_outputs(5643) <= not (a xor b);
    layer6_outputs(5644) <= a or b;
    layer6_outputs(5645) <= not (a xor b);
    layer6_outputs(5646) <= not (a and b);
    layer6_outputs(5647) <= a;
    layer6_outputs(5648) <= not a;
    layer6_outputs(5649) <= not a or b;
    layer6_outputs(5650) <= a and b;
    layer6_outputs(5651) <= a and not b;
    layer6_outputs(5652) <= a xor b;
    layer6_outputs(5653) <= not b or a;
    layer6_outputs(5654) <= not b;
    layer6_outputs(5655) <= a;
    layer6_outputs(5656) <= not a;
    layer6_outputs(5657) <= a;
    layer6_outputs(5658) <= a;
    layer6_outputs(5659) <= a or b;
    layer6_outputs(5660) <= a;
    layer6_outputs(5661) <= not a;
    layer6_outputs(5662) <= 1'b0;
    layer6_outputs(5663) <= b;
    layer6_outputs(5664) <= a xor b;
    layer6_outputs(5665) <= not a or b;
    layer6_outputs(5666) <= not b or a;
    layer6_outputs(5667) <= a and b;
    layer6_outputs(5668) <= a;
    layer6_outputs(5669) <= a;
    layer6_outputs(5670) <= 1'b0;
    layer6_outputs(5671) <= not b;
    layer6_outputs(5672) <= b and not a;
    layer6_outputs(5673) <= a;
    layer6_outputs(5674) <= not (a xor b);
    layer6_outputs(5675) <= 1'b1;
    layer6_outputs(5676) <= not b or a;
    layer6_outputs(5677) <= a;
    layer6_outputs(5678) <= a xor b;
    layer6_outputs(5679) <= a and b;
    layer6_outputs(5680) <= b and not a;
    layer6_outputs(5681) <= not a;
    layer6_outputs(5682) <= a xor b;
    layer6_outputs(5683) <= not (a or b);
    layer6_outputs(5684) <= a or b;
    layer6_outputs(5685) <= not a or b;
    layer6_outputs(5686) <= a xor b;
    layer6_outputs(5687) <= a and not b;
    layer6_outputs(5688) <= a and b;
    layer6_outputs(5689) <= not (a xor b);
    layer6_outputs(5690) <= b;
    layer6_outputs(5691) <= not b;
    layer6_outputs(5692) <= b and not a;
    layer6_outputs(5693) <= b;
    layer6_outputs(5694) <= b and not a;
    layer6_outputs(5695) <= a;
    layer6_outputs(5696) <= a or b;
    layer6_outputs(5697) <= a;
    layer6_outputs(5698) <= not b;
    layer6_outputs(5699) <= not b;
    layer6_outputs(5700) <= not b;
    layer6_outputs(5701) <= a xor b;
    layer6_outputs(5702) <= not (a or b);
    layer6_outputs(5703) <= a or b;
    layer6_outputs(5704) <= a xor b;
    layer6_outputs(5705) <= b and not a;
    layer6_outputs(5706) <= not a;
    layer6_outputs(5707) <= not a;
    layer6_outputs(5708) <= a;
    layer6_outputs(5709) <= 1'b0;
    layer6_outputs(5710) <= not a;
    layer6_outputs(5711) <= b and not a;
    layer6_outputs(5712) <= a xor b;
    layer6_outputs(5713) <= not (a xor b);
    layer6_outputs(5714) <= not a;
    layer6_outputs(5715) <= not a or b;
    layer6_outputs(5716) <= a;
    layer6_outputs(5717) <= a or b;
    layer6_outputs(5718) <= not a;
    layer6_outputs(5719) <= 1'b0;
    layer6_outputs(5720) <= not a;
    layer6_outputs(5721) <= 1'b0;
    layer6_outputs(5722) <= not b;
    layer6_outputs(5723) <= not b or a;
    layer6_outputs(5724) <= b and not a;
    layer6_outputs(5725) <= 1'b1;
    layer6_outputs(5726) <= a or b;
    layer6_outputs(5727) <= not a;
    layer6_outputs(5728) <= not a;
    layer6_outputs(5729) <= a or b;
    layer6_outputs(5730) <= b and not a;
    layer6_outputs(5731) <= not b or a;
    layer6_outputs(5732) <= not (a xor b);
    layer6_outputs(5733) <= not a or b;
    layer6_outputs(5734) <= not b;
    layer6_outputs(5735) <= b;
    layer6_outputs(5736) <= a or b;
    layer6_outputs(5737) <= 1'b1;
    layer6_outputs(5738) <= not a;
    layer6_outputs(5739) <= a or b;
    layer6_outputs(5740) <= b;
    layer6_outputs(5741) <= a or b;
    layer6_outputs(5742) <= a or b;
    layer6_outputs(5743) <= a;
    layer6_outputs(5744) <= b;
    layer6_outputs(5745) <= not a;
    layer6_outputs(5746) <= a and not b;
    layer6_outputs(5747) <= not b;
    layer6_outputs(5748) <= not b;
    layer6_outputs(5749) <= a;
    layer6_outputs(5750) <= a;
    layer6_outputs(5751) <= b;
    layer6_outputs(5752) <= not a or b;
    layer6_outputs(5753) <= not b;
    layer6_outputs(5754) <= not b or a;
    layer6_outputs(5755) <= b;
    layer6_outputs(5756) <= not b or a;
    layer6_outputs(5757) <= not b;
    layer6_outputs(5758) <= not b or a;
    layer6_outputs(5759) <= b and not a;
    layer6_outputs(5760) <= a xor b;
    layer6_outputs(5761) <= not (a and b);
    layer6_outputs(5762) <= a xor b;
    layer6_outputs(5763) <= a and b;
    layer6_outputs(5764) <= a and b;
    layer6_outputs(5765) <= not b;
    layer6_outputs(5766) <= not b;
    layer6_outputs(5767) <= b and not a;
    layer6_outputs(5768) <= not b;
    layer6_outputs(5769) <= a;
    layer6_outputs(5770) <= a;
    layer6_outputs(5771) <= not a;
    layer6_outputs(5772) <= not a;
    layer6_outputs(5773) <= b and not a;
    layer6_outputs(5774) <= a;
    layer6_outputs(5775) <= not a or b;
    layer6_outputs(5776) <= 1'b1;
    layer6_outputs(5777) <= 1'b1;
    layer6_outputs(5778) <= b;
    layer6_outputs(5779) <= not a;
    layer6_outputs(5780) <= 1'b0;
    layer6_outputs(5781) <= not a;
    layer6_outputs(5782) <= b;
    layer6_outputs(5783) <= b;
    layer6_outputs(5784) <= a or b;
    layer6_outputs(5785) <= not (a and b);
    layer6_outputs(5786) <= not a;
    layer6_outputs(5787) <= b and not a;
    layer6_outputs(5788) <= b;
    layer6_outputs(5789) <= not b or a;
    layer6_outputs(5790) <= b and not a;
    layer6_outputs(5791) <= b and not a;
    layer6_outputs(5792) <= a and not b;
    layer6_outputs(5793) <= not b;
    layer6_outputs(5794) <= 1'b0;
    layer6_outputs(5795) <= not (a xor b);
    layer6_outputs(5796) <= a xor b;
    layer6_outputs(5797) <= not b or a;
    layer6_outputs(5798) <= b and not a;
    layer6_outputs(5799) <= not b;
    layer6_outputs(5800) <= not b;
    layer6_outputs(5801) <= a;
    layer6_outputs(5802) <= b and not a;
    layer6_outputs(5803) <= not a;
    layer6_outputs(5804) <= 1'b0;
    layer6_outputs(5805) <= b;
    layer6_outputs(5806) <= not (a or b);
    layer6_outputs(5807) <= not a;
    layer6_outputs(5808) <= not a;
    layer6_outputs(5809) <= a xor b;
    layer6_outputs(5810) <= not a;
    layer6_outputs(5811) <= b;
    layer6_outputs(5812) <= a;
    layer6_outputs(5813) <= not a;
    layer6_outputs(5814) <= not (a or b);
    layer6_outputs(5815) <= not (a and b);
    layer6_outputs(5816) <= not (a or b);
    layer6_outputs(5817) <= not b;
    layer6_outputs(5818) <= a;
    layer6_outputs(5819) <= a and b;
    layer6_outputs(5820) <= a xor b;
    layer6_outputs(5821) <= a;
    layer6_outputs(5822) <= a;
    layer6_outputs(5823) <= a;
    layer6_outputs(5824) <= not b or a;
    layer6_outputs(5825) <= not a;
    layer6_outputs(5826) <= b;
    layer6_outputs(5827) <= a;
    layer6_outputs(5828) <= not b;
    layer6_outputs(5829) <= a;
    layer6_outputs(5830) <= b;
    layer6_outputs(5831) <= a and not b;
    layer6_outputs(5832) <= not (a or b);
    layer6_outputs(5833) <= not b;
    layer6_outputs(5834) <= a or b;
    layer6_outputs(5835) <= a;
    layer6_outputs(5836) <= not a;
    layer6_outputs(5837) <= not b;
    layer6_outputs(5838) <= not b;
    layer6_outputs(5839) <= 1'b0;
    layer6_outputs(5840) <= not a;
    layer6_outputs(5841) <= a;
    layer6_outputs(5842) <= 1'b0;
    layer6_outputs(5843) <= not a or b;
    layer6_outputs(5844) <= not (a xor b);
    layer6_outputs(5845) <= a or b;
    layer6_outputs(5846) <= not b;
    layer6_outputs(5847) <= not b;
    layer6_outputs(5848) <= 1'b1;
    layer6_outputs(5849) <= not a;
    layer6_outputs(5850) <= not a;
    layer6_outputs(5851) <= not (a xor b);
    layer6_outputs(5852) <= b;
    layer6_outputs(5853) <= not (a and b);
    layer6_outputs(5854) <= a;
    layer6_outputs(5855) <= a;
    layer6_outputs(5856) <= 1'b0;
    layer6_outputs(5857) <= a;
    layer6_outputs(5858) <= b;
    layer6_outputs(5859) <= a and b;
    layer6_outputs(5860) <= a and b;
    layer6_outputs(5861) <= not b;
    layer6_outputs(5862) <= b and not a;
    layer6_outputs(5863) <= a and b;
    layer6_outputs(5864) <= not (a xor b);
    layer6_outputs(5865) <= a xor b;
    layer6_outputs(5866) <= a xor b;
    layer6_outputs(5867) <= not a;
    layer6_outputs(5868) <= b and not a;
    layer6_outputs(5869) <= not a;
    layer6_outputs(5870) <= not b;
    layer6_outputs(5871) <= b and not a;
    layer6_outputs(5872) <= b;
    layer6_outputs(5873) <= not (a or b);
    layer6_outputs(5874) <= b and not a;
    layer6_outputs(5875) <= a or b;
    layer6_outputs(5876) <= a;
    layer6_outputs(5877) <= not b;
    layer6_outputs(5878) <= not b;
    layer6_outputs(5879) <= not a or b;
    layer6_outputs(5880) <= not a;
    layer6_outputs(5881) <= b and not a;
    layer6_outputs(5882) <= not b or a;
    layer6_outputs(5883) <= b;
    layer6_outputs(5884) <= not a or b;
    layer6_outputs(5885) <= 1'b0;
    layer6_outputs(5886) <= not (a xor b);
    layer6_outputs(5887) <= a and b;
    layer6_outputs(5888) <= not b or a;
    layer6_outputs(5889) <= b;
    layer6_outputs(5890) <= not (a or b);
    layer6_outputs(5891) <= not (a and b);
    layer6_outputs(5892) <= b;
    layer6_outputs(5893) <= not b or a;
    layer6_outputs(5894) <= b;
    layer6_outputs(5895) <= not a;
    layer6_outputs(5896) <= not b;
    layer6_outputs(5897) <= a xor b;
    layer6_outputs(5898) <= not b or a;
    layer6_outputs(5899) <= not (a xor b);
    layer6_outputs(5900) <= a;
    layer6_outputs(5901) <= not a;
    layer6_outputs(5902) <= not b or a;
    layer6_outputs(5903) <= a and b;
    layer6_outputs(5904) <= not a or b;
    layer6_outputs(5905) <= a;
    layer6_outputs(5906) <= b;
    layer6_outputs(5907) <= a xor b;
    layer6_outputs(5908) <= a and not b;
    layer6_outputs(5909) <= b;
    layer6_outputs(5910) <= a;
    layer6_outputs(5911) <= a and not b;
    layer6_outputs(5912) <= a and b;
    layer6_outputs(5913) <= not (a and b);
    layer6_outputs(5914) <= not (a and b);
    layer6_outputs(5915) <= b;
    layer6_outputs(5916) <= a xor b;
    layer6_outputs(5917) <= not b;
    layer6_outputs(5918) <= not a;
    layer6_outputs(5919) <= a and not b;
    layer6_outputs(5920) <= not (a xor b);
    layer6_outputs(5921) <= a and b;
    layer6_outputs(5922) <= 1'b0;
    layer6_outputs(5923) <= b and not a;
    layer6_outputs(5924) <= not a or b;
    layer6_outputs(5925) <= a and not b;
    layer6_outputs(5926) <= 1'b1;
    layer6_outputs(5927) <= not (a or b);
    layer6_outputs(5928) <= not a;
    layer6_outputs(5929) <= b;
    layer6_outputs(5930) <= 1'b1;
    layer6_outputs(5931) <= not a or b;
    layer6_outputs(5932) <= a or b;
    layer6_outputs(5933) <= not b or a;
    layer6_outputs(5934) <= a or b;
    layer6_outputs(5935) <= not b;
    layer6_outputs(5936) <= 1'b0;
    layer6_outputs(5937) <= b;
    layer6_outputs(5938) <= not b;
    layer6_outputs(5939) <= not a;
    layer6_outputs(5940) <= 1'b1;
    layer6_outputs(5941) <= a;
    layer6_outputs(5942) <= b;
    layer6_outputs(5943) <= not b or a;
    layer6_outputs(5944) <= b and not a;
    layer6_outputs(5945) <= not a;
    layer6_outputs(5946) <= not b;
    layer6_outputs(5947) <= b and not a;
    layer6_outputs(5948) <= a and not b;
    layer6_outputs(5949) <= not (a and b);
    layer6_outputs(5950) <= a xor b;
    layer6_outputs(5951) <= not (a xor b);
    layer6_outputs(5952) <= not (a xor b);
    layer6_outputs(5953) <= not b;
    layer6_outputs(5954) <= not b or a;
    layer6_outputs(5955) <= a or b;
    layer6_outputs(5956) <= a;
    layer6_outputs(5957) <= not b or a;
    layer6_outputs(5958) <= b;
    layer6_outputs(5959) <= b;
    layer6_outputs(5960) <= not (a or b);
    layer6_outputs(5961) <= not b;
    layer6_outputs(5962) <= 1'b1;
    layer6_outputs(5963) <= not b;
    layer6_outputs(5964) <= a and b;
    layer6_outputs(5965) <= a;
    layer6_outputs(5966) <= a xor b;
    layer6_outputs(5967) <= not b;
    layer6_outputs(5968) <= not (a xor b);
    layer6_outputs(5969) <= not b or a;
    layer6_outputs(5970) <= a and b;
    layer6_outputs(5971) <= b;
    layer6_outputs(5972) <= not a;
    layer6_outputs(5973) <= b;
    layer6_outputs(5974) <= a or b;
    layer6_outputs(5975) <= a;
    layer6_outputs(5976) <= a;
    layer6_outputs(5977) <= a;
    layer6_outputs(5978) <= not b;
    layer6_outputs(5979) <= not a;
    layer6_outputs(5980) <= not b;
    layer6_outputs(5981) <= b;
    layer6_outputs(5982) <= not a or b;
    layer6_outputs(5983) <= not (a xor b);
    layer6_outputs(5984) <= not a or b;
    layer6_outputs(5985) <= not a;
    layer6_outputs(5986) <= a or b;
    layer6_outputs(5987) <= b;
    layer6_outputs(5988) <= a and b;
    layer6_outputs(5989) <= 1'b1;
    layer6_outputs(5990) <= not a;
    layer6_outputs(5991) <= b;
    layer6_outputs(5992) <= a xor b;
    layer6_outputs(5993) <= a;
    layer6_outputs(5994) <= b;
    layer6_outputs(5995) <= not a or b;
    layer6_outputs(5996) <= a xor b;
    layer6_outputs(5997) <= not (a xor b);
    layer6_outputs(5998) <= a and b;
    layer6_outputs(5999) <= a xor b;
    layer6_outputs(6000) <= a xor b;
    layer6_outputs(6001) <= not a;
    layer6_outputs(6002) <= a xor b;
    layer6_outputs(6003) <= not b;
    layer6_outputs(6004) <= a and not b;
    layer6_outputs(6005) <= b;
    layer6_outputs(6006) <= a or b;
    layer6_outputs(6007) <= 1'b1;
    layer6_outputs(6008) <= a xor b;
    layer6_outputs(6009) <= a;
    layer6_outputs(6010) <= not a or b;
    layer6_outputs(6011) <= a;
    layer6_outputs(6012) <= a and b;
    layer6_outputs(6013) <= not b;
    layer6_outputs(6014) <= a;
    layer6_outputs(6015) <= not (a or b);
    layer6_outputs(6016) <= not (a xor b);
    layer6_outputs(6017) <= not b;
    layer6_outputs(6018) <= a xor b;
    layer6_outputs(6019) <= b and not a;
    layer6_outputs(6020) <= not (a xor b);
    layer6_outputs(6021) <= not (a xor b);
    layer6_outputs(6022) <= b;
    layer6_outputs(6023) <= 1'b0;
    layer6_outputs(6024) <= a or b;
    layer6_outputs(6025) <= not b or a;
    layer6_outputs(6026) <= not (a xor b);
    layer6_outputs(6027) <= not a;
    layer6_outputs(6028) <= a or b;
    layer6_outputs(6029) <= not a or b;
    layer6_outputs(6030) <= not a;
    layer6_outputs(6031) <= not b;
    layer6_outputs(6032) <= not b;
    layer6_outputs(6033) <= a;
    layer6_outputs(6034) <= not (a and b);
    layer6_outputs(6035) <= not (a and b);
    layer6_outputs(6036) <= not (a xor b);
    layer6_outputs(6037) <= a or b;
    layer6_outputs(6038) <= a and not b;
    layer6_outputs(6039) <= a;
    layer6_outputs(6040) <= not (a and b);
    layer6_outputs(6041) <= not a;
    layer6_outputs(6042) <= not (a or b);
    layer6_outputs(6043) <= not b;
    layer6_outputs(6044) <= a;
    layer6_outputs(6045) <= not b;
    layer6_outputs(6046) <= b and not a;
    layer6_outputs(6047) <= not a or b;
    layer6_outputs(6048) <= b and not a;
    layer6_outputs(6049) <= a and b;
    layer6_outputs(6050) <= not b;
    layer6_outputs(6051) <= b;
    layer6_outputs(6052) <= not (a and b);
    layer6_outputs(6053) <= a;
    layer6_outputs(6054) <= not b or a;
    layer6_outputs(6055) <= b;
    layer6_outputs(6056) <= not b;
    layer6_outputs(6057) <= b;
    layer6_outputs(6058) <= not a or b;
    layer6_outputs(6059) <= not a;
    layer6_outputs(6060) <= a or b;
    layer6_outputs(6061) <= a;
    layer6_outputs(6062) <= not b;
    layer6_outputs(6063) <= b;
    layer6_outputs(6064) <= b and not a;
    layer6_outputs(6065) <= a or b;
    layer6_outputs(6066) <= a xor b;
    layer6_outputs(6067) <= a or b;
    layer6_outputs(6068) <= a and b;
    layer6_outputs(6069) <= not b or a;
    layer6_outputs(6070) <= b and not a;
    layer6_outputs(6071) <= not b;
    layer6_outputs(6072) <= b;
    layer6_outputs(6073) <= not a;
    layer6_outputs(6074) <= a xor b;
    layer6_outputs(6075) <= 1'b0;
    layer6_outputs(6076) <= not b;
    layer6_outputs(6077) <= 1'b1;
    layer6_outputs(6078) <= not b;
    layer6_outputs(6079) <= b;
    layer6_outputs(6080) <= not (a xor b);
    layer6_outputs(6081) <= a xor b;
    layer6_outputs(6082) <= not (a and b);
    layer6_outputs(6083) <= b;
    layer6_outputs(6084) <= not b or a;
    layer6_outputs(6085) <= a;
    layer6_outputs(6086) <= a and b;
    layer6_outputs(6087) <= not b or a;
    layer6_outputs(6088) <= a or b;
    layer6_outputs(6089) <= b and not a;
    layer6_outputs(6090) <= not b or a;
    layer6_outputs(6091) <= not (a or b);
    layer6_outputs(6092) <= b;
    layer6_outputs(6093) <= b and not a;
    layer6_outputs(6094) <= not a;
    layer6_outputs(6095) <= 1'b0;
    layer6_outputs(6096) <= b and not a;
    layer6_outputs(6097) <= b and not a;
    layer6_outputs(6098) <= not a or b;
    layer6_outputs(6099) <= not a;
    layer6_outputs(6100) <= a or b;
    layer6_outputs(6101) <= b;
    layer6_outputs(6102) <= a and not b;
    layer6_outputs(6103) <= not (a xor b);
    layer6_outputs(6104) <= not a;
    layer6_outputs(6105) <= not a or b;
    layer6_outputs(6106) <= 1'b0;
    layer6_outputs(6107) <= not a;
    layer6_outputs(6108) <= b;
    layer6_outputs(6109) <= a;
    layer6_outputs(6110) <= b and not a;
    layer6_outputs(6111) <= not a or b;
    layer6_outputs(6112) <= a or b;
    layer6_outputs(6113) <= not b;
    layer6_outputs(6114) <= not a;
    layer6_outputs(6115) <= b;
    layer6_outputs(6116) <= not (a and b);
    layer6_outputs(6117) <= not (a xor b);
    layer6_outputs(6118) <= a and not b;
    layer6_outputs(6119) <= a xor b;
    layer6_outputs(6120) <= b and not a;
    layer6_outputs(6121) <= not a or b;
    layer6_outputs(6122) <= not a;
    layer6_outputs(6123) <= not a;
    layer6_outputs(6124) <= b;
    layer6_outputs(6125) <= not b;
    layer6_outputs(6126) <= not b;
    layer6_outputs(6127) <= 1'b0;
    layer6_outputs(6128) <= a or b;
    layer6_outputs(6129) <= not a or b;
    layer6_outputs(6130) <= a and not b;
    layer6_outputs(6131) <= 1'b0;
    layer6_outputs(6132) <= a;
    layer6_outputs(6133) <= a and b;
    layer6_outputs(6134) <= 1'b0;
    layer6_outputs(6135) <= not (a and b);
    layer6_outputs(6136) <= b;
    layer6_outputs(6137) <= not a or b;
    layer6_outputs(6138) <= a;
    layer6_outputs(6139) <= not a;
    layer6_outputs(6140) <= not (a or b);
    layer6_outputs(6141) <= not a;
    layer6_outputs(6142) <= a xor b;
    layer6_outputs(6143) <= b and not a;
    layer6_outputs(6144) <= a and b;
    layer6_outputs(6145) <= a and b;
    layer6_outputs(6146) <= a;
    layer6_outputs(6147) <= 1'b1;
    layer6_outputs(6148) <= not b;
    layer6_outputs(6149) <= not (a or b);
    layer6_outputs(6150) <= not (a and b);
    layer6_outputs(6151) <= a;
    layer6_outputs(6152) <= not b or a;
    layer6_outputs(6153) <= a and b;
    layer6_outputs(6154) <= a;
    layer6_outputs(6155) <= not b or a;
    layer6_outputs(6156) <= b;
    layer6_outputs(6157) <= not b or a;
    layer6_outputs(6158) <= b and not a;
    layer6_outputs(6159) <= b and not a;
    layer6_outputs(6160) <= a and not b;
    layer6_outputs(6161) <= b and not a;
    layer6_outputs(6162) <= not (a and b);
    layer6_outputs(6163) <= a;
    layer6_outputs(6164) <= a;
    layer6_outputs(6165) <= a and b;
    layer6_outputs(6166) <= not (a and b);
    layer6_outputs(6167) <= not a;
    layer6_outputs(6168) <= 1'b1;
    layer6_outputs(6169) <= a;
    layer6_outputs(6170) <= a and b;
    layer6_outputs(6171) <= not b or a;
    layer6_outputs(6172) <= not a or b;
    layer6_outputs(6173) <= a;
    layer6_outputs(6174) <= b and not a;
    layer6_outputs(6175) <= not (a xor b);
    layer6_outputs(6176) <= not a or b;
    layer6_outputs(6177) <= not (a or b);
    layer6_outputs(6178) <= not b;
    layer6_outputs(6179) <= not (a or b);
    layer6_outputs(6180) <= not b;
    layer6_outputs(6181) <= a and not b;
    layer6_outputs(6182) <= a and not b;
    layer6_outputs(6183) <= not a;
    layer6_outputs(6184) <= not b;
    layer6_outputs(6185) <= not a or b;
    layer6_outputs(6186) <= not (a xor b);
    layer6_outputs(6187) <= a and b;
    layer6_outputs(6188) <= b and not a;
    layer6_outputs(6189) <= not b;
    layer6_outputs(6190) <= not (a or b);
    layer6_outputs(6191) <= a;
    layer6_outputs(6192) <= not a or b;
    layer6_outputs(6193) <= not a;
    layer6_outputs(6194) <= a;
    layer6_outputs(6195) <= b;
    layer6_outputs(6196) <= not b;
    layer6_outputs(6197) <= not (a xor b);
    layer6_outputs(6198) <= not (a and b);
    layer6_outputs(6199) <= b;
    layer6_outputs(6200) <= a or b;
    layer6_outputs(6201) <= a and b;
    layer6_outputs(6202) <= a;
    layer6_outputs(6203) <= not b;
    layer6_outputs(6204) <= b;
    layer6_outputs(6205) <= not a;
    layer6_outputs(6206) <= a and b;
    layer6_outputs(6207) <= not a or b;
    layer6_outputs(6208) <= not b;
    layer6_outputs(6209) <= a and not b;
    layer6_outputs(6210) <= a;
    layer6_outputs(6211) <= not b;
    layer6_outputs(6212) <= not a or b;
    layer6_outputs(6213) <= not (a xor b);
    layer6_outputs(6214) <= not (a xor b);
    layer6_outputs(6215) <= not (a or b);
    layer6_outputs(6216) <= not (a or b);
    layer6_outputs(6217) <= a or b;
    layer6_outputs(6218) <= not (a and b);
    layer6_outputs(6219) <= a;
    layer6_outputs(6220) <= not (a xor b);
    layer6_outputs(6221) <= a and not b;
    layer6_outputs(6222) <= not b or a;
    layer6_outputs(6223) <= b;
    layer6_outputs(6224) <= not b or a;
    layer6_outputs(6225) <= not a;
    layer6_outputs(6226) <= b;
    layer6_outputs(6227) <= not b;
    layer6_outputs(6228) <= not (a xor b);
    layer6_outputs(6229) <= a or b;
    layer6_outputs(6230) <= not b;
    layer6_outputs(6231) <= a or b;
    layer6_outputs(6232) <= not (a and b);
    layer6_outputs(6233) <= b;
    layer6_outputs(6234) <= not (a or b);
    layer6_outputs(6235) <= not a;
    layer6_outputs(6236) <= a;
    layer6_outputs(6237) <= not a;
    layer6_outputs(6238) <= a and b;
    layer6_outputs(6239) <= a or b;
    layer6_outputs(6240) <= not b;
    layer6_outputs(6241) <= not b or a;
    layer6_outputs(6242) <= not a or b;
    layer6_outputs(6243) <= a;
    layer6_outputs(6244) <= not a;
    layer6_outputs(6245) <= not b;
    layer6_outputs(6246) <= a or b;
    layer6_outputs(6247) <= b and not a;
    layer6_outputs(6248) <= a;
    layer6_outputs(6249) <= not (a xor b);
    layer6_outputs(6250) <= b;
    layer6_outputs(6251) <= not (a or b);
    layer6_outputs(6252) <= not (a or b);
    layer6_outputs(6253) <= not b;
    layer6_outputs(6254) <= b and not a;
    layer6_outputs(6255) <= a;
    layer6_outputs(6256) <= a;
    layer6_outputs(6257) <= not (a and b);
    layer6_outputs(6258) <= a;
    layer6_outputs(6259) <= a;
    layer6_outputs(6260) <= not (a or b);
    layer6_outputs(6261) <= not a;
    layer6_outputs(6262) <= b;
    layer6_outputs(6263) <= a;
    layer6_outputs(6264) <= not b or a;
    layer6_outputs(6265) <= not a or b;
    layer6_outputs(6266) <= not (a or b);
    layer6_outputs(6267) <= not (a and b);
    layer6_outputs(6268) <= b;
    layer6_outputs(6269) <= not a;
    layer6_outputs(6270) <= not a;
    layer6_outputs(6271) <= b;
    layer6_outputs(6272) <= a;
    layer6_outputs(6273) <= 1'b0;
    layer6_outputs(6274) <= a and not b;
    layer6_outputs(6275) <= not (a xor b);
    layer6_outputs(6276) <= a and not b;
    layer6_outputs(6277) <= not (a xor b);
    layer6_outputs(6278) <= b;
    layer6_outputs(6279) <= not b;
    layer6_outputs(6280) <= b and not a;
    layer6_outputs(6281) <= a;
    layer6_outputs(6282) <= b;
    layer6_outputs(6283) <= b;
    layer6_outputs(6284) <= not (a or b);
    layer6_outputs(6285) <= b and not a;
    layer6_outputs(6286) <= not (a and b);
    layer6_outputs(6287) <= a;
    layer6_outputs(6288) <= not a;
    layer6_outputs(6289) <= not (a and b);
    layer6_outputs(6290) <= b and not a;
    layer6_outputs(6291) <= a or b;
    layer6_outputs(6292) <= b;
    layer6_outputs(6293) <= not a;
    layer6_outputs(6294) <= a xor b;
    layer6_outputs(6295) <= a or b;
    layer6_outputs(6296) <= b;
    layer6_outputs(6297) <= a and not b;
    layer6_outputs(6298) <= a and not b;
    layer6_outputs(6299) <= not a;
    layer6_outputs(6300) <= not (a xor b);
    layer6_outputs(6301) <= not (a or b);
    layer6_outputs(6302) <= not (a and b);
    layer6_outputs(6303) <= a xor b;
    layer6_outputs(6304) <= a;
    layer6_outputs(6305) <= b;
    layer6_outputs(6306) <= a;
    layer6_outputs(6307) <= a xor b;
    layer6_outputs(6308) <= not a;
    layer6_outputs(6309) <= a and b;
    layer6_outputs(6310) <= b and not a;
    layer6_outputs(6311) <= not a;
    layer6_outputs(6312) <= b;
    layer6_outputs(6313) <= not a;
    layer6_outputs(6314) <= a or b;
    layer6_outputs(6315) <= a and b;
    layer6_outputs(6316) <= not (a and b);
    layer6_outputs(6317) <= a or b;
    layer6_outputs(6318) <= not (a xor b);
    layer6_outputs(6319) <= not a;
    layer6_outputs(6320) <= not (a and b);
    layer6_outputs(6321) <= not (a or b);
    layer6_outputs(6322) <= not b;
    layer6_outputs(6323) <= not a;
    layer6_outputs(6324) <= not b;
    layer6_outputs(6325) <= not (a and b);
    layer6_outputs(6326) <= a and b;
    layer6_outputs(6327) <= not (a xor b);
    layer6_outputs(6328) <= a xor b;
    layer6_outputs(6329) <= not b;
    layer6_outputs(6330) <= 1'b0;
    layer6_outputs(6331) <= b;
    layer6_outputs(6332) <= a and b;
    layer6_outputs(6333) <= b;
    layer6_outputs(6334) <= b;
    layer6_outputs(6335) <= not (a and b);
    layer6_outputs(6336) <= not b;
    layer6_outputs(6337) <= a and not b;
    layer6_outputs(6338) <= a;
    layer6_outputs(6339) <= a;
    layer6_outputs(6340) <= 1'b1;
    layer6_outputs(6341) <= b;
    layer6_outputs(6342) <= 1'b0;
    layer6_outputs(6343) <= not (a xor b);
    layer6_outputs(6344) <= not b or a;
    layer6_outputs(6345) <= a;
    layer6_outputs(6346) <= not a;
    layer6_outputs(6347) <= a;
    layer6_outputs(6348) <= not (a and b);
    layer6_outputs(6349) <= not a;
    layer6_outputs(6350) <= not b or a;
    layer6_outputs(6351) <= a and not b;
    layer6_outputs(6352) <= 1'b0;
    layer6_outputs(6353) <= 1'b1;
    layer6_outputs(6354) <= a and b;
    layer6_outputs(6355) <= not a;
    layer6_outputs(6356) <= not a;
    layer6_outputs(6357) <= a xor b;
    layer6_outputs(6358) <= a or b;
    layer6_outputs(6359) <= 1'b1;
    layer6_outputs(6360) <= a and not b;
    layer6_outputs(6361) <= a or b;
    layer6_outputs(6362) <= a;
    layer6_outputs(6363) <= not b or a;
    layer6_outputs(6364) <= b;
    layer6_outputs(6365) <= b and not a;
    layer6_outputs(6366) <= not a;
    layer6_outputs(6367) <= b;
    layer6_outputs(6368) <= a or b;
    layer6_outputs(6369) <= a and not b;
    layer6_outputs(6370) <= b;
    layer6_outputs(6371) <= not b;
    layer6_outputs(6372) <= not b;
    layer6_outputs(6373) <= b;
    layer6_outputs(6374) <= a or b;
    layer6_outputs(6375) <= a and not b;
    layer6_outputs(6376) <= b;
    layer6_outputs(6377) <= a or b;
    layer6_outputs(6378) <= b;
    layer6_outputs(6379) <= b;
    layer6_outputs(6380) <= not a;
    layer6_outputs(6381) <= not b or a;
    layer6_outputs(6382) <= not b;
    layer6_outputs(6383) <= not (a or b);
    layer6_outputs(6384) <= not b or a;
    layer6_outputs(6385) <= a or b;
    layer6_outputs(6386) <= b and not a;
    layer6_outputs(6387) <= b;
    layer6_outputs(6388) <= a xor b;
    layer6_outputs(6389) <= not (a xor b);
    layer6_outputs(6390) <= b;
    layer6_outputs(6391) <= not (a xor b);
    layer6_outputs(6392) <= not a;
    layer6_outputs(6393) <= b;
    layer6_outputs(6394) <= not (a or b);
    layer6_outputs(6395) <= not (a xor b);
    layer6_outputs(6396) <= not b;
    layer6_outputs(6397) <= not (a xor b);
    layer6_outputs(6398) <= b;
    layer6_outputs(6399) <= 1'b0;
    layer6_outputs(6400) <= a or b;
    layer6_outputs(6401) <= a and not b;
    layer6_outputs(6402) <= not (a and b);
    layer6_outputs(6403) <= a and b;
    layer6_outputs(6404) <= b;
    layer6_outputs(6405) <= not b or a;
    layer6_outputs(6406) <= not a or b;
    layer6_outputs(6407) <= a;
    layer6_outputs(6408) <= not (a xor b);
    layer6_outputs(6409) <= a;
    layer6_outputs(6410) <= a and b;
    layer6_outputs(6411) <= 1'b0;
    layer6_outputs(6412) <= not (a or b);
    layer6_outputs(6413) <= not a;
    layer6_outputs(6414) <= b and not a;
    layer6_outputs(6415) <= a and b;
    layer6_outputs(6416) <= not b;
    layer6_outputs(6417) <= not a;
    layer6_outputs(6418) <= not a or b;
    layer6_outputs(6419) <= not b or a;
    layer6_outputs(6420) <= a;
    layer6_outputs(6421) <= b and not a;
    layer6_outputs(6422) <= not (a and b);
    layer6_outputs(6423) <= not b;
    layer6_outputs(6424) <= not a;
    layer6_outputs(6425) <= not a;
    layer6_outputs(6426) <= not (a xor b);
    layer6_outputs(6427) <= not (a xor b);
    layer6_outputs(6428) <= not b;
    layer6_outputs(6429) <= b;
    layer6_outputs(6430) <= b and not a;
    layer6_outputs(6431) <= not (a or b);
    layer6_outputs(6432) <= b and not a;
    layer6_outputs(6433) <= a and b;
    layer6_outputs(6434) <= 1'b0;
    layer6_outputs(6435) <= not a;
    layer6_outputs(6436) <= not b;
    layer6_outputs(6437) <= a and b;
    layer6_outputs(6438) <= a or b;
    layer6_outputs(6439) <= not a;
    layer6_outputs(6440) <= b and not a;
    layer6_outputs(6441) <= b;
    layer6_outputs(6442) <= not a;
    layer6_outputs(6443) <= not a;
    layer6_outputs(6444) <= not b or a;
    layer6_outputs(6445) <= not b or a;
    layer6_outputs(6446) <= 1'b0;
    layer6_outputs(6447) <= b;
    layer6_outputs(6448) <= not b or a;
    layer6_outputs(6449) <= b;
    layer6_outputs(6450) <= a;
    layer6_outputs(6451) <= not a or b;
    layer6_outputs(6452) <= not a;
    layer6_outputs(6453) <= not b;
    layer6_outputs(6454) <= a;
    layer6_outputs(6455) <= b;
    layer6_outputs(6456) <= not b;
    layer6_outputs(6457) <= b;
    layer6_outputs(6458) <= not (a and b);
    layer6_outputs(6459) <= not b;
    layer6_outputs(6460) <= a and b;
    layer6_outputs(6461) <= a;
    layer6_outputs(6462) <= b and not a;
    layer6_outputs(6463) <= a and b;
    layer6_outputs(6464) <= not (a and b);
    layer6_outputs(6465) <= not b;
    layer6_outputs(6466) <= a or b;
    layer6_outputs(6467) <= b;
    layer6_outputs(6468) <= b;
    layer6_outputs(6469) <= not a;
    layer6_outputs(6470) <= not a;
    layer6_outputs(6471) <= b;
    layer6_outputs(6472) <= not a or b;
    layer6_outputs(6473) <= not (a xor b);
    layer6_outputs(6474) <= a;
    layer6_outputs(6475) <= not (a or b);
    layer6_outputs(6476) <= a xor b;
    layer6_outputs(6477) <= a and b;
    layer6_outputs(6478) <= a xor b;
    layer6_outputs(6479) <= not b or a;
    layer6_outputs(6480) <= b and not a;
    layer6_outputs(6481) <= not (a xor b);
    layer6_outputs(6482) <= not a;
    layer6_outputs(6483) <= not b or a;
    layer6_outputs(6484) <= a;
    layer6_outputs(6485) <= a or b;
    layer6_outputs(6486) <= a;
    layer6_outputs(6487) <= not a or b;
    layer6_outputs(6488) <= not b;
    layer6_outputs(6489) <= not b;
    layer6_outputs(6490) <= not b or a;
    layer6_outputs(6491) <= not a;
    layer6_outputs(6492) <= a and b;
    layer6_outputs(6493) <= a xor b;
    layer6_outputs(6494) <= not a;
    layer6_outputs(6495) <= not a;
    layer6_outputs(6496) <= not a;
    layer6_outputs(6497) <= a and not b;
    layer6_outputs(6498) <= not (a and b);
    layer6_outputs(6499) <= a;
    layer6_outputs(6500) <= b and not a;
    layer6_outputs(6501) <= a xor b;
    layer6_outputs(6502) <= a or b;
    layer6_outputs(6503) <= b;
    layer6_outputs(6504) <= a or b;
    layer6_outputs(6505) <= a and b;
    layer6_outputs(6506) <= a and b;
    layer6_outputs(6507) <= not (a xor b);
    layer6_outputs(6508) <= not b;
    layer6_outputs(6509) <= not b;
    layer6_outputs(6510) <= b;
    layer6_outputs(6511) <= 1'b1;
    layer6_outputs(6512) <= not (a xor b);
    layer6_outputs(6513) <= b;
    layer6_outputs(6514) <= not (a and b);
    layer6_outputs(6515) <= b;
    layer6_outputs(6516) <= not (a or b);
    layer6_outputs(6517) <= a xor b;
    layer6_outputs(6518) <= a;
    layer6_outputs(6519) <= not (a xor b);
    layer6_outputs(6520) <= not b;
    layer6_outputs(6521) <= a;
    layer6_outputs(6522) <= not a;
    layer6_outputs(6523) <= a;
    layer6_outputs(6524) <= a or b;
    layer6_outputs(6525) <= a and b;
    layer6_outputs(6526) <= not (a or b);
    layer6_outputs(6527) <= not (a xor b);
    layer6_outputs(6528) <= b;
    layer6_outputs(6529) <= b and not a;
    layer6_outputs(6530) <= not a;
    layer6_outputs(6531) <= b;
    layer6_outputs(6532) <= a xor b;
    layer6_outputs(6533) <= not a;
    layer6_outputs(6534) <= not a or b;
    layer6_outputs(6535) <= a or b;
    layer6_outputs(6536) <= not b;
    layer6_outputs(6537) <= not (a xor b);
    layer6_outputs(6538) <= not (a xor b);
    layer6_outputs(6539) <= not (a xor b);
    layer6_outputs(6540) <= not b;
    layer6_outputs(6541) <= b and not a;
    layer6_outputs(6542) <= a xor b;
    layer6_outputs(6543) <= a xor b;
    layer6_outputs(6544) <= not a;
    layer6_outputs(6545) <= a and not b;
    layer6_outputs(6546) <= a and b;
    layer6_outputs(6547) <= 1'b0;
    layer6_outputs(6548) <= not b;
    layer6_outputs(6549) <= not (a and b);
    layer6_outputs(6550) <= b and not a;
    layer6_outputs(6551) <= not a or b;
    layer6_outputs(6552) <= a;
    layer6_outputs(6553) <= a;
    layer6_outputs(6554) <= b and not a;
    layer6_outputs(6555) <= a or b;
    layer6_outputs(6556) <= not a;
    layer6_outputs(6557) <= not (a or b);
    layer6_outputs(6558) <= not a or b;
    layer6_outputs(6559) <= a and b;
    layer6_outputs(6560) <= not a;
    layer6_outputs(6561) <= not b or a;
    layer6_outputs(6562) <= a;
    layer6_outputs(6563) <= a and b;
    layer6_outputs(6564) <= not a;
    layer6_outputs(6565) <= a;
    layer6_outputs(6566) <= a;
    layer6_outputs(6567) <= not b;
    layer6_outputs(6568) <= not a;
    layer6_outputs(6569) <= not a;
    layer6_outputs(6570) <= a and not b;
    layer6_outputs(6571) <= not b;
    layer6_outputs(6572) <= a or b;
    layer6_outputs(6573) <= not a;
    layer6_outputs(6574) <= not a;
    layer6_outputs(6575) <= a xor b;
    layer6_outputs(6576) <= not (a or b);
    layer6_outputs(6577) <= b and not a;
    layer6_outputs(6578) <= a and b;
    layer6_outputs(6579) <= not (a or b);
    layer6_outputs(6580) <= not a;
    layer6_outputs(6581) <= not (a and b);
    layer6_outputs(6582) <= not (a and b);
    layer6_outputs(6583) <= not a or b;
    layer6_outputs(6584) <= 1'b1;
    layer6_outputs(6585) <= not (a xor b);
    layer6_outputs(6586) <= b and not a;
    layer6_outputs(6587) <= b and not a;
    layer6_outputs(6588) <= not (a and b);
    layer6_outputs(6589) <= not a;
    layer6_outputs(6590) <= not (a and b);
    layer6_outputs(6591) <= not b;
    layer6_outputs(6592) <= not a;
    layer6_outputs(6593) <= a and b;
    layer6_outputs(6594) <= a and b;
    layer6_outputs(6595) <= a;
    layer6_outputs(6596) <= not (a xor b);
    layer6_outputs(6597) <= b and not a;
    layer6_outputs(6598) <= a xor b;
    layer6_outputs(6599) <= not a;
    layer6_outputs(6600) <= not b;
    layer6_outputs(6601) <= a and b;
    layer6_outputs(6602) <= a and not b;
    layer6_outputs(6603) <= not b;
    layer6_outputs(6604) <= b;
    layer6_outputs(6605) <= a;
    layer6_outputs(6606) <= 1'b0;
    layer6_outputs(6607) <= not (a and b);
    layer6_outputs(6608) <= b;
    layer6_outputs(6609) <= a and not b;
    layer6_outputs(6610) <= a;
    layer6_outputs(6611) <= not b or a;
    layer6_outputs(6612) <= a and not b;
    layer6_outputs(6613) <= not a;
    layer6_outputs(6614) <= 1'b1;
    layer6_outputs(6615) <= a xor b;
    layer6_outputs(6616) <= b and not a;
    layer6_outputs(6617) <= not (a and b);
    layer6_outputs(6618) <= b;
    layer6_outputs(6619) <= not (a or b);
    layer6_outputs(6620) <= a and b;
    layer6_outputs(6621) <= not a;
    layer6_outputs(6622) <= not (a and b);
    layer6_outputs(6623) <= not a;
    layer6_outputs(6624) <= b;
    layer6_outputs(6625) <= not (a and b);
    layer6_outputs(6626) <= a;
    layer6_outputs(6627) <= not (a xor b);
    layer6_outputs(6628) <= not b;
    layer6_outputs(6629) <= a and b;
    layer6_outputs(6630) <= not a or b;
    layer6_outputs(6631) <= b;
    layer6_outputs(6632) <= not b;
    layer6_outputs(6633) <= a xor b;
    layer6_outputs(6634) <= a and not b;
    layer6_outputs(6635) <= not a or b;
    layer6_outputs(6636) <= a and b;
    layer6_outputs(6637) <= b;
    layer6_outputs(6638) <= not (a or b);
    layer6_outputs(6639) <= a and b;
    layer6_outputs(6640) <= not (a and b);
    layer6_outputs(6641) <= not (a xor b);
    layer6_outputs(6642) <= not (a or b);
    layer6_outputs(6643) <= not b;
    layer6_outputs(6644) <= not a;
    layer6_outputs(6645) <= not a;
    layer6_outputs(6646) <= a;
    layer6_outputs(6647) <= not a;
    layer6_outputs(6648) <= a;
    layer6_outputs(6649) <= not (a and b);
    layer6_outputs(6650) <= not a;
    layer6_outputs(6651) <= 1'b0;
    layer6_outputs(6652) <= a and b;
    layer6_outputs(6653) <= a;
    layer6_outputs(6654) <= b and not a;
    layer6_outputs(6655) <= a and not b;
    layer6_outputs(6656) <= not a;
    layer6_outputs(6657) <= not (a or b);
    layer6_outputs(6658) <= a and b;
    layer6_outputs(6659) <= a xor b;
    layer6_outputs(6660) <= b;
    layer6_outputs(6661) <= not a or b;
    layer6_outputs(6662) <= 1'b0;
    layer6_outputs(6663) <= not a;
    layer6_outputs(6664) <= a;
    layer6_outputs(6665) <= a and not b;
    layer6_outputs(6666) <= a or b;
    layer6_outputs(6667) <= not a or b;
    layer6_outputs(6668) <= b and not a;
    layer6_outputs(6669) <= a and b;
    layer6_outputs(6670) <= not (a and b);
    layer6_outputs(6671) <= not a;
    layer6_outputs(6672) <= not b or a;
    layer6_outputs(6673) <= b;
    layer6_outputs(6674) <= b and not a;
    layer6_outputs(6675) <= not b or a;
    layer6_outputs(6676) <= a xor b;
    layer6_outputs(6677) <= a and not b;
    layer6_outputs(6678) <= not a;
    layer6_outputs(6679) <= not (a and b);
    layer6_outputs(6680) <= b;
    layer6_outputs(6681) <= not b;
    layer6_outputs(6682) <= not (a or b);
    layer6_outputs(6683) <= a and not b;
    layer6_outputs(6684) <= not a or b;
    layer6_outputs(6685) <= not a or b;
    layer6_outputs(6686) <= a;
    layer6_outputs(6687) <= not b;
    layer6_outputs(6688) <= b;
    layer6_outputs(6689) <= not (a or b);
    layer6_outputs(6690) <= not a;
    layer6_outputs(6691) <= a or b;
    layer6_outputs(6692) <= not a;
    layer6_outputs(6693) <= not (a and b);
    layer6_outputs(6694) <= not (a xor b);
    layer6_outputs(6695) <= not a;
    layer6_outputs(6696) <= 1'b1;
    layer6_outputs(6697) <= 1'b0;
    layer6_outputs(6698) <= not a or b;
    layer6_outputs(6699) <= not a or b;
    layer6_outputs(6700) <= a;
    layer6_outputs(6701) <= not (a and b);
    layer6_outputs(6702) <= a and b;
    layer6_outputs(6703) <= not (a xor b);
    layer6_outputs(6704) <= not b or a;
    layer6_outputs(6705) <= b and not a;
    layer6_outputs(6706) <= a and b;
    layer6_outputs(6707) <= not a;
    layer6_outputs(6708) <= b and not a;
    layer6_outputs(6709) <= b;
    layer6_outputs(6710) <= not a;
    layer6_outputs(6711) <= not (a xor b);
    layer6_outputs(6712) <= not a;
    layer6_outputs(6713) <= 1'b1;
    layer6_outputs(6714) <= not a;
    layer6_outputs(6715) <= not b;
    layer6_outputs(6716) <= not b;
    layer6_outputs(6717) <= b;
    layer6_outputs(6718) <= not (a and b);
    layer6_outputs(6719) <= not a;
    layer6_outputs(6720) <= not b or a;
    layer6_outputs(6721) <= not (a or b);
    layer6_outputs(6722) <= not a;
    layer6_outputs(6723) <= not (a and b);
    layer6_outputs(6724) <= b;
    layer6_outputs(6725) <= b;
    layer6_outputs(6726) <= a xor b;
    layer6_outputs(6727) <= b;
    layer6_outputs(6728) <= b;
    layer6_outputs(6729) <= not a;
    layer6_outputs(6730) <= not b;
    layer6_outputs(6731) <= not a or b;
    layer6_outputs(6732) <= not a;
    layer6_outputs(6733) <= a and b;
    layer6_outputs(6734) <= b;
    layer6_outputs(6735) <= a and not b;
    layer6_outputs(6736) <= a and b;
    layer6_outputs(6737) <= a and not b;
    layer6_outputs(6738) <= not (a or b);
    layer6_outputs(6739) <= a;
    layer6_outputs(6740) <= 1'b0;
    layer6_outputs(6741) <= not b;
    layer6_outputs(6742) <= a and not b;
    layer6_outputs(6743) <= 1'b0;
    layer6_outputs(6744) <= b;
    layer6_outputs(6745) <= not (a and b);
    layer6_outputs(6746) <= not (a xor b);
    layer6_outputs(6747) <= not a or b;
    layer6_outputs(6748) <= b;
    layer6_outputs(6749) <= a xor b;
    layer6_outputs(6750) <= not (a and b);
    layer6_outputs(6751) <= not a;
    layer6_outputs(6752) <= b;
    layer6_outputs(6753) <= not (a xor b);
    layer6_outputs(6754) <= not (a or b);
    layer6_outputs(6755) <= not a or b;
    layer6_outputs(6756) <= a and b;
    layer6_outputs(6757) <= not (a or b);
    layer6_outputs(6758) <= not b;
    layer6_outputs(6759) <= a and not b;
    layer6_outputs(6760) <= not a;
    layer6_outputs(6761) <= a and not b;
    layer6_outputs(6762) <= a or b;
    layer6_outputs(6763) <= a and b;
    layer6_outputs(6764) <= not b;
    layer6_outputs(6765) <= not (a xor b);
    layer6_outputs(6766) <= not (a or b);
    layer6_outputs(6767) <= a xor b;
    layer6_outputs(6768) <= a;
    layer6_outputs(6769) <= not a;
    layer6_outputs(6770) <= b and not a;
    layer6_outputs(6771) <= a xor b;
    layer6_outputs(6772) <= a and not b;
    layer6_outputs(6773) <= a xor b;
    layer6_outputs(6774) <= a or b;
    layer6_outputs(6775) <= not a;
    layer6_outputs(6776) <= b and not a;
    layer6_outputs(6777) <= a xor b;
    layer6_outputs(6778) <= not (a or b);
    layer6_outputs(6779) <= b and not a;
    layer6_outputs(6780) <= not (a or b);
    layer6_outputs(6781) <= not b;
    layer6_outputs(6782) <= not b or a;
    layer6_outputs(6783) <= 1'b1;
    layer6_outputs(6784) <= a;
    layer6_outputs(6785) <= not b;
    layer6_outputs(6786) <= b;
    layer6_outputs(6787) <= not a;
    layer6_outputs(6788) <= not a;
    layer6_outputs(6789) <= not b;
    layer6_outputs(6790) <= a;
    layer6_outputs(6791) <= not b or a;
    layer6_outputs(6792) <= b and not a;
    layer6_outputs(6793) <= a and b;
    layer6_outputs(6794) <= a;
    layer6_outputs(6795) <= a and not b;
    layer6_outputs(6796) <= a or b;
    layer6_outputs(6797) <= b;
    layer6_outputs(6798) <= a or b;
    layer6_outputs(6799) <= a;
    layer6_outputs(6800) <= not b or a;
    layer6_outputs(6801) <= b;
    layer6_outputs(6802) <= not (a xor b);
    layer6_outputs(6803) <= b and not a;
    layer6_outputs(6804) <= not (a or b);
    layer6_outputs(6805) <= a or b;
    layer6_outputs(6806) <= a and not b;
    layer6_outputs(6807) <= 1'b0;
    layer6_outputs(6808) <= b;
    layer6_outputs(6809) <= 1'b0;
    layer6_outputs(6810) <= a;
    layer6_outputs(6811) <= b;
    layer6_outputs(6812) <= not a or b;
    layer6_outputs(6813) <= b;
    layer6_outputs(6814) <= b and not a;
    layer6_outputs(6815) <= not a;
    layer6_outputs(6816) <= not a or b;
    layer6_outputs(6817) <= not a or b;
    layer6_outputs(6818) <= not (a xor b);
    layer6_outputs(6819) <= not b;
    layer6_outputs(6820) <= b;
    layer6_outputs(6821) <= a or b;
    layer6_outputs(6822) <= not b or a;
    layer6_outputs(6823) <= not a or b;
    layer6_outputs(6824) <= a or b;
    layer6_outputs(6825) <= b;
    layer6_outputs(6826) <= 1'b0;
    layer6_outputs(6827) <= not a or b;
    layer6_outputs(6828) <= not b;
    layer6_outputs(6829) <= not a;
    layer6_outputs(6830) <= a and b;
    layer6_outputs(6831) <= a or b;
    layer6_outputs(6832) <= not a;
    layer6_outputs(6833) <= b;
    layer6_outputs(6834) <= a and not b;
    layer6_outputs(6835) <= a;
    layer6_outputs(6836) <= not b;
    layer6_outputs(6837) <= not b;
    layer6_outputs(6838) <= not (a and b);
    layer6_outputs(6839) <= a;
    layer6_outputs(6840) <= not b;
    layer6_outputs(6841) <= not (a and b);
    layer6_outputs(6842) <= b;
    layer6_outputs(6843) <= not a;
    layer6_outputs(6844) <= a and b;
    layer6_outputs(6845) <= not (a or b);
    layer6_outputs(6846) <= a or b;
    layer6_outputs(6847) <= b;
    layer6_outputs(6848) <= not a;
    layer6_outputs(6849) <= a or b;
    layer6_outputs(6850) <= not (a and b);
    layer6_outputs(6851) <= a and b;
    layer6_outputs(6852) <= b;
    layer6_outputs(6853) <= b and not a;
    layer6_outputs(6854) <= not b or a;
    layer6_outputs(6855) <= not (a xor b);
    layer6_outputs(6856) <= not b;
    layer6_outputs(6857) <= not a or b;
    layer6_outputs(6858) <= not (a xor b);
    layer6_outputs(6859) <= not b;
    layer6_outputs(6860) <= not b or a;
    layer6_outputs(6861) <= not (a or b);
    layer6_outputs(6862) <= a and not b;
    layer6_outputs(6863) <= a xor b;
    layer6_outputs(6864) <= not a;
    layer6_outputs(6865) <= not a;
    layer6_outputs(6866) <= a and not b;
    layer6_outputs(6867) <= a and b;
    layer6_outputs(6868) <= a;
    layer6_outputs(6869) <= not b;
    layer6_outputs(6870) <= b;
    layer6_outputs(6871) <= not a or b;
    layer6_outputs(6872) <= b;
    layer6_outputs(6873) <= not a or b;
    layer6_outputs(6874) <= 1'b0;
    layer6_outputs(6875) <= not a;
    layer6_outputs(6876) <= 1'b0;
    layer6_outputs(6877) <= not b or a;
    layer6_outputs(6878) <= not a;
    layer6_outputs(6879) <= not (a xor b);
    layer6_outputs(6880) <= b and not a;
    layer6_outputs(6881) <= b and not a;
    layer6_outputs(6882) <= b;
    layer6_outputs(6883) <= not (a and b);
    layer6_outputs(6884) <= a and not b;
    layer6_outputs(6885) <= a;
    layer6_outputs(6886) <= a;
    layer6_outputs(6887) <= not a;
    layer6_outputs(6888) <= b;
    layer6_outputs(6889) <= a xor b;
    layer6_outputs(6890) <= a or b;
    layer6_outputs(6891) <= 1'b0;
    layer6_outputs(6892) <= a xor b;
    layer6_outputs(6893) <= not (a and b);
    layer6_outputs(6894) <= not a;
    layer6_outputs(6895) <= a and not b;
    layer6_outputs(6896) <= b;
    layer6_outputs(6897) <= 1'b1;
    layer6_outputs(6898) <= a xor b;
    layer6_outputs(6899) <= not (a and b);
    layer6_outputs(6900) <= b;
    layer6_outputs(6901) <= not (a or b);
    layer6_outputs(6902) <= not a;
    layer6_outputs(6903) <= not a;
    layer6_outputs(6904) <= not (a and b);
    layer6_outputs(6905) <= not (a and b);
    layer6_outputs(6906) <= not a;
    layer6_outputs(6907) <= a;
    layer6_outputs(6908) <= a and b;
    layer6_outputs(6909) <= not a or b;
    layer6_outputs(6910) <= not a or b;
    layer6_outputs(6911) <= not a;
    layer6_outputs(6912) <= not b;
    layer6_outputs(6913) <= not b or a;
    layer6_outputs(6914) <= not b;
    layer6_outputs(6915) <= not b;
    layer6_outputs(6916) <= 1'b1;
    layer6_outputs(6917) <= not (a or b);
    layer6_outputs(6918) <= b;
    layer6_outputs(6919) <= a and b;
    layer6_outputs(6920) <= not b;
    layer6_outputs(6921) <= a;
    layer6_outputs(6922) <= 1'b1;
    layer6_outputs(6923) <= a;
    layer6_outputs(6924) <= not b;
    layer6_outputs(6925) <= a;
    layer6_outputs(6926) <= a or b;
    layer6_outputs(6927) <= not b;
    layer6_outputs(6928) <= not (a and b);
    layer6_outputs(6929) <= not b or a;
    layer6_outputs(6930) <= a and b;
    layer6_outputs(6931) <= not a;
    layer6_outputs(6932) <= not a or b;
    layer6_outputs(6933) <= not (a and b);
    layer6_outputs(6934) <= not b;
    layer6_outputs(6935) <= a and b;
    layer6_outputs(6936) <= b and not a;
    layer6_outputs(6937) <= not (a and b);
    layer6_outputs(6938) <= not a;
    layer6_outputs(6939) <= not b;
    layer6_outputs(6940) <= not (a xor b);
    layer6_outputs(6941) <= b;
    layer6_outputs(6942) <= not (a and b);
    layer6_outputs(6943) <= not b;
    layer6_outputs(6944) <= a xor b;
    layer6_outputs(6945) <= not (a or b);
    layer6_outputs(6946) <= not a or b;
    layer6_outputs(6947) <= b and not a;
    layer6_outputs(6948) <= not b or a;
    layer6_outputs(6949) <= not a;
    layer6_outputs(6950) <= a;
    layer6_outputs(6951) <= not b;
    layer6_outputs(6952) <= not a;
    layer6_outputs(6953) <= a or b;
    layer6_outputs(6954) <= a;
    layer6_outputs(6955) <= not a;
    layer6_outputs(6956) <= not (a and b);
    layer6_outputs(6957) <= not (a and b);
    layer6_outputs(6958) <= not (a or b);
    layer6_outputs(6959) <= not (a or b);
    layer6_outputs(6960) <= b and not a;
    layer6_outputs(6961) <= not (a xor b);
    layer6_outputs(6962) <= not a or b;
    layer6_outputs(6963) <= not b;
    layer6_outputs(6964) <= not b;
    layer6_outputs(6965) <= not b;
    layer6_outputs(6966) <= not a;
    layer6_outputs(6967) <= a and b;
    layer6_outputs(6968) <= not b;
    layer6_outputs(6969) <= not a;
    layer6_outputs(6970) <= not b;
    layer6_outputs(6971) <= b;
    layer6_outputs(6972) <= b and not a;
    layer6_outputs(6973) <= not b;
    layer6_outputs(6974) <= not b;
    layer6_outputs(6975) <= not (a xor b);
    layer6_outputs(6976) <= not (a and b);
    layer6_outputs(6977) <= a and not b;
    layer6_outputs(6978) <= not b;
    layer6_outputs(6979) <= not b;
    layer6_outputs(6980) <= b;
    layer6_outputs(6981) <= not (a or b);
    layer6_outputs(6982) <= a;
    layer6_outputs(6983) <= not (a or b);
    layer6_outputs(6984) <= not a;
    layer6_outputs(6985) <= a xor b;
    layer6_outputs(6986) <= not b or a;
    layer6_outputs(6987) <= not a or b;
    layer6_outputs(6988) <= a and b;
    layer6_outputs(6989) <= b and not a;
    layer6_outputs(6990) <= a and not b;
    layer6_outputs(6991) <= not b or a;
    layer6_outputs(6992) <= not (a or b);
    layer6_outputs(6993) <= b;
    layer6_outputs(6994) <= not a;
    layer6_outputs(6995) <= not (a and b);
    layer6_outputs(6996) <= b;
    layer6_outputs(6997) <= not b or a;
    layer6_outputs(6998) <= b and not a;
    layer6_outputs(6999) <= not (a and b);
    layer6_outputs(7000) <= not a;
    layer6_outputs(7001) <= a and b;
    layer6_outputs(7002) <= a;
    layer6_outputs(7003) <= not (a and b);
    layer6_outputs(7004) <= a xor b;
    layer6_outputs(7005) <= b;
    layer6_outputs(7006) <= a and b;
    layer6_outputs(7007) <= a;
    layer6_outputs(7008) <= not (a or b);
    layer6_outputs(7009) <= not a or b;
    layer6_outputs(7010) <= not b or a;
    layer6_outputs(7011) <= a;
    layer6_outputs(7012) <= not (a and b);
    layer6_outputs(7013) <= not (a or b);
    layer6_outputs(7014) <= a and not b;
    layer6_outputs(7015) <= a xor b;
    layer6_outputs(7016) <= b and not a;
    layer6_outputs(7017) <= a and b;
    layer6_outputs(7018) <= a xor b;
    layer6_outputs(7019) <= a;
    layer6_outputs(7020) <= 1'b1;
    layer6_outputs(7021) <= a and not b;
    layer6_outputs(7022) <= b;
    layer6_outputs(7023) <= b;
    layer6_outputs(7024) <= not b;
    layer6_outputs(7025) <= a or b;
    layer6_outputs(7026) <= a or b;
    layer6_outputs(7027) <= a or b;
    layer6_outputs(7028) <= a;
    layer6_outputs(7029) <= not b or a;
    layer6_outputs(7030) <= not (a or b);
    layer6_outputs(7031) <= not b;
    layer6_outputs(7032) <= not (a or b);
    layer6_outputs(7033) <= a and not b;
    layer6_outputs(7034) <= not (a xor b);
    layer6_outputs(7035) <= a and b;
    layer6_outputs(7036) <= a xor b;
    layer6_outputs(7037) <= not b;
    layer6_outputs(7038) <= a or b;
    layer6_outputs(7039) <= not b or a;
    layer6_outputs(7040) <= not b;
    layer6_outputs(7041) <= not (a and b);
    layer6_outputs(7042) <= not (a and b);
    layer6_outputs(7043) <= a and b;
    layer6_outputs(7044) <= b;
    layer6_outputs(7045) <= a;
    layer6_outputs(7046) <= not a;
    layer6_outputs(7047) <= b and not a;
    layer6_outputs(7048) <= not a;
    layer6_outputs(7049) <= not (a xor b);
    layer6_outputs(7050) <= not b;
    layer6_outputs(7051) <= b;
    layer6_outputs(7052) <= not a or b;
    layer6_outputs(7053) <= 1'b0;
    layer6_outputs(7054) <= b;
    layer6_outputs(7055) <= b;
    layer6_outputs(7056) <= b and not a;
    layer6_outputs(7057) <= b and not a;
    layer6_outputs(7058) <= not (a or b);
    layer6_outputs(7059) <= a xor b;
    layer6_outputs(7060) <= not a;
    layer6_outputs(7061) <= not (a xor b);
    layer6_outputs(7062) <= b and not a;
    layer6_outputs(7063) <= b;
    layer6_outputs(7064) <= not a;
    layer6_outputs(7065) <= a and b;
    layer6_outputs(7066) <= a or b;
    layer6_outputs(7067) <= not b or a;
    layer6_outputs(7068) <= not (a or b);
    layer6_outputs(7069) <= not a;
    layer6_outputs(7070) <= not b or a;
    layer6_outputs(7071) <= a and b;
    layer6_outputs(7072) <= not a;
    layer6_outputs(7073) <= not b;
    layer6_outputs(7074) <= b and not a;
    layer6_outputs(7075) <= not b or a;
    layer6_outputs(7076) <= a or b;
    layer6_outputs(7077) <= b and not a;
    layer6_outputs(7078) <= not (a xor b);
    layer6_outputs(7079) <= a xor b;
    layer6_outputs(7080) <= b;
    layer6_outputs(7081) <= b;
    layer6_outputs(7082) <= a;
    layer6_outputs(7083) <= not (a xor b);
    layer6_outputs(7084) <= a;
    layer6_outputs(7085) <= a xor b;
    layer6_outputs(7086) <= a;
    layer6_outputs(7087) <= a or b;
    layer6_outputs(7088) <= not b;
    layer6_outputs(7089) <= not b;
    layer6_outputs(7090) <= a and not b;
    layer6_outputs(7091) <= not a;
    layer6_outputs(7092) <= a;
    layer6_outputs(7093) <= not (a xor b);
    layer6_outputs(7094) <= not b or a;
    layer6_outputs(7095) <= a;
    layer6_outputs(7096) <= a xor b;
    layer6_outputs(7097) <= not a;
    layer6_outputs(7098) <= a and not b;
    layer6_outputs(7099) <= not b;
    layer6_outputs(7100) <= a and not b;
    layer6_outputs(7101) <= a xor b;
    layer6_outputs(7102) <= a and b;
    layer6_outputs(7103) <= not (a or b);
    layer6_outputs(7104) <= a;
    layer6_outputs(7105) <= not (a and b);
    layer6_outputs(7106) <= b;
    layer6_outputs(7107) <= a and b;
    layer6_outputs(7108) <= a xor b;
    layer6_outputs(7109) <= not b;
    layer6_outputs(7110) <= b and not a;
    layer6_outputs(7111) <= a;
    layer6_outputs(7112) <= not a;
    layer6_outputs(7113) <= a;
    layer6_outputs(7114) <= not a;
    layer6_outputs(7115) <= not b or a;
    layer6_outputs(7116) <= not a;
    layer6_outputs(7117) <= 1'b1;
    layer6_outputs(7118) <= a and not b;
    layer6_outputs(7119) <= not (a or b);
    layer6_outputs(7120) <= a and b;
    layer6_outputs(7121) <= not a;
    layer6_outputs(7122) <= a;
    layer6_outputs(7123) <= not b;
    layer6_outputs(7124) <= not a;
    layer6_outputs(7125) <= a;
    layer6_outputs(7126) <= a;
    layer6_outputs(7127) <= not b;
    layer6_outputs(7128) <= not b or a;
    layer6_outputs(7129) <= not b;
    layer6_outputs(7130) <= not (a and b);
    layer6_outputs(7131) <= a and not b;
    layer6_outputs(7132) <= not (a or b);
    layer6_outputs(7133) <= a or b;
    layer6_outputs(7134) <= not a;
    layer6_outputs(7135) <= b;
    layer6_outputs(7136) <= a xor b;
    layer6_outputs(7137) <= b;
    layer6_outputs(7138) <= not (a or b);
    layer6_outputs(7139) <= not b or a;
    layer6_outputs(7140) <= not (a xor b);
    layer6_outputs(7141) <= a and b;
    layer6_outputs(7142) <= not b;
    layer6_outputs(7143) <= a;
    layer6_outputs(7144) <= b and not a;
    layer6_outputs(7145) <= a;
    layer6_outputs(7146) <= b and not a;
    layer6_outputs(7147) <= not b;
    layer6_outputs(7148) <= b;
    layer6_outputs(7149) <= not (a xor b);
    layer6_outputs(7150) <= a xor b;
    layer6_outputs(7151) <= b;
    layer6_outputs(7152) <= not b;
    layer6_outputs(7153) <= 1'b1;
    layer6_outputs(7154) <= a and not b;
    layer6_outputs(7155) <= not (a and b);
    layer6_outputs(7156) <= not a;
    layer6_outputs(7157) <= not a;
    layer6_outputs(7158) <= not b;
    layer6_outputs(7159) <= not (a xor b);
    layer6_outputs(7160) <= a and not b;
    layer6_outputs(7161) <= not a;
    layer6_outputs(7162) <= not b;
    layer6_outputs(7163) <= not a;
    layer6_outputs(7164) <= not (a and b);
    layer6_outputs(7165) <= not b;
    layer6_outputs(7166) <= not (a and b);
    layer6_outputs(7167) <= not b;
    layer6_outputs(7168) <= not b;
    layer6_outputs(7169) <= b and not a;
    layer6_outputs(7170) <= not b;
    layer6_outputs(7171) <= b;
    layer6_outputs(7172) <= b;
    layer6_outputs(7173) <= b;
    layer6_outputs(7174) <= b and not a;
    layer6_outputs(7175) <= a;
    layer6_outputs(7176) <= b;
    layer6_outputs(7177) <= a and b;
    layer6_outputs(7178) <= not b;
    layer6_outputs(7179) <= b;
    layer6_outputs(7180) <= not (a xor b);
    layer6_outputs(7181) <= a;
    layer6_outputs(7182) <= not a or b;
    layer6_outputs(7183) <= not (a xor b);
    layer6_outputs(7184) <= not b;
    layer6_outputs(7185) <= not (a xor b);
    layer6_outputs(7186) <= b;
    layer6_outputs(7187) <= b and not a;
    layer6_outputs(7188) <= a;
    layer6_outputs(7189) <= not (a and b);
    layer6_outputs(7190) <= a and not b;
    layer6_outputs(7191) <= a;
    layer6_outputs(7192) <= not a;
    layer6_outputs(7193) <= not a;
    layer6_outputs(7194) <= not a;
    layer6_outputs(7195) <= not (a and b);
    layer6_outputs(7196) <= a;
    layer6_outputs(7197) <= a or b;
    layer6_outputs(7198) <= b;
    layer6_outputs(7199) <= not a;
    layer6_outputs(7200) <= not b or a;
    layer6_outputs(7201) <= not (a or b);
    layer6_outputs(7202) <= not b;
    layer6_outputs(7203) <= not a;
    layer6_outputs(7204) <= a and not b;
    layer6_outputs(7205) <= a and not b;
    layer6_outputs(7206) <= a;
    layer6_outputs(7207) <= not b or a;
    layer6_outputs(7208) <= not b or a;
    layer6_outputs(7209) <= not (a xor b);
    layer6_outputs(7210) <= not b;
    layer6_outputs(7211) <= not b or a;
    layer6_outputs(7212) <= not (a xor b);
    layer6_outputs(7213) <= not a;
    layer6_outputs(7214) <= a or b;
    layer6_outputs(7215) <= not (a or b);
    layer6_outputs(7216) <= not b;
    layer6_outputs(7217) <= a and not b;
    layer6_outputs(7218) <= a;
    layer6_outputs(7219) <= not b;
    layer6_outputs(7220) <= not a or b;
    layer6_outputs(7221) <= a or b;
    layer6_outputs(7222) <= not a;
    layer6_outputs(7223) <= 1'b0;
    layer6_outputs(7224) <= b;
    layer6_outputs(7225) <= not a;
    layer6_outputs(7226) <= not (a xor b);
    layer6_outputs(7227) <= a or b;
    layer6_outputs(7228) <= a xor b;
    layer6_outputs(7229) <= a or b;
    layer6_outputs(7230) <= not a or b;
    layer6_outputs(7231) <= a;
    layer6_outputs(7232) <= b;
    layer6_outputs(7233) <= b;
    layer6_outputs(7234) <= not b;
    layer6_outputs(7235) <= not (a and b);
    layer6_outputs(7236) <= b and not a;
    layer6_outputs(7237) <= b;
    layer6_outputs(7238) <= b and not a;
    layer6_outputs(7239) <= not a;
    layer6_outputs(7240) <= a xor b;
    layer6_outputs(7241) <= not a;
    layer6_outputs(7242) <= not a or b;
    layer6_outputs(7243) <= not (a xor b);
    layer6_outputs(7244) <= 1'b1;
    layer6_outputs(7245) <= a and not b;
    layer6_outputs(7246) <= not a;
    layer6_outputs(7247) <= a and not b;
    layer6_outputs(7248) <= a xor b;
    layer6_outputs(7249) <= a and b;
    layer6_outputs(7250) <= not (a and b);
    layer6_outputs(7251) <= b;
    layer6_outputs(7252) <= not (a and b);
    layer6_outputs(7253) <= not a;
    layer6_outputs(7254) <= a;
    layer6_outputs(7255) <= a and b;
    layer6_outputs(7256) <= a or b;
    layer6_outputs(7257) <= a;
    layer6_outputs(7258) <= 1'b0;
    layer6_outputs(7259) <= a and b;
    layer6_outputs(7260) <= a;
    layer6_outputs(7261) <= b;
    layer6_outputs(7262) <= not (a and b);
    layer6_outputs(7263) <= a and b;
    layer6_outputs(7264) <= a and not b;
    layer6_outputs(7265) <= not b;
    layer6_outputs(7266) <= a;
    layer6_outputs(7267) <= a or b;
    layer6_outputs(7268) <= not a;
    layer6_outputs(7269) <= 1'b0;
    layer6_outputs(7270) <= a xor b;
    layer6_outputs(7271) <= a and b;
    layer6_outputs(7272) <= a and b;
    layer6_outputs(7273) <= a;
    layer6_outputs(7274) <= b and not a;
    layer6_outputs(7275) <= b;
    layer6_outputs(7276) <= not a;
    layer6_outputs(7277) <= a or b;
    layer6_outputs(7278) <= not a;
    layer6_outputs(7279) <= a xor b;
    layer6_outputs(7280) <= not a;
    layer6_outputs(7281) <= b and not a;
    layer6_outputs(7282) <= b;
    layer6_outputs(7283) <= b and not a;
    layer6_outputs(7284) <= b;
    layer6_outputs(7285) <= b;
    layer6_outputs(7286) <= a or b;
    layer6_outputs(7287) <= 1'b0;
    layer6_outputs(7288) <= not (a or b);
    layer6_outputs(7289) <= not (a or b);
    layer6_outputs(7290) <= not a;
    layer6_outputs(7291) <= not a;
    layer6_outputs(7292) <= not a;
    layer6_outputs(7293) <= not b;
    layer6_outputs(7294) <= not (a or b);
    layer6_outputs(7295) <= a;
    layer6_outputs(7296) <= b and not a;
    layer6_outputs(7297) <= a;
    layer6_outputs(7298) <= not b;
    layer6_outputs(7299) <= not b or a;
    layer6_outputs(7300) <= not (a xor b);
    layer6_outputs(7301) <= not (a xor b);
    layer6_outputs(7302) <= b;
    layer6_outputs(7303) <= not a or b;
    layer6_outputs(7304) <= not (a xor b);
    layer6_outputs(7305) <= b;
    layer6_outputs(7306) <= not b;
    layer6_outputs(7307) <= a and not b;
    layer6_outputs(7308) <= not a or b;
    layer6_outputs(7309) <= not (a xor b);
    layer6_outputs(7310) <= b;
    layer6_outputs(7311) <= not (a xor b);
    layer6_outputs(7312) <= not a;
    layer6_outputs(7313) <= not (a and b);
    layer6_outputs(7314) <= not (a xor b);
    layer6_outputs(7315) <= a xor b;
    layer6_outputs(7316) <= not b;
    layer6_outputs(7317) <= a and not b;
    layer6_outputs(7318) <= not a or b;
    layer6_outputs(7319) <= not b or a;
    layer6_outputs(7320) <= not (a and b);
    layer6_outputs(7321) <= 1'b0;
    layer6_outputs(7322) <= b and not a;
    layer6_outputs(7323) <= a and not b;
    layer6_outputs(7324) <= not a;
    layer6_outputs(7325) <= b;
    layer6_outputs(7326) <= not (a and b);
    layer6_outputs(7327) <= a and b;
    layer6_outputs(7328) <= a;
    layer6_outputs(7329) <= b and not a;
    layer6_outputs(7330) <= not b;
    layer6_outputs(7331) <= not a or b;
    layer6_outputs(7332) <= not a;
    layer6_outputs(7333) <= b;
    layer6_outputs(7334) <= a;
    layer6_outputs(7335) <= b;
    layer6_outputs(7336) <= a xor b;
    layer6_outputs(7337) <= not a;
    layer6_outputs(7338) <= not (a and b);
    layer6_outputs(7339) <= not b or a;
    layer6_outputs(7340) <= b;
    layer6_outputs(7341) <= not a or b;
    layer6_outputs(7342) <= not (a or b);
    layer6_outputs(7343) <= not b or a;
    layer6_outputs(7344) <= not (a xor b);
    layer6_outputs(7345) <= not (a and b);
    layer6_outputs(7346) <= a and not b;
    layer6_outputs(7347) <= 1'b0;
    layer6_outputs(7348) <= not b;
    layer6_outputs(7349) <= a xor b;
    layer6_outputs(7350) <= b and not a;
    layer6_outputs(7351) <= not (a and b);
    layer6_outputs(7352) <= not (a and b);
    layer6_outputs(7353) <= not a;
    layer6_outputs(7354) <= b;
    layer6_outputs(7355) <= not a;
    layer6_outputs(7356) <= not b;
    layer6_outputs(7357) <= a and b;
    layer6_outputs(7358) <= not (a and b);
    layer6_outputs(7359) <= not b;
    layer6_outputs(7360) <= not (a xor b);
    layer6_outputs(7361) <= not (a or b);
    layer6_outputs(7362) <= b;
    layer6_outputs(7363) <= a and not b;
    layer6_outputs(7364) <= b and not a;
    layer6_outputs(7365) <= not a or b;
    layer6_outputs(7366) <= b;
    layer6_outputs(7367) <= not a or b;
    layer6_outputs(7368) <= a xor b;
    layer6_outputs(7369) <= not a;
    layer6_outputs(7370) <= 1'b0;
    layer6_outputs(7371) <= a xor b;
    layer6_outputs(7372) <= 1'b1;
    layer6_outputs(7373) <= a or b;
    layer6_outputs(7374) <= b and not a;
    layer6_outputs(7375) <= not a;
    layer6_outputs(7376) <= a and b;
    layer6_outputs(7377) <= b and not a;
    layer6_outputs(7378) <= not b or a;
    layer6_outputs(7379) <= not b or a;
    layer6_outputs(7380) <= a and not b;
    layer6_outputs(7381) <= 1'b0;
    layer6_outputs(7382) <= not a or b;
    layer6_outputs(7383) <= a and b;
    layer6_outputs(7384) <= b;
    layer6_outputs(7385) <= not a;
    layer6_outputs(7386) <= a;
    layer6_outputs(7387) <= b and not a;
    layer6_outputs(7388) <= not a;
    layer6_outputs(7389) <= 1'b0;
    layer6_outputs(7390) <= not a;
    layer6_outputs(7391) <= b and not a;
    layer6_outputs(7392) <= not b or a;
    layer6_outputs(7393) <= not a or b;
    layer6_outputs(7394) <= not (a or b);
    layer6_outputs(7395) <= not a;
    layer6_outputs(7396) <= not (a xor b);
    layer6_outputs(7397) <= not b;
    layer6_outputs(7398) <= b;
    layer6_outputs(7399) <= b;
    layer6_outputs(7400) <= not a;
    layer6_outputs(7401) <= b and not a;
    layer6_outputs(7402) <= 1'b1;
    layer6_outputs(7403) <= b;
    layer6_outputs(7404) <= a xor b;
    layer6_outputs(7405) <= b and not a;
    layer6_outputs(7406) <= a xor b;
    layer6_outputs(7407) <= b and not a;
    layer6_outputs(7408) <= not a or b;
    layer6_outputs(7409) <= a or b;
    layer6_outputs(7410) <= b;
    layer6_outputs(7411) <= a and b;
    layer6_outputs(7412) <= b;
    layer6_outputs(7413) <= a or b;
    layer6_outputs(7414) <= not (a and b);
    layer6_outputs(7415) <= not (a or b);
    layer6_outputs(7416) <= a and not b;
    layer6_outputs(7417) <= a and b;
    layer6_outputs(7418) <= b;
    layer6_outputs(7419) <= b;
    layer6_outputs(7420) <= not (a and b);
    layer6_outputs(7421) <= not a or b;
    layer6_outputs(7422) <= not b or a;
    layer6_outputs(7423) <= not (a or b);
    layer6_outputs(7424) <= a and b;
    layer6_outputs(7425) <= not (a xor b);
    layer6_outputs(7426) <= not (a xor b);
    layer6_outputs(7427) <= not b;
    layer6_outputs(7428) <= not b or a;
    layer6_outputs(7429) <= not a;
    layer6_outputs(7430) <= not b or a;
    layer6_outputs(7431) <= not b;
    layer6_outputs(7432) <= a and b;
    layer6_outputs(7433) <= a xor b;
    layer6_outputs(7434) <= a and b;
    layer6_outputs(7435) <= b and not a;
    layer6_outputs(7436) <= not a;
    layer6_outputs(7437) <= a;
    layer6_outputs(7438) <= not (a and b);
    layer6_outputs(7439) <= 1'b0;
    layer6_outputs(7440) <= b;
    layer6_outputs(7441) <= b and not a;
    layer6_outputs(7442) <= a xor b;
    layer6_outputs(7443) <= b;
    layer6_outputs(7444) <= a;
    layer6_outputs(7445) <= b;
    layer6_outputs(7446) <= b and not a;
    layer6_outputs(7447) <= a and b;
    layer6_outputs(7448) <= not b;
    layer6_outputs(7449) <= not (a and b);
    layer6_outputs(7450) <= not a;
    layer6_outputs(7451) <= a xor b;
    layer6_outputs(7452) <= b;
    layer6_outputs(7453) <= not b or a;
    layer6_outputs(7454) <= not b;
    layer6_outputs(7455) <= a and not b;
    layer6_outputs(7456) <= not a;
    layer6_outputs(7457) <= not (a xor b);
    layer6_outputs(7458) <= not b;
    layer6_outputs(7459) <= not a or b;
    layer6_outputs(7460) <= a xor b;
    layer6_outputs(7461) <= a xor b;
    layer6_outputs(7462) <= a xor b;
    layer6_outputs(7463) <= a and not b;
    layer6_outputs(7464) <= not b;
    layer6_outputs(7465) <= a or b;
    layer6_outputs(7466) <= 1'b0;
    layer6_outputs(7467) <= a xor b;
    layer6_outputs(7468) <= not b;
    layer6_outputs(7469) <= not b;
    layer6_outputs(7470) <= a and b;
    layer6_outputs(7471) <= not b;
    layer6_outputs(7472) <= b;
    layer6_outputs(7473) <= b and not a;
    layer6_outputs(7474) <= not (a and b);
    layer6_outputs(7475) <= a;
    layer6_outputs(7476) <= not (a or b);
    layer6_outputs(7477) <= a and not b;
    layer6_outputs(7478) <= not b;
    layer6_outputs(7479) <= a and not b;
    layer6_outputs(7480) <= a;
    layer6_outputs(7481) <= not (a or b);
    layer6_outputs(7482) <= a;
    layer6_outputs(7483) <= a and b;
    layer6_outputs(7484) <= a;
    layer6_outputs(7485) <= b;
    layer6_outputs(7486) <= not b;
    layer6_outputs(7487) <= b;
    layer6_outputs(7488) <= not (a xor b);
    layer6_outputs(7489) <= not a or b;
    layer6_outputs(7490) <= a and not b;
    layer6_outputs(7491) <= a and not b;
    layer6_outputs(7492) <= not a;
    layer6_outputs(7493) <= b;
    layer6_outputs(7494) <= a;
    layer6_outputs(7495) <= not a;
    layer6_outputs(7496) <= not b or a;
    layer6_outputs(7497) <= b and not a;
    layer6_outputs(7498) <= b and not a;
    layer6_outputs(7499) <= not (a or b);
    layer6_outputs(7500) <= b and not a;
    layer6_outputs(7501) <= not a;
    layer6_outputs(7502) <= b and not a;
    layer6_outputs(7503) <= not a or b;
    layer6_outputs(7504) <= not b or a;
    layer6_outputs(7505) <= not a or b;
    layer6_outputs(7506) <= not (a and b);
    layer6_outputs(7507) <= b;
    layer6_outputs(7508) <= not a;
    layer6_outputs(7509) <= b and not a;
    layer6_outputs(7510) <= 1'b1;
    layer6_outputs(7511) <= a;
    layer6_outputs(7512) <= a;
    layer6_outputs(7513) <= b;
    layer6_outputs(7514) <= a or b;
    layer6_outputs(7515) <= 1'b0;
    layer6_outputs(7516) <= not (a xor b);
    layer6_outputs(7517) <= not a or b;
    layer6_outputs(7518) <= a xor b;
    layer6_outputs(7519) <= 1'b0;
    layer6_outputs(7520) <= b;
    layer6_outputs(7521) <= 1'b1;
    layer6_outputs(7522) <= b and not a;
    layer6_outputs(7523) <= 1'b1;
    layer6_outputs(7524) <= a;
    layer6_outputs(7525) <= not (a and b);
    layer6_outputs(7526) <= a or b;
    layer6_outputs(7527) <= not (a and b);
    layer6_outputs(7528) <= a;
    layer6_outputs(7529) <= b;
    layer6_outputs(7530) <= b and not a;
    layer6_outputs(7531) <= not a;
    layer6_outputs(7532) <= not a or b;
    layer6_outputs(7533) <= not b;
    layer6_outputs(7534) <= not b or a;
    layer6_outputs(7535) <= a and not b;
    layer6_outputs(7536) <= a xor b;
    layer6_outputs(7537) <= a and b;
    layer6_outputs(7538) <= b;
    layer6_outputs(7539) <= 1'b0;
    layer6_outputs(7540) <= a;
    layer6_outputs(7541) <= not (a xor b);
    layer6_outputs(7542) <= not b;
    layer6_outputs(7543) <= b;
    layer6_outputs(7544) <= not a or b;
    layer6_outputs(7545) <= b;
    layer6_outputs(7546) <= a xor b;
    layer6_outputs(7547) <= not (a or b);
    layer6_outputs(7548) <= b and not a;
    layer6_outputs(7549) <= a;
    layer6_outputs(7550) <= not a;
    layer6_outputs(7551) <= a xor b;
    layer6_outputs(7552) <= not (a xor b);
    layer6_outputs(7553) <= not b;
    layer6_outputs(7554) <= not (a or b);
    layer6_outputs(7555) <= not (a and b);
    layer6_outputs(7556) <= not b or a;
    layer6_outputs(7557) <= not (a and b);
    layer6_outputs(7558) <= a;
    layer6_outputs(7559) <= not b or a;
    layer6_outputs(7560) <= not a;
    layer6_outputs(7561) <= not (a and b);
    layer6_outputs(7562) <= not b;
    layer6_outputs(7563) <= b;
    layer6_outputs(7564) <= not (a and b);
    layer6_outputs(7565) <= a;
    layer6_outputs(7566) <= b and not a;
    layer6_outputs(7567) <= not (a and b);
    layer6_outputs(7568) <= b;
    layer6_outputs(7569) <= not (a or b);
    layer6_outputs(7570) <= not a;
    layer6_outputs(7571) <= not a;
    layer6_outputs(7572) <= not a or b;
    layer6_outputs(7573) <= a xor b;
    layer6_outputs(7574) <= 1'b0;
    layer6_outputs(7575) <= b;
    layer6_outputs(7576) <= not b;
    layer6_outputs(7577) <= not b;
    layer6_outputs(7578) <= b;
    layer6_outputs(7579) <= not (a or b);
    layer6_outputs(7580) <= a;
    layer6_outputs(7581) <= a and not b;
    layer6_outputs(7582) <= not (a xor b);
    layer6_outputs(7583) <= not a or b;
    layer6_outputs(7584) <= a xor b;
    layer6_outputs(7585) <= not b;
    layer6_outputs(7586) <= a and b;
    layer6_outputs(7587) <= b;
    layer6_outputs(7588) <= not b;
    layer6_outputs(7589) <= a and not b;
    layer6_outputs(7590) <= a xor b;
    layer6_outputs(7591) <= b;
    layer6_outputs(7592) <= not a;
    layer6_outputs(7593) <= not a or b;
    layer6_outputs(7594) <= not a;
    layer6_outputs(7595) <= a;
    layer6_outputs(7596) <= b;
    layer6_outputs(7597) <= not b;
    layer6_outputs(7598) <= a;
    layer6_outputs(7599) <= not (a and b);
    layer6_outputs(7600) <= not (a and b);
    layer6_outputs(7601) <= a;
    layer6_outputs(7602) <= not a;
    layer6_outputs(7603) <= not (a or b);
    layer6_outputs(7604) <= a or b;
    layer6_outputs(7605) <= a and b;
    layer6_outputs(7606) <= a;
    layer6_outputs(7607) <= a;
    layer6_outputs(7608) <= not a;
    layer6_outputs(7609) <= a and not b;
    layer6_outputs(7610) <= a;
    layer6_outputs(7611) <= a xor b;
    layer6_outputs(7612) <= b;
    layer6_outputs(7613) <= a and b;
    layer6_outputs(7614) <= not a;
    layer6_outputs(7615) <= b;
    layer6_outputs(7616) <= not b;
    layer6_outputs(7617) <= not (a or b);
    layer6_outputs(7618) <= b and not a;
    layer6_outputs(7619) <= not (a xor b);
    layer6_outputs(7620) <= not b;
    layer6_outputs(7621) <= a and not b;
    layer6_outputs(7622) <= b and not a;
    layer6_outputs(7623) <= not (a and b);
    layer6_outputs(7624) <= not b or a;
    layer6_outputs(7625) <= not a or b;
    layer6_outputs(7626) <= not b or a;
    layer6_outputs(7627) <= not (a or b);
    layer6_outputs(7628) <= not b or a;
    layer6_outputs(7629) <= b;
    layer6_outputs(7630) <= not a;
    layer6_outputs(7631) <= b and not a;
    layer6_outputs(7632) <= a or b;
    layer6_outputs(7633) <= a;
    layer6_outputs(7634) <= not (a xor b);
    layer6_outputs(7635) <= a;
    layer6_outputs(7636) <= not a;
    layer6_outputs(7637) <= a;
    layer6_outputs(7638) <= not (a and b);
    layer6_outputs(7639) <= not b;
    layer6_outputs(7640) <= not a;
    layer6_outputs(7641) <= not b;
    layer6_outputs(7642) <= not a or b;
    layer6_outputs(7643) <= a and not b;
    layer6_outputs(7644) <= not a or b;
    layer6_outputs(7645) <= not (a and b);
    layer6_outputs(7646) <= not (a or b);
    layer6_outputs(7647) <= not a or b;
    layer6_outputs(7648) <= a;
    layer6_outputs(7649) <= not b;
    layer6_outputs(7650) <= a or b;
    layer6_outputs(7651) <= not (a or b);
    layer6_outputs(7652) <= a or b;
    layer6_outputs(7653) <= not (a xor b);
    layer6_outputs(7654) <= not a or b;
    layer6_outputs(7655) <= b;
    layer6_outputs(7656) <= b and not a;
    layer6_outputs(7657) <= not b or a;
    layer6_outputs(7658) <= not b or a;
    layer6_outputs(7659) <= a and b;
    layer6_outputs(7660) <= a;
    layer6_outputs(7661) <= not b;
    layer6_outputs(7662) <= b;
    layer6_outputs(7663) <= a and not b;
    layer6_outputs(7664) <= not b or a;
    layer6_outputs(7665) <= b and not a;
    layer6_outputs(7666) <= not a;
    layer6_outputs(7667) <= a and not b;
    layer6_outputs(7668) <= a and not b;
    layer6_outputs(7669) <= not b;
    layer6_outputs(7670) <= not a or b;
    layer6_outputs(7671) <= not a;
    layer6_outputs(7672) <= a or b;
    layer6_outputs(7673) <= a and b;
    layer6_outputs(7674) <= a and not b;
    layer6_outputs(7675) <= a or b;
    layer6_outputs(7676) <= a xor b;
    layer6_outputs(7677) <= not a or b;
    layer6_outputs(7678) <= not a or b;
    layer6_outputs(7679) <= not a or b;
    layer6_outputs(7680) <= not a or b;
    layer6_outputs(7681) <= not (a and b);
    layer6_outputs(7682) <= not a or b;
    layer6_outputs(7683) <= not b;
    layer6_outputs(7684) <= b;
    layer6_outputs(7685) <= b;
    layer6_outputs(7686) <= not (a and b);
    layer6_outputs(7687) <= a and b;
    layer6_outputs(7688) <= b;
    layer6_outputs(7689) <= a and b;
    layer6_outputs(7690) <= b;
    layer6_outputs(7691) <= b and not a;
    layer6_outputs(7692) <= not (a and b);
    layer6_outputs(7693) <= not a;
    layer6_outputs(7694) <= a;
    layer6_outputs(7695) <= a;
    layer6_outputs(7696) <= a and b;
    layer6_outputs(7697) <= not b;
    layer6_outputs(7698) <= a xor b;
    layer6_outputs(7699) <= not b or a;
    layer6_outputs(7700) <= not b;
    layer6_outputs(7701) <= not (a xor b);
    layer6_outputs(7702) <= b;
    layer6_outputs(7703) <= a and b;
    layer6_outputs(7704) <= not (a xor b);
    layer6_outputs(7705) <= b;
    layer6_outputs(7706) <= b and not a;
    layer6_outputs(7707) <= a;
    layer6_outputs(7708) <= b;
    layer6_outputs(7709) <= a and b;
    layer6_outputs(7710) <= not (a xor b);
    layer6_outputs(7711) <= b and not a;
    layer6_outputs(7712) <= a or b;
    layer6_outputs(7713) <= a or b;
    layer6_outputs(7714) <= b;
    layer6_outputs(7715) <= a or b;
    layer6_outputs(7716) <= not b;
    layer6_outputs(7717) <= a and not b;
    layer6_outputs(7718) <= not b;
    layer6_outputs(7719) <= b;
    layer6_outputs(7720) <= a;
    layer6_outputs(7721) <= not (a and b);
    layer6_outputs(7722) <= a or b;
    layer6_outputs(7723) <= a xor b;
    layer6_outputs(7724) <= not a or b;
    layer6_outputs(7725) <= not a;
    layer6_outputs(7726) <= not b or a;
    layer6_outputs(7727) <= a and not b;
    layer6_outputs(7728) <= 1'b0;
    layer6_outputs(7729) <= b;
    layer6_outputs(7730) <= a and b;
    layer6_outputs(7731) <= not b;
    layer6_outputs(7732) <= not (a or b);
    layer6_outputs(7733) <= a xor b;
    layer6_outputs(7734) <= a;
    layer6_outputs(7735) <= a;
    layer6_outputs(7736) <= b;
    layer6_outputs(7737) <= b and not a;
    layer6_outputs(7738) <= b;
    layer6_outputs(7739) <= 1'b1;
    layer6_outputs(7740) <= a and b;
    layer6_outputs(7741) <= not a;
    layer6_outputs(7742) <= a xor b;
    layer6_outputs(7743) <= a or b;
    layer6_outputs(7744) <= b and not a;
    layer6_outputs(7745) <= a xor b;
    layer6_outputs(7746) <= b and not a;
    layer6_outputs(7747) <= not b;
    layer6_outputs(7748) <= a and not b;
    layer6_outputs(7749) <= not (a or b);
    layer6_outputs(7750) <= not a;
    layer6_outputs(7751) <= b;
    layer6_outputs(7752) <= a;
    layer6_outputs(7753) <= not a;
    layer6_outputs(7754) <= a or b;
    layer6_outputs(7755) <= a xor b;
    layer6_outputs(7756) <= b;
    layer6_outputs(7757) <= b;
    layer6_outputs(7758) <= a and b;
    layer6_outputs(7759) <= 1'b1;
    layer6_outputs(7760) <= not a;
    layer6_outputs(7761) <= not (a or b);
    layer6_outputs(7762) <= not b;
    layer6_outputs(7763) <= b and not a;
    layer6_outputs(7764) <= a;
    layer6_outputs(7765) <= a or b;
    layer6_outputs(7766) <= b;
    layer6_outputs(7767) <= a or b;
    layer6_outputs(7768) <= b;
    layer6_outputs(7769) <= a and not b;
    layer6_outputs(7770) <= 1'b1;
    layer6_outputs(7771) <= not (a or b);
    layer6_outputs(7772) <= not b;
    layer6_outputs(7773) <= b;
    layer6_outputs(7774) <= a xor b;
    layer6_outputs(7775) <= not b;
    layer6_outputs(7776) <= not a;
    layer6_outputs(7777) <= not (a and b);
    layer6_outputs(7778) <= not b;
    layer6_outputs(7779) <= a;
    layer6_outputs(7780) <= not b;
    layer6_outputs(7781) <= 1'b0;
    layer6_outputs(7782) <= not b or a;
    layer6_outputs(7783) <= a;
    layer6_outputs(7784) <= a xor b;
    layer6_outputs(7785) <= b and not a;
    layer6_outputs(7786) <= b;
    layer6_outputs(7787) <= a xor b;
    layer6_outputs(7788) <= b;
    layer6_outputs(7789) <= a;
    layer6_outputs(7790) <= not (a and b);
    layer6_outputs(7791) <= not (a and b);
    layer6_outputs(7792) <= a or b;
    layer6_outputs(7793) <= a and b;
    layer6_outputs(7794) <= not b or a;
    layer6_outputs(7795) <= not a or b;
    layer6_outputs(7796) <= a and not b;
    layer6_outputs(7797) <= not (a or b);
    layer6_outputs(7798) <= a or b;
    layer6_outputs(7799) <= a and not b;
    layer6_outputs(7800) <= b;
    layer6_outputs(7801) <= not b;
    layer6_outputs(7802) <= not a;
    layer6_outputs(7803) <= b and not a;
    layer6_outputs(7804) <= not (a xor b);
    layer6_outputs(7805) <= a and b;
    layer6_outputs(7806) <= not a;
    layer6_outputs(7807) <= a or b;
    layer6_outputs(7808) <= a xor b;
    layer6_outputs(7809) <= a;
    layer6_outputs(7810) <= 1'b0;
    layer6_outputs(7811) <= not (a and b);
    layer6_outputs(7812) <= not b;
    layer6_outputs(7813) <= not (a xor b);
    layer6_outputs(7814) <= a xor b;
    layer6_outputs(7815) <= a;
    layer6_outputs(7816) <= a xor b;
    layer6_outputs(7817) <= not (a xor b);
    layer6_outputs(7818) <= not (a or b);
    layer6_outputs(7819) <= b;
    layer6_outputs(7820) <= not a;
    layer6_outputs(7821) <= not (a xor b);
    layer6_outputs(7822) <= not b or a;
    layer6_outputs(7823) <= b;
    layer6_outputs(7824) <= not a or b;
    layer6_outputs(7825) <= b and not a;
    layer6_outputs(7826) <= not b;
    layer6_outputs(7827) <= b and not a;
    layer6_outputs(7828) <= a and not b;
    layer6_outputs(7829) <= a and not b;
    layer6_outputs(7830) <= a or b;
    layer6_outputs(7831) <= 1'b0;
    layer6_outputs(7832) <= b;
    layer6_outputs(7833) <= b;
    layer6_outputs(7834) <= b and not a;
    layer6_outputs(7835) <= a;
    layer6_outputs(7836) <= 1'b1;
    layer6_outputs(7837) <= not b;
    layer6_outputs(7838) <= not b or a;
    layer6_outputs(7839) <= not (a xor b);
    layer6_outputs(7840) <= not a;
    layer6_outputs(7841) <= b;
    layer6_outputs(7842) <= a;
    layer6_outputs(7843) <= not (a or b);
    layer6_outputs(7844) <= not b or a;
    layer6_outputs(7845) <= a;
    layer6_outputs(7846) <= a and not b;
    layer6_outputs(7847) <= a xor b;
    layer6_outputs(7848) <= not a;
    layer6_outputs(7849) <= a or b;
    layer6_outputs(7850) <= not a or b;
    layer6_outputs(7851) <= not (a or b);
    layer6_outputs(7852) <= not (a and b);
    layer6_outputs(7853) <= not b or a;
    layer6_outputs(7854) <= not b;
    layer6_outputs(7855) <= b;
    layer6_outputs(7856) <= not a;
    layer6_outputs(7857) <= 1'b1;
    layer6_outputs(7858) <= a;
    layer6_outputs(7859) <= not (a and b);
    layer6_outputs(7860) <= b;
    layer6_outputs(7861) <= b;
    layer6_outputs(7862) <= not a;
    layer6_outputs(7863) <= not (a xor b);
    layer6_outputs(7864) <= not a;
    layer6_outputs(7865) <= not a or b;
    layer6_outputs(7866) <= b and not a;
    layer6_outputs(7867) <= not (a or b);
    layer6_outputs(7868) <= not a;
    layer6_outputs(7869) <= not b or a;
    layer6_outputs(7870) <= not a;
    layer6_outputs(7871) <= a and not b;
    layer6_outputs(7872) <= not b or a;
    layer6_outputs(7873) <= a or b;
    layer6_outputs(7874) <= not b;
    layer6_outputs(7875) <= b;
    layer6_outputs(7876) <= not (a or b);
    layer6_outputs(7877) <= b;
    layer6_outputs(7878) <= 1'b0;
    layer6_outputs(7879) <= 1'b0;
    layer6_outputs(7880) <= a and b;
    layer6_outputs(7881) <= not a or b;
    layer6_outputs(7882) <= not a or b;
    layer6_outputs(7883) <= a xor b;
    layer6_outputs(7884) <= 1'b0;
    layer6_outputs(7885) <= a or b;
    layer6_outputs(7886) <= b;
    layer6_outputs(7887) <= b;
    layer6_outputs(7888) <= a and b;
    layer6_outputs(7889) <= a and b;
    layer6_outputs(7890) <= not (a xor b);
    layer6_outputs(7891) <= not b or a;
    layer6_outputs(7892) <= a xor b;
    layer6_outputs(7893) <= not b;
    layer6_outputs(7894) <= not b or a;
    layer6_outputs(7895) <= not (a or b);
    layer6_outputs(7896) <= a;
    layer6_outputs(7897) <= not a;
    layer6_outputs(7898) <= b;
    layer6_outputs(7899) <= a;
    layer6_outputs(7900) <= not b;
    layer6_outputs(7901) <= b;
    layer6_outputs(7902) <= b and not a;
    layer6_outputs(7903) <= not a;
    layer6_outputs(7904) <= not b;
    layer6_outputs(7905) <= b and not a;
    layer6_outputs(7906) <= not b or a;
    layer6_outputs(7907) <= not (a and b);
    layer6_outputs(7908) <= a xor b;
    layer6_outputs(7909) <= a;
    layer6_outputs(7910) <= not a;
    layer6_outputs(7911) <= a or b;
    layer6_outputs(7912) <= not a;
    layer6_outputs(7913) <= not b;
    layer6_outputs(7914) <= not (a and b);
    layer6_outputs(7915) <= not b;
    layer6_outputs(7916) <= not b;
    layer6_outputs(7917) <= not (a or b);
    layer6_outputs(7918) <= b;
    layer6_outputs(7919) <= a and not b;
    layer6_outputs(7920) <= a;
    layer6_outputs(7921) <= a or b;
    layer6_outputs(7922) <= b;
    layer6_outputs(7923) <= 1'b1;
    layer6_outputs(7924) <= not b;
    layer6_outputs(7925) <= not (a and b);
    layer6_outputs(7926) <= 1'b0;
    layer6_outputs(7927) <= not a;
    layer6_outputs(7928) <= not a;
    layer6_outputs(7929) <= not (a or b);
    layer6_outputs(7930) <= not a;
    layer6_outputs(7931) <= b and not a;
    layer6_outputs(7932) <= a or b;
    layer6_outputs(7933) <= a;
    layer6_outputs(7934) <= a;
    layer6_outputs(7935) <= not a or b;
    layer6_outputs(7936) <= not b;
    layer6_outputs(7937) <= not (a and b);
    layer6_outputs(7938) <= a or b;
    layer6_outputs(7939) <= not b;
    layer6_outputs(7940) <= a and b;
    layer6_outputs(7941) <= not (a and b);
    layer6_outputs(7942) <= b;
    layer6_outputs(7943) <= not a or b;
    layer6_outputs(7944) <= a xor b;
    layer6_outputs(7945) <= not b;
    layer6_outputs(7946) <= 1'b0;
    layer6_outputs(7947) <= b;
    layer6_outputs(7948) <= a or b;
    layer6_outputs(7949) <= a or b;
    layer6_outputs(7950) <= a;
    layer6_outputs(7951) <= a and not b;
    layer6_outputs(7952) <= not (a xor b);
    layer6_outputs(7953) <= a and b;
    layer6_outputs(7954) <= a and b;
    layer6_outputs(7955) <= a and not b;
    layer6_outputs(7956) <= a and not b;
    layer6_outputs(7957) <= not b or a;
    layer6_outputs(7958) <= not a or b;
    layer6_outputs(7959) <= a xor b;
    layer6_outputs(7960) <= not b or a;
    layer6_outputs(7961) <= a and b;
    layer6_outputs(7962) <= a or b;
    layer6_outputs(7963) <= not (a or b);
    layer6_outputs(7964) <= a xor b;
    layer6_outputs(7965) <= not (a and b);
    layer6_outputs(7966) <= not (a or b);
    layer6_outputs(7967) <= a;
    layer6_outputs(7968) <= not b or a;
    layer6_outputs(7969) <= a;
    layer6_outputs(7970) <= not a;
    layer6_outputs(7971) <= b and not a;
    layer6_outputs(7972) <= a or b;
    layer6_outputs(7973) <= a;
    layer6_outputs(7974) <= 1'b0;
    layer6_outputs(7975) <= b and not a;
    layer6_outputs(7976) <= a and b;
    layer6_outputs(7977) <= not b or a;
    layer6_outputs(7978) <= not b;
    layer6_outputs(7979) <= a;
    layer6_outputs(7980) <= b;
    layer6_outputs(7981) <= a;
    layer6_outputs(7982) <= 1'b0;
    layer6_outputs(7983) <= not (a xor b);
    layer6_outputs(7984) <= not b or a;
    layer6_outputs(7985) <= not a;
    layer6_outputs(7986) <= not a or b;
    layer6_outputs(7987) <= not (a and b);
    layer6_outputs(7988) <= not b;
    layer6_outputs(7989) <= b;
    layer6_outputs(7990) <= b;
    layer6_outputs(7991) <= a or b;
    layer6_outputs(7992) <= not a;
    layer6_outputs(7993) <= not (a xor b);
    layer6_outputs(7994) <= a xor b;
    layer6_outputs(7995) <= a;
    layer6_outputs(7996) <= a;
    layer6_outputs(7997) <= b;
    layer6_outputs(7998) <= not (a or b);
    layer6_outputs(7999) <= a and b;
    layer6_outputs(8000) <= not (a or b);
    layer6_outputs(8001) <= a and not b;
    layer6_outputs(8002) <= not b;
    layer6_outputs(8003) <= not (a xor b);
    layer6_outputs(8004) <= not (a and b);
    layer6_outputs(8005) <= a and not b;
    layer6_outputs(8006) <= a;
    layer6_outputs(8007) <= a or b;
    layer6_outputs(8008) <= b;
    layer6_outputs(8009) <= not b;
    layer6_outputs(8010) <= not a or b;
    layer6_outputs(8011) <= a;
    layer6_outputs(8012) <= b;
    layer6_outputs(8013) <= not a;
    layer6_outputs(8014) <= a or b;
    layer6_outputs(8015) <= a and b;
    layer6_outputs(8016) <= a xor b;
    layer6_outputs(8017) <= not b;
    layer6_outputs(8018) <= a and b;
    layer6_outputs(8019) <= a and b;
    layer6_outputs(8020) <= a or b;
    layer6_outputs(8021) <= a and b;
    layer6_outputs(8022) <= not a;
    layer6_outputs(8023) <= b and not a;
    layer6_outputs(8024) <= not (a xor b);
    layer6_outputs(8025) <= 1'b0;
    layer6_outputs(8026) <= a xor b;
    layer6_outputs(8027) <= not a;
    layer6_outputs(8028) <= not b or a;
    layer6_outputs(8029) <= not a;
    layer6_outputs(8030) <= a and not b;
    layer6_outputs(8031) <= not a or b;
    layer6_outputs(8032) <= not b or a;
    layer6_outputs(8033) <= a and b;
    layer6_outputs(8034) <= a or b;
    layer6_outputs(8035) <= not b;
    layer6_outputs(8036) <= not (a xor b);
    layer6_outputs(8037) <= not b;
    layer6_outputs(8038) <= b and not a;
    layer6_outputs(8039) <= b;
    layer6_outputs(8040) <= b;
    layer6_outputs(8041) <= not (a and b);
    layer6_outputs(8042) <= b and not a;
    layer6_outputs(8043) <= b;
    layer6_outputs(8044) <= not a;
    layer6_outputs(8045) <= not a;
    layer6_outputs(8046) <= b;
    layer6_outputs(8047) <= not b;
    layer6_outputs(8048) <= b;
    layer6_outputs(8049) <= not a or b;
    layer6_outputs(8050) <= not a or b;
    layer6_outputs(8051) <= not (a and b);
    layer6_outputs(8052) <= a;
    layer6_outputs(8053) <= not (a and b);
    layer6_outputs(8054) <= not a or b;
    layer6_outputs(8055) <= not (a and b);
    layer6_outputs(8056) <= not (a or b);
    layer6_outputs(8057) <= a xor b;
    layer6_outputs(8058) <= a or b;
    layer6_outputs(8059) <= not a or b;
    layer6_outputs(8060) <= not b;
    layer6_outputs(8061) <= not (a or b);
    layer6_outputs(8062) <= a and not b;
    layer6_outputs(8063) <= not a;
    layer6_outputs(8064) <= not b;
    layer6_outputs(8065) <= 1'b1;
    layer6_outputs(8066) <= a;
    layer6_outputs(8067) <= a;
    layer6_outputs(8068) <= b;
    layer6_outputs(8069) <= not b or a;
    layer6_outputs(8070) <= not a;
    layer6_outputs(8071) <= a or b;
    layer6_outputs(8072) <= not b or a;
    layer6_outputs(8073) <= not a;
    layer6_outputs(8074) <= not (a and b);
    layer6_outputs(8075) <= not a or b;
    layer6_outputs(8076) <= a;
    layer6_outputs(8077) <= a and not b;
    layer6_outputs(8078) <= a and b;
    layer6_outputs(8079) <= a xor b;
    layer6_outputs(8080) <= not (a or b);
    layer6_outputs(8081) <= not b;
    layer6_outputs(8082) <= a and b;
    layer6_outputs(8083) <= b;
    layer6_outputs(8084) <= a and not b;
    layer6_outputs(8085) <= b and not a;
    layer6_outputs(8086) <= not b;
    layer6_outputs(8087) <= not b;
    layer6_outputs(8088) <= b;
    layer6_outputs(8089) <= not a;
    layer6_outputs(8090) <= a;
    layer6_outputs(8091) <= not (a and b);
    layer6_outputs(8092) <= a and not b;
    layer6_outputs(8093) <= a and b;
    layer6_outputs(8094) <= not (a and b);
    layer6_outputs(8095) <= not b;
    layer6_outputs(8096) <= not b;
    layer6_outputs(8097) <= not b or a;
    layer6_outputs(8098) <= a;
    layer6_outputs(8099) <= not a or b;
    layer6_outputs(8100) <= b;
    layer6_outputs(8101) <= b;
    layer6_outputs(8102) <= b;
    layer6_outputs(8103) <= b;
    layer6_outputs(8104) <= not a or b;
    layer6_outputs(8105) <= a and b;
    layer6_outputs(8106) <= b;
    layer6_outputs(8107) <= b;
    layer6_outputs(8108) <= a and not b;
    layer6_outputs(8109) <= not a or b;
    layer6_outputs(8110) <= b;
    layer6_outputs(8111) <= not a or b;
    layer6_outputs(8112) <= b and not a;
    layer6_outputs(8113) <= a;
    layer6_outputs(8114) <= 1'b1;
    layer6_outputs(8115) <= a and b;
    layer6_outputs(8116) <= 1'b0;
    layer6_outputs(8117) <= not (a or b);
    layer6_outputs(8118) <= not (a xor b);
    layer6_outputs(8119) <= a;
    layer6_outputs(8120) <= not b or a;
    layer6_outputs(8121) <= not (a or b);
    layer6_outputs(8122) <= b;
    layer6_outputs(8123) <= not b or a;
    layer6_outputs(8124) <= a xor b;
    layer6_outputs(8125) <= a or b;
    layer6_outputs(8126) <= not b or a;
    layer6_outputs(8127) <= not a;
    layer6_outputs(8128) <= 1'b1;
    layer6_outputs(8129) <= not a;
    layer6_outputs(8130) <= not a;
    layer6_outputs(8131) <= a;
    layer6_outputs(8132) <= a xor b;
    layer6_outputs(8133) <= not b or a;
    layer6_outputs(8134) <= a and not b;
    layer6_outputs(8135) <= a xor b;
    layer6_outputs(8136) <= a xor b;
    layer6_outputs(8137) <= not b;
    layer6_outputs(8138) <= b;
    layer6_outputs(8139) <= a xor b;
    layer6_outputs(8140) <= not a or b;
    layer6_outputs(8141) <= a and not b;
    layer6_outputs(8142) <= not a;
    layer6_outputs(8143) <= a and not b;
    layer6_outputs(8144) <= 1'b0;
    layer6_outputs(8145) <= not b;
    layer6_outputs(8146) <= not a or b;
    layer6_outputs(8147) <= not b;
    layer6_outputs(8148) <= not b;
    layer6_outputs(8149) <= b and not a;
    layer6_outputs(8150) <= not b;
    layer6_outputs(8151) <= not (a or b);
    layer6_outputs(8152) <= a and not b;
    layer6_outputs(8153) <= not b or a;
    layer6_outputs(8154) <= not b;
    layer6_outputs(8155) <= a;
    layer6_outputs(8156) <= a;
    layer6_outputs(8157) <= not (a or b);
    layer6_outputs(8158) <= 1'b0;
    layer6_outputs(8159) <= not (a and b);
    layer6_outputs(8160) <= b and not a;
    layer6_outputs(8161) <= not b;
    layer6_outputs(8162) <= b and not a;
    layer6_outputs(8163) <= not b or a;
    layer6_outputs(8164) <= not a or b;
    layer6_outputs(8165) <= not b or a;
    layer6_outputs(8166) <= not b or a;
    layer6_outputs(8167) <= not b or a;
    layer6_outputs(8168) <= a or b;
    layer6_outputs(8169) <= not (a or b);
    layer6_outputs(8170) <= not (a and b);
    layer6_outputs(8171) <= a;
    layer6_outputs(8172) <= not (a or b);
    layer6_outputs(8173) <= b;
    layer6_outputs(8174) <= a xor b;
    layer6_outputs(8175) <= a or b;
    layer6_outputs(8176) <= a or b;
    layer6_outputs(8177) <= not (a xor b);
    layer6_outputs(8178) <= a xor b;
    layer6_outputs(8179) <= not a;
    layer6_outputs(8180) <= 1'b0;
    layer6_outputs(8181) <= not (a xor b);
    layer6_outputs(8182) <= not b or a;
    layer6_outputs(8183) <= not b;
    layer6_outputs(8184) <= not a or b;
    layer6_outputs(8185) <= a xor b;
    layer6_outputs(8186) <= not b;
    layer6_outputs(8187) <= a;
    layer6_outputs(8188) <= not b or a;
    layer6_outputs(8189) <= b;
    layer6_outputs(8190) <= not b;
    layer6_outputs(8191) <= b and not a;
    layer6_outputs(8192) <= not b;
    layer6_outputs(8193) <= not a;
    layer6_outputs(8194) <= a or b;
    layer6_outputs(8195) <= not (a and b);
    layer6_outputs(8196) <= b and not a;
    layer6_outputs(8197) <= not b;
    layer6_outputs(8198) <= not b;
    layer6_outputs(8199) <= not b;
    layer6_outputs(8200) <= 1'b1;
    layer6_outputs(8201) <= not (a xor b);
    layer6_outputs(8202) <= b and not a;
    layer6_outputs(8203) <= a or b;
    layer6_outputs(8204) <= a or b;
    layer6_outputs(8205) <= not a or b;
    layer6_outputs(8206) <= not b;
    layer6_outputs(8207) <= b;
    layer6_outputs(8208) <= b;
    layer6_outputs(8209) <= not b or a;
    layer6_outputs(8210) <= a and b;
    layer6_outputs(8211) <= not b;
    layer6_outputs(8212) <= not (a xor b);
    layer6_outputs(8213) <= a;
    layer6_outputs(8214) <= b;
    layer6_outputs(8215) <= not (a xor b);
    layer6_outputs(8216) <= b;
    layer6_outputs(8217) <= a;
    layer6_outputs(8218) <= 1'b0;
    layer6_outputs(8219) <= not b;
    layer6_outputs(8220) <= not a or b;
    layer6_outputs(8221) <= a and not b;
    layer6_outputs(8222) <= not (a and b);
    layer6_outputs(8223) <= b and not a;
    layer6_outputs(8224) <= a;
    layer6_outputs(8225) <= not a or b;
    layer6_outputs(8226) <= a xor b;
    layer6_outputs(8227) <= not (a and b);
    layer6_outputs(8228) <= not (a and b);
    layer6_outputs(8229) <= not b;
    layer6_outputs(8230) <= not a or b;
    layer6_outputs(8231) <= not (a and b);
    layer6_outputs(8232) <= not (a and b);
    layer6_outputs(8233) <= not a;
    layer6_outputs(8234) <= not (a and b);
    layer6_outputs(8235) <= not (a and b);
    layer6_outputs(8236) <= a or b;
    layer6_outputs(8237) <= b and not a;
    layer6_outputs(8238) <= not (a and b);
    layer6_outputs(8239) <= not (a or b);
    layer6_outputs(8240) <= not b;
    layer6_outputs(8241) <= not b;
    layer6_outputs(8242) <= b and not a;
    layer6_outputs(8243) <= not b;
    layer6_outputs(8244) <= a xor b;
    layer6_outputs(8245) <= a and b;
    layer6_outputs(8246) <= a xor b;
    layer6_outputs(8247) <= not a;
    layer6_outputs(8248) <= a xor b;
    layer6_outputs(8249) <= a and b;
    layer6_outputs(8250) <= not (a and b);
    layer6_outputs(8251) <= not a;
    layer6_outputs(8252) <= b;
    layer6_outputs(8253) <= a;
    layer6_outputs(8254) <= a or b;
    layer6_outputs(8255) <= not a or b;
    layer6_outputs(8256) <= b and not a;
    layer6_outputs(8257) <= a;
    layer6_outputs(8258) <= not b;
    layer6_outputs(8259) <= not b or a;
    layer6_outputs(8260) <= 1'b0;
    layer6_outputs(8261) <= not (a and b);
    layer6_outputs(8262) <= 1'b1;
    layer6_outputs(8263) <= a;
    layer6_outputs(8264) <= 1'b0;
    layer6_outputs(8265) <= not a or b;
    layer6_outputs(8266) <= 1'b1;
    layer6_outputs(8267) <= not (a xor b);
    layer6_outputs(8268) <= b;
    layer6_outputs(8269) <= not b or a;
    layer6_outputs(8270) <= not b;
    layer6_outputs(8271) <= a and not b;
    layer6_outputs(8272) <= a or b;
    layer6_outputs(8273) <= not a;
    layer6_outputs(8274) <= a and not b;
    layer6_outputs(8275) <= a and b;
    layer6_outputs(8276) <= a or b;
    layer6_outputs(8277) <= a;
    layer6_outputs(8278) <= a xor b;
    layer6_outputs(8279) <= a;
    layer6_outputs(8280) <= not (a xor b);
    layer6_outputs(8281) <= not b;
    layer6_outputs(8282) <= b and not a;
    layer6_outputs(8283) <= not b;
    layer6_outputs(8284) <= b;
    layer6_outputs(8285) <= b;
    layer6_outputs(8286) <= 1'b0;
    layer6_outputs(8287) <= b;
    layer6_outputs(8288) <= a;
    layer6_outputs(8289) <= a;
    layer6_outputs(8290) <= b;
    layer6_outputs(8291) <= not a or b;
    layer6_outputs(8292) <= not b or a;
    layer6_outputs(8293) <= b;
    layer6_outputs(8294) <= not a or b;
    layer6_outputs(8295) <= a;
    layer6_outputs(8296) <= a and not b;
    layer6_outputs(8297) <= a xor b;
    layer6_outputs(8298) <= b;
    layer6_outputs(8299) <= not (a or b);
    layer6_outputs(8300) <= a;
    layer6_outputs(8301) <= a or b;
    layer6_outputs(8302) <= a and not b;
    layer6_outputs(8303) <= b and not a;
    layer6_outputs(8304) <= 1'b0;
    layer6_outputs(8305) <= a;
    layer6_outputs(8306) <= not b or a;
    layer6_outputs(8307) <= not a;
    layer6_outputs(8308) <= a and not b;
    layer6_outputs(8309) <= a or b;
    layer6_outputs(8310) <= not (a xor b);
    layer6_outputs(8311) <= b and not a;
    layer6_outputs(8312) <= a or b;
    layer6_outputs(8313) <= a;
    layer6_outputs(8314) <= not b or a;
    layer6_outputs(8315) <= a;
    layer6_outputs(8316) <= a;
    layer6_outputs(8317) <= a xor b;
    layer6_outputs(8318) <= b and not a;
    layer6_outputs(8319) <= a or b;
    layer6_outputs(8320) <= b;
    layer6_outputs(8321) <= not (a xor b);
    layer6_outputs(8322) <= 1'b1;
    layer6_outputs(8323) <= not a or b;
    layer6_outputs(8324) <= 1'b1;
    layer6_outputs(8325) <= a xor b;
    layer6_outputs(8326) <= 1'b0;
    layer6_outputs(8327) <= b;
    layer6_outputs(8328) <= not b;
    layer6_outputs(8329) <= a;
    layer6_outputs(8330) <= not a;
    layer6_outputs(8331) <= b;
    layer6_outputs(8332) <= not b;
    layer6_outputs(8333) <= a;
    layer6_outputs(8334) <= b and not a;
    layer6_outputs(8335) <= b;
    layer6_outputs(8336) <= not b;
    layer6_outputs(8337) <= a;
    layer6_outputs(8338) <= not (a or b);
    layer6_outputs(8339) <= not b or a;
    layer6_outputs(8340) <= a or b;
    layer6_outputs(8341) <= b and not a;
    layer6_outputs(8342) <= a or b;
    layer6_outputs(8343) <= not (a xor b);
    layer6_outputs(8344) <= not a;
    layer6_outputs(8345) <= a and b;
    layer6_outputs(8346) <= not b or a;
    layer6_outputs(8347) <= b;
    layer6_outputs(8348) <= a;
    layer6_outputs(8349) <= b and not a;
    layer6_outputs(8350) <= a xor b;
    layer6_outputs(8351) <= not a;
    layer6_outputs(8352) <= a;
    layer6_outputs(8353) <= b;
    layer6_outputs(8354) <= a;
    layer6_outputs(8355) <= a or b;
    layer6_outputs(8356) <= a xor b;
    layer6_outputs(8357) <= not (a and b);
    layer6_outputs(8358) <= a and not b;
    layer6_outputs(8359) <= not a;
    layer6_outputs(8360) <= a;
    layer6_outputs(8361) <= not a;
    layer6_outputs(8362) <= 1'b0;
    layer6_outputs(8363) <= not (a and b);
    layer6_outputs(8364) <= not b;
    layer6_outputs(8365) <= b and not a;
    layer6_outputs(8366) <= a and not b;
    layer6_outputs(8367) <= a and not b;
    layer6_outputs(8368) <= not b or a;
    layer6_outputs(8369) <= not b or a;
    layer6_outputs(8370) <= a or b;
    layer6_outputs(8371) <= b and not a;
    layer6_outputs(8372) <= b;
    layer6_outputs(8373) <= not a or b;
    layer6_outputs(8374) <= b;
    layer6_outputs(8375) <= a and not b;
    layer6_outputs(8376) <= b;
    layer6_outputs(8377) <= not a;
    layer6_outputs(8378) <= not b or a;
    layer6_outputs(8379) <= a and not b;
    layer6_outputs(8380) <= not a;
    layer6_outputs(8381) <= not b or a;
    layer6_outputs(8382) <= a xor b;
    layer6_outputs(8383) <= not a or b;
    layer6_outputs(8384) <= a and b;
    layer6_outputs(8385) <= not (a or b);
    layer6_outputs(8386) <= not b or a;
    layer6_outputs(8387) <= a and not b;
    layer6_outputs(8388) <= not b;
    layer6_outputs(8389) <= not b or a;
    layer6_outputs(8390) <= not (a and b);
    layer6_outputs(8391) <= not b or a;
    layer6_outputs(8392) <= a and not b;
    layer6_outputs(8393) <= not b or a;
    layer6_outputs(8394) <= b;
    layer6_outputs(8395) <= not a;
    layer6_outputs(8396) <= not a;
    layer6_outputs(8397) <= not (a and b);
    layer6_outputs(8398) <= a and not b;
    layer6_outputs(8399) <= not b;
    layer6_outputs(8400) <= not b;
    layer6_outputs(8401) <= a xor b;
    layer6_outputs(8402) <= not a;
    layer6_outputs(8403) <= a and b;
    layer6_outputs(8404) <= not a;
    layer6_outputs(8405) <= a and b;
    layer6_outputs(8406) <= not a or b;
    layer6_outputs(8407) <= not (a xor b);
    layer6_outputs(8408) <= a and not b;
    layer6_outputs(8409) <= not (a and b);
    layer6_outputs(8410) <= a and not b;
    layer6_outputs(8411) <= a xor b;
    layer6_outputs(8412) <= b and not a;
    layer6_outputs(8413) <= not b or a;
    layer6_outputs(8414) <= not b or a;
    layer6_outputs(8415) <= not a;
    layer6_outputs(8416) <= not (a and b);
    layer6_outputs(8417) <= not b;
    layer6_outputs(8418) <= a xor b;
    layer6_outputs(8419) <= not b;
    layer6_outputs(8420) <= a;
    layer6_outputs(8421) <= not a;
    layer6_outputs(8422) <= not a;
    layer6_outputs(8423) <= b;
    layer6_outputs(8424) <= a and b;
    layer6_outputs(8425) <= 1'b1;
    layer6_outputs(8426) <= not a or b;
    layer6_outputs(8427) <= not b;
    layer6_outputs(8428) <= a;
    layer6_outputs(8429) <= a and b;
    layer6_outputs(8430) <= 1'b0;
    layer6_outputs(8431) <= not (a and b);
    layer6_outputs(8432) <= a;
    layer6_outputs(8433) <= a and b;
    layer6_outputs(8434) <= a and b;
    layer6_outputs(8435) <= a and not b;
    layer6_outputs(8436) <= b;
    layer6_outputs(8437) <= not (a xor b);
    layer6_outputs(8438) <= not (a xor b);
    layer6_outputs(8439) <= a;
    layer6_outputs(8440) <= a xor b;
    layer6_outputs(8441) <= not a;
    layer6_outputs(8442) <= a or b;
    layer6_outputs(8443) <= 1'b0;
    layer6_outputs(8444) <= not a;
    layer6_outputs(8445) <= a and b;
    layer6_outputs(8446) <= a;
    layer6_outputs(8447) <= 1'b0;
    layer6_outputs(8448) <= not (a or b);
    layer6_outputs(8449) <= not b or a;
    layer6_outputs(8450) <= b;
    layer6_outputs(8451) <= not a or b;
    layer6_outputs(8452) <= not a;
    layer6_outputs(8453) <= not b;
    layer6_outputs(8454) <= not b;
    layer6_outputs(8455) <= 1'b0;
    layer6_outputs(8456) <= not b;
    layer6_outputs(8457) <= not b or a;
    layer6_outputs(8458) <= b and not a;
    layer6_outputs(8459) <= a or b;
    layer6_outputs(8460) <= not a;
    layer6_outputs(8461) <= a or b;
    layer6_outputs(8462) <= a xor b;
    layer6_outputs(8463) <= not b or a;
    layer6_outputs(8464) <= a;
    layer6_outputs(8465) <= not b;
    layer6_outputs(8466) <= 1'b1;
    layer6_outputs(8467) <= b;
    layer6_outputs(8468) <= not (a or b);
    layer6_outputs(8469) <= b;
    layer6_outputs(8470) <= a and b;
    layer6_outputs(8471) <= a;
    layer6_outputs(8472) <= a;
    layer6_outputs(8473) <= a xor b;
    layer6_outputs(8474) <= a;
    layer6_outputs(8475) <= b;
    layer6_outputs(8476) <= a;
    layer6_outputs(8477) <= not (a or b);
    layer6_outputs(8478) <= a;
    layer6_outputs(8479) <= not (a or b);
    layer6_outputs(8480) <= a;
    layer6_outputs(8481) <= not a;
    layer6_outputs(8482) <= not b or a;
    layer6_outputs(8483) <= a xor b;
    layer6_outputs(8484) <= not b or a;
    layer6_outputs(8485) <= a and not b;
    layer6_outputs(8486) <= not b;
    layer6_outputs(8487) <= not (a or b);
    layer6_outputs(8488) <= not a or b;
    layer6_outputs(8489) <= b and not a;
    layer6_outputs(8490) <= 1'b0;
    layer6_outputs(8491) <= a and b;
    layer6_outputs(8492) <= a;
    layer6_outputs(8493) <= a or b;
    layer6_outputs(8494) <= not a or b;
    layer6_outputs(8495) <= not (a xor b);
    layer6_outputs(8496) <= b;
    layer6_outputs(8497) <= a and b;
    layer6_outputs(8498) <= not b or a;
    layer6_outputs(8499) <= a and b;
    layer6_outputs(8500) <= b;
    layer6_outputs(8501) <= b;
    layer6_outputs(8502) <= a xor b;
    layer6_outputs(8503) <= a;
    layer6_outputs(8504) <= b;
    layer6_outputs(8505) <= not a;
    layer6_outputs(8506) <= a;
    layer6_outputs(8507) <= not a or b;
    layer6_outputs(8508) <= a and not b;
    layer6_outputs(8509) <= not (a or b);
    layer6_outputs(8510) <= not a;
    layer6_outputs(8511) <= not (a and b);
    layer6_outputs(8512) <= not b;
    layer6_outputs(8513) <= not b;
    layer6_outputs(8514) <= not (a or b);
    layer6_outputs(8515) <= 1'b0;
    layer6_outputs(8516) <= 1'b1;
    layer6_outputs(8517) <= b and not a;
    layer6_outputs(8518) <= not a;
    layer6_outputs(8519) <= not (a and b);
    layer6_outputs(8520) <= a or b;
    layer6_outputs(8521) <= not (a xor b);
    layer6_outputs(8522) <= a xor b;
    layer6_outputs(8523) <= a or b;
    layer6_outputs(8524) <= a;
    layer6_outputs(8525) <= not b;
    layer6_outputs(8526) <= not a;
    layer6_outputs(8527) <= not b;
    layer6_outputs(8528) <= b;
    layer6_outputs(8529) <= not (a or b);
    layer6_outputs(8530) <= a or b;
    layer6_outputs(8531) <= b;
    layer6_outputs(8532) <= 1'b1;
    layer6_outputs(8533) <= a;
    layer6_outputs(8534) <= b and not a;
    layer6_outputs(8535) <= not b;
    layer6_outputs(8536) <= a or b;
    layer6_outputs(8537) <= a xor b;
    layer6_outputs(8538) <= a or b;
    layer6_outputs(8539) <= a;
    layer6_outputs(8540) <= not a;
    layer6_outputs(8541) <= a xor b;
    layer6_outputs(8542) <= not (a and b);
    layer6_outputs(8543) <= not (a or b);
    layer6_outputs(8544) <= a xor b;
    layer6_outputs(8545) <= not b;
    layer6_outputs(8546) <= not a;
    layer6_outputs(8547) <= not a or b;
    layer6_outputs(8548) <= not a;
    layer6_outputs(8549) <= not (a and b);
    layer6_outputs(8550) <= a;
    layer6_outputs(8551) <= not (a and b);
    layer6_outputs(8552) <= not a;
    layer6_outputs(8553) <= a or b;
    layer6_outputs(8554) <= not a;
    layer6_outputs(8555) <= a and not b;
    layer6_outputs(8556) <= a;
    layer6_outputs(8557) <= b;
    layer6_outputs(8558) <= not a;
    layer6_outputs(8559) <= not b;
    layer6_outputs(8560) <= b;
    layer6_outputs(8561) <= not b;
    layer6_outputs(8562) <= not b;
    layer6_outputs(8563) <= b;
    layer6_outputs(8564) <= not (a and b);
    layer6_outputs(8565) <= a xor b;
    layer6_outputs(8566) <= a;
    layer6_outputs(8567) <= not a or b;
    layer6_outputs(8568) <= b and not a;
    layer6_outputs(8569) <= a and b;
    layer6_outputs(8570) <= b;
    layer6_outputs(8571) <= b;
    layer6_outputs(8572) <= a;
    layer6_outputs(8573) <= not (a or b);
    layer6_outputs(8574) <= b;
    layer6_outputs(8575) <= not b;
    layer6_outputs(8576) <= a or b;
    layer6_outputs(8577) <= not b or a;
    layer6_outputs(8578) <= not a;
    layer6_outputs(8579) <= a and b;
    layer6_outputs(8580) <= a;
    layer6_outputs(8581) <= a;
    layer6_outputs(8582) <= not (a and b);
    layer6_outputs(8583) <= not b;
    layer6_outputs(8584) <= a and not b;
    layer6_outputs(8585) <= a;
    layer6_outputs(8586) <= b;
    layer6_outputs(8587) <= a and not b;
    layer6_outputs(8588) <= not b or a;
    layer6_outputs(8589) <= a;
    layer6_outputs(8590) <= not (a xor b);
    layer6_outputs(8591) <= a and not b;
    layer6_outputs(8592) <= not (a or b);
    layer6_outputs(8593) <= not (a and b);
    layer6_outputs(8594) <= not (a xor b);
    layer6_outputs(8595) <= not a;
    layer6_outputs(8596) <= a and not b;
    layer6_outputs(8597) <= a;
    layer6_outputs(8598) <= not a;
    layer6_outputs(8599) <= not (a and b);
    layer6_outputs(8600) <= a;
    layer6_outputs(8601) <= a and not b;
    layer6_outputs(8602) <= not b;
    layer6_outputs(8603) <= b and not a;
    layer6_outputs(8604) <= not a;
    layer6_outputs(8605) <= a;
    layer6_outputs(8606) <= b and not a;
    layer6_outputs(8607) <= b;
    layer6_outputs(8608) <= b and not a;
    layer6_outputs(8609) <= a or b;
    layer6_outputs(8610) <= a xor b;
    layer6_outputs(8611) <= a xor b;
    layer6_outputs(8612) <= b and not a;
    layer6_outputs(8613) <= not (a or b);
    layer6_outputs(8614) <= 1'b1;
    layer6_outputs(8615) <= not a;
    layer6_outputs(8616) <= b;
    layer6_outputs(8617) <= a or b;
    layer6_outputs(8618) <= b;
    layer6_outputs(8619) <= a and b;
    layer6_outputs(8620) <= a and not b;
    layer6_outputs(8621) <= b;
    layer6_outputs(8622) <= not (a xor b);
    layer6_outputs(8623) <= not a;
    layer6_outputs(8624) <= b;
    layer6_outputs(8625) <= b;
    layer6_outputs(8626) <= a;
    layer6_outputs(8627) <= a;
    layer6_outputs(8628) <= a;
    layer6_outputs(8629) <= not (a xor b);
    layer6_outputs(8630) <= a xor b;
    layer6_outputs(8631) <= b;
    layer6_outputs(8632) <= a and not b;
    layer6_outputs(8633) <= not a or b;
    layer6_outputs(8634) <= not a;
    layer6_outputs(8635) <= a xor b;
    layer6_outputs(8636) <= a;
    layer6_outputs(8637) <= a or b;
    layer6_outputs(8638) <= not a;
    layer6_outputs(8639) <= 1'b1;
    layer6_outputs(8640) <= a;
    layer6_outputs(8641) <= not b;
    layer6_outputs(8642) <= not a or b;
    layer6_outputs(8643) <= not b or a;
    layer6_outputs(8644) <= not b;
    layer6_outputs(8645) <= b;
    layer6_outputs(8646) <= not a;
    layer6_outputs(8647) <= b and not a;
    layer6_outputs(8648) <= not (a or b);
    layer6_outputs(8649) <= a and b;
    layer6_outputs(8650) <= a xor b;
    layer6_outputs(8651) <= b;
    layer6_outputs(8652) <= not b or a;
    layer6_outputs(8653) <= a and not b;
    layer6_outputs(8654) <= a and b;
    layer6_outputs(8655) <= not (a and b);
    layer6_outputs(8656) <= not (a or b);
    layer6_outputs(8657) <= a;
    layer6_outputs(8658) <= a;
    layer6_outputs(8659) <= b;
    layer6_outputs(8660) <= not a;
    layer6_outputs(8661) <= a or b;
    layer6_outputs(8662) <= a and not b;
    layer6_outputs(8663) <= not (a and b);
    layer6_outputs(8664) <= not a;
    layer6_outputs(8665) <= not b;
    layer6_outputs(8666) <= not a;
    layer6_outputs(8667) <= not b;
    layer6_outputs(8668) <= b and not a;
    layer6_outputs(8669) <= a and not b;
    layer6_outputs(8670) <= b;
    layer6_outputs(8671) <= a;
    layer6_outputs(8672) <= not b;
    layer6_outputs(8673) <= not b;
    layer6_outputs(8674) <= not a or b;
    layer6_outputs(8675) <= not a or b;
    layer6_outputs(8676) <= a and b;
    layer6_outputs(8677) <= not (a or b);
    layer6_outputs(8678) <= b;
    layer6_outputs(8679) <= not a;
    layer6_outputs(8680) <= a;
    layer6_outputs(8681) <= a;
    layer6_outputs(8682) <= a;
    layer6_outputs(8683) <= b;
    layer6_outputs(8684) <= a;
    layer6_outputs(8685) <= not b;
    layer6_outputs(8686) <= not a;
    layer6_outputs(8687) <= not a;
    layer6_outputs(8688) <= a;
    layer6_outputs(8689) <= b and not a;
    layer6_outputs(8690) <= not (a xor b);
    layer6_outputs(8691) <= not (a and b);
    layer6_outputs(8692) <= not b;
    layer6_outputs(8693) <= a and not b;
    layer6_outputs(8694) <= a;
    layer6_outputs(8695) <= 1'b0;
    layer6_outputs(8696) <= b and not a;
    layer6_outputs(8697) <= b;
    layer6_outputs(8698) <= a and b;
    layer6_outputs(8699) <= b;
    layer6_outputs(8700) <= a and b;
    layer6_outputs(8701) <= b;
    layer6_outputs(8702) <= a and not b;
    layer6_outputs(8703) <= not (a or b);
    layer6_outputs(8704) <= b;
    layer6_outputs(8705) <= b;
    layer6_outputs(8706) <= not (a or b);
    layer6_outputs(8707) <= a or b;
    layer6_outputs(8708) <= not a;
    layer6_outputs(8709) <= not (a or b);
    layer6_outputs(8710) <= 1'b0;
    layer6_outputs(8711) <= a;
    layer6_outputs(8712) <= b;
    layer6_outputs(8713) <= 1'b0;
    layer6_outputs(8714) <= a and not b;
    layer6_outputs(8715) <= not (a xor b);
    layer6_outputs(8716) <= b and not a;
    layer6_outputs(8717) <= b;
    layer6_outputs(8718) <= not b or a;
    layer6_outputs(8719) <= a xor b;
    layer6_outputs(8720) <= b;
    layer6_outputs(8721) <= not a or b;
    layer6_outputs(8722) <= not a;
    layer6_outputs(8723) <= a and b;
    layer6_outputs(8724) <= 1'b1;
    layer6_outputs(8725) <= not (a xor b);
    layer6_outputs(8726) <= not a;
    layer6_outputs(8727) <= not b or a;
    layer6_outputs(8728) <= not (a or b);
    layer6_outputs(8729) <= a and b;
    layer6_outputs(8730) <= not a;
    layer6_outputs(8731) <= a and b;
    layer6_outputs(8732) <= a;
    layer6_outputs(8733) <= not a or b;
    layer6_outputs(8734) <= a;
    layer6_outputs(8735) <= not a or b;
    layer6_outputs(8736) <= a;
    layer6_outputs(8737) <= not b or a;
    layer6_outputs(8738) <= not a or b;
    layer6_outputs(8739) <= b;
    layer6_outputs(8740) <= not a or b;
    layer6_outputs(8741) <= a and not b;
    layer6_outputs(8742) <= not a;
    layer6_outputs(8743) <= b;
    layer6_outputs(8744) <= not b or a;
    layer6_outputs(8745) <= a or b;
    layer6_outputs(8746) <= a and b;
    layer6_outputs(8747) <= not (a and b);
    layer6_outputs(8748) <= a xor b;
    layer6_outputs(8749) <= not (a xor b);
    layer6_outputs(8750) <= not b;
    layer6_outputs(8751) <= not b;
    layer6_outputs(8752) <= a or b;
    layer6_outputs(8753) <= not (a xor b);
    layer6_outputs(8754) <= not b;
    layer6_outputs(8755) <= a;
    layer6_outputs(8756) <= a;
    layer6_outputs(8757) <= not a;
    layer6_outputs(8758) <= not a;
    layer6_outputs(8759) <= b and not a;
    layer6_outputs(8760) <= not b or a;
    layer6_outputs(8761) <= not b;
    layer6_outputs(8762) <= a and not b;
    layer6_outputs(8763) <= not a;
    layer6_outputs(8764) <= b;
    layer6_outputs(8765) <= not a;
    layer6_outputs(8766) <= not b;
    layer6_outputs(8767) <= 1'b1;
    layer6_outputs(8768) <= a and b;
    layer6_outputs(8769) <= not b;
    layer6_outputs(8770) <= b;
    layer6_outputs(8771) <= a and b;
    layer6_outputs(8772) <= not (a and b);
    layer6_outputs(8773) <= a xor b;
    layer6_outputs(8774) <= a;
    layer6_outputs(8775) <= 1'b0;
    layer6_outputs(8776) <= not b;
    layer6_outputs(8777) <= a and b;
    layer6_outputs(8778) <= not (a and b);
    layer6_outputs(8779) <= not a;
    layer6_outputs(8780) <= not a;
    layer6_outputs(8781) <= not b;
    layer6_outputs(8782) <= not b or a;
    layer6_outputs(8783) <= not a;
    layer6_outputs(8784) <= b;
    layer6_outputs(8785) <= b;
    layer6_outputs(8786) <= not a;
    layer6_outputs(8787) <= not b;
    layer6_outputs(8788) <= a xor b;
    layer6_outputs(8789) <= b;
    layer6_outputs(8790) <= not (a or b);
    layer6_outputs(8791) <= a;
    layer6_outputs(8792) <= not a;
    layer6_outputs(8793) <= 1'b0;
    layer6_outputs(8794) <= not (a or b);
    layer6_outputs(8795) <= b;
    layer6_outputs(8796) <= not b or a;
    layer6_outputs(8797) <= not (a or b);
    layer6_outputs(8798) <= not b or a;
    layer6_outputs(8799) <= not b;
    layer6_outputs(8800) <= 1'b0;
    layer6_outputs(8801) <= not b;
    layer6_outputs(8802) <= not (a and b);
    layer6_outputs(8803) <= b and not a;
    layer6_outputs(8804) <= not b;
    layer6_outputs(8805) <= not a or b;
    layer6_outputs(8806) <= not (a and b);
    layer6_outputs(8807) <= a;
    layer6_outputs(8808) <= not b;
    layer6_outputs(8809) <= not a;
    layer6_outputs(8810) <= b;
    layer6_outputs(8811) <= b;
    layer6_outputs(8812) <= a;
    layer6_outputs(8813) <= a or b;
    layer6_outputs(8814) <= not (a xor b);
    layer6_outputs(8815) <= b;
    layer6_outputs(8816) <= a and b;
    layer6_outputs(8817) <= not (a and b);
    layer6_outputs(8818) <= b and not a;
    layer6_outputs(8819) <= not a;
    layer6_outputs(8820) <= a;
    layer6_outputs(8821) <= not b or a;
    layer6_outputs(8822) <= a and b;
    layer6_outputs(8823) <= b;
    layer6_outputs(8824) <= not (a or b);
    layer6_outputs(8825) <= a or b;
    layer6_outputs(8826) <= not b or a;
    layer6_outputs(8827) <= a and b;
    layer6_outputs(8828) <= not a;
    layer6_outputs(8829) <= not (a and b);
    layer6_outputs(8830) <= 1'b0;
    layer6_outputs(8831) <= not a;
    layer6_outputs(8832) <= not (a and b);
    layer6_outputs(8833) <= not (a or b);
    layer6_outputs(8834) <= not a;
    layer6_outputs(8835) <= not (a or b);
    layer6_outputs(8836) <= not (a and b);
    layer6_outputs(8837) <= a and b;
    layer6_outputs(8838) <= a and b;
    layer6_outputs(8839) <= a xor b;
    layer6_outputs(8840) <= a xor b;
    layer6_outputs(8841) <= a or b;
    layer6_outputs(8842) <= a or b;
    layer6_outputs(8843) <= b and not a;
    layer6_outputs(8844) <= a;
    layer6_outputs(8845) <= not b;
    layer6_outputs(8846) <= not b;
    layer6_outputs(8847) <= not a;
    layer6_outputs(8848) <= not (a or b);
    layer6_outputs(8849) <= a;
    layer6_outputs(8850) <= b and not a;
    layer6_outputs(8851) <= not a;
    layer6_outputs(8852) <= not a;
    layer6_outputs(8853) <= b;
    layer6_outputs(8854) <= a and not b;
    layer6_outputs(8855) <= b;
    layer6_outputs(8856) <= a;
    layer6_outputs(8857) <= not (a xor b);
    layer6_outputs(8858) <= not b;
    layer6_outputs(8859) <= not b or a;
    layer6_outputs(8860) <= not (a and b);
    layer6_outputs(8861) <= a;
    layer6_outputs(8862) <= a xor b;
    layer6_outputs(8863) <= b;
    layer6_outputs(8864) <= not (a or b);
    layer6_outputs(8865) <= not a;
    layer6_outputs(8866) <= not b or a;
    layer6_outputs(8867) <= 1'b1;
    layer6_outputs(8868) <= not a;
    layer6_outputs(8869) <= not a;
    layer6_outputs(8870) <= not (a or b);
    layer6_outputs(8871) <= b;
    layer6_outputs(8872) <= b;
    layer6_outputs(8873) <= not (a and b);
    layer6_outputs(8874) <= not b;
    layer6_outputs(8875) <= b;
    layer6_outputs(8876) <= not b;
    layer6_outputs(8877) <= b and not a;
    layer6_outputs(8878) <= b;
    layer6_outputs(8879) <= not a;
    layer6_outputs(8880) <= not (a xor b);
    layer6_outputs(8881) <= 1'b0;
    layer6_outputs(8882) <= a;
    layer6_outputs(8883) <= a xor b;
    layer6_outputs(8884) <= a;
    layer6_outputs(8885) <= a and not b;
    layer6_outputs(8886) <= not (a or b);
    layer6_outputs(8887) <= not a or b;
    layer6_outputs(8888) <= a;
    layer6_outputs(8889) <= a and b;
    layer6_outputs(8890) <= not b;
    layer6_outputs(8891) <= b;
    layer6_outputs(8892) <= not (a xor b);
    layer6_outputs(8893) <= a;
    layer6_outputs(8894) <= not a;
    layer6_outputs(8895) <= a xor b;
    layer6_outputs(8896) <= not a;
    layer6_outputs(8897) <= not a;
    layer6_outputs(8898) <= b;
    layer6_outputs(8899) <= a or b;
    layer6_outputs(8900) <= not a;
    layer6_outputs(8901) <= b and not a;
    layer6_outputs(8902) <= b;
    layer6_outputs(8903) <= b;
    layer6_outputs(8904) <= a xor b;
    layer6_outputs(8905) <= b and not a;
    layer6_outputs(8906) <= not b;
    layer6_outputs(8907) <= a;
    layer6_outputs(8908) <= b;
    layer6_outputs(8909) <= not (a or b);
    layer6_outputs(8910) <= not a or b;
    layer6_outputs(8911) <= not (a or b);
    layer6_outputs(8912) <= not b;
    layer6_outputs(8913) <= b;
    layer6_outputs(8914) <= a;
    layer6_outputs(8915) <= 1'b0;
    layer6_outputs(8916) <= not a or b;
    layer6_outputs(8917) <= not a;
    layer6_outputs(8918) <= not a;
    layer6_outputs(8919) <= b and not a;
    layer6_outputs(8920) <= not (a and b);
    layer6_outputs(8921) <= not (a xor b);
    layer6_outputs(8922) <= b and not a;
    layer6_outputs(8923) <= a or b;
    layer6_outputs(8924) <= a;
    layer6_outputs(8925) <= a and b;
    layer6_outputs(8926) <= not (a or b);
    layer6_outputs(8927) <= a or b;
    layer6_outputs(8928) <= a;
    layer6_outputs(8929) <= a and not b;
    layer6_outputs(8930) <= not a;
    layer6_outputs(8931) <= b and not a;
    layer6_outputs(8932) <= a;
    layer6_outputs(8933) <= not b;
    layer6_outputs(8934) <= 1'b0;
    layer6_outputs(8935) <= not b or a;
    layer6_outputs(8936) <= b;
    layer6_outputs(8937) <= not a;
    layer6_outputs(8938) <= a;
    layer6_outputs(8939) <= b;
    layer6_outputs(8940) <= not b or a;
    layer6_outputs(8941) <= a;
    layer6_outputs(8942) <= b;
    layer6_outputs(8943) <= b;
    layer6_outputs(8944) <= a and b;
    layer6_outputs(8945) <= a and b;
    layer6_outputs(8946) <= not b;
    layer6_outputs(8947) <= a and not b;
    layer6_outputs(8948) <= b and not a;
    layer6_outputs(8949) <= a;
    layer6_outputs(8950) <= a and b;
    layer6_outputs(8951) <= not a or b;
    layer6_outputs(8952) <= b;
    layer6_outputs(8953) <= a and not b;
    layer6_outputs(8954) <= a and b;
    layer6_outputs(8955) <= not (a and b);
    layer6_outputs(8956) <= a xor b;
    layer6_outputs(8957) <= a;
    layer6_outputs(8958) <= a and not b;
    layer6_outputs(8959) <= not a or b;
    layer6_outputs(8960) <= a and b;
    layer6_outputs(8961) <= a and b;
    layer6_outputs(8962) <= not a or b;
    layer6_outputs(8963) <= a and b;
    layer6_outputs(8964) <= not a;
    layer6_outputs(8965) <= b and not a;
    layer6_outputs(8966) <= b;
    layer6_outputs(8967) <= not a;
    layer6_outputs(8968) <= b and not a;
    layer6_outputs(8969) <= a;
    layer6_outputs(8970) <= a xor b;
    layer6_outputs(8971) <= not a;
    layer6_outputs(8972) <= a and b;
    layer6_outputs(8973) <= a;
    layer6_outputs(8974) <= not (a xor b);
    layer6_outputs(8975) <= a and not b;
    layer6_outputs(8976) <= not b or a;
    layer6_outputs(8977) <= not b;
    layer6_outputs(8978) <= not b;
    layer6_outputs(8979) <= not (a xor b);
    layer6_outputs(8980) <= not b;
    layer6_outputs(8981) <= 1'b1;
    layer6_outputs(8982) <= a or b;
    layer6_outputs(8983) <= 1'b0;
    layer6_outputs(8984) <= not b or a;
    layer6_outputs(8985) <= 1'b1;
    layer6_outputs(8986) <= not (a or b);
    layer6_outputs(8987) <= not a or b;
    layer6_outputs(8988) <= a;
    layer6_outputs(8989) <= not a;
    layer6_outputs(8990) <= a and not b;
    layer6_outputs(8991) <= a;
    layer6_outputs(8992) <= a xor b;
    layer6_outputs(8993) <= not a;
    layer6_outputs(8994) <= not b;
    layer6_outputs(8995) <= b;
    layer6_outputs(8996) <= 1'b1;
    layer6_outputs(8997) <= not b;
    layer6_outputs(8998) <= a;
    layer6_outputs(8999) <= not b;
    layer6_outputs(9000) <= a;
    layer6_outputs(9001) <= not a or b;
    layer6_outputs(9002) <= not (a or b);
    layer6_outputs(9003) <= a;
    layer6_outputs(9004) <= not (a xor b);
    layer6_outputs(9005) <= not a or b;
    layer6_outputs(9006) <= not a;
    layer6_outputs(9007) <= not a;
    layer6_outputs(9008) <= a or b;
    layer6_outputs(9009) <= a and not b;
    layer6_outputs(9010) <= a;
    layer6_outputs(9011) <= not (a xor b);
    layer6_outputs(9012) <= not a;
    layer6_outputs(9013) <= not b;
    layer6_outputs(9014) <= a xor b;
    layer6_outputs(9015) <= not b;
    layer6_outputs(9016) <= not b;
    layer6_outputs(9017) <= 1'b0;
    layer6_outputs(9018) <= not b;
    layer6_outputs(9019) <= 1'b0;
    layer6_outputs(9020) <= b and not a;
    layer6_outputs(9021) <= b and not a;
    layer6_outputs(9022) <= a;
    layer6_outputs(9023) <= not b;
    layer6_outputs(9024) <= a;
    layer6_outputs(9025) <= not (a or b);
    layer6_outputs(9026) <= not (a xor b);
    layer6_outputs(9027) <= a or b;
    layer6_outputs(9028) <= not a;
    layer6_outputs(9029) <= b;
    layer6_outputs(9030) <= b;
    layer6_outputs(9031) <= a xor b;
    layer6_outputs(9032) <= not b or a;
    layer6_outputs(9033) <= not a or b;
    layer6_outputs(9034) <= a or b;
    layer6_outputs(9035) <= not (a xor b);
    layer6_outputs(9036) <= not b;
    layer6_outputs(9037) <= b;
    layer6_outputs(9038) <= a;
    layer6_outputs(9039) <= not b;
    layer6_outputs(9040) <= a;
    layer6_outputs(9041) <= not (a xor b);
    layer6_outputs(9042) <= not (a xor b);
    layer6_outputs(9043) <= not (a or b);
    layer6_outputs(9044) <= not b;
    layer6_outputs(9045) <= a and b;
    layer6_outputs(9046) <= b;
    layer6_outputs(9047) <= a and not b;
    layer6_outputs(9048) <= a and b;
    layer6_outputs(9049) <= not (a or b);
    layer6_outputs(9050) <= a;
    layer6_outputs(9051) <= a;
    layer6_outputs(9052) <= a;
    layer6_outputs(9053) <= not (a or b);
    layer6_outputs(9054) <= a and b;
    layer6_outputs(9055) <= a and not b;
    layer6_outputs(9056) <= not b;
    layer6_outputs(9057) <= not b or a;
    layer6_outputs(9058) <= b;
    layer6_outputs(9059) <= a;
    layer6_outputs(9060) <= not (a or b);
    layer6_outputs(9061) <= not a;
    layer6_outputs(9062) <= a xor b;
    layer6_outputs(9063) <= b and not a;
    layer6_outputs(9064) <= a and not b;
    layer6_outputs(9065) <= a and b;
    layer6_outputs(9066) <= a;
    layer6_outputs(9067) <= 1'b1;
    layer6_outputs(9068) <= not a or b;
    layer6_outputs(9069) <= not b or a;
    layer6_outputs(9070) <= not a;
    layer6_outputs(9071) <= not a;
    layer6_outputs(9072) <= not b;
    layer6_outputs(9073) <= a;
    layer6_outputs(9074) <= not b;
    layer6_outputs(9075) <= not a or b;
    layer6_outputs(9076) <= a xor b;
    layer6_outputs(9077) <= a;
    layer6_outputs(9078) <= not b;
    layer6_outputs(9079) <= 1'b1;
    layer6_outputs(9080) <= not (a xor b);
    layer6_outputs(9081) <= not (a and b);
    layer6_outputs(9082) <= b and not a;
    layer6_outputs(9083) <= not a or b;
    layer6_outputs(9084) <= not (a and b);
    layer6_outputs(9085) <= b;
    layer6_outputs(9086) <= a;
    layer6_outputs(9087) <= b and not a;
    layer6_outputs(9088) <= 1'b1;
    layer6_outputs(9089) <= not b;
    layer6_outputs(9090) <= not a;
    layer6_outputs(9091) <= a xor b;
    layer6_outputs(9092) <= not a;
    layer6_outputs(9093) <= not a;
    layer6_outputs(9094) <= a and b;
    layer6_outputs(9095) <= a or b;
    layer6_outputs(9096) <= a;
    layer6_outputs(9097) <= a xor b;
    layer6_outputs(9098) <= not b;
    layer6_outputs(9099) <= not b or a;
    layer6_outputs(9100) <= not b or a;
    layer6_outputs(9101) <= not b;
    layer6_outputs(9102) <= a and not b;
    layer6_outputs(9103) <= not b or a;
    layer6_outputs(9104) <= not (a xor b);
    layer6_outputs(9105) <= not b;
    layer6_outputs(9106) <= a xor b;
    layer6_outputs(9107) <= not b or a;
    layer6_outputs(9108) <= not (a xor b);
    layer6_outputs(9109) <= not b or a;
    layer6_outputs(9110) <= not (a and b);
    layer6_outputs(9111) <= not (a or b);
    layer6_outputs(9112) <= not b;
    layer6_outputs(9113) <= a;
    layer6_outputs(9114) <= a or b;
    layer6_outputs(9115) <= not b;
    layer6_outputs(9116) <= a and not b;
    layer6_outputs(9117) <= a and b;
    layer6_outputs(9118) <= not (a xor b);
    layer6_outputs(9119) <= a xor b;
    layer6_outputs(9120) <= a xor b;
    layer6_outputs(9121) <= a or b;
    layer6_outputs(9122) <= not a;
    layer6_outputs(9123) <= b;
    layer6_outputs(9124) <= b;
    layer6_outputs(9125) <= 1'b0;
    layer6_outputs(9126) <= a;
    layer6_outputs(9127) <= not b;
    layer6_outputs(9128) <= a and b;
    layer6_outputs(9129) <= a and b;
    layer6_outputs(9130) <= not (a and b);
    layer6_outputs(9131) <= a;
    layer6_outputs(9132) <= not a;
    layer6_outputs(9133) <= not (a and b);
    layer6_outputs(9134) <= a and not b;
    layer6_outputs(9135) <= not b;
    layer6_outputs(9136) <= not (a or b);
    layer6_outputs(9137) <= a xor b;
    layer6_outputs(9138) <= a;
    layer6_outputs(9139) <= b;
    layer6_outputs(9140) <= not a or b;
    layer6_outputs(9141) <= not b;
    layer6_outputs(9142) <= not b;
    layer6_outputs(9143) <= a;
    layer6_outputs(9144) <= not a or b;
    layer6_outputs(9145) <= not a;
    layer6_outputs(9146) <= not a or b;
    layer6_outputs(9147) <= not (a xor b);
    layer6_outputs(9148) <= a;
    layer6_outputs(9149) <= not a or b;
    layer6_outputs(9150) <= a;
    layer6_outputs(9151) <= not b or a;
    layer6_outputs(9152) <= b;
    layer6_outputs(9153) <= not (a or b);
    layer6_outputs(9154) <= a;
    layer6_outputs(9155) <= not a or b;
    layer6_outputs(9156) <= not (a and b);
    layer6_outputs(9157) <= b;
    layer6_outputs(9158) <= a;
    layer6_outputs(9159) <= a;
    layer6_outputs(9160) <= a;
    layer6_outputs(9161) <= not a or b;
    layer6_outputs(9162) <= b;
    layer6_outputs(9163) <= not (a or b);
    layer6_outputs(9164) <= not (a and b);
    layer6_outputs(9165) <= not (a xor b);
    layer6_outputs(9166) <= a;
    layer6_outputs(9167) <= not a or b;
    layer6_outputs(9168) <= not a;
    layer6_outputs(9169) <= a;
    layer6_outputs(9170) <= not a;
    layer6_outputs(9171) <= b;
    layer6_outputs(9172) <= a and not b;
    layer6_outputs(9173) <= b;
    layer6_outputs(9174) <= b;
    layer6_outputs(9175) <= a or b;
    layer6_outputs(9176) <= not b;
    layer6_outputs(9177) <= a xor b;
    layer6_outputs(9178) <= b;
    layer6_outputs(9179) <= b and not a;
    layer6_outputs(9180) <= 1'b1;
    layer6_outputs(9181) <= 1'b0;
    layer6_outputs(9182) <= b and not a;
    layer6_outputs(9183) <= not b or a;
    layer6_outputs(9184) <= not a;
    layer6_outputs(9185) <= not (a xor b);
    layer6_outputs(9186) <= a or b;
    layer6_outputs(9187) <= not (a or b);
    layer6_outputs(9188) <= a;
    layer6_outputs(9189) <= a;
    layer6_outputs(9190) <= not a or b;
    layer6_outputs(9191) <= not b;
    layer6_outputs(9192) <= 1'b0;
    layer6_outputs(9193) <= not b;
    layer6_outputs(9194) <= not b;
    layer6_outputs(9195) <= not b;
    layer6_outputs(9196) <= not (a and b);
    layer6_outputs(9197) <= not b;
    layer6_outputs(9198) <= a and b;
    layer6_outputs(9199) <= not b or a;
    layer6_outputs(9200) <= 1'b1;
    layer6_outputs(9201) <= not b;
    layer6_outputs(9202) <= not a;
    layer6_outputs(9203) <= a and b;
    layer6_outputs(9204) <= b;
    layer6_outputs(9205) <= not b or a;
    layer6_outputs(9206) <= not b;
    layer6_outputs(9207) <= b;
    layer6_outputs(9208) <= not b or a;
    layer6_outputs(9209) <= b;
    layer6_outputs(9210) <= b;
    layer6_outputs(9211) <= a and not b;
    layer6_outputs(9212) <= a and b;
    layer6_outputs(9213) <= not b;
    layer6_outputs(9214) <= not b or a;
    layer6_outputs(9215) <= not b;
    layer6_outputs(9216) <= b;
    layer6_outputs(9217) <= b and not a;
    layer6_outputs(9218) <= b;
    layer6_outputs(9219) <= 1'b0;
    layer6_outputs(9220) <= not a or b;
    layer6_outputs(9221) <= not b or a;
    layer6_outputs(9222) <= a and b;
    layer6_outputs(9223) <= a;
    layer6_outputs(9224) <= not (a and b);
    layer6_outputs(9225) <= a;
    layer6_outputs(9226) <= a and not b;
    layer6_outputs(9227) <= a and not b;
    layer6_outputs(9228) <= not b;
    layer6_outputs(9229) <= b;
    layer6_outputs(9230) <= not a;
    layer6_outputs(9231) <= 1'b0;
    layer6_outputs(9232) <= a;
    layer6_outputs(9233) <= not b;
    layer6_outputs(9234) <= not b or a;
    layer6_outputs(9235) <= not a;
    layer6_outputs(9236) <= not (a xor b);
    layer6_outputs(9237) <= not (a and b);
    layer6_outputs(9238) <= not b;
    layer6_outputs(9239) <= not b;
    layer6_outputs(9240) <= not b;
    layer6_outputs(9241) <= 1'b1;
    layer6_outputs(9242) <= a or b;
    layer6_outputs(9243) <= 1'b0;
    layer6_outputs(9244) <= not a;
    layer6_outputs(9245) <= not b;
    layer6_outputs(9246) <= not b;
    layer6_outputs(9247) <= not a;
    layer6_outputs(9248) <= not (a xor b);
    layer6_outputs(9249) <= a xor b;
    layer6_outputs(9250) <= not b;
    layer6_outputs(9251) <= a and b;
    layer6_outputs(9252) <= 1'b0;
    layer6_outputs(9253) <= a xor b;
    layer6_outputs(9254) <= b;
    layer6_outputs(9255) <= not (a and b);
    layer6_outputs(9256) <= not a or b;
    layer6_outputs(9257) <= 1'b0;
    layer6_outputs(9258) <= not b or a;
    layer6_outputs(9259) <= a xor b;
    layer6_outputs(9260) <= b and not a;
    layer6_outputs(9261) <= b;
    layer6_outputs(9262) <= a and b;
    layer6_outputs(9263) <= not a;
    layer6_outputs(9264) <= a xor b;
    layer6_outputs(9265) <= a and not b;
    layer6_outputs(9266) <= a and b;
    layer6_outputs(9267) <= a and b;
    layer6_outputs(9268) <= a;
    layer6_outputs(9269) <= a;
    layer6_outputs(9270) <= a;
    layer6_outputs(9271) <= 1'b0;
    layer6_outputs(9272) <= b and not a;
    layer6_outputs(9273) <= not b;
    layer6_outputs(9274) <= not a;
    layer6_outputs(9275) <= not (a or b);
    layer6_outputs(9276) <= not (a xor b);
    layer6_outputs(9277) <= a and b;
    layer6_outputs(9278) <= not (a or b);
    layer6_outputs(9279) <= not (a or b);
    layer6_outputs(9280) <= a and b;
    layer6_outputs(9281) <= not (a xor b);
    layer6_outputs(9282) <= a or b;
    layer6_outputs(9283) <= not b;
    layer6_outputs(9284) <= not a;
    layer6_outputs(9285) <= not b or a;
    layer6_outputs(9286) <= a or b;
    layer6_outputs(9287) <= not (a or b);
    layer6_outputs(9288) <= not b;
    layer6_outputs(9289) <= a xor b;
    layer6_outputs(9290) <= 1'b0;
    layer6_outputs(9291) <= a and b;
    layer6_outputs(9292) <= b;
    layer6_outputs(9293) <= not a;
    layer6_outputs(9294) <= a;
    layer6_outputs(9295) <= not (a or b);
    layer6_outputs(9296) <= not b;
    layer6_outputs(9297) <= not (a and b);
    layer6_outputs(9298) <= a and not b;
    layer6_outputs(9299) <= b;
    layer6_outputs(9300) <= not b;
    layer6_outputs(9301) <= a and not b;
    layer6_outputs(9302) <= a xor b;
    layer6_outputs(9303) <= not a or b;
    layer6_outputs(9304) <= not (a or b);
    layer6_outputs(9305) <= b and not a;
    layer6_outputs(9306) <= a xor b;
    layer6_outputs(9307) <= not b;
    layer6_outputs(9308) <= not b;
    layer6_outputs(9309) <= 1'b0;
    layer6_outputs(9310) <= not (a xor b);
    layer6_outputs(9311) <= not a;
    layer6_outputs(9312) <= not b;
    layer6_outputs(9313) <= a and not b;
    layer6_outputs(9314) <= not b or a;
    layer6_outputs(9315) <= b and not a;
    layer6_outputs(9316) <= 1'b1;
    layer6_outputs(9317) <= not a;
    layer6_outputs(9318) <= not (a xor b);
    layer6_outputs(9319) <= not (a or b);
    layer6_outputs(9320) <= a;
    layer6_outputs(9321) <= not b or a;
    layer6_outputs(9322) <= not b;
    layer6_outputs(9323) <= not (a xor b);
    layer6_outputs(9324) <= not a;
    layer6_outputs(9325) <= not a;
    layer6_outputs(9326) <= a;
    layer6_outputs(9327) <= not b;
    layer6_outputs(9328) <= not b;
    layer6_outputs(9329) <= a xor b;
    layer6_outputs(9330) <= b and not a;
    layer6_outputs(9331) <= a xor b;
    layer6_outputs(9332) <= a;
    layer6_outputs(9333) <= not b or a;
    layer6_outputs(9334) <= a or b;
    layer6_outputs(9335) <= not (a or b);
    layer6_outputs(9336) <= not a;
    layer6_outputs(9337) <= b and not a;
    layer6_outputs(9338) <= not b;
    layer6_outputs(9339) <= not (a or b);
    layer6_outputs(9340) <= not (a xor b);
    layer6_outputs(9341) <= not b;
    layer6_outputs(9342) <= not (a xor b);
    layer6_outputs(9343) <= a and not b;
    layer6_outputs(9344) <= 1'b0;
    layer6_outputs(9345) <= not b;
    layer6_outputs(9346) <= 1'b1;
    layer6_outputs(9347) <= not a;
    layer6_outputs(9348) <= b;
    layer6_outputs(9349) <= 1'b0;
    layer6_outputs(9350) <= b and not a;
    layer6_outputs(9351) <= not b;
    layer6_outputs(9352) <= not (a xor b);
    layer6_outputs(9353) <= not (a and b);
    layer6_outputs(9354) <= a xor b;
    layer6_outputs(9355) <= b;
    layer6_outputs(9356) <= not a;
    layer6_outputs(9357) <= not (a or b);
    layer6_outputs(9358) <= b;
    layer6_outputs(9359) <= not a or b;
    layer6_outputs(9360) <= not b or a;
    layer6_outputs(9361) <= not a;
    layer6_outputs(9362) <= a xor b;
    layer6_outputs(9363) <= not b;
    layer6_outputs(9364) <= not (a or b);
    layer6_outputs(9365) <= b;
    layer6_outputs(9366) <= not b or a;
    layer6_outputs(9367) <= not a;
    layer6_outputs(9368) <= not b;
    layer6_outputs(9369) <= b;
    layer6_outputs(9370) <= not b;
    layer6_outputs(9371) <= not a or b;
    layer6_outputs(9372) <= not a;
    layer6_outputs(9373) <= b;
    layer6_outputs(9374) <= not b;
    layer6_outputs(9375) <= not (a and b);
    layer6_outputs(9376) <= b and not a;
    layer6_outputs(9377) <= a and not b;
    layer6_outputs(9378) <= a;
    layer6_outputs(9379) <= b;
    layer6_outputs(9380) <= b;
    layer6_outputs(9381) <= not b or a;
    layer6_outputs(9382) <= 1'b0;
    layer6_outputs(9383) <= a xor b;
    layer6_outputs(9384) <= a;
    layer6_outputs(9385) <= not a;
    layer6_outputs(9386) <= not a or b;
    layer6_outputs(9387) <= not (a and b);
    layer6_outputs(9388) <= not a or b;
    layer6_outputs(9389) <= not a;
    layer6_outputs(9390) <= a and b;
    layer6_outputs(9391) <= a;
    layer6_outputs(9392) <= not b or a;
    layer6_outputs(9393) <= not (a and b);
    layer6_outputs(9394) <= b and not a;
    layer6_outputs(9395) <= not b;
    layer6_outputs(9396) <= a;
    layer6_outputs(9397) <= not (a or b);
    layer6_outputs(9398) <= not (a xor b);
    layer6_outputs(9399) <= not (a or b);
    layer6_outputs(9400) <= not a or b;
    layer6_outputs(9401) <= not a or b;
    layer6_outputs(9402) <= not b;
    layer6_outputs(9403) <= not (a and b);
    layer6_outputs(9404) <= a and not b;
    layer6_outputs(9405) <= not (a xor b);
    layer6_outputs(9406) <= not a;
    layer6_outputs(9407) <= a;
    layer6_outputs(9408) <= not a;
    layer6_outputs(9409) <= a and not b;
    layer6_outputs(9410) <= a;
    layer6_outputs(9411) <= not b;
    layer6_outputs(9412) <= not a;
    layer6_outputs(9413) <= b;
    layer6_outputs(9414) <= not b or a;
    layer6_outputs(9415) <= a xor b;
    layer6_outputs(9416) <= not (a or b);
    layer6_outputs(9417) <= not b;
    layer6_outputs(9418) <= not a;
    layer6_outputs(9419) <= a xor b;
    layer6_outputs(9420) <= not (a or b);
    layer6_outputs(9421) <= a xor b;
    layer6_outputs(9422) <= not b or a;
    layer6_outputs(9423) <= not b or a;
    layer6_outputs(9424) <= not (a or b);
    layer6_outputs(9425) <= not (a xor b);
    layer6_outputs(9426) <= b;
    layer6_outputs(9427) <= not (a and b);
    layer6_outputs(9428) <= b and not a;
    layer6_outputs(9429) <= not a or b;
    layer6_outputs(9430) <= b;
    layer6_outputs(9431) <= not a;
    layer6_outputs(9432) <= a and b;
    layer6_outputs(9433) <= a and b;
    layer6_outputs(9434) <= not b or a;
    layer6_outputs(9435) <= a or b;
    layer6_outputs(9436) <= not b;
    layer6_outputs(9437) <= a and b;
    layer6_outputs(9438) <= not (a xor b);
    layer6_outputs(9439) <= not b;
    layer6_outputs(9440) <= 1'b0;
    layer6_outputs(9441) <= a or b;
    layer6_outputs(9442) <= not a;
    layer6_outputs(9443) <= a and not b;
    layer6_outputs(9444) <= not a;
    layer6_outputs(9445) <= b;
    layer6_outputs(9446) <= not b;
    layer6_outputs(9447) <= not a or b;
    layer6_outputs(9448) <= not b or a;
    layer6_outputs(9449) <= not (a or b);
    layer6_outputs(9450) <= not (a xor b);
    layer6_outputs(9451) <= not (a and b);
    layer6_outputs(9452) <= not a or b;
    layer6_outputs(9453) <= 1'b0;
    layer6_outputs(9454) <= a xor b;
    layer6_outputs(9455) <= not a or b;
    layer6_outputs(9456) <= not a;
    layer6_outputs(9457) <= not b;
    layer6_outputs(9458) <= b and not a;
    layer6_outputs(9459) <= not b or a;
    layer6_outputs(9460) <= not (a xor b);
    layer6_outputs(9461) <= b and not a;
    layer6_outputs(9462) <= not (a xor b);
    layer6_outputs(9463) <= not a;
    layer6_outputs(9464) <= not a;
    layer6_outputs(9465) <= b;
    layer6_outputs(9466) <= b and not a;
    layer6_outputs(9467) <= not a or b;
    layer6_outputs(9468) <= not (a or b);
    layer6_outputs(9469) <= not b or a;
    layer6_outputs(9470) <= not (a or b);
    layer6_outputs(9471) <= b;
    layer6_outputs(9472) <= not b;
    layer6_outputs(9473) <= a;
    layer6_outputs(9474) <= b;
    layer6_outputs(9475) <= a;
    layer6_outputs(9476) <= b;
    layer6_outputs(9477) <= 1'b1;
    layer6_outputs(9478) <= b;
    layer6_outputs(9479) <= b and not a;
    layer6_outputs(9480) <= not a;
    layer6_outputs(9481) <= not a or b;
    layer6_outputs(9482) <= a and not b;
    layer6_outputs(9483) <= a;
    layer6_outputs(9484) <= b and not a;
    layer6_outputs(9485) <= a xor b;
    layer6_outputs(9486) <= b;
    layer6_outputs(9487) <= not a;
    layer6_outputs(9488) <= 1'b0;
    layer6_outputs(9489) <= not a or b;
    layer6_outputs(9490) <= not b;
    layer6_outputs(9491) <= b and not a;
    layer6_outputs(9492) <= b and not a;
    layer6_outputs(9493) <= not b or a;
    layer6_outputs(9494) <= not a;
    layer6_outputs(9495) <= not (a and b);
    layer6_outputs(9496) <= not a;
    layer6_outputs(9497) <= a or b;
    layer6_outputs(9498) <= not b or a;
    layer6_outputs(9499) <= not b;
    layer6_outputs(9500) <= a and b;
    layer6_outputs(9501) <= not b or a;
    layer6_outputs(9502) <= not a;
    layer6_outputs(9503) <= not b;
    layer6_outputs(9504) <= not (a and b);
    layer6_outputs(9505) <= b and not a;
    layer6_outputs(9506) <= not a;
    layer6_outputs(9507) <= not b;
    layer6_outputs(9508) <= a and not b;
    layer6_outputs(9509) <= a;
    layer6_outputs(9510) <= a;
    layer6_outputs(9511) <= a xor b;
    layer6_outputs(9512) <= b;
    layer6_outputs(9513) <= 1'b1;
    layer6_outputs(9514) <= a;
    layer6_outputs(9515) <= a;
    layer6_outputs(9516) <= not b;
    layer6_outputs(9517) <= not a;
    layer6_outputs(9518) <= not a;
    layer6_outputs(9519) <= not b or a;
    layer6_outputs(9520) <= a xor b;
    layer6_outputs(9521) <= not (a xor b);
    layer6_outputs(9522) <= a;
    layer6_outputs(9523) <= a and b;
    layer6_outputs(9524) <= not (a and b);
    layer6_outputs(9525) <= not (a xor b);
    layer6_outputs(9526) <= not (a xor b);
    layer6_outputs(9527) <= not b or a;
    layer6_outputs(9528) <= a and b;
    layer6_outputs(9529) <= a xor b;
    layer6_outputs(9530) <= b;
    layer6_outputs(9531) <= not a;
    layer6_outputs(9532) <= a and not b;
    layer6_outputs(9533) <= b;
    layer6_outputs(9534) <= a;
    layer6_outputs(9535) <= a xor b;
    layer6_outputs(9536) <= not b;
    layer6_outputs(9537) <= not (a and b);
    layer6_outputs(9538) <= b;
    layer6_outputs(9539) <= b;
    layer6_outputs(9540) <= not (a and b);
    layer6_outputs(9541) <= a and b;
    layer6_outputs(9542) <= a and not b;
    layer6_outputs(9543) <= not a;
    layer6_outputs(9544) <= not b;
    layer6_outputs(9545) <= not b;
    layer6_outputs(9546) <= a;
    layer6_outputs(9547) <= a and not b;
    layer6_outputs(9548) <= a and not b;
    layer6_outputs(9549) <= b;
    layer6_outputs(9550) <= not b;
    layer6_outputs(9551) <= not a;
    layer6_outputs(9552) <= b;
    layer6_outputs(9553) <= 1'b0;
    layer6_outputs(9554) <= not b;
    layer6_outputs(9555) <= not (a or b);
    layer6_outputs(9556) <= b and not a;
    layer6_outputs(9557) <= a xor b;
    layer6_outputs(9558) <= a;
    layer6_outputs(9559) <= not b;
    layer6_outputs(9560) <= not (a or b);
    layer6_outputs(9561) <= b and not a;
    layer6_outputs(9562) <= not b or a;
    layer6_outputs(9563) <= 1'b1;
    layer6_outputs(9564) <= a or b;
    layer6_outputs(9565) <= b;
    layer6_outputs(9566) <= not a;
    layer6_outputs(9567) <= not (a or b);
    layer6_outputs(9568) <= not a;
    layer6_outputs(9569) <= not b;
    layer6_outputs(9570) <= not b or a;
    layer6_outputs(9571) <= not a;
    layer6_outputs(9572) <= a and b;
    layer6_outputs(9573) <= b;
    layer6_outputs(9574) <= a and not b;
    layer6_outputs(9575) <= not b;
    layer6_outputs(9576) <= a and b;
    layer6_outputs(9577) <= not a;
    layer6_outputs(9578) <= a xor b;
    layer6_outputs(9579) <= 1'b0;
    layer6_outputs(9580) <= b;
    layer6_outputs(9581) <= not b or a;
    layer6_outputs(9582) <= 1'b0;
    layer6_outputs(9583) <= b and not a;
    layer6_outputs(9584) <= a and b;
    layer6_outputs(9585) <= b;
    layer6_outputs(9586) <= not b;
    layer6_outputs(9587) <= not b or a;
    layer6_outputs(9588) <= a;
    layer6_outputs(9589) <= a or b;
    layer6_outputs(9590) <= a or b;
    layer6_outputs(9591) <= b and not a;
    layer6_outputs(9592) <= a or b;
    layer6_outputs(9593) <= not (a or b);
    layer6_outputs(9594) <= not a or b;
    layer6_outputs(9595) <= not b or a;
    layer6_outputs(9596) <= b and not a;
    layer6_outputs(9597) <= not (a or b);
    layer6_outputs(9598) <= a;
    layer6_outputs(9599) <= not a or b;
    layer6_outputs(9600) <= 1'b0;
    layer6_outputs(9601) <= b;
    layer6_outputs(9602) <= not a;
    layer6_outputs(9603) <= a;
    layer6_outputs(9604) <= a and b;
    layer6_outputs(9605) <= not (a and b);
    layer6_outputs(9606) <= a;
    layer6_outputs(9607) <= not (a or b);
    layer6_outputs(9608) <= b and not a;
    layer6_outputs(9609) <= a and not b;
    layer6_outputs(9610) <= not (a xor b);
    layer6_outputs(9611) <= not (a and b);
    layer6_outputs(9612) <= b;
    layer6_outputs(9613) <= b;
    layer6_outputs(9614) <= a and b;
    layer6_outputs(9615) <= a or b;
    layer6_outputs(9616) <= not (a and b);
    layer6_outputs(9617) <= not b;
    layer6_outputs(9618) <= b;
    layer6_outputs(9619) <= a and b;
    layer6_outputs(9620) <= 1'b0;
    layer6_outputs(9621) <= a or b;
    layer6_outputs(9622) <= a xor b;
    layer6_outputs(9623) <= not b or a;
    layer6_outputs(9624) <= b and not a;
    layer6_outputs(9625) <= not a;
    layer6_outputs(9626) <= not (a and b);
    layer6_outputs(9627) <= a and b;
    layer6_outputs(9628) <= not (a and b);
    layer6_outputs(9629) <= not b;
    layer6_outputs(9630) <= b and not a;
    layer6_outputs(9631) <= a and not b;
    layer6_outputs(9632) <= a and b;
    layer6_outputs(9633) <= not (a and b);
    layer6_outputs(9634) <= not a or b;
    layer6_outputs(9635) <= not (a xor b);
    layer6_outputs(9636) <= a;
    layer6_outputs(9637) <= 1'b1;
    layer6_outputs(9638) <= not b or a;
    layer6_outputs(9639) <= not (a and b);
    layer6_outputs(9640) <= a and not b;
    layer6_outputs(9641) <= not (a and b);
    layer6_outputs(9642) <= b;
    layer6_outputs(9643) <= a and not b;
    layer6_outputs(9644) <= a;
    layer6_outputs(9645) <= a and b;
    layer6_outputs(9646) <= not (a xor b);
    layer6_outputs(9647) <= not a;
    layer6_outputs(9648) <= a;
    layer6_outputs(9649) <= not b or a;
    layer6_outputs(9650) <= not b;
    layer6_outputs(9651) <= not b;
    layer6_outputs(9652) <= not b;
    layer6_outputs(9653) <= not (a xor b);
    layer6_outputs(9654) <= b and not a;
    layer6_outputs(9655) <= not a;
    layer6_outputs(9656) <= a xor b;
    layer6_outputs(9657) <= not a;
    layer6_outputs(9658) <= not (a and b);
    layer6_outputs(9659) <= not a or b;
    layer6_outputs(9660) <= 1'b1;
    layer6_outputs(9661) <= 1'b1;
    layer6_outputs(9662) <= b;
    layer6_outputs(9663) <= not a;
    layer6_outputs(9664) <= not (a xor b);
    layer6_outputs(9665) <= a or b;
    layer6_outputs(9666) <= not b;
    layer6_outputs(9667) <= not b or a;
    layer6_outputs(9668) <= not a or b;
    layer6_outputs(9669) <= a and not b;
    layer6_outputs(9670) <= not a;
    layer6_outputs(9671) <= not b or a;
    layer6_outputs(9672) <= a and not b;
    layer6_outputs(9673) <= a;
    layer6_outputs(9674) <= a and not b;
    layer6_outputs(9675) <= not a;
    layer6_outputs(9676) <= not a or b;
    layer6_outputs(9677) <= not (a and b);
    layer6_outputs(9678) <= a or b;
    layer6_outputs(9679) <= not a or b;
    layer6_outputs(9680) <= a xor b;
    layer6_outputs(9681) <= not (a xor b);
    layer6_outputs(9682) <= a;
    layer6_outputs(9683) <= a and not b;
    layer6_outputs(9684) <= not (a and b);
    layer6_outputs(9685) <= a;
    layer6_outputs(9686) <= b and not a;
    layer6_outputs(9687) <= a and b;
    layer6_outputs(9688) <= not a;
    layer6_outputs(9689) <= not b;
    layer6_outputs(9690) <= not a;
    layer6_outputs(9691) <= a;
    layer6_outputs(9692) <= not (a and b);
    layer6_outputs(9693) <= not a or b;
    layer6_outputs(9694) <= not b;
    layer6_outputs(9695) <= a xor b;
    layer6_outputs(9696) <= a or b;
    layer6_outputs(9697) <= b;
    layer6_outputs(9698) <= not b or a;
    layer6_outputs(9699) <= not a;
    layer6_outputs(9700) <= not a;
    layer6_outputs(9701) <= a;
    layer6_outputs(9702) <= a;
    layer6_outputs(9703) <= not b;
    layer6_outputs(9704) <= a;
    layer6_outputs(9705) <= not a;
    layer6_outputs(9706) <= not a;
    layer6_outputs(9707) <= 1'b1;
    layer6_outputs(9708) <= a;
    layer6_outputs(9709) <= b and not a;
    layer6_outputs(9710) <= 1'b0;
    layer6_outputs(9711) <= not (a and b);
    layer6_outputs(9712) <= not (a and b);
    layer6_outputs(9713) <= a and not b;
    layer6_outputs(9714) <= not (a or b);
    layer6_outputs(9715) <= not (a xor b);
    layer6_outputs(9716) <= a or b;
    layer6_outputs(9717) <= not b;
    layer6_outputs(9718) <= b;
    layer6_outputs(9719) <= not b;
    layer6_outputs(9720) <= not a;
    layer6_outputs(9721) <= not a;
    layer6_outputs(9722) <= b;
    layer6_outputs(9723) <= b;
    layer6_outputs(9724) <= not (a and b);
    layer6_outputs(9725) <= 1'b1;
    layer6_outputs(9726) <= not b;
    layer6_outputs(9727) <= a and not b;
    layer6_outputs(9728) <= a;
    layer6_outputs(9729) <= a;
    layer6_outputs(9730) <= not (a or b);
    layer6_outputs(9731) <= b;
    layer6_outputs(9732) <= a;
    layer6_outputs(9733) <= a and not b;
    layer6_outputs(9734) <= not b;
    layer6_outputs(9735) <= not (a or b);
    layer6_outputs(9736) <= not a;
    layer6_outputs(9737) <= b;
    layer6_outputs(9738) <= b;
    layer6_outputs(9739) <= a or b;
    layer6_outputs(9740) <= 1'b1;
    layer6_outputs(9741) <= not (a or b);
    layer6_outputs(9742) <= b and not a;
    layer6_outputs(9743) <= b;
    layer6_outputs(9744) <= b and not a;
    layer6_outputs(9745) <= not b or a;
    layer6_outputs(9746) <= a;
    layer6_outputs(9747) <= not (a or b);
    layer6_outputs(9748) <= not (a or b);
    layer6_outputs(9749) <= not a;
    layer6_outputs(9750) <= b;
    layer6_outputs(9751) <= a xor b;
    layer6_outputs(9752) <= not (a and b);
    layer6_outputs(9753) <= b and not a;
    layer6_outputs(9754) <= not b;
    layer6_outputs(9755) <= not (a xor b);
    layer6_outputs(9756) <= not a;
    layer6_outputs(9757) <= b and not a;
    layer6_outputs(9758) <= not b;
    layer6_outputs(9759) <= not a;
    layer6_outputs(9760) <= a;
    layer6_outputs(9761) <= not b or a;
    layer6_outputs(9762) <= not (a and b);
    layer6_outputs(9763) <= not a or b;
    layer6_outputs(9764) <= a and not b;
    layer6_outputs(9765) <= a xor b;
    layer6_outputs(9766) <= 1'b1;
    layer6_outputs(9767) <= not a;
    layer6_outputs(9768) <= not b;
    layer6_outputs(9769) <= a and not b;
    layer6_outputs(9770) <= a xor b;
    layer6_outputs(9771) <= a xor b;
    layer6_outputs(9772) <= a xor b;
    layer6_outputs(9773) <= b;
    layer6_outputs(9774) <= a;
    layer6_outputs(9775) <= not a or b;
    layer6_outputs(9776) <= a or b;
    layer6_outputs(9777) <= b;
    layer6_outputs(9778) <= not a;
    layer6_outputs(9779) <= not a;
    layer6_outputs(9780) <= not b or a;
    layer6_outputs(9781) <= not (a or b);
    layer6_outputs(9782) <= not (a and b);
    layer6_outputs(9783) <= a or b;
    layer6_outputs(9784) <= b and not a;
    layer6_outputs(9785) <= not (a or b);
    layer6_outputs(9786) <= b;
    layer6_outputs(9787) <= a;
    layer6_outputs(9788) <= a and not b;
    layer6_outputs(9789) <= not b;
    layer6_outputs(9790) <= a or b;
    layer6_outputs(9791) <= a;
    layer6_outputs(9792) <= not a or b;
    layer6_outputs(9793) <= a;
    layer6_outputs(9794) <= b;
    layer6_outputs(9795) <= not a or b;
    layer6_outputs(9796) <= 1'b0;
    layer6_outputs(9797) <= a or b;
    layer6_outputs(9798) <= b and not a;
    layer6_outputs(9799) <= not (a and b);
    layer6_outputs(9800) <= not (a or b);
    layer6_outputs(9801) <= not (a xor b);
    layer6_outputs(9802) <= not b or a;
    layer6_outputs(9803) <= a xor b;
    layer6_outputs(9804) <= not a or b;
    layer6_outputs(9805) <= not a or b;
    layer6_outputs(9806) <= not a;
    layer6_outputs(9807) <= not (a xor b);
    layer6_outputs(9808) <= not a;
    layer6_outputs(9809) <= not a or b;
    layer6_outputs(9810) <= not a;
    layer6_outputs(9811) <= b and not a;
    layer6_outputs(9812) <= not (a or b);
    layer6_outputs(9813) <= not a or b;
    layer6_outputs(9814) <= not a;
    layer6_outputs(9815) <= a or b;
    layer6_outputs(9816) <= a and b;
    layer6_outputs(9817) <= b;
    layer6_outputs(9818) <= not (a and b);
    layer6_outputs(9819) <= a and not b;
    layer6_outputs(9820) <= a and b;
    layer6_outputs(9821) <= 1'b1;
    layer6_outputs(9822) <= a and b;
    layer6_outputs(9823) <= not b;
    layer6_outputs(9824) <= a and not b;
    layer6_outputs(9825) <= a and not b;
    layer6_outputs(9826) <= not a;
    layer6_outputs(9827) <= a;
    layer6_outputs(9828) <= b;
    layer6_outputs(9829) <= not b;
    layer6_outputs(9830) <= b and not a;
    layer6_outputs(9831) <= b;
    layer6_outputs(9832) <= 1'b0;
    layer6_outputs(9833) <= not (a xor b);
    layer6_outputs(9834) <= not a;
    layer6_outputs(9835) <= not a;
    layer6_outputs(9836) <= a and not b;
    layer6_outputs(9837) <= not b;
    layer6_outputs(9838) <= a and b;
    layer6_outputs(9839) <= not (a xor b);
    layer6_outputs(9840) <= a;
    layer6_outputs(9841) <= not a;
    layer6_outputs(9842) <= b;
    layer6_outputs(9843) <= b and not a;
    layer6_outputs(9844) <= not (a or b);
    layer6_outputs(9845) <= b;
    layer6_outputs(9846) <= not (a and b);
    layer6_outputs(9847) <= not b;
    layer6_outputs(9848) <= not a;
    layer6_outputs(9849) <= not b;
    layer6_outputs(9850) <= not a or b;
    layer6_outputs(9851) <= not b;
    layer6_outputs(9852) <= b and not a;
    layer6_outputs(9853) <= not b or a;
    layer6_outputs(9854) <= b and not a;
    layer6_outputs(9855) <= not b or a;
    layer6_outputs(9856) <= not b or a;
    layer6_outputs(9857) <= a and not b;
    layer6_outputs(9858) <= b;
    layer6_outputs(9859) <= not (a xor b);
    layer6_outputs(9860) <= b;
    layer6_outputs(9861) <= a and not b;
    layer6_outputs(9862) <= not (a and b);
    layer6_outputs(9863) <= b;
    layer6_outputs(9864) <= not (a and b);
    layer6_outputs(9865) <= a and not b;
    layer6_outputs(9866) <= not b;
    layer6_outputs(9867) <= b;
    layer6_outputs(9868) <= a and not b;
    layer6_outputs(9869) <= not (a xor b);
    layer6_outputs(9870) <= not a;
    layer6_outputs(9871) <= not a;
    layer6_outputs(9872) <= not (a and b);
    layer6_outputs(9873) <= not b;
    layer6_outputs(9874) <= not b;
    layer6_outputs(9875) <= not b or a;
    layer6_outputs(9876) <= not b;
    layer6_outputs(9877) <= b and not a;
    layer6_outputs(9878) <= not (a xor b);
    layer6_outputs(9879) <= not a;
    layer6_outputs(9880) <= a;
    layer6_outputs(9881) <= a and not b;
    layer6_outputs(9882) <= a or b;
    layer6_outputs(9883) <= a;
    layer6_outputs(9884) <= a and b;
    layer6_outputs(9885) <= 1'b0;
    layer6_outputs(9886) <= a xor b;
    layer6_outputs(9887) <= not a or b;
    layer6_outputs(9888) <= b;
    layer6_outputs(9889) <= not (a or b);
    layer6_outputs(9890) <= not a;
    layer6_outputs(9891) <= 1'b1;
    layer6_outputs(9892) <= a and not b;
    layer6_outputs(9893) <= not b;
    layer6_outputs(9894) <= a or b;
    layer6_outputs(9895) <= a;
    layer6_outputs(9896) <= not b;
    layer6_outputs(9897) <= a and b;
    layer6_outputs(9898) <= a;
    layer6_outputs(9899) <= not (a xor b);
    layer6_outputs(9900) <= a or b;
    layer6_outputs(9901) <= 1'b1;
    layer6_outputs(9902) <= not a;
    layer6_outputs(9903) <= not a;
    layer6_outputs(9904) <= a;
    layer6_outputs(9905) <= not (a or b);
    layer6_outputs(9906) <= not a;
    layer6_outputs(9907) <= a and not b;
    layer6_outputs(9908) <= a;
    layer6_outputs(9909) <= a and b;
    layer6_outputs(9910) <= b;
    layer6_outputs(9911) <= not b or a;
    layer6_outputs(9912) <= not (a xor b);
    layer6_outputs(9913) <= a or b;
    layer6_outputs(9914) <= not b;
    layer6_outputs(9915) <= a xor b;
    layer6_outputs(9916) <= a or b;
    layer6_outputs(9917) <= a and not b;
    layer6_outputs(9918) <= b;
    layer6_outputs(9919) <= a and b;
    layer6_outputs(9920) <= b;
    layer6_outputs(9921) <= a;
    layer6_outputs(9922) <= not a;
    layer6_outputs(9923) <= a;
    layer6_outputs(9924) <= not a;
    layer6_outputs(9925) <= not a;
    layer6_outputs(9926) <= not b;
    layer6_outputs(9927) <= a or b;
    layer6_outputs(9928) <= a and b;
    layer6_outputs(9929) <= b;
    layer6_outputs(9930) <= not a;
    layer6_outputs(9931) <= 1'b0;
    layer6_outputs(9932) <= not a or b;
    layer6_outputs(9933) <= b;
    layer6_outputs(9934) <= b;
    layer6_outputs(9935) <= b;
    layer6_outputs(9936) <= b;
    layer6_outputs(9937) <= a and not b;
    layer6_outputs(9938) <= not b;
    layer6_outputs(9939) <= b;
    layer6_outputs(9940) <= b;
    layer6_outputs(9941) <= not (a or b);
    layer6_outputs(9942) <= not a;
    layer6_outputs(9943) <= a and not b;
    layer6_outputs(9944) <= a xor b;
    layer6_outputs(9945) <= b;
    layer6_outputs(9946) <= not (a and b);
    layer6_outputs(9947) <= a and b;
    layer6_outputs(9948) <= not a;
    layer6_outputs(9949) <= not a;
    layer6_outputs(9950) <= 1'b0;
    layer6_outputs(9951) <= not (a xor b);
    layer6_outputs(9952) <= b;
    layer6_outputs(9953) <= 1'b0;
    layer6_outputs(9954) <= not (a and b);
    layer6_outputs(9955) <= b;
    layer6_outputs(9956) <= a xor b;
    layer6_outputs(9957) <= b;
    layer6_outputs(9958) <= a;
    layer6_outputs(9959) <= a or b;
    layer6_outputs(9960) <= a and not b;
    layer6_outputs(9961) <= a or b;
    layer6_outputs(9962) <= not (a and b);
    layer6_outputs(9963) <= not b;
    layer6_outputs(9964) <= not b;
    layer6_outputs(9965) <= b and not a;
    layer6_outputs(9966) <= a or b;
    layer6_outputs(9967) <= a and b;
    layer6_outputs(9968) <= a;
    layer6_outputs(9969) <= a and not b;
    layer6_outputs(9970) <= not (a or b);
    layer6_outputs(9971) <= a and not b;
    layer6_outputs(9972) <= not b or a;
    layer6_outputs(9973) <= not a or b;
    layer6_outputs(9974) <= not (a or b);
    layer6_outputs(9975) <= b;
    layer6_outputs(9976) <= not a;
    layer6_outputs(9977) <= not (a and b);
    layer6_outputs(9978) <= not a or b;
    layer6_outputs(9979) <= 1'b1;
    layer6_outputs(9980) <= b;
    layer6_outputs(9981) <= not b or a;
    layer6_outputs(9982) <= a;
    layer6_outputs(9983) <= not a or b;
    layer6_outputs(9984) <= a or b;
    layer6_outputs(9985) <= 1'b0;
    layer6_outputs(9986) <= not b;
    layer6_outputs(9987) <= a xor b;
    layer6_outputs(9988) <= b and not a;
    layer6_outputs(9989) <= b and not a;
    layer6_outputs(9990) <= a xor b;
    layer6_outputs(9991) <= 1'b0;
    layer6_outputs(9992) <= not b or a;
    layer6_outputs(9993) <= b;
    layer6_outputs(9994) <= a;
    layer6_outputs(9995) <= not b or a;
    layer6_outputs(9996) <= not (a or b);
    layer6_outputs(9997) <= not (a xor b);
    layer6_outputs(9998) <= a xor b;
    layer6_outputs(9999) <= not b;
    layer6_outputs(10000) <= not a;
    layer6_outputs(10001) <= not (a xor b);
    layer6_outputs(10002) <= a and b;
    layer6_outputs(10003) <= not b;
    layer6_outputs(10004) <= not a;
    layer6_outputs(10005) <= a and not b;
    layer6_outputs(10006) <= a and b;
    layer6_outputs(10007) <= a xor b;
    layer6_outputs(10008) <= 1'b1;
    layer6_outputs(10009) <= not b;
    layer6_outputs(10010) <= a and b;
    layer6_outputs(10011) <= a and not b;
    layer6_outputs(10012) <= a and not b;
    layer6_outputs(10013) <= not a;
    layer6_outputs(10014) <= not (a and b);
    layer6_outputs(10015) <= not (a and b);
    layer6_outputs(10016) <= a and b;
    layer6_outputs(10017) <= a and not b;
    layer6_outputs(10018) <= b;
    layer6_outputs(10019) <= not b;
    layer6_outputs(10020) <= not (a and b);
    layer6_outputs(10021) <= 1'b1;
    layer6_outputs(10022) <= a;
    layer6_outputs(10023) <= not a;
    layer6_outputs(10024) <= a and not b;
    layer6_outputs(10025) <= a and b;
    layer6_outputs(10026) <= a;
    layer6_outputs(10027) <= b and not a;
    layer6_outputs(10028) <= not b;
    layer6_outputs(10029) <= not (a xor b);
    layer6_outputs(10030) <= b;
    layer6_outputs(10031) <= not b;
    layer6_outputs(10032) <= b and not a;
    layer6_outputs(10033) <= a or b;
    layer6_outputs(10034) <= not a;
    layer6_outputs(10035) <= not b;
    layer6_outputs(10036) <= not (a and b);
    layer6_outputs(10037) <= a and not b;
    layer6_outputs(10038) <= 1'b1;
    layer6_outputs(10039) <= a xor b;
    layer6_outputs(10040) <= a and not b;
    layer6_outputs(10041) <= not a or b;
    layer6_outputs(10042) <= not b;
    layer6_outputs(10043) <= b;
    layer6_outputs(10044) <= b and not a;
    layer6_outputs(10045) <= a;
    layer6_outputs(10046) <= not (a and b);
    layer6_outputs(10047) <= 1'b1;
    layer6_outputs(10048) <= not b or a;
    layer6_outputs(10049) <= not b;
    layer6_outputs(10050) <= not (a and b);
    layer6_outputs(10051) <= a;
    layer6_outputs(10052) <= b and not a;
    layer6_outputs(10053) <= a;
    layer6_outputs(10054) <= b;
    layer6_outputs(10055) <= not a;
    layer6_outputs(10056) <= a and not b;
    layer6_outputs(10057) <= not (a and b);
    layer6_outputs(10058) <= not a;
    layer6_outputs(10059) <= a or b;
    layer6_outputs(10060) <= not (a xor b);
    layer6_outputs(10061) <= not b;
    layer6_outputs(10062) <= not a or b;
    layer6_outputs(10063) <= not (a or b);
    layer6_outputs(10064) <= not (a xor b);
    layer6_outputs(10065) <= not (a and b);
    layer6_outputs(10066) <= not a;
    layer6_outputs(10067) <= not a or b;
    layer6_outputs(10068) <= a xor b;
    layer6_outputs(10069) <= a and not b;
    layer6_outputs(10070) <= a;
    layer6_outputs(10071) <= not b;
    layer6_outputs(10072) <= b;
    layer6_outputs(10073) <= not (a and b);
    layer6_outputs(10074) <= not a;
    layer6_outputs(10075) <= not (a xor b);
    layer6_outputs(10076) <= a or b;
    layer6_outputs(10077) <= not b or a;
    layer6_outputs(10078) <= a and not b;
    layer6_outputs(10079) <= not b;
    layer6_outputs(10080) <= not b;
    layer6_outputs(10081) <= not a;
    layer6_outputs(10082) <= a;
    layer6_outputs(10083) <= a xor b;
    layer6_outputs(10084) <= a or b;
    layer6_outputs(10085) <= b;
    layer6_outputs(10086) <= not a or b;
    layer6_outputs(10087) <= a and b;
    layer6_outputs(10088) <= 1'b1;
    layer6_outputs(10089) <= not (a xor b);
    layer6_outputs(10090) <= a or b;
    layer6_outputs(10091) <= not a or b;
    layer6_outputs(10092) <= a and not b;
    layer6_outputs(10093) <= b;
    layer6_outputs(10094) <= not (a or b);
    layer6_outputs(10095) <= not a;
    layer6_outputs(10096) <= not b or a;
    layer6_outputs(10097) <= not (a or b);
    layer6_outputs(10098) <= b;
    layer6_outputs(10099) <= b;
    layer6_outputs(10100) <= b and not a;
    layer6_outputs(10101) <= a;
    layer6_outputs(10102) <= a or b;
    layer6_outputs(10103) <= a and not b;
    layer6_outputs(10104) <= not a;
    layer6_outputs(10105) <= not a;
    layer6_outputs(10106) <= a;
    layer6_outputs(10107) <= not a or b;
    layer6_outputs(10108) <= not b;
    layer6_outputs(10109) <= a;
    layer6_outputs(10110) <= not (a or b);
    layer6_outputs(10111) <= not b;
    layer6_outputs(10112) <= b;
    layer6_outputs(10113) <= not b;
    layer6_outputs(10114) <= 1'b0;
    layer6_outputs(10115) <= not b or a;
    layer6_outputs(10116) <= not b or a;
    layer6_outputs(10117) <= a;
    layer6_outputs(10118) <= not (a xor b);
    layer6_outputs(10119) <= a and b;
    layer6_outputs(10120) <= not (a xor b);
    layer6_outputs(10121) <= a;
    layer6_outputs(10122) <= a and not b;
    layer6_outputs(10123) <= a;
    layer6_outputs(10124) <= a or b;
    layer6_outputs(10125) <= a and not b;
    layer6_outputs(10126) <= not b;
    layer6_outputs(10127) <= not (a xor b);
    layer6_outputs(10128) <= a and b;
    layer6_outputs(10129) <= a and not b;
    layer6_outputs(10130) <= b;
    layer6_outputs(10131) <= not a;
    layer6_outputs(10132) <= not a;
    layer6_outputs(10133) <= a;
    layer6_outputs(10134) <= a and not b;
    layer6_outputs(10135) <= a or b;
    layer6_outputs(10136) <= a or b;
    layer6_outputs(10137) <= not (a and b);
    layer6_outputs(10138) <= 1'b1;
    layer6_outputs(10139) <= b;
    layer6_outputs(10140) <= not b or a;
    layer6_outputs(10141) <= not b;
    layer6_outputs(10142) <= b and not a;
    layer6_outputs(10143) <= b;
    layer6_outputs(10144) <= b and not a;
    layer6_outputs(10145) <= 1'b0;
    layer6_outputs(10146) <= a;
    layer6_outputs(10147) <= a and b;
    layer6_outputs(10148) <= not a;
    layer6_outputs(10149) <= b;
    layer6_outputs(10150) <= not (a and b);
    layer6_outputs(10151) <= a;
    layer6_outputs(10152) <= a xor b;
    layer6_outputs(10153) <= not (a xor b);
    layer6_outputs(10154) <= not b;
    layer6_outputs(10155) <= not (a and b);
    layer6_outputs(10156) <= b and not a;
    layer6_outputs(10157) <= not (a and b);
    layer6_outputs(10158) <= not (a and b);
    layer6_outputs(10159) <= not (a and b);
    layer6_outputs(10160) <= a and b;
    layer6_outputs(10161) <= not a or b;
    layer6_outputs(10162) <= not a;
    layer6_outputs(10163) <= a xor b;
    layer6_outputs(10164) <= a and not b;
    layer6_outputs(10165) <= a xor b;
    layer6_outputs(10166) <= a;
    layer6_outputs(10167) <= not a;
    layer6_outputs(10168) <= not b or a;
    layer6_outputs(10169) <= not b;
    layer6_outputs(10170) <= b;
    layer6_outputs(10171) <= a;
    layer6_outputs(10172) <= not b;
    layer6_outputs(10173) <= not (a and b);
    layer6_outputs(10174) <= a;
    layer6_outputs(10175) <= a;
    layer6_outputs(10176) <= 1'b0;
    layer6_outputs(10177) <= a;
    layer6_outputs(10178) <= not a;
    layer6_outputs(10179) <= a;
    layer6_outputs(10180) <= a;
    layer6_outputs(10181) <= a or b;
    layer6_outputs(10182) <= 1'b1;
    layer6_outputs(10183) <= not b or a;
    layer6_outputs(10184) <= not a or b;
    layer6_outputs(10185) <= a xor b;
    layer6_outputs(10186) <= a xor b;
    layer6_outputs(10187) <= not a or b;
    layer6_outputs(10188) <= a or b;
    layer6_outputs(10189) <= a xor b;
    layer6_outputs(10190) <= a;
    layer6_outputs(10191) <= b;
    layer6_outputs(10192) <= a and b;
    layer6_outputs(10193) <= a and not b;
    layer6_outputs(10194) <= b and not a;
    layer6_outputs(10195) <= not b or a;
    layer6_outputs(10196) <= b;
    layer6_outputs(10197) <= a and not b;
    layer6_outputs(10198) <= not (a and b);
    layer6_outputs(10199) <= not (a and b);
    layer6_outputs(10200) <= a and not b;
    layer6_outputs(10201) <= a and b;
    layer6_outputs(10202) <= not a;
    layer6_outputs(10203) <= not b;
    layer6_outputs(10204) <= not a;
    layer6_outputs(10205) <= not a;
    layer6_outputs(10206) <= a;
    layer6_outputs(10207) <= a xor b;
    layer6_outputs(10208) <= a or b;
    layer6_outputs(10209) <= not (a and b);
    layer6_outputs(10210) <= 1'b1;
    layer6_outputs(10211) <= a;
    layer6_outputs(10212) <= a;
    layer6_outputs(10213) <= a and not b;
    layer6_outputs(10214) <= b;
    layer6_outputs(10215) <= not b;
    layer6_outputs(10216) <= a and not b;
    layer6_outputs(10217) <= not a;
    layer6_outputs(10218) <= not a;
    layer6_outputs(10219) <= not (a and b);
    layer6_outputs(10220) <= b;
    layer6_outputs(10221) <= a;
    layer6_outputs(10222) <= a or b;
    layer6_outputs(10223) <= 1'b0;
    layer6_outputs(10224) <= not a;
    layer6_outputs(10225) <= not a;
    layer6_outputs(10226) <= not a;
    layer6_outputs(10227) <= b;
    layer6_outputs(10228) <= not b or a;
    layer6_outputs(10229) <= not b;
    layer6_outputs(10230) <= b;
    layer6_outputs(10231) <= not b;
    layer6_outputs(10232) <= a and b;
    layer6_outputs(10233) <= not b or a;
    layer6_outputs(10234) <= a;
    layer6_outputs(10235) <= a and b;
    layer6_outputs(10236) <= not a;
    layer6_outputs(10237) <= not b;
    layer6_outputs(10238) <= b;
    layer6_outputs(10239) <= not (a xor b);
    layer7_outputs(0) <= not b or a;
    layer7_outputs(1) <= a;
    layer7_outputs(2) <= a;
    layer7_outputs(3) <= not a or b;
    layer7_outputs(4) <= a and not b;
    layer7_outputs(5) <= a and b;
    layer7_outputs(6) <= not a or b;
    layer7_outputs(7) <= b and not a;
    layer7_outputs(8) <= not a;
    layer7_outputs(9) <= a and b;
    layer7_outputs(10) <= 1'b0;
    layer7_outputs(11) <= b and not a;
    layer7_outputs(12) <= a xor b;
    layer7_outputs(13) <= not a or b;
    layer7_outputs(14) <= not (a xor b);
    layer7_outputs(15) <= a;
    layer7_outputs(16) <= a;
    layer7_outputs(17) <= not b;
    layer7_outputs(18) <= a and not b;
    layer7_outputs(19) <= not b or a;
    layer7_outputs(20) <= a;
    layer7_outputs(21) <= 1'b1;
    layer7_outputs(22) <= not (a and b);
    layer7_outputs(23) <= not a;
    layer7_outputs(24) <= not a or b;
    layer7_outputs(25) <= not b;
    layer7_outputs(26) <= b;
    layer7_outputs(27) <= not (a or b);
    layer7_outputs(28) <= 1'b1;
    layer7_outputs(29) <= not a;
    layer7_outputs(30) <= not b;
    layer7_outputs(31) <= b and not a;
    layer7_outputs(32) <= not b or a;
    layer7_outputs(33) <= not (a and b);
    layer7_outputs(34) <= not (a xor b);
    layer7_outputs(35) <= not (a xor b);
    layer7_outputs(36) <= a xor b;
    layer7_outputs(37) <= a xor b;
    layer7_outputs(38) <= not (a xor b);
    layer7_outputs(39) <= a and not b;
    layer7_outputs(40) <= not (a xor b);
    layer7_outputs(41) <= a and not b;
    layer7_outputs(42) <= not b;
    layer7_outputs(43) <= not (a or b);
    layer7_outputs(44) <= not a;
    layer7_outputs(45) <= not a;
    layer7_outputs(46) <= a or b;
    layer7_outputs(47) <= not b;
    layer7_outputs(48) <= a;
    layer7_outputs(49) <= not b;
    layer7_outputs(50) <= not b;
    layer7_outputs(51) <= a and b;
    layer7_outputs(52) <= b and not a;
    layer7_outputs(53) <= b;
    layer7_outputs(54) <= not a;
    layer7_outputs(55) <= b and not a;
    layer7_outputs(56) <= not a;
    layer7_outputs(57) <= a and b;
    layer7_outputs(58) <= not a or b;
    layer7_outputs(59) <= a and not b;
    layer7_outputs(60) <= b and not a;
    layer7_outputs(61) <= not (a xor b);
    layer7_outputs(62) <= not b or a;
    layer7_outputs(63) <= not a;
    layer7_outputs(64) <= not a or b;
    layer7_outputs(65) <= a and b;
    layer7_outputs(66) <= not (a and b);
    layer7_outputs(67) <= not b or a;
    layer7_outputs(68) <= not (a xor b);
    layer7_outputs(69) <= b and not a;
    layer7_outputs(70) <= a and not b;
    layer7_outputs(71) <= a;
    layer7_outputs(72) <= a xor b;
    layer7_outputs(73) <= a;
    layer7_outputs(74) <= a;
    layer7_outputs(75) <= a;
    layer7_outputs(76) <= not (a xor b);
    layer7_outputs(77) <= a;
    layer7_outputs(78) <= not a;
    layer7_outputs(79) <= not b;
    layer7_outputs(80) <= b;
    layer7_outputs(81) <= not b;
    layer7_outputs(82) <= a xor b;
    layer7_outputs(83) <= a and not b;
    layer7_outputs(84) <= b;
    layer7_outputs(85) <= b;
    layer7_outputs(86) <= not b;
    layer7_outputs(87) <= a xor b;
    layer7_outputs(88) <= not (a and b);
    layer7_outputs(89) <= not (a or b);
    layer7_outputs(90) <= a and not b;
    layer7_outputs(91) <= not b;
    layer7_outputs(92) <= a;
    layer7_outputs(93) <= not (a and b);
    layer7_outputs(94) <= not a;
    layer7_outputs(95) <= not b;
    layer7_outputs(96) <= a and not b;
    layer7_outputs(97) <= not a;
    layer7_outputs(98) <= b and not a;
    layer7_outputs(99) <= a xor b;
    layer7_outputs(100) <= a or b;
    layer7_outputs(101) <= not a;
    layer7_outputs(102) <= b and not a;
    layer7_outputs(103) <= b;
    layer7_outputs(104) <= a;
    layer7_outputs(105) <= b;
    layer7_outputs(106) <= not b;
    layer7_outputs(107) <= b and not a;
    layer7_outputs(108) <= not a;
    layer7_outputs(109) <= b;
    layer7_outputs(110) <= b;
    layer7_outputs(111) <= not (a xor b);
    layer7_outputs(112) <= a;
    layer7_outputs(113) <= a xor b;
    layer7_outputs(114) <= not a or b;
    layer7_outputs(115) <= a or b;
    layer7_outputs(116) <= b and not a;
    layer7_outputs(117) <= not b or a;
    layer7_outputs(118) <= a;
    layer7_outputs(119) <= not (a or b);
    layer7_outputs(120) <= b and not a;
    layer7_outputs(121) <= a;
    layer7_outputs(122) <= not b;
    layer7_outputs(123) <= not a;
    layer7_outputs(124) <= not (a xor b);
    layer7_outputs(125) <= a xor b;
    layer7_outputs(126) <= b and not a;
    layer7_outputs(127) <= not b;
    layer7_outputs(128) <= not (a or b);
    layer7_outputs(129) <= not a;
    layer7_outputs(130) <= a xor b;
    layer7_outputs(131) <= a and not b;
    layer7_outputs(132) <= a and not b;
    layer7_outputs(133) <= b;
    layer7_outputs(134) <= a;
    layer7_outputs(135) <= not a;
    layer7_outputs(136) <= not b or a;
    layer7_outputs(137) <= a xor b;
    layer7_outputs(138) <= not (a xor b);
    layer7_outputs(139) <= not (a xor b);
    layer7_outputs(140) <= not (a xor b);
    layer7_outputs(141) <= a and b;
    layer7_outputs(142) <= a and b;
    layer7_outputs(143) <= not (a and b);
    layer7_outputs(144) <= not a;
    layer7_outputs(145) <= not b;
    layer7_outputs(146) <= not (a xor b);
    layer7_outputs(147) <= a;
    layer7_outputs(148) <= not (a and b);
    layer7_outputs(149) <= not (a xor b);
    layer7_outputs(150) <= a and b;
    layer7_outputs(151) <= not b;
    layer7_outputs(152) <= a and not b;
    layer7_outputs(153) <= a and b;
    layer7_outputs(154) <= b;
    layer7_outputs(155) <= a and b;
    layer7_outputs(156) <= a or b;
    layer7_outputs(157) <= not b;
    layer7_outputs(158) <= not (a xor b);
    layer7_outputs(159) <= not a;
    layer7_outputs(160) <= a;
    layer7_outputs(161) <= not (a or b);
    layer7_outputs(162) <= not a;
    layer7_outputs(163) <= not (a xor b);
    layer7_outputs(164) <= a;
    layer7_outputs(165) <= not a or b;
    layer7_outputs(166) <= a or b;
    layer7_outputs(167) <= not (a or b);
    layer7_outputs(168) <= not a;
    layer7_outputs(169) <= a;
    layer7_outputs(170) <= a xor b;
    layer7_outputs(171) <= a and b;
    layer7_outputs(172) <= not a;
    layer7_outputs(173) <= not (a or b);
    layer7_outputs(174) <= a xor b;
    layer7_outputs(175) <= a xor b;
    layer7_outputs(176) <= not a or b;
    layer7_outputs(177) <= a xor b;
    layer7_outputs(178) <= not (a xor b);
    layer7_outputs(179) <= not b;
    layer7_outputs(180) <= not (a xor b);
    layer7_outputs(181) <= not b;
    layer7_outputs(182) <= a xor b;
    layer7_outputs(183) <= not (a xor b);
    layer7_outputs(184) <= a and b;
    layer7_outputs(185) <= a;
    layer7_outputs(186) <= a xor b;
    layer7_outputs(187) <= a xor b;
    layer7_outputs(188) <= b and not a;
    layer7_outputs(189) <= not a;
    layer7_outputs(190) <= not (a and b);
    layer7_outputs(191) <= not (a or b);
    layer7_outputs(192) <= not (a or b);
    layer7_outputs(193) <= a;
    layer7_outputs(194) <= b;
    layer7_outputs(195) <= not (a and b);
    layer7_outputs(196) <= not b or a;
    layer7_outputs(197) <= a;
    layer7_outputs(198) <= not a;
    layer7_outputs(199) <= not a;
    layer7_outputs(200) <= not a;
    layer7_outputs(201) <= not b;
    layer7_outputs(202) <= not a;
    layer7_outputs(203) <= not a;
    layer7_outputs(204) <= a or b;
    layer7_outputs(205) <= a and b;
    layer7_outputs(206) <= not (a xor b);
    layer7_outputs(207) <= a;
    layer7_outputs(208) <= not (a and b);
    layer7_outputs(209) <= not (a and b);
    layer7_outputs(210) <= not b or a;
    layer7_outputs(211) <= not (a and b);
    layer7_outputs(212) <= a or b;
    layer7_outputs(213) <= a;
    layer7_outputs(214) <= a;
    layer7_outputs(215) <= not (a and b);
    layer7_outputs(216) <= not (a or b);
    layer7_outputs(217) <= not b;
    layer7_outputs(218) <= a and not b;
    layer7_outputs(219) <= a and not b;
    layer7_outputs(220) <= a xor b;
    layer7_outputs(221) <= b;
    layer7_outputs(222) <= b;
    layer7_outputs(223) <= a xor b;
    layer7_outputs(224) <= a xor b;
    layer7_outputs(225) <= not a;
    layer7_outputs(226) <= not (a or b);
    layer7_outputs(227) <= a and not b;
    layer7_outputs(228) <= not (a or b);
    layer7_outputs(229) <= not b;
    layer7_outputs(230) <= b and not a;
    layer7_outputs(231) <= b and not a;
    layer7_outputs(232) <= a xor b;
    layer7_outputs(233) <= a;
    layer7_outputs(234) <= b and not a;
    layer7_outputs(235) <= not a;
    layer7_outputs(236) <= not (a or b);
    layer7_outputs(237) <= not b or a;
    layer7_outputs(238) <= a xor b;
    layer7_outputs(239) <= a xor b;
    layer7_outputs(240) <= b and not a;
    layer7_outputs(241) <= not b;
    layer7_outputs(242) <= a and not b;
    layer7_outputs(243) <= not (a xor b);
    layer7_outputs(244) <= a or b;
    layer7_outputs(245) <= not (a and b);
    layer7_outputs(246) <= not b or a;
    layer7_outputs(247) <= 1'b0;
    layer7_outputs(248) <= not b or a;
    layer7_outputs(249) <= b and not a;
    layer7_outputs(250) <= not a;
    layer7_outputs(251) <= a;
    layer7_outputs(252) <= not a;
    layer7_outputs(253) <= a and not b;
    layer7_outputs(254) <= b and not a;
    layer7_outputs(255) <= not a;
    layer7_outputs(256) <= 1'b1;
    layer7_outputs(257) <= not a;
    layer7_outputs(258) <= b;
    layer7_outputs(259) <= a and not b;
    layer7_outputs(260) <= b;
    layer7_outputs(261) <= a;
    layer7_outputs(262) <= not b;
    layer7_outputs(263) <= not a or b;
    layer7_outputs(264) <= b;
    layer7_outputs(265) <= not b;
    layer7_outputs(266) <= a and b;
    layer7_outputs(267) <= not a;
    layer7_outputs(268) <= a xor b;
    layer7_outputs(269) <= a and not b;
    layer7_outputs(270) <= not (a or b);
    layer7_outputs(271) <= a or b;
    layer7_outputs(272) <= not b;
    layer7_outputs(273) <= not a;
    layer7_outputs(274) <= not a;
    layer7_outputs(275) <= not b;
    layer7_outputs(276) <= a xor b;
    layer7_outputs(277) <= 1'b0;
    layer7_outputs(278) <= a xor b;
    layer7_outputs(279) <= a and not b;
    layer7_outputs(280) <= a;
    layer7_outputs(281) <= not a or b;
    layer7_outputs(282) <= a xor b;
    layer7_outputs(283) <= not (a xor b);
    layer7_outputs(284) <= a xor b;
    layer7_outputs(285) <= b and not a;
    layer7_outputs(286) <= not (a xor b);
    layer7_outputs(287) <= not (a or b);
    layer7_outputs(288) <= b and not a;
    layer7_outputs(289) <= b;
    layer7_outputs(290) <= b;
    layer7_outputs(291) <= a and b;
    layer7_outputs(292) <= a and b;
    layer7_outputs(293) <= not (a and b);
    layer7_outputs(294) <= a or b;
    layer7_outputs(295) <= a;
    layer7_outputs(296) <= not a;
    layer7_outputs(297) <= a and b;
    layer7_outputs(298) <= a;
    layer7_outputs(299) <= b and not a;
    layer7_outputs(300) <= a xor b;
    layer7_outputs(301) <= a;
    layer7_outputs(302) <= not (a or b);
    layer7_outputs(303) <= not (a and b);
    layer7_outputs(304) <= b;
    layer7_outputs(305) <= not a;
    layer7_outputs(306) <= a xor b;
    layer7_outputs(307) <= not (a or b);
    layer7_outputs(308) <= b;
    layer7_outputs(309) <= a and b;
    layer7_outputs(310) <= a and b;
    layer7_outputs(311) <= not a;
    layer7_outputs(312) <= a or b;
    layer7_outputs(313) <= a xor b;
    layer7_outputs(314) <= not a or b;
    layer7_outputs(315) <= not a;
    layer7_outputs(316) <= a xor b;
    layer7_outputs(317) <= b;
    layer7_outputs(318) <= not a;
    layer7_outputs(319) <= not b;
    layer7_outputs(320) <= not a;
    layer7_outputs(321) <= not (a and b);
    layer7_outputs(322) <= a;
    layer7_outputs(323) <= b and not a;
    layer7_outputs(324) <= b and not a;
    layer7_outputs(325) <= not b;
    layer7_outputs(326) <= not b;
    layer7_outputs(327) <= not a;
    layer7_outputs(328) <= not (a xor b);
    layer7_outputs(329) <= not a or b;
    layer7_outputs(330) <= a;
    layer7_outputs(331) <= b;
    layer7_outputs(332) <= not a;
    layer7_outputs(333) <= a;
    layer7_outputs(334) <= a;
    layer7_outputs(335) <= a xor b;
    layer7_outputs(336) <= a;
    layer7_outputs(337) <= a and not b;
    layer7_outputs(338) <= a;
    layer7_outputs(339) <= not a;
    layer7_outputs(340) <= not (a and b);
    layer7_outputs(341) <= b and not a;
    layer7_outputs(342) <= not (a xor b);
    layer7_outputs(343) <= not a;
    layer7_outputs(344) <= not (a and b);
    layer7_outputs(345) <= not a;
    layer7_outputs(346) <= not b or a;
    layer7_outputs(347) <= not (a xor b);
    layer7_outputs(348) <= a;
    layer7_outputs(349) <= not (a and b);
    layer7_outputs(350) <= not (a or b);
    layer7_outputs(351) <= a and not b;
    layer7_outputs(352) <= not (a xor b);
    layer7_outputs(353) <= not a;
    layer7_outputs(354) <= a xor b;
    layer7_outputs(355) <= a xor b;
    layer7_outputs(356) <= a and b;
    layer7_outputs(357) <= not b;
    layer7_outputs(358) <= b;
    layer7_outputs(359) <= not (a and b);
    layer7_outputs(360) <= not b;
    layer7_outputs(361) <= not b;
    layer7_outputs(362) <= a and not b;
    layer7_outputs(363) <= not a;
    layer7_outputs(364) <= not (a or b);
    layer7_outputs(365) <= not b;
    layer7_outputs(366) <= not (a xor b);
    layer7_outputs(367) <= not (a xor b);
    layer7_outputs(368) <= not a;
    layer7_outputs(369) <= not (a xor b);
    layer7_outputs(370) <= a and b;
    layer7_outputs(371) <= b;
    layer7_outputs(372) <= not a or b;
    layer7_outputs(373) <= not b;
    layer7_outputs(374) <= a;
    layer7_outputs(375) <= not (a xor b);
    layer7_outputs(376) <= not a;
    layer7_outputs(377) <= not a;
    layer7_outputs(378) <= a;
    layer7_outputs(379) <= not a;
    layer7_outputs(380) <= not (a or b);
    layer7_outputs(381) <= not a;
    layer7_outputs(382) <= b and not a;
    layer7_outputs(383) <= not a;
    layer7_outputs(384) <= not a;
    layer7_outputs(385) <= not b;
    layer7_outputs(386) <= not b;
    layer7_outputs(387) <= b;
    layer7_outputs(388) <= not b;
    layer7_outputs(389) <= a and not b;
    layer7_outputs(390) <= a xor b;
    layer7_outputs(391) <= not a;
    layer7_outputs(392) <= b and not a;
    layer7_outputs(393) <= not b;
    layer7_outputs(394) <= not (a xor b);
    layer7_outputs(395) <= a or b;
    layer7_outputs(396) <= b;
    layer7_outputs(397) <= a or b;
    layer7_outputs(398) <= not a or b;
    layer7_outputs(399) <= b;
    layer7_outputs(400) <= b;
    layer7_outputs(401) <= not a;
    layer7_outputs(402) <= b and not a;
    layer7_outputs(403) <= not b;
    layer7_outputs(404) <= not b;
    layer7_outputs(405) <= not (a or b);
    layer7_outputs(406) <= b and not a;
    layer7_outputs(407) <= not b or a;
    layer7_outputs(408) <= a xor b;
    layer7_outputs(409) <= b and not a;
    layer7_outputs(410) <= a and b;
    layer7_outputs(411) <= not (a xor b);
    layer7_outputs(412) <= not b;
    layer7_outputs(413) <= not b or a;
    layer7_outputs(414) <= not a;
    layer7_outputs(415) <= a and b;
    layer7_outputs(416) <= a and b;
    layer7_outputs(417) <= not b or a;
    layer7_outputs(418) <= a and b;
    layer7_outputs(419) <= a and b;
    layer7_outputs(420) <= not b or a;
    layer7_outputs(421) <= not a or b;
    layer7_outputs(422) <= not a;
    layer7_outputs(423) <= not a;
    layer7_outputs(424) <= not b;
    layer7_outputs(425) <= a xor b;
    layer7_outputs(426) <= not b;
    layer7_outputs(427) <= not a;
    layer7_outputs(428) <= not a or b;
    layer7_outputs(429) <= a and b;
    layer7_outputs(430) <= not (a xor b);
    layer7_outputs(431) <= b and not a;
    layer7_outputs(432) <= a xor b;
    layer7_outputs(433) <= a;
    layer7_outputs(434) <= b and not a;
    layer7_outputs(435) <= not a;
    layer7_outputs(436) <= not b or a;
    layer7_outputs(437) <= not (a xor b);
    layer7_outputs(438) <= not a or b;
    layer7_outputs(439) <= a and b;
    layer7_outputs(440) <= a;
    layer7_outputs(441) <= not (a or b);
    layer7_outputs(442) <= a xor b;
    layer7_outputs(443) <= a;
    layer7_outputs(444) <= a and b;
    layer7_outputs(445) <= a and b;
    layer7_outputs(446) <= not b;
    layer7_outputs(447) <= not a;
    layer7_outputs(448) <= a and b;
    layer7_outputs(449) <= a;
    layer7_outputs(450) <= not (a or b);
    layer7_outputs(451) <= not (a xor b);
    layer7_outputs(452) <= b and not a;
    layer7_outputs(453) <= a and not b;
    layer7_outputs(454) <= a xor b;
    layer7_outputs(455) <= b and not a;
    layer7_outputs(456) <= not a;
    layer7_outputs(457) <= a or b;
    layer7_outputs(458) <= 1'b1;
    layer7_outputs(459) <= b;
    layer7_outputs(460) <= a;
    layer7_outputs(461) <= a xor b;
    layer7_outputs(462) <= a;
    layer7_outputs(463) <= a;
    layer7_outputs(464) <= b;
    layer7_outputs(465) <= a;
    layer7_outputs(466) <= a and not b;
    layer7_outputs(467) <= a and not b;
    layer7_outputs(468) <= a and not b;
    layer7_outputs(469) <= not a;
    layer7_outputs(470) <= a or b;
    layer7_outputs(471) <= a or b;
    layer7_outputs(472) <= b;
    layer7_outputs(473) <= b;
    layer7_outputs(474) <= not b;
    layer7_outputs(475) <= a or b;
    layer7_outputs(476) <= not a;
    layer7_outputs(477) <= b;
    layer7_outputs(478) <= not (a xor b);
    layer7_outputs(479) <= not (a xor b);
    layer7_outputs(480) <= not b;
    layer7_outputs(481) <= not a or b;
    layer7_outputs(482) <= not a;
    layer7_outputs(483) <= a and b;
    layer7_outputs(484) <= a xor b;
    layer7_outputs(485) <= a xor b;
    layer7_outputs(486) <= a and not b;
    layer7_outputs(487) <= a;
    layer7_outputs(488) <= not a or b;
    layer7_outputs(489) <= not b;
    layer7_outputs(490) <= a;
    layer7_outputs(491) <= a;
    layer7_outputs(492) <= not b;
    layer7_outputs(493) <= not a;
    layer7_outputs(494) <= b;
    layer7_outputs(495) <= not b;
    layer7_outputs(496) <= not a;
    layer7_outputs(497) <= not a;
    layer7_outputs(498) <= a;
    layer7_outputs(499) <= not (a and b);
    layer7_outputs(500) <= not a;
    layer7_outputs(501) <= not (a xor b);
    layer7_outputs(502) <= b and not a;
    layer7_outputs(503) <= not b;
    layer7_outputs(504) <= not b or a;
    layer7_outputs(505) <= not (a and b);
    layer7_outputs(506) <= b and not a;
    layer7_outputs(507) <= not (a xor b);
    layer7_outputs(508) <= a and b;
    layer7_outputs(509) <= b;
    layer7_outputs(510) <= b;
    layer7_outputs(511) <= a and b;
    layer7_outputs(512) <= not (a xor b);
    layer7_outputs(513) <= not b;
    layer7_outputs(514) <= a xor b;
    layer7_outputs(515) <= not b;
    layer7_outputs(516) <= b;
    layer7_outputs(517) <= a;
    layer7_outputs(518) <= a xor b;
    layer7_outputs(519) <= not a;
    layer7_outputs(520) <= a xor b;
    layer7_outputs(521) <= a;
    layer7_outputs(522) <= a or b;
    layer7_outputs(523) <= not b;
    layer7_outputs(524) <= b;
    layer7_outputs(525) <= not (a or b);
    layer7_outputs(526) <= not a;
    layer7_outputs(527) <= not b;
    layer7_outputs(528) <= not a or b;
    layer7_outputs(529) <= a or b;
    layer7_outputs(530) <= a xor b;
    layer7_outputs(531) <= b;
    layer7_outputs(532) <= not a or b;
    layer7_outputs(533) <= a;
    layer7_outputs(534) <= not (a or b);
    layer7_outputs(535) <= not a;
    layer7_outputs(536) <= not b or a;
    layer7_outputs(537) <= not a;
    layer7_outputs(538) <= b;
    layer7_outputs(539) <= b;
    layer7_outputs(540) <= a and not b;
    layer7_outputs(541) <= a xor b;
    layer7_outputs(542) <= not a;
    layer7_outputs(543) <= a xor b;
    layer7_outputs(544) <= not a;
    layer7_outputs(545) <= not b or a;
    layer7_outputs(546) <= not b;
    layer7_outputs(547) <= b and not a;
    layer7_outputs(548) <= a and not b;
    layer7_outputs(549) <= not a or b;
    layer7_outputs(550) <= not (a and b);
    layer7_outputs(551) <= a;
    layer7_outputs(552) <= not b or a;
    layer7_outputs(553) <= a;
    layer7_outputs(554) <= a or b;
    layer7_outputs(555) <= b;
    layer7_outputs(556) <= a and b;
    layer7_outputs(557) <= not b;
    layer7_outputs(558) <= b;
    layer7_outputs(559) <= a xor b;
    layer7_outputs(560) <= not (a xor b);
    layer7_outputs(561) <= not (a xor b);
    layer7_outputs(562) <= b and not a;
    layer7_outputs(563) <= b;
    layer7_outputs(564) <= not (a xor b);
    layer7_outputs(565) <= a and not b;
    layer7_outputs(566) <= not a;
    layer7_outputs(567) <= a xor b;
    layer7_outputs(568) <= not a;
    layer7_outputs(569) <= not a;
    layer7_outputs(570) <= a and b;
    layer7_outputs(571) <= a xor b;
    layer7_outputs(572) <= not a;
    layer7_outputs(573) <= not (a xor b);
    layer7_outputs(574) <= not b;
    layer7_outputs(575) <= a and not b;
    layer7_outputs(576) <= a;
    layer7_outputs(577) <= not a;
    layer7_outputs(578) <= a;
    layer7_outputs(579) <= a or b;
    layer7_outputs(580) <= b;
    layer7_outputs(581) <= not a;
    layer7_outputs(582) <= not (a xor b);
    layer7_outputs(583) <= not b;
    layer7_outputs(584) <= b and not a;
    layer7_outputs(585) <= a and not b;
    layer7_outputs(586) <= not (a xor b);
    layer7_outputs(587) <= not b or a;
    layer7_outputs(588) <= not a;
    layer7_outputs(589) <= not a;
    layer7_outputs(590) <= not a or b;
    layer7_outputs(591) <= not b or a;
    layer7_outputs(592) <= not b;
    layer7_outputs(593) <= not b or a;
    layer7_outputs(594) <= not (a or b);
    layer7_outputs(595) <= b and not a;
    layer7_outputs(596) <= not (a and b);
    layer7_outputs(597) <= not (a and b);
    layer7_outputs(598) <= a and b;
    layer7_outputs(599) <= not b or a;
    layer7_outputs(600) <= not b;
    layer7_outputs(601) <= not a;
    layer7_outputs(602) <= a xor b;
    layer7_outputs(603) <= a and b;
    layer7_outputs(604) <= not b;
    layer7_outputs(605) <= not (a and b);
    layer7_outputs(606) <= not a;
    layer7_outputs(607) <= b;
    layer7_outputs(608) <= a xor b;
    layer7_outputs(609) <= not (a or b);
    layer7_outputs(610) <= not a;
    layer7_outputs(611) <= a xor b;
    layer7_outputs(612) <= not a;
    layer7_outputs(613) <= a;
    layer7_outputs(614) <= not (a xor b);
    layer7_outputs(615) <= not a;
    layer7_outputs(616) <= not (a and b);
    layer7_outputs(617) <= b;
    layer7_outputs(618) <= not (a or b);
    layer7_outputs(619) <= not (a or b);
    layer7_outputs(620) <= not a or b;
    layer7_outputs(621) <= not b;
    layer7_outputs(622) <= a;
    layer7_outputs(623) <= not a;
    layer7_outputs(624) <= b;
    layer7_outputs(625) <= not b or a;
    layer7_outputs(626) <= a;
    layer7_outputs(627) <= b;
    layer7_outputs(628) <= not a;
    layer7_outputs(629) <= a;
    layer7_outputs(630) <= not b;
    layer7_outputs(631) <= not (a xor b);
    layer7_outputs(632) <= not b;
    layer7_outputs(633) <= not a;
    layer7_outputs(634) <= b and not a;
    layer7_outputs(635) <= 1'b0;
    layer7_outputs(636) <= a or b;
    layer7_outputs(637) <= not b or a;
    layer7_outputs(638) <= 1'b0;
    layer7_outputs(639) <= a;
    layer7_outputs(640) <= a or b;
    layer7_outputs(641) <= a xor b;
    layer7_outputs(642) <= 1'b1;
    layer7_outputs(643) <= not (a and b);
    layer7_outputs(644) <= a;
    layer7_outputs(645) <= a and not b;
    layer7_outputs(646) <= 1'b0;
    layer7_outputs(647) <= not a;
    layer7_outputs(648) <= a and b;
    layer7_outputs(649) <= b;
    layer7_outputs(650) <= b;
    layer7_outputs(651) <= b and not a;
    layer7_outputs(652) <= b;
    layer7_outputs(653) <= not (a xor b);
    layer7_outputs(654) <= not a or b;
    layer7_outputs(655) <= a xor b;
    layer7_outputs(656) <= not a;
    layer7_outputs(657) <= not (a or b);
    layer7_outputs(658) <= a xor b;
    layer7_outputs(659) <= not (a xor b);
    layer7_outputs(660) <= not (a and b);
    layer7_outputs(661) <= b;
    layer7_outputs(662) <= not (a and b);
    layer7_outputs(663) <= a or b;
    layer7_outputs(664) <= b and not a;
    layer7_outputs(665) <= a xor b;
    layer7_outputs(666) <= a or b;
    layer7_outputs(667) <= a xor b;
    layer7_outputs(668) <= a or b;
    layer7_outputs(669) <= a xor b;
    layer7_outputs(670) <= a and not b;
    layer7_outputs(671) <= a xor b;
    layer7_outputs(672) <= not b or a;
    layer7_outputs(673) <= a and not b;
    layer7_outputs(674) <= b;
    layer7_outputs(675) <= not a;
    layer7_outputs(676) <= not (a or b);
    layer7_outputs(677) <= not a or b;
    layer7_outputs(678) <= a or b;
    layer7_outputs(679) <= a and b;
    layer7_outputs(680) <= not (a or b);
    layer7_outputs(681) <= not (a xor b);
    layer7_outputs(682) <= not a;
    layer7_outputs(683) <= b;
    layer7_outputs(684) <= not (a and b);
    layer7_outputs(685) <= a and b;
    layer7_outputs(686) <= not b or a;
    layer7_outputs(687) <= a and b;
    layer7_outputs(688) <= a and b;
    layer7_outputs(689) <= a and b;
    layer7_outputs(690) <= a and b;
    layer7_outputs(691) <= not a;
    layer7_outputs(692) <= not b or a;
    layer7_outputs(693) <= not (a or b);
    layer7_outputs(694) <= not a;
    layer7_outputs(695) <= b;
    layer7_outputs(696) <= not a;
    layer7_outputs(697) <= b;
    layer7_outputs(698) <= a or b;
    layer7_outputs(699) <= a xor b;
    layer7_outputs(700) <= not a;
    layer7_outputs(701) <= not (a xor b);
    layer7_outputs(702) <= not (a or b);
    layer7_outputs(703) <= not b;
    layer7_outputs(704) <= a xor b;
    layer7_outputs(705) <= not a;
    layer7_outputs(706) <= a and b;
    layer7_outputs(707) <= a and not b;
    layer7_outputs(708) <= a;
    layer7_outputs(709) <= not b;
    layer7_outputs(710) <= b and not a;
    layer7_outputs(711) <= not a;
    layer7_outputs(712) <= not b;
    layer7_outputs(713) <= a xor b;
    layer7_outputs(714) <= not (a or b);
    layer7_outputs(715) <= not a;
    layer7_outputs(716) <= b and not a;
    layer7_outputs(717) <= a or b;
    layer7_outputs(718) <= a;
    layer7_outputs(719) <= not b;
    layer7_outputs(720) <= not (a xor b);
    layer7_outputs(721) <= not (a and b);
    layer7_outputs(722) <= b;
    layer7_outputs(723) <= not b or a;
    layer7_outputs(724) <= a and not b;
    layer7_outputs(725) <= not b;
    layer7_outputs(726) <= not b;
    layer7_outputs(727) <= a and not b;
    layer7_outputs(728) <= a or b;
    layer7_outputs(729) <= a xor b;
    layer7_outputs(730) <= not a or b;
    layer7_outputs(731) <= not (a and b);
    layer7_outputs(732) <= a and not b;
    layer7_outputs(733) <= a;
    layer7_outputs(734) <= not (a xor b);
    layer7_outputs(735) <= a;
    layer7_outputs(736) <= not (a xor b);
    layer7_outputs(737) <= a and b;
    layer7_outputs(738) <= b and not a;
    layer7_outputs(739) <= not (a xor b);
    layer7_outputs(740) <= not (a and b);
    layer7_outputs(741) <= not (a xor b);
    layer7_outputs(742) <= b;
    layer7_outputs(743) <= not a;
    layer7_outputs(744) <= a or b;
    layer7_outputs(745) <= a xor b;
    layer7_outputs(746) <= not (a or b);
    layer7_outputs(747) <= not b or a;
    layer7_outputs(748) <= a;
    layer7_outputs(749) <= a or b;
    layer7_outputs(750) <= a xor b;
    layer7_outputs(751) <= not b or a;
    layer7_outputs(752) <= a;
    layer7_outputs(753) <= a;
    layer7_outputs(754) <= not b;
    layer7_outputs(755) <= not (a or b);
    layer7_outputs(756) <= not a;
    layer7_outputs(757) <= a and b;
    layer7_outputs(758) <= a;
    layer7_outputs(759) <= a;
    layer7_outputs(760) <= a;
    layer7_outputs(761) <= not b;
    layer7_outputs(762) <= b;
    layer7_outputs(763) <= not a or b;
    layer7_outputs(764) <= not (a or b);
    layer7_outputs(765) <= not (a and b);
    layer7_outputs(766) <= a xor b;
    layer7_outputs(767) <= b;
    layer7_outputs(768) <= not b or a;
    layer7_outputs(769) <= b;
    layer7_outputs(770) <= not b;
    layer7_outputs(771) <= not b or a;
    layer7_outputs(772) <= b;
    layer7_outputs(773) <= not (a xor b);
    layer7_outputs(774) <= a;
    layer7_outputs(775) <= not b;
    layer7_outputs(776) <= not b;
    layer7_outputs(777) <= not (a xor b);
    layer7_outputs(778) <= a;
    layer7_outputs(779) <= a;
    layer7_outputs(780) <= not (a xor b);
    layer7_outputs(781) <= a xor b;
    layer7_outputs(782) <= b and not a;
    layer7_outputs(783) <= not (a or b);
    layer7_outputs(784) <= a and not b;
    layer7_outputs(785) <= not a or b;
    layer7_outputs(786) <= a xor b;
    layer7_outputs(787) <= not b;
    layer7_outputs(788) <= a and b;
    layer7_outputs(789) <= a;
    layer7_outputs(790) <= not (a or b);
    layer7_outputs(791) <= a;
    layer7_outputs(792) <= not (a xor b);
    layer7_outputs(793) <= b and not a;
    layer7_outputs(794) <= a;
    layer7_outputs(795) <= not b or a;
    layer7_outputs(796) <= not b;
    layer7_outputs(797) <= not (a xor b);
    layer7_outputs(798) <= not b;
    layer7_outputs(799) <= not b;
    layer7_outputs(800) <= not a or b;
    layer7_outputs(801) <= a xor b;
    layer7_outputs(802) <= not (a and b);
    layer7_outputs(803) <= not a;
    layer7_outputs(804) <= a;
    layer7_outputs(805) <= not a;
    layer7_outputs(806) <= not (a xor b);
    layer7_outputs(807) <= not a or b;
    layer7_outputs(808) <= not a;
    layer7_outputs(809) <= b and not a;
    layer7_outputs(810) <= a or b;
    layer7_outputs(811) <= not (a xor b);
    layer7_outputs(812) <= not b;
    layer7_outputs(813) <= a;
    layer7_outputs(814) <= not a;
    layer7_outputs(815) <= not b;
    layer7_outputs(816) <= not b;
    layer7_outputs(817) <= not (a and b);
    layer7_outputs(818) <= a xor b;
    layer7_outputs(819) <= b;
    layer7_outputs(820) <= a and not b;
    layer7_outputs(821) <= not b or a;
    layer7_outputs(822) <= a;
    layer7_outputs(823) <= not (a and b);
    layer7_outputs(824) <= not b;
    layer7_outputs(825) <= a and not b;
    layer7_outputs(826) <= not b;
    layer7_outputs(827) <= not a;
    layer7_outputs(828) <= not (a and b);
    layer7_outputs(829) <= b;
    layer7_outputs(830) <= b and not a;
    layer7_outputs(831) <= not b;
    layer7_outputs(832) <= a and not b;
    layer7_outputs(833) <= a and not b;
    layer7_outputs(834) <= a xor b;
    layer7_outputs(835) <= b;
    layer7_outputs(836) <= not b or a;
    layer7_outputs(837) <= a or b;
    layer7_outputs(838) <= a;
    layer7_outputs(839) <= not b;
    layer7_outputs(840) <= not b;
    layer7_outputs(841) <= not b;
    layer7_outputs(842) <= b;
    layer7_outputs(843) <= 1'b0;
    layer7_outputs(844) <= not (a xor b);
    layer7_outputs(845) <= b;
    layer7_outputs(846) <= a and not b;
    layer7_outputs(847) <= a;
    layer7_outputs(848) <= not b;
    layer7_outputs(849) <= not b;
    layer7_outputs(850) <= not a;
    layer7_outputs(851) <= a xor b;
    layer7_outputs(852) <= not b;
    layer7_outputs(853) <= b and not a;
    layer7_outputs(854) <= a xor b;
    layer7_outputs(855) <= a xor b;
    layer7_outputs(856) <= not (a xor b);
    layer7_outputs(857) <= not a;
    layer7_outputs(858) <= a or b;
    layer7_outputs(859) <= not a or b;
    layer7_outputs(860) <= not (a and b);
    layer7_outputs(861) <= not b;
    layer7_outputs(862) <= 1'b0;
    layer7_outputs(863) <= not b or a;
    layer7_outputs(864) <= a;
    layer7_outputs(865) <= b;
    layer7_outputs(866) <= not a;
    layer7_outputs(867) <= a and b;
    layer7_outputs(868) <= a;
    layer7_outputs(869) <= not b;
    layer7_outputs(870) <= not b;
    layer7_outputs(871) <= b;
    layer7_outputs(872) <= not (a and b);
    layer7_outputs(873) <= a or b;
    layer7_outputs(874) <= a;
    layer7_outputs(875) <= not a;
    layer7_outputs(876) <= b;
    layer7_outputs(877) <= b and not a;
    layer7_outputs(878) <= 1'b0;
    layer7_outputs(879) <= a xor b;
    layer7_outputs(880) <= not b;
    layer7_outputs(881) <= a or b;
    layer7_outputs(882) <= a;
    layer7_outputs(883) <= b and not a;
    layer7_outputs(884) <= a xor b;
    layer7_outputs(885) <= not b;
    layer7_outputs(886) <= 1'b0;
    layer7_outputs(887) <= b and not a;
    layer7_outputs(888) <= not (a xor b);
    layer7_outputs(889) <= not b;
    layer7_outputs(890) <= not (a or b);
    layer7_outputs(891) <= not (a xor b);
    layer7_outputs(892) <= not a or b;
    layer7_outputs(893) <= not a;
    layer7_outputs(894) <= not a;
    layer7_outputs(895) <= 1'b1;
    layer7_outputs(896) <= not (a xor b);
    layer7_outputs(897) <= a and not b;
    layer7_outputs(898) <= b and not a;
    layer7_outputs(899) <= a;
    layer7_outputs(900) <= b and not a;
    layer7_outputs(901) <= a and not b;
    layer7_outputs(902) <= a;
    layer7_outputs(903) <= b and not a;
    layer7_outputs(904) <= not b or a;
    layer7_outputs(905) <= a xor b;
    layer7_outputs(906) <= a;
    layer7_outputs(907) <= a xor b;
    layer7_outputs(908) <= a;
    layer7_outputs(909) <= not (a xor b);
    layer7_outputs(910) <= not (a and b);
    layer7_outputs(911) <= not b;
    layer7_outputs(912) <= a and not b;
    layer7_outputs(913) <= a xor b;
    layer7_outputs(914) <= not a;
    layer7_outputs(915) <= not a;
    layer7_outputs(916) <= not b;
    layer7_outputs(917) <= not a;
    layer7_outputs(918) <= b;
    layer7_outputs(919) <= a;
    layer7_outputs(920) <= 1'b0;
    layer7_outputs(921) <= not (a and b);
    layer7_outputs(922) <= a;
    layer7_outputs(923) <= not b;
    layer7_outputs(924) <= not (a or b);
    layer7_outputs(925) <= not a;
    layer7_outputs(926) <= not a or b;
    layer7_outputs(927) <= not b or a;
    layer7_outputs(928) <= b;
    layer7_outputs(929) <= a;
    layer7_outputs(930) <= 1'b0;
    layer7_outputs(931) <= b;
    layer7_outputs(932) <= not a or b;
    layer7_outputs(933) <= not a;
    layer7_outputs(934) <= not b;
    layer7_outputs(935) <= a xor b;
    layer7_outputs(936) <= not b or a;
    layer7_outputs(937) <= 1'b0;
    layer7_outputs(938) <= a;
    layer7_outputs(939) <= not (a or b);
    layer7_outputs(940) <= a and b;
    layer7_outputs(941) <= not (a xor b);
    layer7_outputs(942) <= a xor b;
    layer7_outputs(943) <= not a;
    layer7_outputs(944) <= not (a xor b);
    layer7_outputs(945) <= not b;
    layer7_outputs(946) <= not a or b;
    layer7_outputs(947) <= not b;
    layer7_outputs(948) <= 1'b1;
    layer7_outputs(949) <= not b or a;
    layer7_outputs(950) <= not b;
    layer7_outputs(951) <= 1'b1;
    layer7_outputs(952) <= a and not b;
    layer7_outputs(953) <= a or b;
    layer7_outputs(954) <= a or b;
    layer7_outputs(955) <= b and not a;
    layer7_outputs(956) <= not (a xor b);
    layer7_outputs(957) <= a;
    layer7_outputs(958) <= a xor b;
    layer7_outputs(959) <= not a;
    layer7_outputs(960) <= not a or b;
    layer7_outputs(961) <= not b;
    layer7_outputs(962) <= a or b;
    layer7_outputs(963) <= a xor b;
    layer7_outputs(964) <= a;
    layer7_outputs(965) <= a or b;
    layer7_outputs(966) <= b and not a;
    layer7_outputs(967) <= not (a or b);
    layer7_outputs(968) <= a and not b;
    layer7_outputs(969) <= not a;
    layer7_outputs(970) <= a xor b;
    layer7_outputs(971) <= b;
    layer7_outputs(972) <= a;
    layer7_outputs(973) <= a;
    layer7_outputs(974) <= not a or b;
    layer7_outputs(975) <= not b;
    layer7_outputs(976) <= a;
    layer7_outputs(977) <= b;
    layer7_outputs(978) <= not (a xor b);
    layer7_outputs(979) <= a;
    layer7_outputs(980) <= not a or b;
    layer7_outputs(981) <= b;
    layer7_outputs(982) <= a xor b;
    layer7_outputs(983) <= not b;
    layer7_outputs(984) <= b;
    layer7_outputs(985) <= a;
    layer7_outputs(986) <= b;
    layer7_outputs(987) <= a;
    layer7_outputs(988) <= not a;
    layer7_outputs(989) <= a;
    layer7_outputs(990) <= a;
    layer7_outputs(991) <= 1'b1;
    layer7_outputs(992) <= not (a xor b);
    layer7_outputs(993) <= a xor b;
    layer7_outputs(994) <= not a;
    layer7_outputs(995) <= not (a xor b);
    layer7_outputs(996) <= not a;
    layer7_outputs(997) <= not b;
    layer7_outputs(998) <= not b;
    layer7_outputs(999) <= not b;
    layer7_outputs(1000) <= b;
    layer7_outputs(1001) <= not a;
    layer7_outputs(1002) <= a or b;
    layer7_outputs(1003) <= b;
    layer7_outputs(1004) <= not a;
    layer7_outputs(1005) <= a;
    layer7_outputs(1006) <= a;
    layer7_outputs(1007) <= not b;
    layer7_outputs(1008) <= not a or b;
    layer7_outputs(1009) <= not a or b;
    layer7_outputs(1010) <= a and b;
    layer7_outputs(1011) <= not b;
    layer7_outputs(1012) <= a;
    layer7_outputs(1013) <= b;
    layer7_outputs(1014) <= a;
    layer7_outputs(1015) <= a;
    layer7_outputs(1016) <= b;
    layer7_outputs(1017) <= not b or a;
    layer7_outputs(1018) <= a xor b;
    layer7_outputs(1019) <= a xor b;
    layer7_outputs(1020) <= a;
    layer7_outputs(1021) <= b;
    layer7_outputs(1022) <= not (a xor b);
    layer7_outputs(1023) <= not (a and b);
    layer7_outputs(1024) <= not a or b;
    layer7_outputs(1025) <= a xor b;
    layer7_outputs(1026) <= not b or a;
    layer7_outputs(1027) <= a and not b;
    layer7_outputs(1028) <= not b;
    layer7_outputs(1029) <= not (a and b);
    layer7_outputs(1030) <= not (a xor b);
    layer7_outputs(1031) <= b;
    layer7_outputs(1032) <= a and b;
    layer7_outputs(1033) <= not a;
    layer7_outputs(1034) <= not a;
    layer7_outputs(1035) <= b;
    layer7_outputs(1036) <= not a or b;
    layer7_outputs(1037) <= 1'b0;
    layer7_outputs(1038) <= not (a or b);
    layer7_outputs(1039) <= b and not a;
    layer7_outputs(1040) <= not a;
    layer7_outputs(1041) <= a;
    layer7_outputs(1042) <= not b;
    layer7_outputs(1043) <= b;
    layer7_outputs(1044) <= a;
    layer7_outputs(1045) <= a;
    layer7_outputs(1046) <= b and not a;
    layer7_outputs(1047) <= not b;
    layer7_outputs(1048) <= b and not a;
    layer7_outputs(1049) <= not b;
    layer7_outputs(1050) <= b;
    layer7_outputs(1051) <= b and not a;
    layer7_outputs(1052) <= b;
    layer7_outputs(1053) <= a;
    layer7_outputs(1054) <= b and not a;
    layer7_outputs(1055) <= not a;
    layer7_outputs(1056) <= a and not b;
    layer7_outputs(1057) <= a;
    layer7_outputs(1058) <= not a;
    layer7_outputs(1059) <= a;
    layer7_outputs(1060) <= not a;
    layer7_outputs(1061) <= a xor b;
    layer7_outputs(1062) <= a and not b;
    layer7_outputs(1063) <= not a or b;
    layer7_outputs(1064) <= not a or b;
    layer7_outputs(1065) <= a xor b;
    layer7_outputs(1066) <= not (a or b);
    layer7_outputs(1067) <= not a or b;
    layer7_outputs(1068) <= b and not a;
    layer7_outputs(1069) <= not a;
    layer7_outputs(1070) <= not b;
    layer7_outputs(1071) <= not a;
    layer7_outputs(1072) <= not (a xor b);
    layer7_outputs(1073) <= not b;
    layer7_outputs(1074) <= not a;
    layer7_outputs(1075) <= b;
    layer7_outputs(1076) <= b;
    layer7_outputs(1077) <= a;
    layer7_outputs(1078) <= not b;
    layer7_outputs(1079) <= not a;
    layer7_outputs(1080) <= a and not b;
    layer7_outputs(1081) <= a;
    layer7_outputs(1082) <= not b;
    layer7_outputs(1083) <= not (a xor b);
    layer7_outputs(1084) <= a;
    layer7_outputs(1085) <= not (a xor b);
    layer7_outputs(1086) <= not b;
    layer7_outputs(1087) <= not b;
    layer7_outputs(1088) <= a and not b;
    layer7_outputs(1089) <= a;
    layer7_outputs(1090) <= a and b;
    layer7_outputs(1091) <= b;
    layer7_outputs(1092) <= a or b;
    layer7_outputs(1093) <= 1'b0;
    layer7_outputs(1094) <= not b;
    layer7_outputs(1095) <= a;
    layer7_outputs(1096) <= b;
    layer7_outputs(1097) <= a and not b;
    layer7_outputs(1098) <= b;
    layer7_outputs(1099) <= not a or b;
    layer7_outputs(1100) <= not a or b;
    layer7_outputs(1101) <= a;
    layer7_outputs(1102) <= not (a xor b);
    layer7_outputs(1103) <= a and not b;
    layer7_outputs(1104) <= not b;
    layer7_outputs(1105) <= not b or a;
    layer7_outputs(1106) <= not a;
    layer7_outputs(1107) <= b and not a;
    layer7_outputs(1108) <= a xor b;
    layer7_outputs(1109) <= a;
    layer7_outputs(1110) <= a;
    layer7_outputs(1111) <= not b;
    layer7_outputs(1112) <= not b or a;
    layer7_outputs(1113) <= not a or b;
    layer7_outputs(1114) <= not a;
    layer7_outputs(1115) <= not a;
    layer7_outputs(1116) <= a and not b;
    layer7_outputs(1117) <= b;
    layer7_outputs(1118) <= b;
    layer7_outputs(1119) <= not (a and b);
    layer7_outputs(1120) <= b;
    layer7_outputs(1121) <= a and b;
    layer7_outputs(1122) <= not b;
    layer7_outputs(1123) <= not a;
    layer7_outputs(1124) <= not (a xor b);
    layer7_outputs(1125) <= not (a xor b);
    layer7_outputs(1126) <= not a;
    layer7_outputs(1127) <= a;
    layer7_outputs(1128) <= a xor b;
    layer7_outputs(1129) <= a and not b;
    layer7_outputs(1130) <= not (a xor b);
    layer7_outputs(1131) <= not b;
    layer7_outputs(1132) <= not a;
    layer7_outputs(1133) <= a and b;
    layer7_outputs(1134) <= not a;
    layer7_outputs(1135) <= not b or a;
    layer7_outputs(1136) <= not (a and b);
    layer7_outputs(1137) <= not a;
    layer7_outputs(1138) <= b;
    layer7_outputs(1139) <= a or b;
    layer7_outputs(1140) <= a xor b;
    layer7_outputs(1141) <= not b or a;
    layer7_outputs(1142) <= not (a or b);
    layer7_outputs(1143) <= not (a xor b);
    layer7_outputs(1144) <= b;
    layer7_outputs(1145) <= not (a xor b);
    layer7_outputs(1146) <= a xor b;
    layer7_outputs(1147) <= not b or a;
    layer7_outputs(1148) <= not (a xor b);
    layer7_outputs(1149) <= a and not b;
    layer7_outputs(1150) <= not b;
    layer7_outputs(1151) <= a;
    layer7_outputs(1152) <= b;
    layer7_outputs(1153) <= not b;
    layer7_outputs(1154) <= a and not b;
    layer7_outputs(1155) <= not b or a;
    layer7_outputs(1156) <= not (a and b);
    layer7_outputs(1157) <= 1'b0;
    layer7_outputs(1158) <= a xor b;
    layer7_outputs(1159) <= a and not b;
    layer7_outputs(1160) <= not b;
    layer7_outputs(1161) <= not (a xor b);
    layer7_outputs(1162) <= not a;
    layer7_outputs(1163) <= not (a or b);
    layer7_outputs(1164) <= a or b;
    layer7_outputs(1165) <= b;
    layer7_outputs(1166) <= not b;
    layer7_outputs(1167) <= not a;
    layer7_outputs(1168) <= not b or a;
    layer7_outputs(1169) <= a;
    layer7_outputs(1170) <= a xor b;
    layer7_outputs(1171) <= a and not b;
    layer7_outputs(1172) <= not a;
    layer7_outputs(1173) <= not (a xor b);
    layer7_outputs(1174) <= not b or a;
    layer7_outputs(1175) <= a;
    layer7_outputs(1176) <= a xor b;
    layer7_outputs(1177) <= b and not a;
    layer7_outputs(1178) <= not (a and b);
    layer7_outputs(1179) <= a or b;
    layer7_outputs(1180) <= b;
    layer7_outputs(1181) <= not a or b;
    layer7_outputs(1182) <= a;
    layer7_outputs(1183) <= a and b;
    layer7_outputs(1184) <= 1'b1;
    layer7_outputs(1185) <= not a;
    layer7_outputs(1186) <= not a;
    layer7_outputs(1187) <= a xor b;
    layer7_outputs(1188) <= not b;
    layer7_outputs(1189) <= b;
    layer7_outputs(1190) <= not a;
    layer7_outputs(1191) <= a;
    layer7_outputs(1192) <= b;
    layer7_outputs(1193) <= a;
    layer7_outputs(1194) <= a or b;
    layer7_outputs(1195) <= a xor b;
    layer7_outputs(1196) <= a;
    layer7_outputs(1197) <= not b or a;
    layer7_outputs(1198) <= not (a or b);
    layer7_outputs(1199) <= a;
    layer7_outputs(1200) <= a and not b;
    layer7_outputs(1201) <= not b or a;
    layer7_outputs(1202) <= a xor b;
    layer7_outputs(1203) <= not a or b;
    layer7_outputs(1204) <= not b;
    layer7_outputs(1205) <= a xor b;
    layer7_outputs(1206) <= a;
    layer7_outputs(1207) <= not b;
    layer7_outputs(1208) <= a and not b;
    layer7_outputs(1209) <= a or b;
    layer7_outputs(1210) <= a and b;
    layer7_outputs(1211) <= a xor b;
    layer7_outputs(1212) <= a and b;
    layer7_outputs(1213) <= not b;
    layer7_outputs(1214) <= b and not a;
    layer7_outputs(1215) <= a xor b;
    layer7_outputs(1216) <= not (a or b);
    layer7_outputs(1217) <= b;
    layer7_outputs(1218) <= not (a and b);
    layer7_outputs(1219) <= not a or b;
    layer7_outputs(1220) <= a or b;
    layer7_outputs(1221) <= a and b;
    layer7_outputs(1222) <= a xor b;
    layer7_outputs(1223) <= a and not b;
    layer7_outputs(1224) <= a and not b;
    layer7_outputs(1225) <= a and b;
    layer7_outputs(1226) <= not (a or b);
    layer7_outputs(1227) <= a or b;
    layer7_outputs(1228) <= a;
    layer7_outputs(1229) <= 1'b0;
    layer7_outputs(1230) <= a and b;
    layer7_outputs(1231) <= a or b;
    layer7_outputs(1232) <= not b;
    layer7_outputs(1233) <= b;
    layer7_outputs(1234) <= a and b;
    layer7_outputs(1235) <= not (a xor b);
    layer7_outputs(1236) <= not (a or b);
    layer7_outputs(1237) <= not b;
    layer7_outputs(1238) <= b;
    layer7_outputs(1239) <= b;
    layer7_outputs(1240) <= not b;
    layer7_outputs(1241) <= a;
    layer7_outputs(1242) <= not a;
    layer7_outputs(1243) <= not (a or b);
    layer7_outputs(1244) <= not (a or b);
    layer7_outputs(1245) <= b;
    layer7_outputs(1246) <= b and not a;
    layer7_outputs(1247) <= not a;
    layer7_outputs(1248) <= not a or b;
    layer7_outputs(1249) <= not a or b;
    layer7_outputs(1250) <= not (a and b);
    layer7_outputs(1251) <= not a;
    layer7_outputs(1252) <= not a;
    layer7_outputs(1253) <= a;
    layer7_outputs(1254) <= b;
    layer7_outputs(1255) <= a xor b;
    layer7_outputs(1256) <= not a or b;
    layer7_outputs(1257) <= a;
    layer7_outputs(1258) <= not b;
    layer7_outputs(1259) <= not (a and b);
    layer7_outputs(1260) <= not (a xor b);
    layer7_outputs(1261) <= a;
    layer7_outputs(1262) <= not a or b;
    layer7_outputs(1263) <= not b or a;
    layer7_outputs(1264) <= a xor b;
    layer7_outputs(1265) <= not a;
    layer7_outputs(1266) <= a and not b;
    layer7_outputs(1267) <= a or b;
    layer7_outputs(1268) <= not a;
    layer7_outputs(1269) <= a xor b;
    layer7_outputs(1270) <= a xor b;
    layer7_outputs(1271) <= not a;
    layer7_outputs(1272) <= a;
    layer7_outputs(1273) <= a and not b;
    layer7_outputs(1274) <= not b;
    layer7_outputs(1275) <= a or b;
    layer7_outputs(1276) <= not (a and b);
    layer7_outputs(1277) <= a and b;
    layer7_outputs(1278) <= a xor b;
    layer7_outputs(1279) <= b;
    layer7_outputs(1280) <= 1'b1;
    layer7_outputs(1281) <= a and b;
    layer7_outputs(1282) <= a or b;
    layer7_outputs(1283) <= a or b;
    layer7_outputs(1284) <= a;
    layer7_outputs(1285) <= not a;
    layer7_outputs(1286) <= b;
    layer7_outputs(1287) <= not (a and b);
    layer7_outputs(1288) <= not b;
    layer7_outputs(1289) <= a or b;
    layer7_outputs(1290) <= a xor b;
    layer7_outputs(1291) <= a xor b;
    layer7_outputs(1292) <= b and not a;
    layer7_outputs(1293) <= not b;
    layer7_outputs(1294) <= not (a or b);
    layer7_outputs(1295) <= not (a xor b);
    layer7_outputs(1296) <= b;
    layer7_outputs(1297) <= not (a or b);
    layer7_outputs(1298) <= not b;
    layer7_outputs(1299) <= not b;
    layer7_outputs(1300) <= not a;
    layer7_outputs(1301) <= b;
    layer7_outputs(1302) <= b;
    layer7_outputs(1303) <= a xor b;
    layer7_outputs(1304) <= a;
    layer7_outputs(1305) <= not b or a;
    layer7_outputs(1306) <= a and not b;
    layer7_outputs(1307) <= a;
    layer7_outputs(1308) <= not b or a;
    layer7_outputs(1309) <= not (a and b);
    layer7_outputs(1310) <= not b or a;
    layer7_outputs(1311) <= not a;
    layer7_outputs(1312) <= not b or a;
    layer7_outputs(1313) <= b;
    layer7_outputs(1314) <= a xor b;
    layer7_outputs(1315) <= a;
    layer7_outputs(1316) <= b;
    layer7_outputs(1317) <= not b or a;
    layer7_outputs(1318) <= not (a and b);
    layer7_outputs(1319) <= a and b;
    layer7_outputs(1320) <= not b;
    layer7_outputs(1321) <= a and b;
    layer7_outputs(1322) <= a xor b;
    layer7_outputs(1323) <= b;
    layer7_outputs(1324) <= 1'b0;
    layer7_outputs(1325) <= not a or b;
    layer7_outputs(1326) <= a;
    layer7_outputs(1327) <= not a;
    layer7_outputs(1328) <= a and b;
    layer7_outputs(1329) <= not a;
    layer7_outputs(1330) <= not b;
    layer7_outputs(1331) <= not (a and b);
    layer7_outputs(1332) <= not (a and b);
    layer7_outputs(1333) <= a xor b;
    layer7_outputs(1334) <= a and b;
    layer7_outputs(1335) <= a xor b;
    layer7_outputs(1336) <= b and not a;
    layer7_outputs(1337) <= not (a xor b);
    layer7_outputs(1338) <= not (a xor b);
    layer7_outputs(1339) <= b and not a;
    layer7_outputs(1340) <= a and not b;
    layer7_outputs(1341) <= not a or b;
    layer7_outputs(1342) <= 1'b1;
    layer7_outputs(1343) <= b;
    layer7_outputs(1344) <= not a;
    layer7_outputs(1345) <= a xor b;
    layer7_outputs(1346) <= b;
    layer7_outputs(1347) <= b;
    layer7_outputs(1348) <= not a;
    layer7_outputs(1349) <= a;
    layer7_outputs(1350) <= a and b;
    layer7_outputs(1351) <= not (a or b);
    layer7_outputs(1352) <= b and not a;
    layer7_outputs(1353) <= a;
    layer7_outputs(1354) <= 1'b1;
    layer7_outputs(1355) <= not b;
    layer7_outputs(1356) <= a;
    layer7_outputs(1357) <= a;
    layer7_outputs(1358) <= not (a xor b);
    layer7_outputs(1359) <= not a;
    layer7_outputs(1360) <= not a or b;
    layer7_outputs(1361) <= a or b;
    layer7_outputs(1362) <= a xor b;
    layer7_outputs(1363) <= not a;
    layer7_outputs(1364) <= b;
    layer7_outputs(1365) <= not b;
    layer7_outputs(1366) <= a or b;
    layer7_outputs(1367) <= not (a or b);
    layer7_outputs(1368) <= a;
    layer7_outputs(1369) <= a;
    layer7_outputs(1370) <= not a;
    layer7_outputs(1371) <= not (a xor b);
    layer7_outputs(1372) <= not (a or b);
    layer7_outputs(1373) <= not a;
    layer7_outputs(1374) <= a xor b;
    layer7_outputs(1375) <= not a;
    layer7_outputs(1376) <= b;
    layer7_outputs(1377) <= not b;
    layer7_outputs(1378) <= a xor b;
    layer7_outputs(1379) <= not a;
    layer7_outputs(1380) <= a or b;
    layer7_outputs(1381) <= a;
    layer7_outputs(1382) <= not b;
    layer7_outputs(1383) <= a and b;
    layer7_outputs(1384) <= b;
    layer7_outputs(1385) <= not b or a;
    layer7_outputs(1386) <= not (a or b);
    layer7_outputs(1387) <= not b;
    layer7_outputs(1388) <= b;
    layer7_outputs(1389) <= a xor b;
    layer7_outputs(1390) <= a;
    layer7_outputs(1391) <= a xor b;
    layer7_outputs(1392) <= not a or b;
    layer7_outputs(1393) <= not (a xor b);
    layer7_outputs(1394) <= not a;
    layer7_outputs(1395) <= not (a xor b);
    layer7_outputs(1396) <= a;
    layer7_outputs(1397) <= not b;
    layer7_outputs(1398) <= 1'b0;
    layer7_outputs(1399) <= not b;
    layer7_outputs(1400) <= a or b;
    layer7_outputs(1401) <= b;
    layer7_outputs(1402) <= a xor b;
    layer7_outputs(1403) <= a xor b;
    layer7_outputs(1404) <= not b;
    layer7_outputs(1405) <= not b;
    layer7_outputs(1406) <= not (a and b);
    layer7_outputs(1407) <= not (a and b);
    layer7_outputs(1408) <= not a;
    layer7_outputs(1409) <= b;
    layer7_outputs(1410) <= not (a xor b);
    layer7_outputs(1411) <= not a;
    layer7_outputs(1412) <= not a;
    layer7_outputs(1413) <= 1'b0;
    layer7_outputs(1414) <= a or b;
    layer7_outputs(1415) <= a xor b;
    layer7_outputs(1416) <= not (a or b);
    layer7_outputs(1417) <= not b;
    layer7_outputs(1418) <= not (a and b);
    layer7_outputs(1419) <= b;
    layer7_outputs(1420) <= not a;
    layer7_outputs(1421) <= not b;
    layer7_outputs(1422) <= not b;
    layer7_outputs(1423) <= a;
    layer7_outputs(1424) <= not (a and b);
    layer7_outputs(1425) <= not b;
    layer7_outputs(1426) <= not b;
    layer7_outputs(1427) <= not b;
    layer7_outputs(1428) <= a xor b;
    layer7_outputs(1429) <= not a;
    layer7_outputs(1430) <= a xor b;
    layer7_outputs(1431) <= a or b;
    layer7_outputs(1432) <= not a or b;
    layer7_outputs(1433) <= not (a and b);
    layer7_outputs(1434) <= not a;
    layer7_outputs(1435) <= a or b;
    layer7_outputs(1436) <= a or b;
    layer7_outputs(1437) <= a or b;
    layer7_outputs(1438) <= b;
    layer7_outputs(1439) <= not (a and b);
    layer7_outputs(1440) <= not a;
    layer7_outputs(1441) <= a or b;
    layer7_outputs(1442) <= b;
    layer7_outputs(1443) <= a or b;
    layer7_outputs(1444) <= a or b;
    layer7_outputs(1445) <= not (a or b);
    layer7_outputs(1446) <= not a;
    layer7_outputs(1447) <= a and b;
    layer7_outputs(1448) <= b;
    layer7_outputs(1449) <= b;
    layer7_outputs(1450) <= a xor b;
    layer7_outputs(1451) <= not (a xor b);
    layer7_outputs(1452) <= a and b;
    layer7_outputs(1453) <= not a;
    layer7_outputs(1454) <= not (a xor b);
    layer7_outputs(1455) <= a or b;
    layer7_outputs(1456) <= a;
    layer7_outputs(1457) <= a xor b;
    layer7_outputs(1458) <= a and not b;
    layer7_outputs(1459) <= a and not b;
    layer7_outputs(1460) <= not b or a;
    layer7_outputs(1461) <= not a;
    layer7_outputs(1462) <= a and not b;
    layer7_outputs(1463) <= a;
    layer7_outputs(1464) <= not b;
    layer7_outputs(1465) <= not b;
    layer7_outputs(1466) <= not a or b;
    layer7_outputs(1467) <= a and b;
    layer7_outputs(1468) <= a and b;
    layer7_outputs(1469) <= not (a xor b);
    layer7_outputs(1470) <= not (a and b);
    layer7_outputs(1471) <= b;
    layer7_outputs(1472) <= not a or b;
    layer7_outputs(1473) <= not (a or b);
    layer7_outputs(1474) <= a or b;
    layer7_outputs(1475) <= not (a xor b);
    layer7_outputs(1476) <= not a or b;
    layer7_outputs(1477) <= a;
    layer7_outputs(1478) <= a;
    layer7_outputs(1479) <= not (a or b);
    layer7_outputs(1480) <= b;
    layer7_outputs(1481) <= not (a or b);
    layer7_outputs(1482) <= not (a xor b);
    layer7_outputs(1483) <= a;
    layer7_outputs(1484) <= not a or b;
    layer7_outputs(1485) <= a;
    layer7_outputs(1486) <= not (a and b);
    layer7_outputs(1487) <= not b;
    layer7_outputs(1488) <= not b;
    layer7_outputs(1489) <= not a;
    layer7_outputs(1490) <= a or b;
    layer7_outputs(1491) <= a;
    layer7_outputs(1492) <= a and not b;
    layer7_outputs(1493) <= not (a and b);
    layer7_outputs(1494) <= not b or a;
    layer7_outputs(1495) <= a;
    layer7_outputs(1496) <= not (a xor b);
    layer7_outputs(1497) <= a xor b;
    layer7_outputs(1498) <= not (a or b);
    layer7_outputs(1499) <= a;
    layer7_outputs(1500) <= not b or a;
    layer7_outputs(1501) <= not (a and b);
    layer7_outputs(1502) <= b and not a;
    layer7_outputs(1503) <= a or b;
    layer7_outputs(1504) <= a xor b;
    layer7_outputs(1505) <= b and not a;
    layer7_outputs(1506) <= a xor b;
    layer7_outputs(1507) <= not b or a;
    layer7_outputs(1508) <= a;
    layer7_outputs(1509) <= b;
    layer7_outputs(1510) <= not a or b;
    layer7_outputs(1511) <= a;
    layer7_outputs(1512) <= a;
    layer7_outputs(1513) <= not b or a;
    layer7_outputs(1514) <= not b;
    layer7_outputs(1515) <= b and not a;
    layer7_outputs(1516) <= a xor b;
    layer7_outputs(1517) <= a;
    layer7_outputs(1518) <= a;
    layer7_outputs(1519) <= a xor b;
    layer7_outputs(1520) <= not (a xor b);
    layer7_outputs(1521) <= not (a xor b);
    layer7_outputs(1522) <= not b;
    layer7_outputs(1523) <= b;
    layer7_outputs(1524) <= not (a or b);
    layer7_outputs(1525) <= not (a or b);
    layer7_outputs(1526) <= 1'b1;
    layer7_outputs(1527) <= a xor b;
    layer7_outputs(1528) <= a or b;
    layer7_outputs(1529) <= not b or a;
    layer7_outputs(1530) <= not b or a;
    layer7_outputs(1531) <= not (a and b);
    layer7_outputs(1532) <= b and not a;
    layer7_outputs(1533) <= not b or a;
    layer7_outputs(1534) <= a xor b;
    layer7_outputs(1535) <= not (a xor b);
    layer7_outputs(1536) <= not (a and b);
    layer7_outputs(1537) <= a and not b;
    layer7_outputs(1538) <= a and b;
    layer7_outputs(1539) <= not a;
    layer7_outputs(1540) <= not (a xor b);
    layer7_outputs(1541) <= not b;
    layer7_outputs(1542) <= a xor b;
    layer7_outputs(1543) <= a or b;
    layer7_outputs(1544) <= not a;
    layer7_outputs(1545) <= a or b;
    layer7_outputs(1546) <= not (a or b);
    layer7_outputs(1547) <= b;
    layer7_outputs(1548) <= not a or b;
    layer7_outputs(1549) <= a xor b;
    layer7_outputs(1550) <= a;
    layer7_outputs(1551) <= b and not a;
    layer7_outputs(1552) <= not (a and b);
    layer7_outputs(1553) <= a or b;
    layer7_outputs(1554) <= not a;
    layer7_outputs(1555) <= not a;
    layer7_outputs(1556) <= a;
    layer7_outputs(1557) <= a;
    layer7_outputs(1558) <= a and b;
    layer7_outputs(1559) <= not (a xor b);
    layer7_outputs(1560) <= not (a and b);
    layer7_outputs(1561) <= a;
    layer7_outputs(1562) <= a and b;
    layer7_outputs(1563) <= not a;
    layer7_outputs(1564) <= a xor b;
    layer7_outputs(1565) <= a and b;
    layer7_outputs(1566) <= not b;
    layer7_outputs(1567) <= a;
    layer7_outputs(1568) <= a;
    layer7_outputs(1569) <= b;
    layer7_outputs(1570) <= b;
    layer7_outputs(1571) <= not b;
    layer7_outputs(1572) <= b;
    layer7_outputs(1573) <= a;
    layer7_outputs(1574) <= not b;
    layer7_outputs(1575) <= not a;
    layer7_outputs(1576) <= b;
    layer7_outputs(1577) <= not (a and b);
    layer7_outputs(1578) <= a xor b;
    layer7_outputs(1579) <= b;
    layer7_outputs(1580) <= a and b;
    layer7_outputs(1581) <= b;
    layer7_outputs(1582) <= b and not a;
    layer7_outputs(1583) <= a and b;
    layer7_outputs(1584) <= not b;
    layer7_outputs(1585) <= not a;
    layer7_outputs(1586) <= a xor b;
    layer7_outputs(1587) <= not a;
    layer7_outputs(1588) <= not (a or b);
    layer7_outputs(1589) <= a;
    layer7_outputs(1590) <= a;
    layer7_outputs(1591) <= not (a xor b);
    layer7_outputs(1592) <= a;
    layer7_outputs(1593) <= a or b;
    layer7_outputs(1594) <= not b;
    layer7_outputs(1595) <= not b;
    layer7_outputs(1596) <= not a;
    layer7_outputs(1597) <= not a or b;
    layer7_outputs(1598) <= a and b;
    layer7_outputs(1599) <= b;
    layer7_outputs(1600) <= not (a xor b);
    layer7_outputs(1601) <= a and b;
    layer7_outputs(1602) <= not (a xor b);
    layer7_outputs(1603) <= a;
    layer7_outputs(1604) <= not b;
    layer7_outputs(1605) <= a xor b;
    layer7_outputs(1606) <= not (a xor b);
    layer7_outputs(1607) <= a;
    layer7_outputs(1608) <= a;
    layer7_outputs(1609) <= 1'b0;
    layer7_outputs(1610) <= not b;
    layer7_outputs(1611) <= b and not a;
    layer7_outputs(1612) <= 1'b1;
    layer7_outputs(1613) <= b;
    layer7_outputs(1614) <= not a;
    layer7_outputs(1615) <= not (a xor b);
    layer7_outputs(1616) <= a;
    layer7_outputs(1617) <= b;
    layer7_outputs(1618) <= not b or a;
    layer7_outputs(1619) <= b;
    layer7_outputs(1620) <= not (a or b);
    layer7_outputs(1621) <= a xor b;
    layer7_outputs(1622) <= a and not b;
    layer7_outputs(1623) <= 1'b0;
    layer7_outputs(1624) <= b and not a;
    layer7_outputs(1625) <= not a;
    layer7_outputs(1626) <= not a or b;
    layer7_outputs(1627) <= b;
    layer7_outputs(1628) <= not a;
    layer7_outputs(1629) <= a;
    layer7_outputs(1630) <= not a;
    layer7_outputs(1631) <= not b;
    layer7_outputs(1632) <= a and not b;
    layer7_outputs(1633) <= not a or b;
    layer7_outputs(1634) <= b and not a;
    layer7_outputs(1635) <= a xor b;
    layer7_outputs(1636) <= not a or b;
    layer7_outputs(1637) <= not b;
    layer7_outputs(1638) <= not (a xor b);
    layer7_outputs(1639) <= b;
    layer7_outputs(1640) <= not b;
    layer7_outputs(1641) <= not b;
    layer7_outputs(1642) <= a and b;
    layer7_outputs(1643) <= not (a and b);
    layer7_outputs(1644) <= a or b;
    layer7_outputs(1645) <= not a or b;
    layer7_outputs(1646) <= not (a or b);
    layer7_outputs(1647) <= b and not a;
    layer7_outputs(1648) <= a;
    layer7_outputs(1649) <= 1'b0;
    layer7_outputs(1650) <= a xor b;
    layer7_outputs(1651) <= a;
    layer7_outputs(1652) <= not a;
    layer7_outputs(1653) <= not a;
    layer7_outputs(1654) <= not b;
    layer7_outputs(1655) <= not (a and b);
    layer7_outputs(1656) <= a or b;
    layer7_outputs(1657) <= not (a xor b);
    layer7_outputs(1658) <= a;
    layer7_outputs(1659) <= a;
    layer7_outputs(1660) <= b;
    layer7_outputs(1661) <= 1'b1;
    layer7_outputs(1662) <= b;
    layer7_outputs(1663) <= not a or b;
    layer7_outputs(1664) <= a or b;
    layer7_outputs(1665) <= not b;
    layer7_outputs(1666) <= b;
    layer7_outputs(1667) <= not a;
    layer7_outputs(1668) <= b;
    layer7_outputs(1669) <= a xor b;
    layer7_outputs(1670) <= a xor b;
    layer7_outputs(1671) <= b;
    layer7_outputs(1672) <= a and b;
    layer7_outputs(1673) <= b;
    layer7_outputs(1674) <= not a;
    layer7_outputs(1675) <= 1'b0;
    layer7_outputs(1676) <= not b;
    layer7_outputs(1677) <= not (a or b);
    layer7_outputs(1678) <= a and not b;
    layer7_outputs(1679) <= not b or a;
    layer7_outputs(1680) <= not b or a;
    layer7_outputs(1681) <= not (a xor b);
    layer7_outputs(1682) <= not b;
    layer7_outputs(1683) <= a;
    layer7_outputs(1684) <= 1'b1;
    layer7_outputs(1685) <= not (a or b);
    layer7_outputs(1686) <= b;
    layer7_outputs(1687) <= not b or a;
    layer7_outputs(1688) <= not a;
    layer7_outputs(1689) <= not a;
    layer7_outputs(1690) <= not (a or b);
    layer7_outputs(1691) <= not b or a;
    layer7_outputs(1692) <= not a;
    layer7_outputs(1693) <= not b;
    layer7_outputs(1694) <= not b;
    layer7_outputs(1695) <= not b;
    layer7_outputs(1696) <= not b;
    layer7_outputs(1697) <= not a or b;
    layer7_outputs(1698) <= not (a xor b);
    layer7_outputs(1699) <= not (a xor b);
    layer7_outputs(1700) <= not b;
    layer7_outputs(1701) <= 1'b1;
    layer7_outputs(1702) <= b;
    layer7_outputs(1703) <= a or b;
    layer7_outputs(1704) <= a and not b;
    layer7_outputs(1705) <= a;
    layer7_outputs(1706) <= a;
    layer7_outputs(1707) <= b and not a;
    layer7_outputs(1708) <= not a or b;
    layer7_outputs(1709) <= a and b;
    layer7_outputs(1710) <= not a;
    layer7_outputs(1711) <= not (a xor b);
    layer7_outputs(1712) <= a;
    layer7_outputs(1713) <= not (a or b);
    layer7_outputs(1714) <= a;
    layer7_outputs(1715) <= a xor b;
    layer7_outputs(1716) <= not a;
    layer7_outputs(1717) <= not a;
    layer7_outputs(1718) <= a xor b;
    layer7_outputs(1719) <= not (a and b);
    layer7_outputs(1720) <= a and not b;
    layer7_outputs(1721) <= a;
    layer7_outputs(1722) <= b and not a;
    layer7_outputs(1723) <= not a or b;
    layer7_outputs(1724) <= not b;
    layer7_outputs(1725) <= a;
    layer7_outputs(1726) <= a;
    layer7_outputs(1727) <= not b;
    layer7_outputs(1728) <= a;
    layer7_outputs(1729) <= a;
    layer7_outputs(1730) <= not b;
    layer7_outputs(1731) <= not a;
    layer7_outputs(1732) <= a xor b;
    layer7_outputs(1733) <= a and b;
    layer7_outputs(1734) <= not (a and b);
    layer7_outputs(1735) <= not a;
    layer7_outputs(1736) <= not a;
    layer7_outputs(1737) <= b and not a;
    layer7_outputs(1738) <= not b or a;
    layer7_outputs(1739) <= not b or a;
    layer7_outputs(1740) <= b;
    layer7_outputs(1741) <= a and b;
    layer7_outputs(1742) <= a and not b;
    layer7_outputs(1743) <= not b;
    layer7_outputs(1744) <= a;
    layer7_outputs(1745) <= a;
    layer7_outputs(1746) <= b;
    layer7_outputs(1747) <= not a;
    layer7_outputs(1748) <= a;
    layer7_outputs(1749) <= not b;
    layer7_outputs(1750) <= not b or a;
    layer7_outputs(1751) <= a xor b;
    layer7_outputs(1752) <= b and not a;
    layer7_outputs(1753) <= b;
    layer7_outputs(1754) <= a;
    layer7_outputs(1755) <= b;
    layer7_outputs(1756) <= a and b;
    layer7_outputs(1757) <= b;
    layer7_outputs(1758) <= b;
    layer7_outputs(1759) <= a;
    layer7_outputs(1760) <= not a;
    layer7_outputs(1761) <= a xor b;
    layer7_outputs(1762) <= not (a xor b);
    layer7_outputs(1763) <= a xor b;
    layer7_outputs(1764) <= not (a or b);
    layer7_outputs(1765) <= a;
    layer7_outputs(1766) <= not (a and b);
    layer7_outputs(1767) <= a or b;
    layer7_outputs(1768) <= a;
    layer7_outputs(1769) <= a and not b;
    layer7_outputs(1770) <= a and b;
    layer7_outputs(1771) <= not (a xor b);
    layer7_outputs(1772) <= a;
    layer7_outputs(1773) <= 1'b0;
    layer7_outputs(1774) <= not a;
    layer7_outputs(1775) <= not a;
    layer7_outputs(1776) <= b and not a;
    layer7_outputs(1777) <= a;
    layer7_outputs(1778) <= b;
    layer7_outputs(1779) <= b;
    layer7_outputs(1780) <= a;
    layer7_outputs(1781) <= not b;
    layer7_outputs(1782) <= a and b;
    layer7_outputs(1783) <= not b or a;
    layer7_outputs(1784) <= not (a xor b);
    layer7_outputs(1785) <= b;
    layer7_outputs(1786) <= not (a xor b);
    layer7_outputs(1787) <= a and not b;
    layer7_outputs(1788) <= a xor b;
    layer7_outputs(1789) <= a and b;
    layer7_outputs(1790) <= a;
    layer7_outputs(1791) <= not (a and b);
    layer7_outputs(1792) <= not b;
    layer7_outputs(1793) <= b;
    layer7_outputs(1794) <= a;
    layer7_outputs(1795) <= b;
    layer7_outputs(1796) <= not (a xor b);
    layer7_outputs(1797) <= a xor b;
    layer7_outputs(1798) <= a xor b;
    layer7_outputs(1799) <= not (a xor b);
    layer7_outputs(1800) <= a;
    layer7_outputs(1801) <= not (a or b);
    layer7_outputs(1802) <= a and not b;
    layer7_outputs(1803) <= a;
    layer7_outputs(1804) <= not a;
    layer7_outputs(1805) <= not b or a;
    layer7_outputs(1806) <= not a or b;
    layer7_outputs(1807) <= a and not b;
    layer7_outputs(1808) <= a;
    layer7_outputs(1809) <= a;
    layer7_outputs(1810) <= not (a xor b);
    layer7_outputs(1811) <= not b;
    layer7_outputs(1812) <= b;
    layer7_outputs(1813) <= not b;
    layer7_outputs(1814) <= not (a or b);
    layer7_outputs(1815) <= a or b;
    layer7_outputs(1816) <= a;
    layer7_outputs(1817) <= not a;
    layer7_outputs(1818) <= a xor b;
    layer7_outputs(1819) <= b;
    layer7_outputs(1820) <= not a;
    layer7_outputs(1821) <= not (a and b);
    layer7_outputs(1822) <= b;
    layer7_outputs(1823) <= 1'b1;
    layer7_outputs(1824) <= a and b;
    layer7_outputs(1825) <= not a;
    layer7_outputs(1826) <= not (a or b);
    layer7_outputs(1827) <= a xor b;
    layer7_outputs(1828) <= not b or a;
    layer7_outputs(1829) <= not a;
    layer7_outputs(1830) <= b and not a;
    layer7_outputs(1831) <= not a or b;
    layer7_outputs(1832) <= b and not a;
    layer7_outputs(1833) <= b;
    layer7_outputs(1834) <= b;
    layer7_outputs(1835) <= 1'b1;
    layer7_outputs(1836) <= not (a xor b);
    layer7_outputs(1837) <= b;
    layer7_outputs(1838) <= a;
    layer7_outputs(1839) <= not a;
    layer7_outputs(1840) <= not b or a;
    layer7_outputs(1841) <= a and b;
    layer7_outputs(1842) <= not b;
    layer7_outputs(1843) <= not a;
    layer7_outputs(1844) <= a xor b;
    layer7_outputs(1845) <= not (a xor b);
    layer7_outputs(1846) <= 1'b1;
    layer7_outputs(1847) <= b and not a;
    layer7_outputs(1848) <= not (a and b);
    layer7_outputs(1849) <= not (a xor b);
    layer7_outputs(1850) <= a;
    layer7_outputs(1851) <= a;
    layer7_outputs(1852) <= a and not b;
    layer7_outputs(1853) <= a and not b;
    layer7_outputs(1854) <= not (a xor b);
    layer7_outputs(1855) <= not b;
    layer7_outputs(1856) <= a xor b;
    layer7_outputs(1857) <= not b or a;
    layer7_outputs(1858) <= a;
    layer7_outputs(1859) <= a;
    layer7_outputs(1860) <= a;
    layer7_outputs(1861) <= not b;
    layer7_outputs(1862) <= not a;
    layer7_outputs(1863) <= not (a xor b);
    layer7_outputs(1864) <= a xor b;
    layer7_outputs(1865) <= not (a or b);
    layer7_outputs(1866) <= not a;
    layer7_outputs(1867) <= not b;
    layer7_outputs(1868) <= not (a xor b);
    layer7_outputs(1869) <= b;
    layer7_outputs(1870) <= not b;
    layer7_outputs(1871) <= b;
    layer7_outputs(1872) <= a xor b;
    layer7_outputs(1873) <= a and not b;
    layer7_outputs(1874) <= not (a and b);
    layer7_outputs(1875) <= not a;
    layer7_outputs(1876) <= b and not a;
    layer7_outputs(1877) <= not b;
    layer7_outputs(1878) <= a and not b;
    layer7_outputs(1879) <= not b;
    layer7_outputs(1880) <= a;
    layer7_outputs(1881) <= not a;
    layer7_outputs(1882) <= a or b;
    layer7_outputs(1883) <= b and not a;
    layer7_outputs(1884) <= a xor b;
    layer7_outputs(1885) <= b;
    layer7_outputs(1886) <= b;
    layer7_outputs(1887) <= not (a xor b);
    layer7_outputs(1888) <= a and b;
    layer7_outputs(1889) <= not (a and b);
    layer7_outputs(1890) <= b and not a;
    layer7_outputs(1891) <= not a or b;
    layer7_outputs(1892) <= a or b;
    layer7_outputs(1893) <= a and b;
    layer7_outputs(1894) <= a xor b;
    layer7_outputs(1895) <= not a;
    layer7_outputs(1896) <= not a or b;
    layer7_outputs(1897) <= not b;
    layer7_outputs(1898) <= a xor b;
    layer7_outputs(1899) <= not (a or b);
    layer7_outputs(1900) <= a xor b;
    layer7_outputs(1901) <= b;
    layer7_outputs(1902) <= not b or a;
    layer7_outputs(1903) <= a or b;
    layer7_outputs(1904) <= a xor b;
    layer7_outputs(1905) <= b;
    layer7_outputs(1906) <= not b;
    layer7_outputs(1907) <= not (a and b);
    layer7_outputs(1908) <= b and not a;
    layer7_outputs(1909) <= not (a or b);
    layer7_outputs(1910) <= a or b;
    layer7_outputs(1911) <= a and b;
    layer7_outputs(1912) <= a and b;
    layer7_outputs(1913) <= not (a and b);
    layer7_outputs(1914) <= a or b;
    layer7_outputs(1915) <= not a;
    layer7_outputs(1916) <= not b;
    layer7_outputs(1917) <= b;
    layer7_outputs(1918) <= not b or a;
    layer7_outputs(1919) <= a xor b;
    layer7_outputs(1920) <= b;
    layer7_outputs(1921) <= a and b;
    layer7_outputs(1922) <= b;
    layer7_outputs(1923) <= not a;
    layer7_outputs(1924) <= not a;
    layer7_outputs(1925) <= a;
    layer7_outputs(1926) <= not b;
    layer7_outputs(1927) <= a and b;
    layer7_outputs(1928) <= b and not a;
    layer7_outputs(1929) <= not (a or b);
    layer7_outputs(1930) <= not (a and b);
    layer7_outputs(1931) <= b and not a;
    layer7_outputs(1932) <= not b or a;
    layer7_outputs(1933) <= a xor b;
    layer7_outputs(1934) <= not b;
    layer7_outputs(1935) <= a;
    layer7_outputs(1936) <= a;
    layer7_outputs(1937) <= not (a xor b);
    layer7_outputs(1938) <= b;
    layer7_outputs(1939) <= a and not b;
    layer7_outputs(1940) <= not a or b;
    layer7_outputs(1941) <= not (a xor b);
    layer7_outputs(1942) <= not b;
    layer7_outputs(1943) <= not b;
    layer7_outputs(1944) <= not b or a;
    layer7_outputs(1945) <= not a;
    layer7_outputs(1946) <= not (a or b);
    layer7_outputs(1947) <= b;
    layer7_outputs(1948) <= not b;
    layer7_outputs(1949) <= not b or a;
    layer7_outputs(1950) <= not a;
    layer7_outputs(1951) <= a and not b;
    layer7_outputs(1952) <= not (a or b);
    layer7_outputs(1953) <= not b;
    layer7_outputs(1954) <= not b;
    layer7_outputs(1955) <= b;
    layer7_outputs(1956) <= a or b;
    layer7_outputs(1957) <= a and not b;
    layer7_outputs(1958) <= not a;
    layer7_outputs(1959) <= a;
    layer7_outputs(1960) <= a;
    layer7_outputs(1961) <= not b;
    layer7_outputs(1962) <= a or b;
    layer7_outputs(1963) <= b;
    layer7_outputs(1964) <= not (a xor b);
    layer7_outputs(1965) <= a;
    layer7_outputs(1966) <= not a or b;
    layer7_outputs(1967) <= not b;
    layer7_outputs(1968) <= a;
    layer7_outputs(1969) <= a;
    layer7_outputs(1970) <= a and b;
    layer7_outputs(1971) <= b;
    layer7_outputs(1972) <= not b;
    layer7_outputs(1973) <= not (a or b);
    layer7_outputs(1974) <= not (a xor b);
    layer7_outputs(1975) <= a or b;
    layer7_outputs(1976) <= not b;
    layer7_outputs(1977) <= not (a xor b);
    layer7_outputs(1978) <= not b or a;
    layer7_outputs(1979) <= not a;
    layer7_outputs(1980) <= not (a or b);
    layer7_outputs(1981) <= a and b;
    layer7_outputs(1982) <= not b;
    layer7_outputs(1983) <= 1'b0;
    layer7_outputs(1984) <= b;
    layer7_outputs(1985) <= not b;
    layer7_outputs(1986) <= a or b;
    layer7_outputs(1987) <= not (a or b);
    layer7_outputs(1988) <= not a;
    layer7_outputs(1989) <= not (a or b);
    layer7_outputs(1990) <= not b or a;
    layer7_outputs(1991) <= not b or a;
    layer7_outputs(1992) <= not (a or b);
    layer7_outputs(1993) <= a xor b;
    layer7_outputs(1994) <= not b;
    layer7_outputs(1995) <= not (a and b);
    layer7_outputs(1996) <= not (a and b);
    layer7_outputs(1997) <= not (a xor b);
    layer7_outputs(1998) <= b and not a;
    layer7_outputs(1999) <= b and not a;
    layer7_outputs(2000) <= a;
    layer7_outputs(2001) <= a xor b;
    layer7_outputs(2002) <= a or b;
    layer7_outputs(2003) <= not a;
    layer7_outputs(2004) <= a xor b;
    layer7_outputs(2005) <= not b;
    layer7_outputs(2006) <= not (a or b);
    layer7_outputs(2007) <= a and not b;
    layer7_outputs(2008) <= b;
    layer7_outputs(2009) <= not a or b;
    layer7_outputs(2010) <= not (a and b);
    layer7_outputs(2011) <= a and not b;
    layer7_outputs(2012) <= not a or b;
    layer7_outputs(2013) <= b;
    layer7_outputs(2014) <= b and not a;
    layer7_outputs(2015) <= not b or a;
    layer7_outputs(2016) <= a or b;
    layer7_outputs(2017) <= b;
    layer7_outputs(2018) <= b;
    layer7_outputs(2019) <= b and not a;
    layer7_outputs(2020) <= a;
    layer7_outputs(2021) <= not a;
    layer7_outputs(2022) <= not b;
    layer7_outputs(2023) <= b;
    layer7_outputs(2024) <= not a or b;
    layer7_outputs(2025) <= a;
    layer7_outputs(2026) <= not a;
    layer7_outputs(2027) <= not b or a;
    layer7_outputs(2028) <= not b or a;
    layer7_outputs(2029) <= 1'b1;
    layer7_outputs(2030) <= a xor b;
    layer7_outputs(2031) <= a or b;
    layer7_outputs(2032) <= not b;
    layer7_outputs(2033) <= b;
    layer7_outputs(2034) <= not b;
    layer7_outputs(2035) <= not (a and b);
    layer7_outputs(2036) <= a and not b;
    layer7_outputs(2037) <= not (a and b);
    layer7_outputs(2038) <= not a;
    layer7_outputs(2039) <= b;
    layer7_outputs(2040) <= not (a xor b);
    layer7_outputs(2041) <= a;
    layer7_outputs(2042) <= not b;
    layer7_outputs(2043) <= not a or b;
    layer7_outputs(2044) <= a;
    layer7_outputs(2045) <= not a;
    layer7_outputs(2046) <= not b;
    layer7_outputs(2047) <= a;
    layer7_outputs(2048) <= not a or b;
    layer7_outputs(2049) <= a;
    layer7_outputs(2050) <= a xor b;
    layer7_outputs(2051) <= not (a and b);
    layer7_outputs(2052) <= b;
    layer7_outputs(2053) <= a and b;
    layer7_outputs(2054) <= a xor b;
    layer7_outputs(2055) <= a xor b;
    layer7_outputs(2056) <= b and not a;
    layer7_outputs(2057) <= a xor b;
    layer7_outputs(2058) <= b;
    layer7_outputs(2059) <= not (a xor b);
    layer7_outputs(2060) <= b;
    layer7_outputs(2061) <= not b or a;
    layer7_outputs(2062) <= not (a and b);
    layer7_outputs(2063) <= not b;
    layer7_outputs(2064) <= not (a xor b);
    layer7_outputs(2065) <= a or b;
    layer7_outputs(2066) <= a or b;
    layer7_outputs(2067) <= b;
    layer7_outputs(2068) <= a or b;
    layer7_outputs(2069) <= not (a or b);
    layer7_outputs(2070) <= b;
    layer7_outputs(2071) <= a xor b;
    layer7_outputs(2072) <= a;
    layer7_outputs(2073) <= b;
    layer7_outputs(2074) <= a and b;
    layer7_outputs(2075) <= a;
    layer7_outputs(2076) <= a;
    layer7_outputs(2077) <= 1'b0;
    layer7_outputs(2078) <= not a or b;
    layer7_outputs(2079) <= b;
    layer7_outputs(2080) <= not (a and b);
    layer7_outputs(2081) <= not a;
    layer7_outputs(2082) <= not a;
    layer7_outputs(2083) <= a and b;
    layer7_outputs(2084) <= b;
    layer7_outputs(2085) <= b and not a;
    layer7_outputs(2086) <= not b;
    layer7_outputs(2087) <= not b or a;
    layer7_outputs(2088) <= a and not b;
    layer7_outputs(2089) <= b;
    layer7_outputs(2090) <= not b;
    layer7_outputs(2091) <= not (a xor b);
    layer7_outputs(2092) <= a and not b;
    layer7_outputs(2093) <= b;
    layer7_outputs(2094) <= a or b;
    layer7_outputs(2095) <= not b or a;
    layer7_outputs(2096) <= not (a and b);
    layer7_outputs(2097) <= a and not b;
    layer7_outputs(2098) <= a or b;
    layer7_outputs(2099) <= not (a and b);
    layer7_outputs(2100) <= not a;
    layer7_outputs(2101) <= b and not a;
    layer7_outputs(2102) <= not (a or b);
    layer7_outputs(2103) <= not a;
    layer7_outputs(2104) <= a xor b;
    layer7_outputs(2105) <= a or b;
    layer7_outputs(2106) <= not b;
    layer7_outputs(2107) <= 1'b1;
    layer7_outputs(2108) <= a and not b;
    layer7_outputs(2109) <= a;
    layer7_outputs(2110) <= not (a xor b);
    layer7_outputs(2111) <= not a;
    layer7_outputs(2112) <= 1'b1;
    layer7_outputs(2113) <= a and not b;
    layer7_outputs(2114) <= b;
    layer7_outputs(2115) <= not b;
    layer7_outputs(2116) <= a xor b;
    layer7_outputs(2117) <= not b;
    layer7_outputs(2118) <= b;
    layer7_outputs(2119) <= not b or a;
    layer7_outputs(2120) <= b;
    layer7_outputs(2121) <= not b or a;
    layer7_outputs(2122) <= b;
    layer7_outputs(2123) <= not a or b;
    layer7_outputs(2124) <= not b;
    layer7_outputs(2125) <= b and not a;
    layer7_outputs(2126) <= not b or a;
    layer7_outputs(2127) <= b;
    layer7_outputs(2128) <= b;
    layer7_outputs(2129) <= b;
    layer7_outputs(2130) <= not b or a;
    layer7_outputs(2131) <= a;
    layer7_outputs(2132) <= a and b;
    layer7_outputs(2133) <= not b;
    layer7_outputs(2134) <= not a;
    layer7_outputs(2135) <= not (a xor b);
    layer7_outputs(2136) <= b;
    layer7_outputs(2137) <= a;
    layer7_outputs(2138) <= a xor b;
    layer7_outputs(2139) <= not a;
    layer7_outputs(2140) <= b;
    layer7_outputs(2141) <= not (a or b);
    layer7_outputs(2142) <= not a;
    layer7_outputs(2143) <= not a or b;
    layer7_outputs(2144) <= a;
    layer7_outputs(2145) <= not a;
    layer7_outputs(2146) <= a;
    layer7_outputs(2147) <= not (a xor b);
    layer7_outputs(2148) <= not b;
    layer7_outputs(2149) <= a and not b;
    layer7_outputs(2150) <= a;
    layer7_outputs(2151) <= a xor b;
    layer7_outputs(2152) <= b and not a;
    layer7_outputs(2153) <= not (a and b);
    layer7_outputs(2154) <= b;
    layer7_outputs(2155) <= not a or b;
    layer7_outputs(2156) <= not (a xor b);
    layer7_outputs(2157) <= not b;
    layer7_outputs(2158) <= b;
    layer7_outputs(2159) <= not b;
    layer7_outputs(2160) <= b;
    layer7_outputs(2161) <= not (a and b);
    layer7_outputs(2162) <= not a;
    layer7_outputs(2163) <= not a;
    layer7_outputs(2164) <= a and not b;
    layer7_outputs(2165) <= b;
    layer7_outputs(2166) <= not (a and b);
    layer7_outputs(2167) <= a;
    layer7_outputs(2168) <= not (a or b);
    layer7_outputs(2169) <= a;
    layer7_outputs(2170) <= not (a xor b);
    layer7_outputs(2171) <= not b;
    layer7_outputs(2172) <= not a or b;
    layer7_outputs(2173) <= not a;
    layer7_outputs(2174) <= not b or a;
    layer7_outputs(2175) <= a;
    layer7_outputs(2176) <= not b;
    layer7_outputs(2177) <= a and not b;
    layer7_outputs(2178) <= not b;
    layer7_outputs(2179) <= a xor b;
    layer7_outputs(2180) <= not (a and b);
    layer7_outputs(2181) <= a and b;
    layer7_outputs(2182) <= a and not b;
    layer7_outputs(2183) <= b and not a;
    layer7_outputs(2184) <= a and b;
    layer7_outputs(2185) <= a and b;
    layer7_outputs(2186) <= not a;
    layer7_outputs(2187) <= not a;
    layer7_outputs(2188) <= a xor b;
    layer7_outputs(2189) <= not a or b;
    layer7_outputs(2190) <= not a;
    layer7_outputs(2191) <= a;
    layer7_outputs(2192) <= a;
    layer7_outputs(2193) <= b and not a;
    layer7_outputs(2194) <= a;
    layer7_outputs(2195) <= not b;
    layer7_outputs(2196) <= a and not b;
    layer7_outputs(2197) <= not (a or b);
    layer7_outputs(2198) <= not (a xor b);
    layer7_outputs(2199) <= not (a and b);
    layer7_outputs(2200) <= a;
    layer7_outputs(2201) <= a xor b;
    layer7_outputs(2202) <= not a;
    layer7_outputs(2203) <= not (a and b);
    layer7_outputs(2204) <= a or b;
    layer7_outputs(2205) <= 1'b1;
    layer7_outputs(2206) <= not (a and b);
    layer7_outputs(2207) <= not (a xor b);
    layer7_outputs(2208) <= b;
    layer7_outputs(2209) <= not (a xor b);
    layer7_outputs(2210) <= not (a or b);
    layer7_outputs(2211) <= b and not a;
    layer7_outputs(2212) <= not a or b;
    layer7_outputs(2213) <= a and b;
    layer7_outputs(2214) <= not b or a;
    layer7_outputs(2215) <= not (a or b);
    layer7_outputs(2216) <= a xor b;
    layer7_outputs(2217) <= not (a or b);
    layer7_outputs(2218) <= a or b;
    layer7_outputs(2219) <= a or b;
    layer7_outputs(2220) <= not a;
    layer7_outputs(2221) <= b and not a;
    layer7_outputs(2222) <= a;
    layer7_outputs(2223) <= a;
    layer7_outputs(2224) <= not b;
    layer7_outputs(2225) <= not (a or b);
    layer7_outputs(2226) <= b;
    layer7_outputs(2227) <= a and b;
    layer7_outputs(2228) <= a;
    layer7_outputs(2229) <= not b;
    layer7_outputs(2230) <= b;
    layer7_outputs(2231) <= a and not b;
    layer7_outputs(2232) <= a and not b;
    layer7_outputs(2233) <= not (a xor b);
    layer7_outputs(2234) <= a and not b;
    layer7_outputs(2235) <= b and not a;
    layer7_outputs(2236) <= not (a or b);
    layer7_outputs(2237) <= b;
    layer7_outputs(2238) <= a and not b;
    layer7_outputs(2239) <= 1'b1;
    layer7_outputs(2240) <= not (a and b);
    layer7_outputs(2241) <= not a;
    layer7_outputs(2242) <= not a or b;
    layer7_outputs(2243) <= a and b;
    layer7_outputs(2244) <= not a or b;
    layer7_outputs(2245) <= a or b;
    layer7_outputs(2246) <= b;
    layer7_outputs(2247) <= not a or b;
    layer7_outputs(2248) <= not b;
    layer7_outputs(2249) <= not (a and b);
    layer7_outputs(2250) <= not (a and b);
    layer7_outputs(2251) <= b;
    layer7_outputs(2252) <= not (a xor b);
    layer7_outputs(2253) <= not a or b;
    layer7_outputs(2254) <= a;
    layer7_outputs(2255) <= b and not a;
    layer7_outputs(2256) <= not (a and b);
    layer7_outputs(2257) <= b;
    layer7_outputs(2258) <= b and not a;
    layer7_outputs(2259) <= not b or a;
    layer7_outputs(2260) <= a xor b;
    layer7_outputs(2261) <= a;
    layer7_outputs(2262) <= a or b;
    layer7_outputs(2263) <= not (a xor b);
    layer7_outputs(2264) <= b;
    layer7_outputs(2265) <= not (a and b);
    layer7_outputs(2266) <= not a;
    layer7_outputs(2267) <= not a;
    layer7_outputs(2268) <= b;
    layer7_outputs(2269) <= not a;
    layer7_outputs(2270) <= not (a or b);
    layer7_outputs(2271) <= not (a and b);
    layer7_outputs(2272) <= a or b;
    layer7_outputs(2273) <= a xor b;
    layer7_outputs(2274) <= 1'b0;
    layer7_outputs(2275) <= a;
    layer7_outputs(2276) <= b;
    layer7_outputs(2277) <= not (a xor b);
    layer7_outputs(2278) <= not b or a;
    layer7_outputs(2279) <= a xor b;
    layer7_outputs(2280) <= not (a xor b);
    layer7_outputs(2281) <= not (a xor b);
    layer7_outputs(2282) <= b;
    layer7_outputs(2283) <= b;
    layer7_outputs(2284) <= b;
    layer7_outputs(2285) <= not b;
    layer7_outputs(2286) <= a xor b;
    layer7_outputs(2287) <= b;
    layer7_outputs(2288) <= a;
    layer7_outputs(2289) <= a xor b;
    layer7_outputs(2290) <= 1'b1;
    layer7_outputs(2291) <= a xor b;
    layer7_outputs(2292) <= not b;
    layer7_outputs(2293) <= a;
    layer7_outputs(2294) <= not b;
    layer7_outputs(2295) <= b and not a;
    layer7_outputs(2296) <= b;
    layer7_outputs(2297) <= not (a xor b);
    layer7_outputs(2298) <= a xor b;
    layer7_outputs(2299) <= not b or a;
    layer7_outputs(2300) <= a xor b;
    layer7_outputs(2301) <= b;
    layer7_outputs(2302) <= b;
    layer7_outputs(2303) <= not (a xor b);
    layer7_outputs(2304) <= a or b;
    layer7_outputs(2305) <= not b;
    layer7_outputs(2306) <= not b;
    layer7_outputs(2307) <= b and not a;
    layer7_outputs(2308) <= not b;
    layer7_outputs(2309) <= b;
    layer7_outputs(2310) <= b;
    layer7_outputs(2311) <= b;
    layer7_outputs(2312) <= a;
    layer7_outputs(2313) <= a and not b;
    layer7_outputs(2314) <= a and not b;
    layer7_outputs(2315) <= a xor b;
    layer7_outputs(2316) <= a and not b;
    layer7_outputs(2317) <= not (a or b);
    layer7_outputs(2318) <= a and not b;
    layer7_outputs(2319) <= a;
    layer7_outputs(2320) <= a;
    layer7_outputs(2321) <= a xor b;
    layer7_outputs(2322) <= b;
    layer7_outputs(2323) <= not (a xor b);
    layer7_outputs(2324) <= a and b;
    layer7_outputs(2325) <= a and not b;
    layer7_outputs(2326) <= a or b;
    layer7_outputs(2327) <= a;
    layer7_outputs(2328) <= not (a and b);
    layer7_outputs(2329) <= a and b;
    layer7_outputs(2330) <= not a;
    layer7_outputs(2331) <= not a;
    layer7_outputs(2332) <= not b;
    layer7_outputs(2333) <= a;
    layer7_outputs(2334) <= not (a or b);
    layer7_outputs(2335) <= not (a xor b);
    layer7_outputs(2336) <= a or b;
    layer7_outputs(2337) <= not (a xor b);
    layer7_outputs(2338) <= not a;
    layer7_outputs(2339) <= a xor b;
    layer7_outputs(2340) <= not a or b;
    layer7_outputs(2341) <= not a;
    layer7_outputs(2342) <= b and not a;
    layer7_outputs(2343) <= a and not b;
    layer7_outputs(2344) <= not (a or b);
    layer7_outputs(2345) <= not a;
    layer7_outputs(2346) <= not (a or b);
    layer7_outputs(2347) <= not a;
    layer7_outputs(2348) <= not a or b;
    layer7_outputs(2349) <= a and b;
    layer7_outputs(2350) <= 1'b1;
    layer7_outputs(2351) <= not a;
    layer7_outputs(2352) <= not a;
    layer7_outputs(2353) <= not (a xor b);
    layer7_outputs(2354) <= not a or b;
    layer7_outputs(2355) <= not b;
    layer7_outputs(2356) <= a xor b;
    layer7_outputs(2357) <= not b;
    layer7_outputs(2358) <= a xor b;
    layer7_outputs(2359) <= not a or b;
    layer7_outputs(2360) <= a;
    layer7_outputs(2361) <= not b;
    layer7_outputs(2362) <= not b or a;
    layer7_outputs(2363) <= not a;
    layer7_outputs(2364) <= a;
    layer7_outputs(2365) <= not (a and b);
    layer7_outputs(2366) <= a xor b;
    layer7_outputs(2367) <= not b;
    layer7_outputs(2368) <= a;
    layer7_outputs(2369) <= not b or a;
    layer7_outputs(2370) <= a or b;
    layer7_outputs(2371) <= a and not b;
    layer7_outputs(2372) <= b and not a;
    layer7_outputs(2373) <= not (a or b);
    layer7_outputs(2374) <= a;
    layer7_outputs(2375) <= a and not b;
    layer7_outputs(2376) <= a;
    layer7_outputs(2377) <= not (a xor b);
    layer7_outputs(2378) <= a and b;
    layer7_outputs(2379) <= not a;
    layer7_outputs(2380) <= not b or a;
    layer7_outputs(2381) <= not (a or b);
    layer7_outputs(2382) <= not a;
    layer7_outputs(2383) <= b;
    layer7_outputs(2384) <= not (a or b);
    layer7_outputs(2385) <= a and b;
    layer7_outputs(2386) <= a xor b;
    layer7_outputs(2387) <= a;
    layer7_outputs(2388) <= a and not b;
    layer7_outputs(2389) <= not b;
    layer7_outputs(2390) <= not (a and b);
    layer7_outputs(2391) <= a and b;
    layer7_outputs(2392) <= a;
    layer7_outputs(2393) <= not (a or b);
    layer7_outputs(2394) <= not a;
    layer7_outputs(2395) <= b;
    layer7_outputs(2396) <= not (a xor b);
    layer7_outputs(2397) <= a and b;
    layer7_outputs(2398) <= not a;
    layer7_outputs(2399) <= not (a xor b);
    layer7_outputs(2400) <= a xor b;
    layer7_outputs(2401) <= a xor b;
    layer7_outputs(2402) <= not (a xor b);
    layer7_outputs(2403) <= not b or a;
    layer7_outputs(2404) <= b;
    layer7_outputs(2405) <= b;
    layer7_outputs(2406) <= not (a or b);
    layer7_outputs(2407) <= not b;
    layer7_outputs(2408) <= not a;
    layer7_outputs(2409) <= a;
    layer7_outputs(2410) <= not (a xor b);
    layer7_outputs(2411) <= a and not b;
    layer7_outputs(2412) <= not a;
    layer7_outputs(2413) <= not b;
    layer7_outputs(2414) <= a xor b;
    layer7_outputs(2415) <= not (a or b);
    layer7_outputs(2416) <= b and not a;
    layer7_outputs(2417) <= b and not a;
    layer7_outputs(2418) <= b;
    layer7_outputs(2419) <= not (a and b);
    layer7_outputs(2420) <= not b;
    layer7_outputs(2421) <= not a or b;
    layer7_outputs(2422) <= a xor b;
    layer7_outputs(2423) <= b and not a;
    layer7_outputs(2424) <= a xor b;
    layer7_outputs(2425) <= not (a xor b);
    layer7_outputs(2426) <= not a;
    layer7_outputs(2427) <= not (a or b);
    layer7_outputs(2428) <= a;
    layer7_outputs(2429) <= b;
    layer7_outputs(2430) <= a;
    layer7_outputs(2431) <= b;
    layer7_outputs(2432) <= a and b;
    layer7_outputs(2433) <= not a;
    layer7_outputs(2434) <= not b;
    layer7_outputs(2435) <= a or b;
    layer7_outputs(2436) <= b;
    layer7_outputs(2437) <= a;
    layer7_outputs(2438) <= b and not a;
    layer7_outputs(2439) <= not a;
    layer7_outputs(2440) <= a and b;
    layer7_outputs(2441) <= b;
    layer7_outputs(2442) <= a;
    layer7_outputs(2443) <= not b;
    layer7_outputs(2444) <= a and b;
    layer7_outputs(2445) <= not b;
    layer7_outputs(2446) <= b and not a;
    layer7_outputs(2447) <= not b;
    layer7_outputs(2448) <= b;
    layer7_outputs(2449) <= not b;
    layer7_outputs(2450) <= not a;
    layer7_outputs(2451) <= not b;
    layer7_outputs(2452) <= a;
    layer7_outputs(2453) <= not b;
    layer7_outputs(2454) <= not b or a;
    layer7_outputs(2455) <= a or b;
    layer7_outputs(2456) <= a and not b;
    layer7_outputs(2457) <= not a;
    layer7_outputs(2458) <= not a;
    layer7_outputs(2459) <= not a or b;
    layer7_outputs(2460) <= b and not a;
    layer7_outputs(2461) <= 1'b1;
    layer7_outputs(2462) <= b and not a;
    layer7_outputs(2463) <= not a or b;
    layer7_outputs(2464) <= not a or b;
    layer7_outputs(2465) <= a;
    layer7_outputs(2466) <= a and b;
    layer7_outputs(2467) <= not b or a;
    layer7_outputs(2468) <= not (a or b);
    layer7_outputs(2469) <= not a;
    layer7_outputs(2470) <= not a;
    layer7_outputs(2471) <= not a;
    layer7_outputs(2472) <= not b;
    layer7_outputs(2473) <= a or b;
    layer7_outputs(2474) <= b;
    layer7_outputs(2475) <= b and not a;
    layer7_outputs(2476) <= b;
    layer7_outputs(2477) <= b;
    layer7_outputs(2478) <= a and b;
    layer7_outputs(2479) <= not a;
    layer7_outputs(2480) <= b;
    layer7_outputs(2481) <= not a or b;
    layer7_outputs(2482) <= a;
    layer7_outputs(2483) <= a xor b;
    layer7_outputs(2484) <= not a;
    layer7_outputs(2485) <= 1'b1;
    layer7_outputs(2486) <= a xor b;
    layer7_outputs(2487) <= not a or b;
    layer7_outputs(2488) <= b;
    layer7_outputs(2489) <= a;
    layer7_outputs(2490) <= 1'b0;
    layer7_outputs(2491) <= a and not b;
    layer7_outputs(2492) <= b;
    layer7_outputs(2493) <= a xor b;
    layer7_outputs(2494) <= not a or b;
    layer7_outputs(2495) <= a or b;
    layer7_outputs(2496) <= not a;
    layer7_outputs(2497) <= b and not a;
    layer7_outputs(2498) <= a xor b;
    layer7_outputs(2499) <= not b;
    layer7_outputs(2500) <= a or b;
    layer7_outputs(2501) <= not a or b;
    layer7_outputs(2502) <= a and b;
    layer7_outputs(2503) <= not b;
    layer7_outputs(2504) <= a xor b;
    layer7_outputs(2505) <= not b;
    layer7_outputs(2506) <= not b;
    layer7_outputs(2507) <= not a;
    layer7_outputs(2508) <= not a;
    layer7_outputs(2509) <= b;
    layer7_outputs(2510) <= a xor b;
    layer7_outputs(2511) <= 1'b0;
    layer7_outputs(2512) <= b;
    layer7_outputs(2513) <= a or b;
    layer7_outputs(2514) <= b;
    layer7_outputs(2515) <= not a;
    layer7_outputs(2516) <= a xor b;
    layer7_outputs(2517) <= not b;
    layer7_outputs(2518) <= b;
    layer7_outputs(2519) <= b;
    layer7_outputs(2520) <= a;
    layer7_outputs(2521) <= not b;
    layer7_outputs(2522) <= not b;
    layer7_outputs(2523) <= not (a and b);
    layer7_outputs(2524) <= not a;
    layer7_outputs(2525) <= not a or b;
    layer7_outputs(2526) <= a and not b;
    layer7_outputs(2527) <= a;
    layer7_outputs(2528) <= not a or b;
    layer7_outputs(2529) <= not b;
    layer7_outputs(2530) <= b;
    layer7_outputs(2531) <= a;
    layer7_outputs(2532) <= a xor b;
    layer7_outputs(2533) <= b;
    layer7_outputs(2534) <= not a;
    layer7_outputs(2535) <= not (a xor b);
    layer7_outputs(2536) <= 1'b1;
    layer7_outputs(2537) <= a and not b;
    layer7_outputs(2538) <= not a;
    layer7_outputs(2539) <= not b;
    layer7_outputs(2540) <= a;
    layer7_outputs(2541) <= a;
    layer7_outputs(2542) <= b and not a;
    layer7_outputs(2543) <= not a;
    layer7_outputs(2544) <= a;
    layer7_outputs(2545) <= not a;
    layer7_outputs(2546) <= not b;
    layer7_outputs(2547) <= a and not b;
    layer7_outputs(2548) <= a and not b;
    layer7_outputs(2549) <= not (a xor b);
    layer7_outputs(2550) <= not a or b;
    layer7_outputs(2551) <= not a or b;
    layer7_outputs(2552) <= a;
    layer7_outputs(2553) <= a xor b;
    layer7_outputs(2554) <= a or b;
    layer7_outputs(2555) <= a;
    layer7_outputs(2556) <= b;
    layer7_outputs(2557) <= not (a and b);
    layer7_outputs(2558) <= not (a xor b);
    layer7_outputs(2559) <= not (a xor b);
    layer7_outputs(2560) <= a xor b;
    layer7_outputs(2561) <= a;
    layer7_outputs(2562) <= not b or a;
    layer7_outputs(2563) <= not a;
    layer7_outputs(2564) <= not b;
    layer7_outputs(2565) <= b;
    layer7_outputs(2566) <= not (a xor b);
    layer7_outputs(2567) <= a;
    layer7_outputs(2568) <= b and not a;
    layer7_outputs(2569) <= not a;
    layer7_outputs(2570) <= a;
    layer7_outputs(2571) <= a or b;
    layer7_outputs(2572) <= not b;
    layer7_outputs(2573) <= a;
    layer7_outputs(2574) <= a;
    layer7_outputs(2575) <= not (a or b);
    layer7_outputs(2576) <= not a or b;
    layer7_outputs(2577) <= not a;
    layer7_outputs(2578) <= not (a xor b);
    layer7_outputs(2579) <= a xor b;
    layer7_outputs(2580) <= a or b;
    layer7_outputs(2581) <= not a;
    layer7_outputs(2582) <= a and not b;
    layer7_outputs(2583) <= a and not b;
    layer7_outputs(2584) <= b and not a;
    layer7_outputs(2585) <= not b;
    layer7_outputs(2586) <= a and b;
    layer7_outputs(2587) <= a or b;
    layer7_outputs(2588) <= a and b;
    layer7_outputs(2589) <= b;
    layer7_outputs(2590) <= not b;
    layer7_outputs(2591) <= 1'b1;
    layer7_outputs(2592) <= a and b;
    layer7_outputs(2593) <= not b or a;
    layer7_outputs(2594) <= not b;
    layer7_outputs(2595) <= a xor b;
    layer7_outputs(2596) <= b and not a;
    layer7_outputs(2597) <= not (a or b);
    layer7_outputs(2598) <= not a;
    layer7_outputs(2599) <= b;
    layer7_outputs(2600) <= not a or b;
    layer7_outputs(2601) <= a;
    layer7_outputs(2602) <= a xor b;
    layer7_outputs(2603) <= not a;
    layer7_outputs(2604) <= a;
    layer7_outputs(2605) <= b and not a;
    layer7_outputs(2606) <= not b;
    layer7_outputs(2607) <= b;
    layer7_outputs(2608) <= not a;
    layer7_outputs(2609) <= not (a and b);
    layer7_outputs(2610) <= not b;
    layer7_outputs(2611) <= not (a xor b);
    layer7_outputs(2612) <= not (a xor b);
    layer7_outputs(2613) <= a;
    layer7_outputs(2614) <= a or b;
    layer7_outputs(2615) <= not (a or b);
    layer7_outputs(2616) <= a and b;
    layer7_outputs(2617) <= not a or b;
    layer7_outputs(2618) <= not (a xor b);
    layer7_outputs(2619) <= not a;
    layer7_outputs(2620) <= not b;
    layer7_outputs(2621) <= a;
    layer7_outputs(2622) <= a or b;
    layer7_outputs(2623) <= not a or b;
    layer7_outputs(2624) <= not a;
    layer7_outputs(2625) <= 1'b0;
    layer7_outputs(2626) <= not b;
    layer7_outputs(2627) <= not b;
    layer7_outputs(2628) <= not a;
    layer7_outputs(2629) <= a;
    layer7_outputs(2630) <= b;
    layer7_outputs(2631) <= not a;
    layer7_outputs(2632) <= not b or a;
    layer7_outputs(2633) <= not a;
    layer7_outputs(2634) <= not a;
    layer7_outputs(2635) <= 1'b1;
    layer7_outputs(2636) <= b;
    layer7_outputs(2637) <= not a or b;
    layer7_outputs(2638) <= b and not a;
    layer7_outputs(2639) <= b;
    layer7_outputs(2640) <= b;
    layer7_outputs(2641) <= a xor b;
    layer7_outputs(2642) <= not b;
    layer7_outputs(2643) <= not (a or b);
    layer7_outputs(2644) <= a xor b;
    layer7_outputs(2645) <= not a;
    layer7_outputs(2646) <= not a;
    layer7_outputs(2647) <= b;
    layer7_outputs(2648) <= a;
    layer7_outputs(2649) <= a or b;
    layer7_outputs(2650) <= not b;
    layer7_outputs(2651) <= a xor b;
    layer7_outputs(2652) <= not a;
    layer7_outputs(2653) <= a and not b;
    layer7_outputs(2654) <= not b or a;
    layer7_outputs(2655) <= not (a xor b);
    layer7_outputs(2656) <= not a;
    layer7_outputs(2657) <= a or b;
    layer7_outputs(2658) <= not b;
    layer7_outputs(2659) <= not b;
    layer7_outputs(2660) <= not b;
    layer7_outputs(2661) <= not (a xor b);
    layer7_outputs(2662) <= not (a and b);
    layer7_outputs(2663) <= not (a or b);
    layer7_outputs(2664) <= a xor b;
    layer7_outputs(2665) <= b;
    layer7_outputs(2666) <= not b;
    layer7_outputs(2667) <= not a;
    layer7_outputs(2668) <= not (a xor b);
    layer7_outputs(2669) <= b;
    layer7_outputs(2670) <= a;
    layer7_outputs(2671) <= a and b;
    layer7_outputs(2672) <= a and not b;
    layer7_outputs(2673) <= not (a xor b);
    layer7_outputs(2674) <= b;
    layer7_outputs(2675) <= not (a xor b);
    layer7_outputs(2676) <= not a;
    layer7_outputs(2677) <= b;
    layer7_outputs(2678) <= not a;
    layer7_outputs(2679) <= not (a xor b);
    layer7_outputs(2680) <= a;
    layer7_outputs(2681) <= not a or b;
    layer7_outputs(2682) <= b;
    layer7_outputs(2683) <= not (a and b);
    layer7_outputs(2684) <= not b;
    layer7_outputs(2685) <= not a;
    layer7_outputs(2686) <= not a;
    layer7_outputs(2687) <= not a or b;
    layer7_outputs(2688) <= a;
    layer7_outputs(2689) <= a xor b;
    layer7_outputs(2690) <= a xor b;
    layer7_outputs(2691) <= not a;
    layer7_outputs(2692) <= b;
    layer7_outputs(2693) <= not b;
    layer7_outputs(2694) <= b;
    layer7_outputs(2695) <= not a;
    layer7_outputs(2696) <= 1'b0;
    layer7_outputs(2697) <= a;
    layer7_outputs(2698) <= b;
    layer7_outputs(2699) <= not (a xor b);
    layer7_outputs(2700) <= b;
    layer7_outputs(2701) <= a;
    layer7_outputs(2702) <= b;
    layer7_outputs(2703) <= b;
    layer7_outputs(2704) <= b;
    layer7_outputs(2705) <= not b or a;
    layer7_outputs(2706) <= not b;
    layer7_outputs(2707) <= not a;
    layer7_outputs(2708) <= not a or b;
    layer7_outputs(2709) <= not (a and b);
    layer7_outputs(2710) <= a;
    layer7_outputs(2711) <= a and not b;
    layer7_outputs(2712) <= not (a xor b);
    layer7_outputs(2713) <= not a;
    layer7_outputs(2714) <= a;
    layer7_outputs(2715) <= a xor b;
    layer7_outputs(2716) <= a;
    layer7_outputs(2717) <= b;
    layer7_outputs(2718) <= a;
    layer7_outputs(2719) <= b and not a;
    layer7_outputs(2720) <= a or b;
    layer7_outputs(2721) <= b and not a;
    layer7_outputs(2722) <= b and not a;
    layer7_outputs(2723) <= a xor b;
    layer7_outputs(2724) <= 1'b1;
    layer7_outputs(2725) <= not (a xor b);
    layer7_outputs(2726) <= not (a or b);
    layer7_outputs(2727) <= b;
    layer7_outputs(2728) <= not (a xor b);
    layer7_outputs(2729) <= b and not a;
    layer7_outputs(2730) <= not (a or b);
    layer7_outputs(2731) <= b;
    layer7_outputs(2732) <= 1'b1;
    layer7_outputs(2733) <= b;
    layer7_outputs(2734) <= not b or a;
    layer7_outputs(2735) <= not a;
    layer7_outputs(2736) <= a and not b;
    layer7_outputs(2737) <= a;
    layer7_outputs(2738) <= a xor b;
    layer7_outputs(2739) <= b;
    layer7_outputs(2740) <= 1'b1;
    layer7_outputs(2741) <= not (a xor b);
    layer7_outputs(2742) <= a or b;
    layer7_outputs(2743) <= not (a or b);
    layer7_outputs(2744) <= b;
    layer7_outputs(2745) <= not (a xor b);
    layer7_outputs(2746) <= not (a or b);
    layer7_outputs(2747) <= a;
    layer7_outputs(2748) <= not b;
    layer7_outputs(2749) <= not (a xor b);
    layer7_outputs(2750) <= not (a xor b);
    layer7_outputs(2751) <= a and not b;
    layer7_outputs(2752) <= a and b;
    layer7_outputs(2753) <= b;
    layer7_outputs(2754) <= a and b;
    layer7_outputs(2755) <= not a;
    layer7_outputs(2756) <= not a;
    layer7_outputs(2757) <= not a or b;
    layer7_outputs(2758) <= a;
    layer7_outputs(2759) <= not a;
    layer7_outputs(2760) <= b;
    layer7_outputs(2761) <= not b;
    layer7_outputs(2762) <= a;
    layer7_outputs(2763) <= a and b;
    layer7_outputs(2764) <= not b;
    layer7_outputs(2765) <= not (a or b);
    layer7_outputs(2766) <= not a;
    layer7_outputs(2767) <= a or b;
    layer7_outputs(2768) <= not a;
    layer7_outputs(2769) <= a;
    layer7_outputs(2770) <= not (a or b);
    layer7_outputs(2771) <= not (a xor b);
    layer7_outputs(2772) <= a xor b;
    layer7_outputs(2773) <= not b;
    layer7_outputs(2774) <= not (a xor b);
    layer7_outputs(2775) <= b;
    layer7_outputs(2776) <= a and not b;
    layer7_outputs(2777) <= not (a and b);
    layer7_outputs(2778) <= not (a xor b);
    layer7_outputs(2779) <= a;
    layer7_outputs(2780) <= b;
    layer7_outputs(2781) <= a;
    layer7_outputs(2782) <= not b or a;
    layer7_outputs(2783) <= not (a or b);
    layer7_outputs(2784) <= a;
    layer7_outputs(2785) <= b;
    layer7_outputs(2786) <= a xor b;
    layer7_outputs(2787) <= not b;
    layer7_outputs(2788) <= not (a or b);
    layer7_outputs(2789) <= not a;
    layer7_outputs(2790) <= not a;
    layer7_outputs(2791) <= b;
    layer7_outputs(2792) <= a;
    layer7_outputs(2793) <= not b;
    layer7_outputs(2794) <= not a or b;
    layer7_outputs(2795) <= a and not b;
    layer7_outputs(2796) <= not a;
    layer7_outputs(2797) <= a and b;
    layer7_outputs(2798) <= a xor b;
    layer7_outputs(2799) <= not b;
    layer7_outputs(2800) <= not (a or b);
    layer7_outputs(2801) <= b;
    layer7_outputs(2802) <= 1'b0;
    layer7_outputs(2803) <= b;
    layer7_outputs(2804) <= not a or b;
    layer7_outputs(2805) <= not (a and b);
    layer7_outputs(2806) <= not a;
    layer7_outputs(2807) <= not b or a;
    layer7_outputs(2808) <= b and not a;
    layer7_outputs(2809) <= not a or b;
    layer7_outputs(2810) <= not (a xor b);
    layer7_outputs(2811) <= a xor b;
    layer7_outputs(2812) <= not a;
    layer7_outputs(2813) <= not a or b;
    layer7_outputs(2814) <= a or b;
    layer7_outputs(2815) <= a and not b;
    layer7_outputs(2816) <= a;
    layer7_outputs(2817) <= a;
    layer7_outputs(2818) <= b;
    layer7_outputs(2819) <= b;
    layer7_outputs(2820) <= b;
    layer7_outputs(2821) <= not a;
    layer7_outputs(2822) <= not a;
    layer7_outputs(2823) <= a and b;
    layer7_outputs(2824) <= not (a xor b);
    layer7_outputs(2825) <= a xor b;
    layer7_outputs(2826) <= not a or b;
    layer7_outputs(2827) <= a and b;
    layer7_outputs(2828) <= b and not a;
    layer7_outputs(2829) <= not (a xor b);
    layer7_outputs(2830) <= b;
    layer7_outputs(2831) <= not a;
    layer7_outputs(2832) <= not b;
    layer7_outputs(2833) <= a and b;
    layer7_outputs(2834) <= a and b;
    layer7_outputs(2835) <= a or b;
    layer7_outputs(2836) <= not (a xor b);
    layer7_outputs(2837) <= not a;
    layer7_outputs(2838) <= a and b;
    layer7_outputs(2839) <= b and not a;
    layer7_outputs(2840) <= b and not a;
    layer7_outputs(2841) <= not b;
    layer7_outputs(2842) <= a and not b;
    layer7_outputs(2843) <= a or b;
    layer7_outputs(2844) <= b and not a;
    layer7_outputs(2845) <= b;
    layer7_outputs(2846) <= a and not b;
    layer7_outputs(2847) <= not (a or b);
    layer7_outputs(2848) <= not b;
    layer7_outputs(2849) <= not b;
    layer7_outputs(2850) <= not b;
    layer7_outputs(2851) <= not (a xor b);
    layer7_outputs(2852) <= b;
    layer7_outputs(2853) <= a xor b;
    layer7_outputs(2854) <= not a;
    layer7_outputs(2855) <= a and b;
    layer7_outputs(2856) <= not (a and b);
    layer7_outputs(2857) <= a;
    layer7_outputs(2858) <= b;
    layer7_outputs(2859) <= not (a xor b);
    layer7_outputs(2860) <= not b or a;
    layer7_outputs(2861) <= a and b;
    layer7_outputs(2862) <= 1'b0;
    layer7_outputs(2863) <= not b;
    layer7_outputs(2864) <= b and not a;
    layer7_outputs(2865) <= not (a xor b);
    layer7_outputs(2866) <= not b;
    layer7_outputs(2867) <= a xor b;
    layer7_outputs(2868) <= not (a or b);
    layer7_outputs(2869) <= b and not a;
    layer7_outputs(2870) <= a and b;
    layer7_outputs(2871) <= a or b;
    layer7_outputs(2872) <= a or b;
    layer7_outputs(2873) <= 1'b0;
    layer7_outputs(2874) <= a xor b;
    layer7_outputs(2875) <= a and b;
    layer7_outputs(2876) <= not b;
    layer7_outputs(2877) <= not a;
    layer7_outputs(2878) <= a;
    layer7_outputs(2879) <= a;
    layer7_outputs(2880) <= a xor b;
    layer7_outputs(2881) <= not (a and b);
    layer7_outputs(2882) <= a;
    layer7_outputs(2883) <= not (a or b);
    layer7_outputs(2884) <= not (a xor b);
    layer7_outputs(2885) <= a;
    layer7_outputs(2886) <= b and not a;
    layer7_outputs(2887) <= not (a xor b);
    layer7_outputs(2888) <= b;
    layer7_outputs(2889) <= a xor b;
    layer7_outputs(2890) <= b;
    layer7_outputs(2891) <= a or b;
    layer7_outputs(2892) <= a;
    layer7_outputs(2893) <= not b or a;
    layer7_outputs(2894) <= not a;
    layer7_outputs(2895) <= not b or a;
    layer7_outputs(2896) <= a;
    layer7_outputs(2897) <= not b or a;
    layer7_outputs(2898) <= not (a or b);
    layer7_outputs(2899) <= not a or b;
    layer7_outputs(2900) <= not a or b;
    layer7_outputs(2901) <= a or b;
    layer7_outputs(2902) <= not (a xor b);
    layer7_outputs(2903) <= a xor b;
    layer7_outputs(2904) <= 1'b0;
    layer7_outputs(2905) <= not a or b;
    layer7_outputs(2906) <= a and not b;
    layer7_outputs(2907) <= not (a or b);
    layer7_outputs(2908) <= a;
    layer7_outputs(2909) <= a xor b;
    layer7_outputs(2910) <= b;
    layer7_outputs(2911) <= a and not b;
    layer7_outputs(2912) <= a;
    layer7_outputs(2913) <= not a;
    layer7_outputs(2914) <= a xor b;
    layer7_outputs(2915) <= not (a xor b);
    layer7_outputs(2916) <= not b;
    layer7_outputs(2917) <= not a;
    layer7_outputs(2918) <= a xor b;
    layer7_outputs(2919) <= not b;
    layer7_outputs(2920) <= a;
    layer7_outputs(2921) <= b;
    layer7_outputs(2922) <= 1'b1;
    layer7_outputs(2923) <= not b;
    layer7_outputs(2924) <= not b;
    layer7_outputs(2925) <= a and b;
    layer7_outputs(2926) <= a xor b;
    layer7_outputs(2927) <= a and b;
    layer7_outputs(2928) <= not (a or b);
    layer7_outputs(2929) <= a and b;
    layer7_outputs(2930) <= a;
    layer7_outputs(2931) <= not a;
    layer7_outputs(2932) <= not a;
    layer7_outputs(2933) <= not (a xor b);
    layer7_outputs(2934) <= not (a xor b);
    layer7_outputs(2935) <= not b or a;
    layer7_outputs(2936) <= not b;
    layer7_outputs(2937) <= a;
    layer7_outputs(2938) <= a and b;
    layer7_outputs(2939) <= not a or b;
    layer7_outputs(2940) <= not a;
    layer7_outputs(2941) <= a and b;
    layer7_outputs(2942) <= not (a or b);
    layer7_outputs(2943) <= a and not b;
    layer7_outputs(2944) <= not a or b;
    layer7_outputs(2945) <= a and b;
    layer7_outputs(2946) <= a and not b;
    layer7_outputs(2947) <= not a or b;
    layer7_outputs(2948) <= not a or b;
    layer7_outputs(2949) <= b;
    layer7_outputs(2950) <= not (a xor b);
    layer7_outputs(2951) <= not (a and b);
    layer7_outputs(2952) <= a xor b;
    layer7_outputs(2953) <= not a;
    layer7_outputs(2954) <= b;
    layer7_outputs(2955) <= not a or b;
    layer7_outputs(2956) <= a or b;
    layer7_outputs(2957) <= not (a xor b);
    layer7_outputs(2958) <= a xor b;
    layer7_outputs(2959) <= a;
    layer7_outputs(2960) <= not (a and b);
    layer7_outputs(2961) <= a;
    layer7_outputs(2962) <= b;
    layer7_outputs(2963) <= not a;
    layer7_outputs(2964) <= not b;
    layer7_outputs(2965) <= a and b;
    layer7_outputs(2966) <= a;
    layer7_outputs(2967) <= not a;
    layer7_outputs(2968) <= not a;
    layer7_outputs(2969) <= a or b;
    layer7_outputs(2970) <= not b;
    layer7_outputs(2971) <= a and b;
    layer7_outputs(2972) <= not b;
    layer7_outputs(2973) <= a or b;
    layer7_outputs(2974) <= not a;
    layer7_outputs(2975) <= b and not a;
    layer7_outputs(2976) <= not a;
    layer7_outputs(2977) <= not b;
    layer7_outputs(2978) <= b and not a;
    layer7_outputs(2979) <= b;
    layer7_outputs(2980) <= a;
    layer7_outputs(2981) <= not (a xor b);
    layer7_outputs(2982) <= b and not a;
    layer7_outputs(2983) <= a;
    layer7_outputs(2984) <= a xor b;
    layer7_outputs(2985) <= a;
    layer7_outputs(2986) <= a xor b;
    layer7_outputs(2987) <= not b;
    layer7_outputs(2988) <= not b;
    layer7_outputs(2989) <= b;
    layer7_outputs(2990) <= b;
    layer7_outputs(2991) <= not a or b;
    layer7_outputs(2992) <= b and not a;
    layer7_outputs(2993) <= b and not a;
    layer7_outputs(2994) <= not a;
    layer7_outputs(2995) <= not a;
    layer7_outputs(2996) <= a xor b;
    layer7_outputs(2997) <= not (a xor b);
    layer7_outputs(2998) <= a;
    layer7_outputs(2999) <= not (a xor b);
    layer7_outputs(3000) <= not (a xor b);
    layer7_outputs(3001) <= a xor b;
    layer7_outputs(3002) <= a;
    layer7_outputs(3003) <= not a;
    layer7_outputs(3004) <= b;
    layer7_outputs(3005) <= 1'b0;
    layer7_outputs(3006) <= b;
    layer7_outputs(3007) <= a and b;
    layer7_outputs(3008) <= a xor b;
    layer7_outputs(3009) <= b and not a;
    layer7_outputs(3010) <= not (a and b);
    layer7_outputs(3011) <= b;
    layer7_outputs(3012) <= not b;
    layer7_outputs(3013) <= not (a and b);
    layer7_outputs(3014) <= not b;
    layer7_outputs(3015) <= b and not a;
    layer7_outputs(3016) <= a xor b;
    layer7_outputs(3017) <= a;
    layer7_outputs(3018) <= b and not a;
    layer7_outputs(3019) <= not (a xor b);
    layer7_outputs(3020) <= not b;
    layer7_outputs(3021) <= not (a and b);
    layer7_outputs(3022) <= a and not b;
    layer7_outputs(3023) <= a;
    layer7_outputs(3024) <= not (a xor b);
    layer7_outputs(3025) <= a;
    layer7_outputs(3026) <= a;
    layer7_outputs(3027) <= a;
    layer7_outputs(3028) <= a and not b;
    layer7_outputs(3029) <= a and not b;
    layer7_outputs(3030) <= 1'b0;
    layer7_outputs(3031) <= a;
    layer7_outputs(3032) <= 1'b0;
    layer7_outputs(3033) <= not a;
    layer7_outputs(3034) <= not b or a;
    layer7_outputs(3035) <= a;
    layer7_outputs(3036) <= not b;
    layer7_outputs(3037) <= not (a and b);
    layer7_outputs(3038) <= a xor b;
    layer7_outputs(3039) <= b and not a;
    layer7_outputs(3040) <= a;
    layer7_outputs(3041) <= not (a or b);
    layer7_outputs(3042) <= b;
    layer7_outputs(3043) <= not (a and b);
    layer7_outputs(3044) <= not a;
    layer7_outputs(3045) <= a and b;
    layer7_outputs(3046) <= not (a xor b);
    layer7_outputs(3047) <= not (a xor b);
    layer7_outputs(3048) <= not b;
    layer7_outputs(3049) <= not (a xor b);
    layer7_outputs(3050) <= not (a xor b);
    layer7_outputs(3051) <= not (a xor b);
    layer7_outputs(3052) <= a and b;
    layer7_outputs(3053) <= not a;
    layer7_outputs(3054) <= a xor b;
    layer7_outputs(3055) <= a and b;
    layer7_outputs(3056) <= b and not a;
    layer7_outputs(3057) <= not (a xor b);
    layer7_outputs(3058) <= not (a and b);
    layer7_outputs(3059) <= a xor b;
    layer7_outputs(3060) <= not b;
    layer7_outputs(3061) <= a;
    layer7_outputs(3062) <= not a;
    layer7_outputs(3063) <= not a;
    layer7_outputs(3064) <= a;
    layer7_outputs(3065) <= not b;
    layer7_outputs(3066) <= a xor b;
    layer7_outputs(3067) <= not b;
    layer7_outputs(3068) <= not a;
    layer7_outputs(3069) <= not (a xor b);
    layer7_outputs(3070) <= not a or b;
    layer7_outputs(3071) <= a;
    layer7_outputs(3072) <= not b;
    layer7_outputs(3073) <= b;
    layer7_outputs(3074) <= a and not b;
    layer7_outputs(3075) <= not (a and b);
    layer7_outputs(3076) <= not b;
    layer7_outputs(3077) <= a;
    layer7_outputs(3078) <= b and not a;
    layer7_outputs(3079) <= a or b;
    layer7_outputs(3080) <= a or b;
    layer7_outputs(3081) <= b and not a;
    layer7_outputs(3082) <= a;
    layer7_outputs(3083) <= a xor b;
    layer7_outputs(3084) <= not a or b;
    layer7_outputs(3085) <= a and not b;
    layer7_outputs(3086) <= not (a xor b);
    layer7_outputs(3087) <= not (a or b);
    layer7_outputs(3088) <= not (a xor b);
    layer7_outputs(3089) <= not b;
    layer7_outputs(3090) <= a and not b;
    layer7_outputs(3091) <= b;
    layer7_outputs(3092) <= a xor b;
    layer7_outputs(3093) <= not b;
    layer7_outputs(3094) <= not a;
    layer7_outputs(3095) <= not (a xor b);
    layer7_outputs(3096) <= a or b;
    layer7_outputs(3097) <= not (a xor b);
    layer7_outputs(3098) <= a and b;
    layer7_outputs(3099) <= b;
    layer7_outputs(3100) <= a and b;
    layer7_outputs(3101) <= b;
    layer7_outputs(3102) <= not b or a;
    layer7_outputs(3103) <= not b;
    layer7_outputs(3104) <= b;
    layer7_outputs(3105) <= b and not a;
    layer7_outputs(3106) <= b and not a;
    layer7_outputs(3107) <= b;
    layer7_outputs(3108) <= not a;
    layer7_outputs(3109) <= b;
    layer7_outputs(3110) <= not b or a;
    layer7_outputs(3111) <= a xor b;
    layer7_outputs(3112) <= not (a or b);
    layer7_outputs(3113) <= not a;
    layer7_outputs(3114) <= not b;
    layer7_outputs(3115) <= not b;
    layer7_outputs(3116) <= not a;
    layer7_outputs(3117) <= a;
    layer7_outputs(3118) <= b;
    layer7_outputs(3119) <= a xor b;
    layer7_outputs(3120) <= b;
    layer7_outputs(3121) <= not (a xor b);
    layer7_outputs(3122) <= a;
    layer7_outputs(3123) <= b;
    layer7_outputs(3124) <= 1'b0;
    layer7_outputs(3125) <= a;
    layer7_outputs(3126) <= a and b;
    layer7_outputs(3127) <= not (a and b);
    layer7_outputs(3128) <= 1'b0;
    layer7_outputs(3129) <= not b;
    layer7_outputs(3130) <= a;
    layer7_outputs(3131) <= not (a or b);
    layer7_outputs(3132) <= not a;
    layer7_outputs(3133) <= not b;
    layer7_outputs(3134) <= not (a or b);
    layer7_outputs(3135) <= 1'b1;
    layer7_outputs(3136) <= not b or a;
    layer7_outputs(3137) <= not b;
    layer7_outputs(3138) <= b and not a;
    layer7_outputs(3139) <= not a or b;
    layer7_outputs(3140) <= not (a or b);
    layer7_outputs(3141) <= b;
    layer7_outputs(3142) <= not (a and b);
    layer7_outputs(3143) <= b;
    layer7_outputs(3144) <= b and not a;
    layer7_outputs(3145) <= not a or b;
    layer7_outputs(3146) <= not b;
    layer7_outputs(3147) <= not (a and b);
    layer7_outputs(3148) <= a xor b;
    layer7_outputs(3149) <= not (a or b);
    layer7_outputs(3150) <= b;
    layer7_outputs(3151) <= not b;
    layer7_outputs(3152) <= not a or b;
    layer7_outputs(3153) <= not b;
    layer7_outputs(3154) <= b;
    layer7_outputs(3155) <= not b;
    layer7_outputs(3156) <= not (a xor b);
    layer7_outputs(3157) <= a and not b;
    layer7_outputs(3158) <= a xor b;
    layer7_outputs(3159) <= not b;
    layer7_outputs(3160) <= not b or a;
    layer7_outputs(3161) <= a and b;
    layer7_outputs(3162) <= not a;
    layer7_outputs(3163) <= not b;
    layer7_outputs(3164) <= 1'b0;
    layer7_outputs(3165) <= a;
    layer7_outputs(3166) <= a;
    layer7_outputs(3167) <= a and not b;
    layer7_outputs(3168) <= b;
    layer7_outputs(3169) <= b;
    layer7_outputs(3170) <= not b;
    layer7_outputs(3171) <= not (a or b);
    layer7_outputs(3172) <= not a;
    layer7_outputs(3173) <= not a;
    layer7_outputs(3174) <= not a;
    layer7_outputs(3175) <= b;
    layer7_outputs(3176) <= a;
    layer7_outputs(3177) <= 1'b1;
    layer7_outputs(3178) <= b and not a;
    layer7_outputs(3179) <= b;
    layer7_outputs(3180) <= b;
    layer7_outputs(3181) <= not b;
    layer7_outputs(3182) <= a or b;
    layer7_outputs(3183) <= a or b;
    layer7_outputs(3184) <= not b;
    layer7_outputs(3185) <= not (a xor b);
    layer7_outputs(3186) <= a xor b;
    layer7_outputs(3187) <= a xor b;
    layer7_outputs(3188) <= a xor b;
    layer7_outputs(3189) <= not a;
    layer7_outputs(3190) <= not (a or b);
    layer7_outputs(3191) <= not b;
    layer7_outputs(3192) <= a;
    layer7_outputs(3193) <= not b or a;
    layer7_outputs(3194) <= not (a or b);
    layer7_outputs(3195) <= not (a or b);
    layer7_outputs(3196) <= not (a or b);
    layer7_outputs(3197) <= not (a xor b);
    layer7_outputs(3198) <= b;
    layer7_outputs(3199) <= not (a or b);
    layer7_outputs(3200) <= not b;
    layer7_outputs(3201) <= a;
    layer7_outputs(3202) <= b and not a;
    layer7_outputs(3203) <= a or b;
    layer7_outputs(3204) <= b;
    layer7_outputs(3205) <= a and not b;
    layer7_outputs(3206) <= a and b;
    layer7_outputs(3207) <= b;
    layer7_outputs(3208) <= a;
    layer7_outputs(3209) <= b;
    layer7_outputs(3210) <= b and not a;
    layer7_outputs(3211) <= not (a or b);
    layer7_outputs(3212) <= a or b;
    layer7_outputs(3213) <= not (a xor b);
    layer7_outputs(3214) <= a;
    layer7_outputs(3215) <= not (a xor b);
    layer7_outputs(3216) <= not b;
    layer7_outputs(3217) <= not a;
    layer7_outputs(3218) <= a;
    layer7_outputs(3219) <= a;
    layer7_outputs(3220) <= a or b;
    layer7_outputs(3221) <= a or b;
    layer7_outputs(3222) <= a;
    layer7_outputs(3223) <= not b;
    layer7_outputs(3224) <= not b;
    layer7_outputs(3225) <= not b or a;
    layer7_outputs(3226) <= a or b;
    layer7_outputs(3227) <= not (a xor b);
    layer7_outputs(3228) <= a and b;
    layer7_outputs(3229) <= not b;
    layer7_outputs(3230) <= not (a xor b);
    layer7_outputs(3231) <= a xor b;
    layer7_outputs(3232) <= a and b;
    layer7_outputs(3233) <= not a;
    layer7_outputs(3234) <= a and not b;
    layer7_outputs(3235) <= a and b;
    layer7_outputs(3236) <= b and not a;
    layer7_outputs(3237) <= not a;
    layer7_outputs(3238) <= a or b;
    layer7_outputs(3239) <= not (a xor b);
    layer7_outputs(3240) <= b;
    layer7_outputs(3241) <= not a or b;
    layer7_outputs(3242) <= not (a xor b);
    layer7_outputs(3243) <= b;
    layer7_outputs(3244) <= b;
    layer7_outputs(3245) <= 1'b1;
    layer7_outputs(3246) <= not a;
    layer7_outputs(3247) <= not a;
    layer7_outputs(3248) <= not b or a;
    layer7_outputs(3249) <= not (a or b);
    layer7_outputs(3250) <= not b;
    layer7_outputs(3251) <= b;
    layer7_outputs(3252) <= a;
    layer7_outputs(3253) <= not b;
    layer7_outputs(3254) <= a;
    layer7_outputs(3255) <= not (a and b);
    layer7_outputs(3256) <= not (a or b);
    layer7_outputs(3257) <= not b or a;
    layer7_outputs(3258) <= a and not b;
    layer7_outputs(3259) <= a;
    layer7_outputs(3260) <= not b;
    layer7_outputs(3261) <= a and b;
    layer7_outputs(3262) <= not a;
    layer7_outputs(3263) <= b;
    layer7_outputs(3264) <= 1'b0;
    layer7_outputs(3265) <= a or b;
    layer7_outputs(3266) <= a and not b;
    layer7_outputs(3267) <= not (a and b);
    layer7_outputs(3268) <= b;
    layer7_outputs(3269) <= a;
    layer7_outputs(3270) <= not (a xor b);
    layer7_outputs(3271) <= not (a xor b);
    layer7_outputs(3272) <= b and not a;
    layer7_outputs(3273) <= not b;
    layer7_outputs(3274) <= not a or b;
    layer7_outputs(3275) <= a;
    layer7_outputs(3276) <= b;
    layer7_outputs(3277) <= a;
    layer7_outputs(3278) <= a and b;
    layer7_outputs(3279) <= a;
    layer7_outputs(3280) <= a;
    layer7_outputs(3281) <= not a;
    layer7_outputs(3282) <= not (a or b);
    layer7_outputs(3283) <= not b or a;
    layer7_outputs(3284) <= not (a xor b);
    layer7_outputs(3285) <= a or b;
    layer7_outputs(3286) <= not (a xor b);
    layer7_outputs(3287) <= a xor b;
    layer7_outputs(3288) <= a and b;
    layer7_outputs(3289) <= not b or a;
    layer7_outputs(3290) <= a;
    layer7_outputs(3291) <= not a;
    layer7_outputs(3292) <= a and not b;
    layer7_outputs(3293) <= a;
    layer7_outputs(3294) <= b;
    layer7_outputs(3295) <= a and b;
    layer7_outputs(3296) <= b;
    layer7_outputs(3297) <= not a or b;
    layer7_outputs(3298) <= not (a or b);
    layer7_outputs(3299) <= not (a and b);
    layer7_outputs(3300) <= b;
    layer7_outputs(3301) <= b and not a;
    layer7_outputs(3302) <= a and b;
    layer7_outputs(3303) <= a;
    layer7_outputs(3304) <= not a;
    layer7_outputs(3305) <= not a;
    layer7_outputs(3306) <= not b or a;
    layer7_outputs(3307) <= not (a or b);
    layer7_outputs(3308) <= not b;
    layer7_outputs(3309) <= a xor b;
    layer7_outputs(3310) <= a and not b;
    layer7_outputs(3311) <= not b;
    layer7_outputs(3312) <= a and b;
    layer7_outputs(3313) <= b and not a;
    layer7_outputs(3314) <= not a;
    layer7_outputs(3315) <= not a;
    layer7_outputs(3316) <= not b;
    layer7_outputs(3317) <= a;
    layer7_outputs(3318) <= not a;
    layer7_outputs(3319) <= not a;
    layer7_outputs(3320) <= b;
    layer7_outputs(3321) <= not a;
    layer7_outputs(3322) <= a xor b;
    layer7_outputs(3323) <= b and not a;
    layer7_outputs(3324) <= a xor b;
    layer7_outputs(3325) <= b;
    layer7_outputs(3326) <= a and not b;
    layer7_outputs(3327) <= b and not a;
    layer7_outputs(3328) <= a and not b;
    layer7_outputs(3329) <= a;
    layer7_outputs(3330) <= not (a or b);
    layer7_outputs(3331) <= not b or a;
    layer7_outputs(3332) <= b;
    layer7_outputs(3333) <= a and b;
    layer7_outputs(3334) <= not a;
    layer7_outputs(3335) <= b and not a;
    layer7_outputs(3336) <= a and b;
    layer7_outputs(3337) <= not b;
    layer7_outputs(3338) <= not b;
    layer7_outputs(3339) <= a and not b;
    layer7_outputs(3340) <= b;
    layer7_outputs(3341) <= not a;
    layer7_outputs(3342) <= not b;
    layer7_outputs(3343) <= not b or a;
    layer7_outputs(3344) <= a;
    layer7_outputs(3345) <= b;
    layer7_outputs(3346) <= a;
    layer7_outputs(3347) <= not (a and b);
    layer7_outputs(3348) <= a and not b;
    layer7_outputs(3349) <= not (a or b);
    layer7_outputs(3350) <= not a;
    layer7_outputs(3351) <= a and not b;
    layer7_outputs(3352) <= b;
    layer7_outputs(3353) <= a and not b;
    layer7_outputs(3354) <= a;
    layer7_outputs(3355) <= b and not a;
    layer7_outputs(3356) <= b;
    layer7_outputs(3357) <= not a;
    layer7_outputs(3358) <= a or b;
    layer7_outputs(3359) <= b and not a;
    layer7_outputs(3360) <= not (a and b);
    layer7_outputs(3361) <= not b;
    layer7_outputs(3362) <= not (a and b);
    layer7_outputs(3363) <= not (a xor b);
    layer7_outputs(3364) <= not (a and b);
    layer7_outputs(3365) <= not (a and b);
    layer7_outputs(3366) <= not b;
    layer7_outputs(3367) <= b and not a;
    layer7_outputs(3368) <= a xor b;
    layer7_outputs(3369) <= not b;
    layer7_outputs(3370) <= a xor b;
    layer7_outputs(3371) <= a;
    layer7_outputs(3372) <= not a;
    layer7_outputs(3373) <= not (a xor b);
    layer7_outputs(3374) <= a and b;
    layer7_outputs(3375) <= b and not a;
    layer7_outputs(3376) <= b;
    layer7_outputs(3377) <= a and not b;
    layer7_outputs(3378) <= b;
    layer7_outputs(3379) <= a;
    layer7_outputs(3380) <= not b or a;
    layer7_outputs(3381) <= a;
    layer7_outputs(3382) <= a;
    layer7_outputs(3383) <= not b or a;
    layer7_outputs(3384) <= a;
    layer7_outputs(3385) <= 1'b1;
    layer7_outputs(3386) <= not a or b;
    layer7_outputs(3387) <= a xor b;
    layer7_outputs(3388) <= not b;
    layer7_outputs(3389) <= not b;
    layer7_outputs(3390) <= b;
    layer7_outputs(3391) <= not b or a;
    layer7_outputs(3392) <= a;
    layer7_outputs(3393) <= not a;
    layer7_outputs(3394) <= a;
    layer7_outputs(3395) <= 1'b0;
    layer7_outputs(3396) <= a;
    layer7_outputs(3397) <= a and not b;
    layer7_outputs(3398) <= 1'b0;
    layer7_outputs(3399) <= not (a or b);
    layer7_outputs(3400) <= a xor b;
    layer7_outputs(3401) <= not b;
    layer7_outputs(3402) <= b and not a;
    layer7_outputs(3403) <= a;
    layer7_outputs(3404) <= not (a xor b);
    layer7_outputs(3405) <= a or b;
    layer7_outputs(3406) <= b and not a;
    layer7_outputs(3407) <= not b or a;
    layer7_outputs(3408) <= not (a and b);
    layer7_outputs(3409) <= 1'b1;
    layer7_outputs(3410) <= a or b;
    layer7_outputs(3411) <= not (a or b);
    layer7_outputs(3412) <= not b or a;
    layer7_outputs(3413) <= a and not b;
    layer7_outputs(3414) <= a xor b;
    layer7_outputs(3415) <= a xor b;
    layer7_outputs(3416) <= a or b;
    layer7_outputs(3417) <= a and not b;
    layer7_outputs(3418) <= not (a or b);
    layer7_outputs(3419) <= a and b;
    layer7_outputs(3420) <= a or b;
    layer7_outputs(3421) <= not a;
    layer7_outputs(3422) <= b;
    layer7_outputs(3423) <= b;
    layer7_outputs(3424) <= b;
    layer7_outputs(3425) <= a and b;
    layer7_outputs(3426) <= not a or b;
    layer7_outputs(3427) <= a xor b;
    layer7_outputs(3428) <= not (a xor b);
    layer7_outputs(3429) <= a or b;
    layer7_outputs(3430) <= not b;
    layer7_outputs(3431) <= b;
    layer7_outputs(3432) <= not (a xor b);
    layer7_outputs(3433) <= not (a and b);
    layer7_outputs(3434) <= not b or a;
    layer7_outputs(3435) <= a;
    layer7_outputs(3436) <= not a or b;
    layer7_outputs(3437) <= not (a or b);
    layer7_outputs(3438) <= not a;
    layer7_outputs(3439) <= not a;
    layer7_outputs(3440) <= not b;
    layer7_outputs(3441) <= a and b;
    layer7_outputs(3442) <= b and not a;
    layer7_outputs(3443) <= not b;
    layer7_outputs(3444) <= not (a and b);
    layer7_outputs(3445) <= a and not b;
    layer7_outputs(3446) <= a;
    layer7_outputs(3447) <= not a;
    layer7_outputs(3448) <= not (a xor b);
    layer7_outputs(3449) <= not a or b;
    layer7_outputs(3450) <= a;
    layer7_outputs(3451) <= not (a xor b);
    layer7_outputs(3452) <= a xor b;
    layer7_outputs(3453) <= not b;
    layer7_outputs(3454) <= a and b;
    layer7_outputs(3455) <= a xor b;
    layer7_outputs(3456) <= not (a and b);
    layer7_outputs(3457) <= b;
    layer7_outputs(3458) <= b;
    layer7_outputs(3459) <= a;
    layer7_outputs(3460) <= not a;
    layer7_outputs(3461) <= a;
    layer7_outputs(3462) <= a or b;
    layer7_outputs(3463) <= not b or a;
    layer7_outputs(3464) <= not (a xor b);
    layer7_outputs(3465) <= b;
    layer7_outputs(3466) <= b;
    layer7_outputs(3467) <= not b;
    layer7_outputs(3468) <= not a or b;
    layer7_outputs(3469) <= not a or b;
    layer7_outputs(3470) <= not (a and b);
    layer7_outputs(3471) <= a or b;
    layer7_outputs(3472) <= a;
    layer7_outputs(3473) <= not (a xor b);
    layer7_outputs(3474) <= b and not a;
    layer7_outputs(3475) <= a and b;
    layer7_outputs(3476) <= not b;
    layer7_outputs(3477) <= not (a xor b);
    layer7_outputs(3478) <= a or b;
    layer7_outputs(3479) <= not a;
    layer7_outputs(3480) <= not (a and b);
    layer7_outputs(3481) <= a or b;
    layer7_outputs(3482) <= not (a xor b);
    layer7_outputs(3483) <= not a or b;
    layer7_outputs(3484) <= not (a or b);
    layer7_outputs(3485) <= b;
    layer7_outputs(3486) <= a and b;
    layer7_outputs(3487) <= not b;
    layer7_outputs(3488) <= not b;
    layer7_outputs(3489) <= not b or a;
    layer7_outputs(3490) <= not (a or b);
    layer7_outputs(3491) <= a;
    layer7_outputs(3492) <= not (a xor b);
    layer7_outputs(3493) <= not a;
    layer7_outputs(3494) <= not a;
    layer7_outputs(3495) <= not b;
    layer7_outputs(3496) <= b;
    layer7_outputs(3497) <= not a or b;
    layer7_outputs(3498) <= not (a and b);
    layer7_outputs(3499) <= a and not b;
    layer7_outputs(3500) <= not (a xor b);
    layer7_outputs(3501) <= a and not b;
    layer7_outputs(3502) <= not a;
    layer7_outputs(3503) <= not b or a;
    layer7_outputs(3504) <= not a;
    layer7_outputs(3505) <= a xor b;
    layer7_outputs(3506) <= a or b;
    layer7_outputs(3507) <= a or b;
    layer7_outputs(3508) <= b;
    layer7_outputs(3509) <= a;
    layer7_outputs(3510) <= a and not b;
    layer7_outputs(3511) <= not (a or b);
    layer7_outputs(3512) <= not a;
    layer7_outputs(3513) <= not a or b;
    layer7_outputs(3514) <= not b;
    layer7_outputs(3515) <= not (a xor b);
    layer7_outputs(3516) <= a xor b;
    layer7_outputs(3517) <= b;
    layer7_outputs(3518) <= not (a and b);
    layer7_outputs(3519) <= not (a xor b);
    layer7_outputs(3520) <= a;
    layer7_outputs(3521) <= b;
    layer7_outputs(3522) <= not b;
    layer7_outputs(3523) <= b;
    layer7_outputs(3524) <= not (a or b);
    layer7_outputs(3525) <= a xor b;
    layer7_outputs(3526) <= not (a and b);
    layer7_outputs(3527) <= b and not a;
    layer7_outputs(3528) <= b;
    layer7_outputs(3529) <= b and not a;
    layer7_outputs(3530) <= not b;
    layer7_outputs(3531) <= 1'b0;
    layer7_outputs(3532) <= not a;
    layer7_outputs(3533) <= a or b;
    layer7_outputs(3534) <= not (a xor b);
    layer7_outputs(3535) <= a xor b;
    layer7_outputs(3536) <= a and not b;
    layer7_outputs(3537) <= b;
    layer7_outputs(3538) <= not b;
    layer7_outputs(3539) <= a xor b;
    layer7_outputs(3540) <= a;
    layer7_outputs(3541) <= a and not b;
    layer7_outputs(3542) <= not a;
    layer7_outputs(3543) <= b;
    layer7_outputs(3544) <= a;
    layer7_outputs(3545) <= not (a and b);
    layer7_outputs(3546) <= a and not b;
    layer7_outputs(3547) <= not a;
    layer7_outputs(3548) <= not a;
    layer7_outputs(3549) <= b and not a;
    layer7_outputs(3550) <= a;
    layer7_outputs(3551) <= not b;
    layer7_outputs(3552) <= not b;
    layer7_outputs(3553) <= b;
    layer7_outputs(3554) <= not (a and b);
    layer7_outputs(3555) <= not (a xor b);
    layer7_outputs(3556) <= b and not a;
    layer7_outputs(3557) <= b;
    layer7_outputs(3558) <= not a;
    layer7_outputs(3559) <= b;
    layer7_outputs(3560) <= a or b;
    layer7_outputs(3561) <= not a;
    layer7_outputs(3562) <= a and not b;
    layer7_outputs(3563) <= a and b;
    layer7_outputs(3564) <= not b or a;
    layer7_outputs(3565) <= a xor b;
    layer7_outputs(3566) <= not (a xor b);
    layer7_outputs(3567) <= a;
    layer7_outputs(3568) <= a and not b;
    layer7_outputs(3569) <= a and not b;
    layer7_outputs(3570) <= a and b;
    layer7_outputs(3571) <= a;
    layer7_outputs(3572) <= b;
    layer7_outputs(3573) <= a;
    layer7_outputs(3574) <= not b;
    layer7_outputs(3575) <= not a;
    layer7_outputs(3576) <= a;
    layer7_outputs(3577) <= not b;
    layer7_outputs(3578) <= not b or a;
    layer7_outputs(3579) <= a and not b;
    layer7_outputs(3580) <= 1'b0;
    layer7_outputs(3581) <= b and not a;
    layer7_outputs(3582) <= b and not a;
    layer7_outputs(3583) <= not (a or b);
    layer7_outputs(3584) <= a;
    layer7_outputs(3585) <= a and b;
    layer7_outputs(3586) <= a;
    layer7_outputs(3587) <= not (a xor b);
    layer7_outputs(3588) <= not (a xor b);
    layer7_outputs(3589) <= not (a and b);
    layer7_outputs(3590) <= not (a or b);
    layer7_outputs(3591) <= not (a or b);
    layer7_outputs(3592) <= not b;
    layer7_outputs(3593) <= not (a and b);
    layer7_outputs(3594) <= not b;
    layer7_outputs(3595) <= not a or b;
    layer7_outputs(3596) <= not b or a;
    layer7_outputs(3597) <= b;
    layer7_outputs(3598) <= not (a xor b);
    layer7_outputs(3599) <= not a or b;
    layer7_outputs(3600) <= not b;
    layer7_outputs(3601) <= a;
    layer7_outputs(3602) <= a;
    layer7_outputs(3603) <= not (a xor b);
    layer7_outputs(3604) <= a and b;
    layer7_outputs(3605) <= not (a xor b);
    layer7_outputs(3606) <= not a or b;
    layer7_outputs(3607) <= a xor b;
    layer7_outputs(3608) <= not a;
    layer7_outputs(3609) <= a or b;
    layer7_outputs(3610) <= not a or b;
    layer7_outputs(3611) <= not b;
    layer7_outputs(3612) <= a xor b;
    layer7_outputs(3613) <= not a or b;
    layer7_outputs(3614) <= not b;
    layer7_outputs(3615) <= a xor b;
    layer7_outputs(3616) <= not b;
    layer7_outputs(3617) <= not b or a;
    layer7_outputs(3618) <= not a;
    layer7_outputs(3619) <= b;
    layer7_outputs(3620) <= a xor b;
    layer7_outputs(3621) <= b and not a;
    layer7_outputs(3622) <= not b;
    layer7_outputs(3623) <= not a;
    layer7_outputs(3624) <= b;
    layer7_outputs(3625) <= not b;
    layer7_outputs(3626) <= not (a xor b);
    layer7_outputs(3627) <= not b;
    layer7_outputs(3628) <= not (a or b);
    layer7_outputs(3629) <= a xor b;
    layer7_outputs(3630) <= not (a or b);
    layer7_outputs(3631) <= a and not b;
    layer7_outputs(3632) <= a xor b;
    layer7_outputs(3633) <= not (a xor b);
    layer7_outputs(3634) <= a and not b;
    layer7_outputs(3635) <= b;
    layer7_outputs(3636) <= a and b;
    layer7_outputs(3637) <= b;
    layer7_outputs(3638) <= a;
    layer7_outputs(3639) <= a and not b;
    layer7_outputs(3640) <= not (a and b);
    layer7_outputs(3641) <= not a;
    layer7_outputs(3642) <= a xor b;
    layer7_outputs(3643) <= b;
    layer7_outputs(3644) <= b and not a;
    layer7_outputs(3645) <= not a or b;
    layer7_outputs(3646) <= not a;
    layer7_outputs(3647) <= b;
    layer7_outputs(3648) <= a xor b;
    layer7_outputs(3649) <= not (a xor b);
    layer7_outputs(3650) <= not a or b;
    layer7_outputs(3651) <= a;
    layer7_outputs(3652) <= b and not a;
    layer7_outputs(3653) <= a;
    layer7_outputs(3654) <= not (a or b);
    layer7_outputs(3655) <= not (a xor b);
    layer7_outputs(3656) <= not (a xor b);
    layer7_outputs(3657) <= not b;
    layer7_outputs(3658) <= b;
    layer7_outputs(3659) <= not a or b;
    layer7_outputs(3660) <= not b;
    layer7_outputs(3661) <= not b;
    layer7_outputs(3662) <= not b or a;
    layer7_outputs(3663) <= a or b;
    layer7_outputs(3664) <= a or b;
    layer7_outputs(3665) <= not (a xor b);
    layer7_outputs(3666) <= not a or b;
    layer7_outputs(3667) <= not a;
    layer7_outputs(3668) <= a;
    layer7_outputs(3669) <= not b;
    layer7_outputs(3670) <= a and b;
    layer7_outputs(3671) <= not (a xor b);
    layer7_outputs(3672) <= not a;
    layer7_outputs(3673) <= 1'b1;
    layer7_outputs(3674) <= b;
    layer7_outputs(3675) <= not b or a;
    layer7_outputs(3676) <= a and not b;
    layer7_outputs(3677) <= not (a and b);
    layer7_outputs(3678) <= not (a xor b);
    layer7_outputs(3679) <= b;
    layer7_outputs(3680) <= not a or b;
    layer7_outputs(3681) <= 1'b0;
    layer7_outputs(3682) <= not a;
    layer7_outputs(3683) <= b;
    layer7_outputs(3684) <= a and not b;
    layer7_outputs(3685) <= not a or b;
    layer7_outputs(3686) <= not b;
    layer7_outputs(3687) <= a and not b;
    layer7_outputs(3688) <= not (a xor b);
    layer7_outputs(3689) <= not a or b;
    layer7_outputs(3690) <= a and b;
    layer7_outputs(3691) <= not a or b;
    layer7_outputs(3692) <= not (a xor b);
    layer7_outputs(3693) <= a and not b;
    layer7_outputs(3694) <= a and not b;
    layer7_outputs(3695) <= a or b;
    layer7_outputs(3696) <= not (a or b);
    layer7_outputs(3697) <= b;
    layer7_outputs(3698) <= b and not a;
    layer7_outputs(3699) <= a and b;
    layer7_outputs(3700) <= b;
    layer7_outputs(3701) <= a and not b;
    layer7_outputs(3702) <= a and not b;
    layer7_outputs(3703) <= not a;
    layer7_outputs(3704) <= not b;
    layer7_outputs(3705) <= a xor b;
    layer7_outputs(3706) <= b and not a;
    layer7_outputs(3707) <= a xor b;
    layer7_outputs(3708) <= not b;
    layer7_outputs(3709) <= a and not b;
    layer7_outputs(3710) <= b;
    layer7_outputs(3711) <= a and not b;
    layer7_outputs(3712) <= a xor b;
    layer7_outputs(3713) <= not (a xor b);
    layer7_outputs(3714) <= a or b;
    layer7_outputs(3715) <= not a;
    layer7_outputs(3716) <= not b;
    layer7_outputs(3717) <= b;
    layer7_outputs(3718) <= not b or a;
    layer7_outputs(3719) <= not a;
    layer7_outputs(3720) <= a;
    layer7_outputs(3721) <= not a or b;
    layer7_outputs(3722) <= not (a xor b);
    layer7_outputs(3723) <= 1'b0;
    layer7_outputs(3724) <= a xor b;
    layer7_outputs(3725) <= b;
    layer7_outputs(3726) <= not b;
    layer7_outputs(3727) <= a xor b;
    layer7_outputs(3728) <= not b;
    layer7_outputs(3729) <= not a;
    layer7_outputs(3730) <= a and not b;
    layer7_outputs(3731) <= a;
    layer7_outputs(3732) <= not a;
    layer7_outputs(3733) <= not a;
    layer7_outputs(3734) <= not (a xor b);
    layer7_outputs(3735) <= a;
    layer7_outputs(3736) <= not a;
    layer7_outputs(3737) <= a and not b;
    layer7_outputs(3738) <= b;
    layer7_outputs(3739) <= b;
    layer7_outputs(3740) <= not (a xor b);
    layer7_outputs(3741) <= a xor b;
    layer7_outputs(3742) <= a or b;
    layer7_outputs(3743) <= not a or b;
    layer7_outputs(3744) <= a;
    layer7_outputs(3745) <= 1'b0;
    layer7_outputs(3746) <= not b;
    layer7_outputs(3747) <= a and b;
    layer7_outputs(3748) <= a;
    layer7_outputs(3749) <= a or b;
    layer7_outputs(3750) <= not a;
    layer7_outputs(3751) <= not a or b;
    layer7_outputs(3752) <= not b;
    layer7_outputs(3753) <= a;
    layer7_outputs(3754) <= not b or a;
    layer7_outputs(3755) <= a and not b;
    layer7_outputs(3756) <= b;
    layer7_outputs(3757) <= b;
    layer7_outputs(3758) <= not b;
    layer7_outputs(3759) <= a xor b;
    layer7_outputs(3760) <= not a;
    layer7_outputs(3761) <= not a;
    layer7_outputs(3762) <= not b;
    layer7_outputs(3763) <= a;
    layer7_outputs(3764) <= not a;
    layer7_outputs(3765) <= not a or b;
    layer7_outputs(3766) <= not b or a;
    layer7_outputs(3767) <= not (a xor b);
    layer7_outputs(3768) <= b;
    layer7_outputs(3769) <= a and b;
    layer7_outputs(3770) <= not a;
    layer7_outputs(3771) <= a or b;
    layer7_outputs(3772) <= not b;
    layer7_outputs(3773) <= a xor b;
    layer7_outputs(3774) <= not a;
    layer7_outputs(3775) <= b;
    layer7_outputs(3776) <= a xor b;
    layer7_outputs(3777) <= not (a and b);
    layer7_outputs(3778) <= not b;
    layer7_outputs(3779) <= a;
    layer7_outputs(3780) <= not (a xor b);
    layer7_outputs(3781) <= not a;
    layer7_outputs(3782) <= a;
    layer7_outputs(3783) <= a or b;
    layer7_outputs(3784) <= b;
    layer7_outputs(3785) <= a or b;
    layer7_outputs(3786) <= a and b;
    layer7_outputs(3787) <= b;
    layer7_outputs(3788) <= a;
    layer7_outputs(3789) <= not a;
    layer7_outputs(3790) <= a or b;
    layer7_outputs(3791) <= b;
    layer7_outputs(3792) <= not a or b;
    layer7_outputs(3793) <= not b;
    layer7_outputs(3794) <= b;
    layer7_outputs(3795) <= not (a or b);
    layer7_outputs(3796) <= not a;
    layer7_outputs(3797) <= a;
    layer7_outputs(3798) <= not a;
    layer7_outputs(3799) <= b;
    layer7_outputs(3800) <= not a or b;
    layer7_outputs(3801) <= a and not b;
    layer7_outputs(3802) <= a;
    layer7_outputs(3803) <= not (a xor b);
    layer7_outputs(3804) <= a;
    layer7_outputs(3805) <= a or b;
    layer7_outputs(3806) <= a xor b;
    layer7_outputs(3807) <= not a;
    layer7_outputs(3808) <= a and not b;
    layer7_outputs(3809) <= not a or b;
    layer7_outputs(3810) <= a and not b;
    layer7_outputs(3811) <= a;
    layer7_outputs(3812) <= a;
    layer7_outputs(3813) <= b;
    layer7_outputs(3814) <= b and not a;
    layer7_outputs(3815) <= a;
    layer7_outputs(3816) <= not b;
    layer7_outputs(3817) <= not (a and b);
    layer7_outputs(3818) <= not (a and b);
    layer7_outputs(3819) <= a xor b;
    layer7_outputs(3820) <= not a or b;
    layer7_outputs(3821) <= a or b;
    layer7_outputs(3822) <= a xor b;
    layer7_outputs(3823) <= b;
    layer7_outputs(3824) <= b;
    layer7_outputs(3825) <= 1'b0;
    layer7_outputs(3826) <= a or b;
    layer7_outputs(3827) <= not b;
    layer7_outputs(3828) <= not a;
    layer7_outputs(3829) <= b;
    layer7_outputs(3830) <= not (a xor b);
    layer7_outputs(3831) <= not (a or b);
    layer7_outputs(3832) <= a or b;
    layer7_outputs(3833) <= b;
    layer7_outputs(3834) <= a and not b;
    layer7_outputs(3835) <= not (a or b);
    layer7_outputs(3836) <= a;
    layer7_outputs(3837) <= b and not a;
    layer7_outputs(3838) <= not (a and b);
    layer7_outputs(3839) <= a xor b;
    layer7_outputs(3840) <= a xor b;
    layer7_outputs(3841) <= a xor b;
    layer7_outputs(3842) <= not (a and b);
    layer7_outputs(3843) <= a;
    layer7_outputs(3844) <= b;
    layer7_outputs(3845) <= b;
    layer7_outputs(3846) <= a;
    layer7_outputs(3847) <= not a;
    layer7_outputs(3848) <= a xor b;
    layer7_outputs(3849) <= not b or a;
    layer7_outputs(3850) <= a or b;
    layer7_outputs(3851) <= b;
    layer7_outputs(3852) <= not (a xor b);
    layer7_outputs(3853) <= a and b;
    layer7_outputs(3854) <= not (a or b);
    layer7_outputs(3855) <= a and not b;
    layer7_outputs(3856) <= not (a xor b);
    layer7_outputs(3857) <= b;
    layer7_outputs(3858) <= not b;
    layer7_outputs(3859) <= b and not a;
    layer7_outputs(3860) <= a or b;
    layer7_outputs(3861) <= b;
    layer7_outputs(3862) <= b;
    layer7_outputs(3863) <= a or b;
    layer7_outputs(3864) <= b;
    layer7_outputs(3865) <= not (a or b);
    layer7_outputs(3866) <= a and not b;
    layer7_outputs(3867) <= not a;
    layer7_outputs(3868) <= not (a xor b);
    layer7_outputs(3869) <= a and not b;
    layer7_outputs(3870) <= not b;
    layer7_outputs(3871) <= a and not b;
    layer7_outputs(3872) <= not b;
    layer7_outputs(3873) <= b;
    layer7_outputs(3874) <= a xor b;
    layer7_outputs(3875) <= not (a xor b);
    layer7_outputs(3876) <= a and b;
    layer7_outputs(3877) <= b and not a;
    layer7_outputs(3878) <= not b;
    layer7_outputs(3879) <= a xor b;
    layer7_outputs(3880) <= not (a xor b);
    layer7_outputs(3881) <= not a or b;
    layer7_outputs(3882) <= not b;
    layer7_outputs(3883) <= not b or a;
    layer7_outputs(3884) <= a xor b;
    layer7_outputs(3885) <= not (a or b);
    layer7_outputs(3886) <= 1'b1;
    layer7_outputs(3887) <= a xor b;
    layer7_outputs(3888) <= not b;
    layer7_outputs(3889) <= not a or b;
    layer7_outputs(3890) <= b and not a;
    layer7_outputs(3891) <= b;
    layer7_outputs(3892) <= a and not b;
    layer7_outputs(3893) <= b;
    layer7_outputs(3894) <= a xor b;
    layer7_outputs(3895) <= not b;
    layer7_outputs(3896) <= b and not a;
    layer7_outputs(3897) <= not (a or b);
    layer7_outputs(3898) <= not (a or b);
    layer7_outputs(3899) <= a;
    layer7_outputs(3900) <= a;
    layer7_outputs(3901) <= not a;
    layer7_outputs(3902) <= not b;
    layer7_outputs(3903) <= a xor b;
    layer7_outputs(3904) <= not b;
    layer7_outputs(3905) <= a;
    layer7_outputs(3906) <= a and not b;
    layer7_outputs(3907) <= a;
    layer7_outputs(3908) <= a xor b;
    layer7_outputs(3909) <= a xor b;
    layer7_outputs(3910) <= not b or a;
    layer7_outputs(3911) <= not (a and b);
    layer7_outputs(3912) <= not (a xor b);
    layer7_outputs(3913) <= a and not b;
    layer7_outputs(3914) <= a;
    layer7_outputs(3915) <= not a;
    layer7_outputs(3916) <= a xor b;
    layer7_outputs(3917) <= not (a xor b);
    layer7_outputs(3918) <= not b;
    layer7_outputs(3919) <= not (a or b);
    layer7_outputs(3920) <= 1'b0;
    layer7_outputs(3921) <= a xor b;
    layer7_outputs(3922) <= not (a and b);
    layer7_outputs(3923) <= not b or a;
    layer7_outputs(3924) <= 1'b1;
    layer7_outputs(3925) <= b and not a;
    layer7_outputs(3926) <= b;
    layer7_outputs(3927) <= not a;
    layer7_outputs(3928) <= not (a xor b);
    layer7_outputs(3929) <= a and b;
    layer7_outputs(3930) <= b;
    layer7_outputs(3931) <= not a;
    layer7_outputs(3932) <= b and not a;
    layer7_outputs(3933) <= b and not a;
    layer7_outputs(3934) <= not a;
    layer7_outputs(3935) <= a xor b;
    layer7_outputs(3936) <= not (a or b);
    layer7_outputs(3937) <= a or b;
    layer7_outputs(3938) <= a and b;
    layer7_outputs(3939) <= not b;
    layer7_outputs(3940) <= b;
    layer7_outputs(3941) <= b and not a;
    layer7_outputs(3942) <= not (a xor b);
    layer7_outputs(3943) <= not b;
    layer7_outputs(3944) <= not (a and b);
    layer7_outputs(3945) <= a and not b;
    layer7_outputs(3946) <= not b or a;
    layer7_outputs(3947) <= a;
    layer7_outputs(3948) <= not b;
    layer7_outputs(3949) <= b;
    layer7_outputs(3950) <= not b;
    layer7_outputs(3951) <= not b;
    layer7_outputs(3952) <= a xor b;
    layer7_outputs(3953) <= b;
    layer7_outputs(3954) <= not b or a;
    layer7_outputs(3955) <= not a;
    layer7_outputs(3956) <= not (a and b);
    layer7_outputs(3957) <= not (a xor b);
    layer7_outputs(3958) <= not a;
    layer7_outputs(3959) <= b;
    layer7_outputs(3960) <= a and not b;
    layer7_outputs(3961) <= not a or b;
    layer7_outputs(3962) <= not (a xor b);
    layer7_outputs(3963) <= not b or a;
    layer7_outputs(3964) <= 1'b1;
    layer7_outputs(3965) <= b and not a;
    layer7_outputs(3966) <= a and b;
    layer7_outputs(3967) <= a or b;
    layer7_outputs(3968) <= not b or a;
    layer7_outputs(3969) <= not b;
    layer7_outputs(3970) <= not b;
    layer7_outputs(3971) <= not b;
    layer7_outputs(3972) <= not (a or b);
    layer7_outputs(3973) <= a;
    layer7_outputs(3974) <= a xor b;
    layer7_outputs(3975) <= a xor b;
    layer7_outputs(3976) <= a;
    layer7_outputs(3977) <= not (a xor b);
    layer7_outputs(3978) <= b and not a;
    layer7_outputs(3979) <= not a;
    layer7_outputs(3980) <= a;
    layer7_outputs(3981) <= 1'b0;
    layer7_outputs(3982) <= b;
    layer7_outputs(3983) <= not a or b;
    layer7_outputs(3984) <= a and b;
    layer7_outputs(3985) <= a and not b;
    layer7_outputs(3986) <= b and not a;
    layer7_outputs(3987) <= not a;
    layer7_outputs(3988) <= a xor b;
    layer7_outputs(3989) <= b;
    layer7_outputs(3990) <= not a or b;
    layer7_outputs(3991) <= not b or a;
    layer7_outputs(3992) <= not a;
    layer7_outputs(3993) <= not (a or b);
    layer7_outputs(3994) <= a xor b;
    layer7_outputs(3995) <= not b or a;
    layer7_outputs(3996) <= not b;
    layer7_outputs(3997) <= a and b;
    layer7_outputs(3998) <= b;
    layer7_outputs(3999) <= b;
    layer7_outputs(4000) <= not (a xor b);
    layer7_outputs(4001) <= a and b;
    layer7_outputs(4002) <= a and b;
    layer7_outputs(4003) <= b and not a;
    layer7_outputs(4004) <= not a or b;
    layer7_outputs(4005) <= a;
    layer7_outputs(4006) <= not b or a;
    layer7_outputs(4007) <= a or b;
    layer7_outputs(4008) <= not a;
    layer7_outputs(4009) <= not (a and b);
    layer7_outputs(4010) <= not b or a;
    layer7_outputs(4011) <= a xor b;
    layer7_outputs(4012) <= 1'b1;
    layer7_outputs(4013) <= not b;
    layer7_outputs(4014) <= a;
    layer7_outputs(4015) <= not a;
    layer7_outputs(4016) <= not (a or b);
    layer7_outputs(4017) <= a;
    layer7_outputs(4018) <= not b;
    layer7_outputs(4019) <= not b;
    layer7_outputs(4020) <= a and not b;
    layer7_outputs(4021) <= not b;
    layer7_outputs(4022) <= not a;
    layer7_outputs(4023) <= a and not b;
    layer7_outputs(4024) <= a and b;
    layer7_outputs(4025) <= a;
    layer7_outputs(4026) <= not b;
    layer7_outputs(4027) <= a;
    layer7_outputs(4028) <= not b;
    layer7_outputs(4029) <= a xor b;
    layer7_outputs(4030) <= a or b;
    layer7_outputs(4031) <= not (a xor b);
    layer7_outputs(4032) <= b and not a;
    layer7_outputs(4033) <= not b;
    layer7_outputs(4034) <= b;
    layer7_outputs(4035) <= a;
    layer7_outputs(4036) <= 1'b0;
    layer7_outputs(4037) <= a and not b;
    layer7_outputs(4038) <= b;
    layer7_outputs(4039) <= a xor b;
    layer7_outputs(4040) <= a or b;
    layer7_outputs(4041) <= not a;
    layer7_outputs(4042) <= b and not a;
    layer7_outputs(4043) <= a xor b;
    layer7_outputs(4044) <= 1'b0;
    layer7_outputs(4045) <= not a or b;
    layer7_outputs(4046) <= a xor b;
    layer7_outputs(4047) <= not b or a;
    layer7_outputs(4048) <= not b;
    layer7_outputs(4049) <= not a;
    layer7_outputs(4050) <= a and b;
    layer7_outputs(4051) <= not b;
    layer7_outputs(4052) <= 1'b1;
    layer7_outputs(4053) <= a;
    layer7_outputs(4054) <= b;
    layer7_outputs(4055) <= b and not a;
    layer7_outputs(4056) <= not a or b;
    layer7_outputs(4057) <= not b;
    layer7_outputs(4058) <= 1'b1;
    layer7_outputs(4059) <= b;
    layer7_outputs(4060) <= b;
    layer7_outputs(4061) <= b;
    layer7_outputs(4062) <= a and b;
    layer7_outputs(4063) <= not a;
    layer7_outputs(4064) <= b and not a;
    layer7_outputs(4065) <= not (a and b);
    layer7_outputs(4066) <= b;
    layer7_outputs(4067) <= b and not a;
    layer7_outputs(4068) <= a or b;
    layer7_outputs(4069) <= a and not b;
    layer7_outputs(4070) <= a or b;
    layer7_outputs(4071) <= b;
    layer7_outputs(4072) <= not (a xor b);
    layer7_outputs(4073) <= a xor b;
    layer7_outputs(4074) <= not (a or b);
    layer7_outputs(4075) <= not a;
    layer7_outputs(4076) <= a xor b;
    layer7_outputs(4077) <= not (a xor b);
    layer7_outputs(4078) <= a;
    layer7_outputs(4079) <= not (a or b);
    layer7_outputs(4080) <= not (a xor b);
    layer7_outputs(4081) <= b;
    layer7_outputs(4082) <= not (a or b);
    layer7_outputs(4083) <= not b or a;
    layer7_outputs(4084) <= not (a xor b);
    layer7_outputs(4085) <= not a;
    layer7_outputs(4086) <= a and b;
    layer7_outputs(4087) <= a or b;
    layer7_outputs(4088) <= not b;
    layer7_outputs(4089) <= not (a or b);
    layer7_outputs(4090) <= a or b;
    layer7_outputs(4091) <= not (a or b);
    layer7_outputs(4092) <= a;
    layer7_outputs(4093) <= a or b;
    layer7_outputs(4094) <= not b;
    layer7_outputs(4095) <= not a;
    layer7_outputs(4096) <= not a or b;
    layer7_outputs(4097) <= b;
    layer7_outputs(4098) <= not b or a;
    layer7_outputs(4099) <= not (a xor b);
    layer7_outputs(4100) <= not b;
    layer7_outputs(4101) <= a;
    layer7_outputs(4102) <= not b;
    layer7_outputs(4103) <= not a;
    layer7_outputs(4104) <= a;
    layer7_outputs(4105) <= not b;
    layer7_outputs(4106) <= a;
    layer7_outputs(4107) <= not b;
    layer7_outputs(4108) <= not b;
    layer7_outputs(4109) <= not b or a;
    layer7_outputs(4110) <= a;
    layer7_outputs(4111) <= not a or b;
    layer7_outputs(4112) <= a;
    layer7_outputs(4113) <= not b;
    layer7_outputs(4114) <= not a or b;
    layer7_outputs(4115) <= a or b;
    layer7_outputs(4116) <= a and b;
    layer7_outputs(4117) <= not a;
    layer7_outputs(4118) <= not b;
    layer7_outputs(4119) <= not a;
    layer7_outputs(4120) <= b and not a;
    layer7_outputs(4121) <= a and not b;
    layer7_outputs(4122) <= not a;
    layer7_outputs(4123) <= b;
    layer7_outputs(4124) <= a and not b;
    layer7_outputs(4125) <= a xor b;
    layer7_outputs(4126) <= not (a xor b);
    layer7_outputs(4127) <= b;
    layer7_outputs(4128) <= a and b;
    layer7_outputs(4129) <= not (a or b);
    layer7_outputs(4130) <= 1'b1;
    layer7_outputs(4131) <= not (a xor b);
    layer7_outputs(4132) <= not a or b;
    layer7_outputs(4133) <= a or b;
    layer7_outputs(4134) <= not a;
    layer7_outputs(4135) <= b;
    layer7_outputs(4136) <= a xor b;
    layer7_outputs(4137) <= a and b;
    layer7_outputs(4138) <= not a;
    layer7_outputs(4139) <= not (a xor b);
    layer7_outputs(4140) <= not (a xor b);
    layer7_outputs(4141) <= not (a xor b);
    layer7_outputs(4142) <= not (a and b);
    layer7_outputs(4143) <= not a;
    layer7_outputs(4144) <= not b or a;
    layer7_outputs(4145) <= not b;
    layer7_outputs(4146) <= b;
    layer7_outputs(4147) <= 1'b1;
    layer7_outputs(4148) <= not b or a;
    layer7_outputs(4149) <= b;
    layer7_outputs(4150) <= a and not b;
    layer7_outputs(4151) <= a;
    layer7_outputs(4152) <= b;
    layer7_outputs(4153) <= a;
    layer7_outputs(4154) <= not (a xor b);
    layer7_outputs(4155) <= b and not a;
    layer7_outputs(4156) <= not a;
    layer7_outputs(4157) <= b;
    layer7_outputs(4158) <= a or b;
    layer7_outputs(4159) <= a xor b;
    layer7_outputs(4160) <= b;
    layer7_outputs(4161) <= not a;
    layer7_outputs(4162) <= b and not a;
    layer7_outputs(4163) <= not a;
    layer7_outputs(4164) <= a and not b;
    layer7_outputs(4165) <= a;
    layer7_outputs(4166) <= a xor b;
    layer7_outputs(4167) <= not a or b;
    layer7_outputs(4168) <= not a;
    layer7_outputs(4169) <= a;
    layer7_outputs(4170) <= a xor b;
    layer7_outputs(4171) <= a and not b;
    layer7_outputs(4172) <= not (a or b);
    layer7_outputs(4173) <= not a or b;
    layer7_outputs(4174) <= not b or a;
    layer7_outputs(4175) <= not (a xor b);
    layer7_outputs(4176) <= not b or a;
    layer7_outputs(4177) <= b;
    layer7_outputs(4178) <= a or b;
    layer7_outputs(4179) <= a and not b;
    layer7_outputs(4180) <= not (a or b);
    layer7_outputs(4181) <= not (a xor b);
    layer7_outputs(4182) <= a and not b;
    layer7_outputs(4183) <= a and b;
    layer7_outputs(4184) <= not (a xor b);
    layer7_outputs(4185) <= not a;
    layer7_outputs(4186) <= not (a or b);
    layer7_outputs(4187) <= a;
    layer7_outputs(4188) <= not b;
    layer7_outputs(4189) <= a xor b;
    layer7_outputs(4190) <= not a;
    layer7_outputs(4191) <= not (a or b);
    layer7_outputs(4192) <= not (a xor b);
    layer7_outputs(4193) <= not a;
    layer7_outputs(4194) <= b;
    layer7_outputs(4195) <= a or b;
    layer7_outputs(4196) <= a;
    layer7_outputs(4197) <= 1'b0;
    layer7_outputs(4198) <= not a;
    layer7_outputs(4199) <= not (a or b);
    layer7_outputs(4200) <= not b;
    layer7_outputs(4201) <= not a;
    layer7_outputs(4202) <= a and not b;
    layer7_outputs(4203) <= a xor b;
    layer7_outputs(4204) <= not a;
    layer7_outputs(4205) <= a;
    layer7_outputs(4206) <= not b;
    layer7_outputs(4207) <= a or b;
    layer7_outputs(4208) <= a and b;
    layer7_outputs(4209) <= a;
    layer7_outputs(4210) <= b;
    layer7_outputs(4211) <= b and not a;
    layer7_outputs(4212) <= not b;
    layer7_outputs(4213) <= a and b;
    layer7_outputs(4214) <= not b;
    layer7_outputs(4215) <= not (a and b);
    layer7_outputs(4216) <= a;
    layer7_outputs(4217) <= not b;
    layer7_outputs(4218) <= not b or a;
    layer7_outputs(4219) <= a and b;
    layer7_outputs(4220) <= not b;
    layer7_outputs(4221) <= not (a xor b);
    layer7_outputs(4222) <= not (a xor b);
    layer7_outputs(4223) <= not b;
    layer7_outputs(4224) <= b;
    layer7_outputs(4225) <= not (a xor b);
    layer7_outputs(4226) <= b;
    layer7_outputs(4227) <= not a;
    layer7_outputs(4228) <= b;
    layer7_outputs(4229) <= b and not a;
    layer7_outputs(4230) <= a;
    layer7_outputs(4231) <= a and not b;
    layer7_outputs(4232) <= not b;
    layer7_outputs(4233) <= b and not a;
    layer7_outputs(4234) <= a;
    layer7_outputs(4235) <= not (a xor b);
    layer7_outputs(4236) <= not a or b;
    layer7_outputs(4237) <= not a or b;
    layer7_outputs(4238) <= not a;
    layer7_outputs(4239) <= not (a and b);
    layer7_outputs(4240) <= not a or b;
    layer7_outputs(4241) <= a xor b;
    layer7_outputs(4242) <= a;
    layer7_outputs(4243) <= a and b;
    layer7_outputs(4244) <= b and not a;
    layer7_outputs(4245) <= not (a xor b);
    layer7_outputs(4246) <= not b;
    layer7_outputs(4247) <= a xor b;
    layer7_outputs(4248) <= not b;
    layer7_outputs(4249) <= b and not a;
    layer7_outputs(4250) <= not b;
    layer7_outputs(4251) <= a and not b;
    layer7_outputs(4252) <= a;
    layer7_outputs(4253) <= not a;
    layer7_outputs(4254) <= not a or b;
    layer7_outputs(4255) <= not a;
    layer7_outputs(4256) <= not (a and b);
    layer7_outputs(4257) <= a and b;
    layer7_outputs(4258) <= a;
    layer7_outputs(4259) <= not (a and b);
    layer7_outputs(4260) <= a and b;
    layer7_outputs(4261) <= not a or b;
    layer7_outputs(4262) <= not b;
    layer7_outputs(4263) <= not b or a;
    layer7_outputs(4264) <= a;
    layer7_outputs(4265) <= not b;
    layer7_outputs(4266) <= not b;
    layer7_outputs(4267) <= b;
    layer7_outputs(4268) <= not (a and b);
    layer7_outputs(4269) <= b;
    layer7_outputs(4270) <= b and not a;
    layer7_outputs(4271) <= a and not b;
    layer7_outputs(4272) <= not b;
    layer7_outputs(4273) <= not b;
    layer7_outputs(4274) <= not (a and b);
    layer7_outputs(4275) <= b;
    layer7_outputs(4276) <= a and b;
    layer7_outputs(4277) <= 1'b0;
    layer7_outputs(4278) <= not a;
    layer7_outputs(4279) <= a;
    layer7_outputs(4280) <= b and not a;
    layer7_outputs(4281) <= a and b;
    layer7_outputs(4282) <= not a;
    layer7_outputs(4283) <= a;
    layer7_outputs(4284) <= a or b;
    layer7_outputs(4285) <= a xor b;
    layer7_outputs(4286) <= b;
    layer7_outputs(4287) <= a and not b;
    layer7_outputs(4288) <= 1'b0;
    layer7_outputs(4289) <= a and not b;
    layer7_outputs(4290) <= not (a xor b);
    layer7_outputs(4291) <= b and not a;
    layer7_outputs(4292) <= a or b;
    layer7_outputs(4293) <= not a;
    layer7_outputs(4294) <= b;
    layer7_outputs(4295) <= a or b;
    layer7_outputs(4296) <= 1'b0;
    layer7_outputs(4297) <= a xor b;
    layer7_outputs(4298) <= 1'b1;
    layer7_outputs(4299) <= a or b;
    layer7_outputs(4300) <= b;
    layer7_outputs(4301) <= a xor b;
    layer7_outputs(4302) <= not a;
    layer7_outputs(4303) <= a;
    layer7_outputs(4304) <= b;
    layer7_outputs(4305) <= a and b;
    layer7_outputs(4306) <= not (a xor b);
    layer7_outputs(4307) <= b;
    layer7_outputs(4308) <= a or b;
    layer7_outputs(4309) <= a;
    layer7_outputs(4310) <= a and not b;
    layer7_outputs(4311) <= not (a and b);
    layer7_outputs(4312) <= a and b;
    layer7_outputs(4313) <= not b or a;
    layer7_outputs(4314) <= b;
    layer7_outputs(4315) <= not a;
    layer7_outputs(4316) <= not (a xor b);
    layer7_outputs(4317) <= not b or a;
    layer7_outputs(4318) <= not a or b;
    layer7_outputs(4319) <= not a;
    layer7_outputs(4320) <= b;
    layer7_outputs(4321) <= not a;
    layer7_outputs(4322) <= not (a or b);
    layer7_outputs(4323) <= a and not b;
    layer7_outputs(4324) <= a or b;
    layer7_outputs(4325) <= not (a or b);
    layer7_outputs(4326) <= a;
    layer7_outputs(4327) <= a xor b;
    layer7_outputs(4328) <= not (a and b);
    layer7_outputs(4329) <= not a or b;
    layer7_outputs(4330) <= b;
    layer7_outputs(4331) <= not (a xor b);
    layer7_outputs(4332) <= not (a or b);
    layer7_outputs(4333) <= a;
    layer7_outputs(4334) <= a;
    layer7_outputs(4335) <= 1'b0;
    layer7_outputs(4336) <= a and not b;
    layer7_outputs(4337) <= not (a xor b);
    layer7_outputs(4338) <= a;
    layer7_outputs(4339) <= not a;
    layer7_outputs(4340) <= not a;
    layer7_outputs(4341) <= not b;
    layer7_outputs(4342) <= not b;
    layer7_outputs(4343) <= b;
    layer7_outputs(4344) <= not (a or b);
    layer7_outputs(4345) <= a;
    layer7_outputs(4346) <= b;
    layer7_outputs(4347) <= not b or a;
    layer7_outputs(4348) <= not b or a;
    layer7_outputs(4349) <= not (a xor b);
    layer7_outputs(4350) <= a;
    layer7_outputs(4351) <= a or b;
    layer7_outputs(4352) <= not b;
    layer7_outputs(4353) <= a;
    layer7_outputs(4354) <= a and b;
    layer7_outputs(4355) <= not b;
    layer7_outputs(4356) <= b;
    layer7_outputs(4357) <= not (a xor b);
    layer7_outputs(4358) <= b;
    layer7_outputs(4359) <= a and b;
    layer7_outputs(4360) <= a;
    layer7_outputs(4361) <= b;
    layer7_outputs(4362) <= not a;
    layer7_outputs(4363) <= not (a xor b);
    layer7_outputs(4364) <= not (a and b);
    layer7_outputs(4365) <= not (a or b);
    layer7_outputs(4366) <= a xor b;
    layer7_outputs(4367) <= b;
    layer7_outputs(4368) <= a and not b;
    layer7_outputs(4369) <= not (a and b);
    layer7_outputs(4370) <= a;
    layer7_outputs(4371) <= not b;
    layer7_outputs(4372) <= not (a and b);
    layer7_outputs(4373) <= not a;
    layer7_outputs(4374) <= not b or a;
    layer7_outputs(4375) <= b;
    layer7_outputs(4376) <= not b or a;
    layer7_outputs(4377) <= a or b;
    layer7_outputs(4378) <= not b;
    layer7_outputs(4379) <= not b;
    layer7_outputs(4380) <= not a or b;
    layer7_outputs(4381) <= b;
    layer7_outputs(4382) <= b;
    layer7_outputs(4383) <= b;
    layer7_outputs(4384) <= a;
    layer7_outputs(4385) <= not (a or b);
    layer7_outputs(4386) <= not (a xor b);
    layer7_outputs(4387) <= a and not b;
    layer7_outputs(4388) <= not (a xor b);
    layer7_outputs(4389) <= not b;
    layer7_outputs(4390) <= 1'b1;
    layer7_outputs(4391) <= not a;
    layer7_outputs(4392) <= a and b;
    layer7_outputs(4393) <= b;
    layer7_outputs(4394) <= 1'b1;
    layer7_outputs(4395) <= not a or b;
    layer7_outputs(4396) <= not (a xor b);
    layer7_outputs(4397) <= a;
    layer7_outputs(4398) <= not a or b;
    layer7_outputs(4399) <= not (a and b);
    layer7_outputs(4400) <= not a or b;
    layer7_outputs(4401) <= not (a xor b);
    layer7_outputs(4402) <= not b or a;
    layer7_outputs(4403) <= not (a and b);
    layer7_outputs(4404) <= not (a or b);
    layer7_outputs(4405) <= not a or b;
    layer7_outputs(4406) <= a and b;
    layer7_outputs(4407) <= not b;
    layer7_outputs(4408) <= b;
    layer7_outputs(4409) <= not a or b;
    layer7_outputs(4410) <= b;
    layer7_outputs(4411) <= not b;
    layer7_outputs(4412) <= not (a xor b);
    layer7_outputs(4413) <= a;
    layer7_outputs(4414) <= not a;
    layer7_outputs(4415) <= not b;
    layer7_outputs(4416) <= not (a xor b);
    layer7_outputs(4417) <= not a;
    layer7_outputs(4418) <= not b;
    layer7_outputs(4419) <= not (a xor b);
    layer7_outputs(4420) <= not b;
    layer7_outputs(4421) <= a xor b;
    layer7_outputs(4422) <= a xor b;
    layer7_outputs(4423) <= a or b;
    layer7_outputs(4424) <= not (a and b);
    layer7_outputs(4425) <= a xor b;
    layer7_outputs(4426) <= not (a xor b);
    layer7_outputs(4427) <= b and not a;
    layer7_outputs(4428) <= not a or b;
    layer7_outputs(4429) <= not a;
    layer7_outputs(4430) <= not (a xor b);
    layer7_outputs(4431) <= not a or b;
    layer7_outputs(4432) <= a or b;
    layer7_outputs(4433) <= not a;
    layer7_outputs(4434) <= not b;
    layer7_outputs(4435) <= b;
    layer7_outputs(4436) <= a;
    layer7_outputs(4437) <= not b or a;
    layer7_outputs(4438) <= not (a xor b);
    layer7_outputs(4439) <= a xor b;
    layer7_outputs(4440) <= a or b;
    layer7_outputs(4441) <= a xor b;
    layer7_outputs(4442) <= a xor b;
    layer7_outputs(4443) <= b;
    layer7_outputs(4444) <= b;
    layer7_outputs(4445) <= not a;
    layer7_outputs(4446) <= not b;
    layer7_outputs(4447) <= not (a or b);
    layer7_outputs(4448) <= not b;
    layer7_outputs(4449) <= not a;
    layer7_outputs(4450) <= not (a xor b);
    layer7_outputs(4451) <= not b;
    layer7_outputs(4452) <= not b;
    layer7_outputs(4453) <= a or b;
    layer7_outputs(4454) <= a;
    layer7_outputs(4455) <= not (a xor b);
    layer7_outputs(4456) <= not (a xor b);
    layer7_outputs(4457) <= b;
    layer7_outputs(4458) <= not a or b;
    layer7_outputs(4459) <= 1'b0;
    layer7_outputs(4460) <= not (a xor b);
    layer7_outputs(4461) <= not b;
    layer7_outputs(4462) <= a;
    layer7_outputs(4463) <= a xor b;
    layer7_outputs(4464) <= a;
    layer7_outputs(4465) <= not a;
    layer7_outputs(4466) <= b;
    layer7_outputs(4467) <= a or b;
    layer7_outputs(4468) <= a xor b;
    layer7_outputs(4469) <= not (a and b);
    layer7_outputs(4470) <= 1'b1;
    layer7_outputs(4471) <= not a or b;
    layer7_outputs(4472) <= a xor b;
    layer7_outputs(4473) <= a;
    layer7_outputs(4474) <= not b;
    layer7_outputs(4475) <= b;
    layer7_outputs(4476) <= not a;
    layer7_outputs(4477) <= b;
    layer7_outputs(4478) <= not (a or b);
    layer7_outputs(4479) <= not (a xor b);
    layer7_outputs(4480) <= not (a or b);
    layer7_outputs(4481) <= a;
    layer7_outputs(4482) <= a;
    layer7_outputs(4483) <= not a or b;
    layer7_outputs(4484) <= not b or a;
    layer7_outputs(4485) <= not a;
    layer7_outputs(4486) <= b;
    layer7_outputs(4487) <= not a;
    layer7_outputs(4488) <= not a or b;
    layer7_outputs(4489) <= b;
    layer7_outputs(4490) <= not (a and b);
    layer7_outputs(4491) <= not (a xor b);
    layer7_outputs(4492) <= not a or b;
    layer7_outputs(4493) <= a;
    layer7_outputs(4494) <= a and not b;
    layer7_outputs(4495) <= not b;
    layer7_outputs(4496) <= not (a or b);
    layer7_outputs(4497) <= b and not a;
    layer7_outputs(4498) <= not b;
    layer7_outputs(4499) <= a or b;
    layer7_outputs(4500) <= 1'b1;
    layer7_outputs(4501) <= not (a or b);
    layer7_outputs(4502) <= not b or a;
    layer7_outputs(4503) <= not (a xor b);
    layer7_outputs(4504) <= a;
    layer7_outputs(4505) <= not b;
    layer7_outputs(4506) <= a and not b;
    layer7_outputs(4507) <= a xor b;
    layer7_outputs(4508) <= b;
    layer7_outputs(4509) <= not a;
    layer7_outputs(4510) <= b;
    layer7_outputs(4511) <= b;
    layer7_outputs(4512) <= a;
    layer7_outputs(4513) <= not b;
    layer7_outputs(4514) <= a;
    layer7_outputs(4515) <= not (a or b);
    layer7_outputs(4516) <= not a;
    layer7_outputs(4517) <= not b;
    layer7_outputs(4518) <= b and not a;
    layer7_outputs(4519) <= a;
    layer7_outputs(4520) <= not b;
    layer7_outputs(4521) <= a xor b;
    layer7_outputs(4522) <= not (a and b);
    layer7_outputs(4523) <= b;
    layer7_outputs(4524) <= b;
    layer7_outputs(4525) <= not (a and b);
    layer7_outputs(4526) <= not a;
    layer7_outputs(4527) <= b and not a;
    layer7_outputs(4528) <= not a;
    layer7_outputs(4529) <= a and b;
    layer7_outputs(4530) <= not a or b;
    layer7_outputs(4531) <= not (a xor b);
    layer7_outputs(4532) <= b;
    layer7_outputs(4533) <= b;
    layer7_outputs(4534) <= not a;
    layer7_outputs(4535) <= a;
    layer7_outputs(4536) <= not (a and b);
    layer7_outputs(4537) <= a or b;
    layer7_outputs(4538) <= not a or b;
    layer7_outputs(4539) <= a and b;
    layer7_outputs(4540) <= not a;
    layer7_outputs(4541) <= a or b;
    layer7_outputs(4542) <= not (a and b);
    layer7_outputs(4543) <= not a;
    layer7_outputs(4544) <= not (a and b);
    layer7_outputs(4545) <= not a;
    layer7_outputs(4546) <= not (a or b);
    layer7_outputs(4547) <= not a or b;
    layer7_outputs(4548) <= a xor b;
    layer7_outputs(4549) <= not (a xor b);
    layer7_outputs(4550) <= not a or b;
    layer7_outputs(4551) <= not (a xor b);
    layer7_outputs(4552) <= a xor b;
    layer7_outputs(4553) <= b and not a;
    layer7_outputs(4554) <= b and not a;
    layer7_outputs(4555) <= not b or a;
    layer7_outputs(4556) <= b;
    layer7_outputs(4557) <= a;
    layer7_outputs(4558) <= a xor b;
    layer7_outputs(4559) <= a;
    layer7_outputs(4560) <= b and not a;
    layer7_outputs(4561) <= a and b;
    layer7_outputs(4562) <= not b or a;
    layer7_outputs(4563) <= not a;
    layer7_outputs(4564) <= b and not a;
    layer7_outputs(4565) <= not b;
    layer7_outputs(4566) <= not b;
    layer7_outputs(4567) <= not b;
    layer7_outputs(4568) <= a or b;
    layer7_outputs(4569) <= b;
    layer7_outputs(4570) <= not a;
    layer7_outputs(4571) <= not (a and b);
    layer7_outputs(4572) <= not a;
    layer7_outputs(4573) <= not a;
    layer7_outputs(4574) <= b;
    layer7_outputs(4575) <= b;
    layer7_outputs(4576) <= not b;
    layer7_outputs(4577) <= not a or b;
    layer7_outputs(4578) <= not (a xor b);
    layer7_outputs(4579) <= a;
    layer7_outputs(4580) <= not b;
    layer7_outputs(4581) <= not b;
    layer7_outputs(4582) <= not (a or b);
    layer7_outputs(4583) <= a and not b;
    layer7_outputs(4584) <= a;
    layer7_outputs(4585) <= not b;
    layer7_outputs(4586) <= 1'b1;
    layer7_outputs(4587) <= not a;
    layer7_outputs(4588) <= a;
    layer7_outputs(4589) <= b;
    layer7_outputs(4590) <= a;
    layer7_outputs(4591) <= a;
    layer7_outputs(4592) <= a xor b;
    layer7_outputs(4593) <= a or b;
    layer7_outputs(4594) <= not b or a;
    layer7_outputs(4595) <= b;
    layer7_outputs(4596) <= not a;
    layer7_outputs(4597) <= not a;
    layer7_outputs(4598) <= not a;
    layer7_outputs(4599) <= a and not b;
    layer7_outputs(4600) <= a;
    layer7_outputs(4601) <= a xor b;
    layer7_outputs(4602) <= not a;
    layer7_outputs(4603) <= not (a or b);
    layer7_outputs(4604) <= a or b;
    layer7_outputs(4605) <= a;
    layer7_outputs(4606) <= not a;
    layer7_outputs(4607) <= not a;
    layer7_outputs(4608) <= a;
    layer7_outputs(4609) <= a;
    layer7_outputs(4610) <= not a;
    layer7_outputs(4611) <= not a;
    layer7_outputs(4612) <= not b;
    layer7_outputs(4613) <= not (a and b);
    layer7_outputs(4614) <= a xor b;
    layer7_outputs(4615) <= a and not b;
    layer7_outputs(4616) <= a xor b;
    layer7_outputs(4617) <= not b;
    layer7_outputs(4618) <= a;
    layer7_outputs(4619) <= 1'b1;
    layer7_outputs(4620) <= b;
    layer7_outputs(4621) <= 1'b0;
    layer7_outputs(4622) <= a or b;
    layer7_outputs(4623) <= a and not b;
    layer7_outputs(4624) <= not (a and b);
    layer7_outputs(4625) <= not b;
    layer7_outputs(4626) <= not b;
    layer7_outputs(4627) <= a xor b;
    layer7_outputs(4628) <= b;
    layer7_outputs(4629) <= a or b;
    layer7_outputs(4630) <= b;
    layer7_outputs(4631) <= a xor b;
    layer7_outputs(4632) <= not b;
    layer7_outputs(4633) <= a and b;
    layer7_outputs(4634) <= not a;
    layer7_outputs(4635) <= not (a xor b);
    layer7_outputs(4636) <= not a or b;
    layer7_outputs(4637) <= not b;
    layer7_outputs(4638) <= not b;
    layer7_outputs(4639) <= a;
    layer7_outputs(4640) <= not a;
    layer7_outputs(4641) <= a;
    layer7_outputs(4642) <= b;
    layer7_outputs(4643) <= a;
    layer7_outputs(4644) <= not b;
    layer7_outputs(4645) <= a and b;
    layer7_outputs(4646) <= not (a xor b);
    layer7_outputs(4647) <= b;
    layer7_outputs(4648) <= a xor b;
    layer7_outputs(4649) <= not b;
    layer7_outputs(4650) <= not (a and b);
    layer7_outputs(4651) <= not b or a;
    layer7_outputs(4652) <= not (a and b);
    layer7_outputs(4653) <= b;
    layer7_outputs(4654) <= a and b;
    layer7_outputs(4655) <= a and not b;
    layer7_outputs(4656) <= not b;
    layer7_outputs(4657) <= not a;
    layer7_outputs(4658) <= a xor b;
    layer7_outputs(4659) <= not a;
    layer7_outputs(4660) <= b and not a;
    layer7_outputs(4661) <= b and not a;
    layer7_outputs(4662) <= b;
    layer7_outputs(4663) <= not (a xor b);
    layer7_outputs(4664) <= not b or a;
    layer7_outputs(4665) <= a and not b;
    layer7_outputs(4666) <= not b;
    layer7_outputs(4667) <= b and not a;
    layer7_outputs(4668) <= a;
    layer7_outputs(4669) <= b;
    layer7_outputs(4670) <= not b;
    layer7_outputs(4671) <= b and not a;
    layer7_outputs(4672) <= not (a or b);
    layer7_outputs(4673) <= b;
    layer7_outputs(4674) <= not a;
    layer7_outputs(4675) <= not (a or b);
    layer7_outputs(4676) <= not a;
    layer7_outputs(4677) <= not b or a;
    layer7_outputs(4678) <= a and not b;
    layer7_outputs(4679) <= not a or b;
    layer7_outputs(4680) <= not b or a;
    layer7_outputs(4681) <= b;
    layer7_outputs(4682) <= not b or a;
    layer7_outputs(4683) <= not (a xor b);
    layer7_outputs(4684) <= a and not b;
    layer7_outputs(4685) <= a;
    layer7_outputs(4686) <= not a;
    layer7_outputs(4687) <= b;
    layer7_outputs(4688) <= not a;
    layer7_outputs(4689) <= a and b;
    layer7_outputs(4690) <= not a;
    layer7_outputs(4691) <= a xor b;
    layer7_outputs(4692) <= b;
    layer7_outputs(4693) <= a xor b;
    layer7_outputs(4694) <= b and not a;
    layer7_outputs(4695) <= a;
    layer7_outputs(4696) <= not a;
    layer7_outputs(4697) <= not a or b;
    layer7_outputs(4698) <= 1'b0;
    layer7_outputs(4699) <= not b;
    layer7_outputs(4700) <= not b;
    layer7_outputs(4701) <= not a or b;
    layer7_outputs(4702) <= not a or b;
    layer7_outputs(4703) <= not (a xor b);
    layer7_outputs(4704) <= not b;
    layer7_outputs(4705) <= not a;
    layer7_outputs(4706) <= a or b;
    layer7_outputs(4707) <= b;
    layer7_outputs(4708) <= not (a and b);
    layer7_outputs(4709) <= not a or b;
    layer7_outputs(4710) <= a;
    layer7_outputs(4711) <= not b;
    layer7_outputs(4712) <= not (a xor b);
    layer7_outputs(4713) <= a and not b;
    layer7_outputs(4714) <= a xor b;
    layer7_outputs(4715) <= 1'b0;
    layer7_outputs(4716) <= not (a xor b);
    layer7_outputs(4717) <= not a;
    layer7_outputs(4718) <= not a or b;
    layer7_outputs(4719) <= not b;
    layer7_outputs(4720) <= a;
    layer7_outputs(4721) <= not b;
    layer7_outputs(4722) <= not (a xor b);
    layer7_outputs(4723) <= not (a and b);
    layer7_outputs(4724) <= not a;
    layer7_outputs(4725) <= a;
    layer7_outputs(4726) <= a xor b;
    layer7_outputs(4727) <= not (a xor b);
    layer7_outputs(4728) <= b;
    layer7_outputs(4729) <= not a;
    layer7_outputs(4730) <= a and b;
    layer7_outputs(4731) <= not (a or b);
    layer7_outputs(4732) <= a xor b;
    layer7_outputs(4733) <= not a;
    layer7_outputs(4734) <= not b;
    layer7_outputs(4735) <= not b;
    layer7_outputs(4736) <= b and not a;
    layer7_outputs(4737) <= b;
    layer7_outputs(4738) <= not (a and b);
    layer7_outputs(4739) <= not (a xor b);
    layer7_outputs(4740) <= a and not b;
    layer7_outputs(4741) <= b;
    layer7_outputs(4742) <= b;
    layer7_outputs(4743) <= a;
    layer7_outputs(4744) <= a and b;
    layer7_outputs(4745) <= not b or a;
    layer7_outputs(4746) <= not a or b;
    layer7_outputs(4747) <= not (a xor b);
    layer7_outputs(4748) <= not a;
    layer7_outputs(4749) <= not (a and b);
    layer7_outputs(4750) <= a;
    layer7_outputs(4751) <= not b;
    layer7_outputs(4752) <= b;
    layer7_outputs(4753) <= not b;
    layer7_outputs(4754) <= b;
    layer7_outputs(4755) <= not a;
    layer7_outputs(4756) <= a;
    layer7_outputs(4757) <= not a;
    layer7_outputs(4758) <= a xor b;
    layer7_outputs(4759) <= not b;
    layer7_outputs(4760) <= not a;
    layer7_outputs(4761) <= 1'b0;
    layer7_outputs(4762) <= not b;
    layer7_outputs(4763) <= not a;
    layer7_outputs(4764) <= not (a and b);
    layer7_outputs(4765) <= a xor b;
    layer7_outputs(4766) <= a xor b;
    layer7_outputs(4767) <= not a;
    layer7_outputs(4768) <= a and b;
    layer7_outputs(4769) <= a or b;
    layer7_outputs(4770) <= a;
    layer7_outputs(4771) <= b;
    layer7_outputs(4772) <= not (a or b);
    layer7_outputs(4773) <= a or b;
    layer7_outputs(4774) <= a or b;
    layer7_outputs(4775) <= b;
    layer7_outputs(4776) <= not a or b;
    layer7_outputs(4777) <= not a or b;
    layer7_outputs(4778) <= 1'b1;
    layer7_outputs(4779) <= a;
    layer7_outputs(4780) <= a;
    layer7_outputs(4781) <= not a or b;
    layer7_outputs(4782) <= b and not a;
    layer7_outputs(4783) <= a and not b;
    layer7_outputs(4784) <= a xor b;
    layer7_outputs(4785) <= a or b;
    layer7_outputs(4786) <= a and b;
    layer7_outputs(4787) <= not (a xor b);
    layer7_outputs(4788) <= a and b;
    layer7_outputs(4789) <= a xor b;
    layer7_outputs(4790) <= not b;
    layer7_outputs(4791) <= not a;
    layer7_outputs(4792) <= not a;
    layer7_outputs(4793) <= not (a and b);
    layer7_outputs(4794) <= a and not b;
    layer7_outputs(4795) <= a or b;
    layer7_outputs(4796) <= b and not a;
    layer7_outputs(4797) <= a;
    layer7_outputs(4798) <= not (a xor b);
    layer7_outputs(4799) <= a xor b;
    layer7_outputs(4800) <= not b;
    layer7_outputs(4801) <= not (a or b);
    layer7_outputs(4802) <= not a;
    layer7_outputs(4803) <= b;
    layer7_outputs(4804) <= a xor b;
    layer7_outputs(4805) <= a and b;
    layer7_outputs(4806) <= b;
    layer7_outputs(4807) <= not (a xor b);
    layer7_outputs(4808) <= not (a and b);
    layer7_outputs(4809) <= not b or a;
    layer7_outputs(4810) <= b and not a;
    layer7_outputs(4811) <= a;
    layer7_outputs(4812) <= a;
    layer7_outputs(4813) <= a and b;
    layer7_outputs(4814) <= a;
    layer7_outputs(4815) <= a xor b;
    layer7_outputs(4816) <= not a;
    layer7_outputs(4817) <= a;
    layer7_outputs(4818) <= b;
    layer7_outputs(4819) <= not a;
    layer7_outputs(4820) <= not a;
    layer7_outputs(4821) <= a and b;
    layer7_outputs(4822) <= a and b;
    layer7_outputs(4823) <= 1'b1;
    layer7_outputs(4824) <= b and not a;
    layer7_outputs(4825) <= a and not b;
    layer7_outputs(4826) <= a;
    layer7_outputs(4827) <= not a;
    layer7_outputs(4828) <= a and b;
    layer7_outputs(4829) <= not a;
    layer7_outputs(4830) <= not b;
    layer7_outputs(4831) <= b;
    layer7_outputs(4832) <= not b or a;
    layer7_outputs(4833) <= not a;
    layer7_outputs(4834) <= a or b;
    layer7_outputs(4835) <= not b or a;
    layer7_outputs(4836) <= b;
    layer7_outputs(4837) <= not a;
    layer7_outputs(4838) <= not b;
    layer7_outputs(4839) <= a or b;
    layer7_outputs(4840) <= not b;
    layer7_outputs(4841) <= 1'b0;
    layer7_outputs(4842) <= a;
    layer7_outputs(4843) <= b and not a;
    layer7_outputs(4844) <= a and not b;
    layer7_outputs(4845) <= b;
    layer7_outputs(4846) <= b and not a;
    layer7_outputs(4847) <= a and b;
    layer7_outputs(4848) <= a;
    layer7_outputs(4849) <= a xor b;
    layer7_outputs(4850) <= b;
    layer7_outputs(4851) <= a;
    layer7_outputs(4852) <= a or b;
    layer7_outputs(4853) <= 1'b1;
    layer7_outputs(4854) <= not a;
    layer7_outputs(4855) <= not a or b;
    layer7_outputs(4856) <= not (a xor b);
    layer7_outputs(4857) <= not a or b;
    layer7_outputs(4858) <= a xor b;
    layer7_outputs(4859) <= a;
    layer7_outputs(4860) <= 1'b1;
    layer7_outputs(4861) <= not (a or b);
    layer7_outputs(4862) <= not (a xor b);
    layer7_outputs(4863) <= not (a and b);
    layer7_outputs(4864) <= a or b;
    layer7_outputs(4865) <= not b;
    layer7_outputs(4866) <= not a;
    layer7_outputs(4867) <= not a or b;
    layer7_outputs(4868) <= not (a xor b);
    layer7_outputs(4869) <= a;
    layer7_outputs(4870) <= not b;
    layer7_outputs(4871) <= not b;
    layer7_outputs(4872) <= a and not b;
    layer7_outputs(4873) <= not (a xor b);
    layer7_outputs(4874) <= a xor b;
    layer7_outputs(4875) <= not b or a;
    layer7_outputs(4876) <= not a or b;
    layer7_outputs(4877) <= not a;
    layer7_outputs(4878) <= not (a xor b);
    layer7_outputs(4879) <= not (a xor b);
    layer7_outputs(4880) <= not (a xor b);
    layer7_outputs(4881) <= a and not b;
    layer7_outputs(4882) <= a and not b;
    layer7_outputs(4883) <= a and b;
    layer7_outputs(4884) <= b;
    layer7_outputs(4885) <= not b;
    layer7_outputs(4886) <= not (a and b);
    layer7_outputs(4887) <= b and not a;
    layer7_outputs(4888) <= a and not b;
    layer7_outputs(4889) <= not b;
    layer7_outputs(4890) <= not a;
    layer7_outputs(4891) <= a xor b;
    layer7_outputs(4892) <= not (a xor b);
    layer7_outputs(4893) <= not (a or b);
    layer7_outputs(4894) <= a and b;
    layer7_outputs(4895) <= a;
    layer7_outputs(4896) <= not a or b;
    layer7_outputs(4897) <= a;
    layer7_outputs(4898) <= not (a xor b);
    layer7_outputs(4899) <= not a;
    layer7_outputs(4900) <= not a;
    layer7_outputs(4901) <= not a;
    layer7_outputs(4902) <= b;
    layer7_outputs(4903) <= a;
    layer7_outputs(4904) <= not b or a;
    layer7_outputs(4905) <= not (a xor b);
    layer7_outputs(4906) <= not a or b;
    layer7_outputs(4907) <= b;
    layer7_outputs(4908) <= b and not a;
    layer7_outputs(4909) <= a xor b;
    layer7_outputs(4910) <= a xor b;
    layer7_outputs(4911) <= b;
    layer7_outputs(4912) <= b;
    layer7_outputs(4913) <= a;
    layer7_outputs(4914) <= b;
    layer7_outputs(4915) <= not (a or b);
    layer7_outputs(4916) <= not b or a;
    layer7_outputs(4917) <= not (a or b);
    layer7_outputs(4918) <= not (a xor b);
    layer7_outputs(4919) <= not a;
    layer7_outputs(4920) <= not a or b;
    layer7_outputs(4921) <= not a or b;
    layer7_outputs(4922) <= not a;
    layer7_outputs(4923) <= not (a or b);
    layer7_outputs(4924) <= b;
    layer7_outputs(4925) <= not a;
    layer7_outputs(4926) <= a or b;
    layer7_outputs(4927) <= b and not a;
    layer7_outputs(4928) <= not (a and b);
    layer7_outputs(4929) <= not b;
    layer7_outputs(4930) <= b;
    layer7_outputs(4931) <= not b;
    layer7_outputs(4932) <= a;
    layer7_outputs(4933) <= a and b;
    layer7_outputs(4934) <= not a;
    layer7_outputs(4935) <= not a or b;
    layer7_outputs(4936) <= not a or b;
    layer7_outputs(4937) <= a;
    layer7_outputs(4938) <= b;
    layer7_outputs(4939) <= not a;
    layer7_outputs(4940) <= b and not a;
    layer7_outputs(4941) <= not a;
    layer7_outputs(4942) <= a;
    layer7_outputs(4943) <= not a or b;
    layer7_outputs(4944) <= b;
    layer7_outputs(4945) <= not a;
    layer7_outputs(4946) <= not (a xor b);
    layer7_outputs(4947) <= a;
    layer7_outputs(4948) <= not a;
    layer7_outputs(4949) <= not a or b;
    layer7_outputs(4950) <= not a;
    layer7_outputs(4951) <= not a or b;
    layer7_outputs(4952) <= not a or b;
    layer7_outputs(4953) <= not (a and b);
    layer7_outputs(4954) <= b and not a;
    layer7_outputs(4955) <= a xor b;
    layer7_outputs(4956) <= a xor b;
    layer7_outputs(4957) <= not a or b;
    layer7_outputs(4958) <= a;
    layer7_outputs(4959) <= a;
    layer7_outputs(4960) <= a and not b;
    layer7_outputs(4961) <= not (a and b);
    layer7_outputs(4962) <= not (a and b);
    layer7_outputs(4963) <= a;
    layer7_outputs(4964) <= a;
    layer7_outputs(4965) <= not (a and b);
    layer7_outputs(4966) <= not (a and b);
    layer7_outputs(4967) <= a and not b;
    layer7_outputs(4968) <= a;
    layer7_outputs(4969) <= not (a or b);
    layer7_outputs(4970) <= a xor b;
    layer7_outputs(4971) <= not a or b;
    layer7_outputs(4972) <= a;
    layer7_outputs(4973) <= not b;
    layer7_outputs(4974) <= b;
    layer7_outputs(4975) <= b;
    layer7_outputs(4976) <= b and not a;
    layer7_outputs(4977) <= a;
    layer7_outputs(4978) <= b and not a;
    layer7_outputs(4979) <= a and b;
    layer7_outputs(4980) <= b and not a;
    layer7_outputs(4981) <= not a;
    layer7_outputs(4982) <= a and not b;
    layer7_outputs(4983) <= b and not a;
    layer7_outputs(4984) <= not b;
    layer7_outputs(4985) <= a;
    layer7_outputs(4986) <= not b;
    layer7_outputs(4987) <= not a;
    layer7_outputs(4988) <= a;
    layer7_outputs(4989) <= not b or a;
    layer7_outputs(4990) <= a xor b;
    layer7_outputs(4991) <= not (a and b);
    layer7_outputs(4992) <= not b or a;
    layer7_outputs(4993) <= not (a and b);
    layer7_outputs(4994) <= a xor b;
    layer7_outputs(4995) <= not a;
    layer7_outputs(4996) <= not a;
    layer7_outputs(4997) <= b and not a;
    layer7_outputs(4998) <= b and not a;
    layer7_outputs(4999) <= not (a and b);
    layer7_outputs(5000) <= b;
    layer7_outputs(5001) <= b and not a;
    layer7_outputs(5002) <= not (a or b);
    layer7_outputs(5003) <= a and b;
    layer7_outputs(5004) <= not (a or b);
    layer7_outputs(5005) <= b;
    layer7_outputs(5006) <= a;
    layer7_outputs(5007) <= not a or b;
    layer7_outputs(5008) <= b;
    layer7_outputs(5009) <= b and not a;
    layer7_outputs(5010) <= a xor b;
    layer7_outputs(5011) <= a;
    layer7_outputs(5012) <= 1'b1;
    layer7_outputs(5013) <= not (a xor b);
    layer7_outputs(5014) <= a xor b;
    layer7_outputs(5015) <= not (a and b);
    layer7_outputs(5016) <= not a;
    layer7_outputs(5017) <= not (a xor b);
    layer7_outputs(5018) <= 1'b1;
    layer7_outputs(5019) <= not (a and b);
    layer7_outputs(5020) <= a xor b;
    layer7_outputs(5021) <= not a;
    layer7_outputs(5022) <= not b;
    layer7_outputs(5023) <= not b or a;
    layer7_outputs(5024) <= not (a or b);
    layer7_outputs(5025) <= not b or a;
    layer7_outputs(5026) <= a or b;
    layer7_outputs(5027) <= not b or a;
    layer7_outputs(5028) <= not b;
    layer7_outputs(5029) <= a or b;
    layer7_outputs(5030) <= b;
    layer7_outputs(5031) <= not (a xor b);
    layer7_outputs(5032) <= a and not b;
    layer7_outputs(5033) <= b;
    layer7_outputs(5034) <= not b;
    layer7_outputs(5035) <= a or b;
    layer7_outputs(5036) <= not b;
    layer7_outputs(5037) <= not (a and b);
    layer7_outputs(5038) <= a;
    layer7_outputs(5039) <= b;
    layer7_outputs(5040) <= not b or a;
    layer7_outputs(5041) <= not a;
    layer7_outputs(5042) <= not a;
    layer7_outputs(5043) <= b;
    layer7_outputs(5044) <= not (a xor b);
    layer7_outputs(5045) <= not (a xor b);
    layer7_outputs(5046) <= a or b;
    layer7_outputs(5047) <= not a;
    layer7_outputs(5048) <= not b;
    layer7_outputs(5049) <= b;
    layer7_outputs(5050) <= not (a xor b);
    layer7_outputs(5051) <= not (a xor b);
    layer7_outputs(5052) <= a and b;
    layer7_outputs(5053) <= not a;
    layer7_outputs(5054) <= a and not b;
    layer7_outputs(5055) <= not (a or b);
    layer7_outputs(5056) <= not (a or b);
    layer7_outputs(5057) <= a xor b;
    layer7_outputs(5058) <= b;
    layer7_outputs(5059) <= not a or b;
    layer7_outputs(5060) <= not (a xor b);
    layer7_outputs(5061) <= not b;
    layer7_outputs(5062) <= b;
    layer7_outputs(5063) <= not (a xor b);
    layer7_outputs(5064) <= not b;
    layer7_outputs(5065) <= b;
    layer7_outputs(5066) <= not b or a;
    layer7_outputs(5067) <= not (a xor b);
    layer7_outputs(5068) <= not b;
    layer7_outputs(5069) <= b and not a;
    layer7_outputs(5070) <= not (a or b);
    layer7_outputs(5071) <= not a;
    layer7_outputs(5072) <= not (a or b);
    layer7_outputs(5073) <= not a;
    layer7_outputs(5074) <= b;
    layer7_outputs(5075) <= a;
    layer7_outputs(5076) <= b and not a;
    layer7_outputs(5077) <= b;
    layer7_outputs(5078) <= not (a xor b);
    layer7_outputs(5079) <= not a;
    layer7_outputs(5080) <= not a;
    layer7_outputs(5081) <= a and b;
    layer7_outputs(5082) <= a;
    layer7_outputs(5083) <= not b;
    layer7_outputs(5084) <= not (a and b);
    layer7_outputs(5085) <= not a;
    layer7_outputs(5086) <= not (a xor b);
    layer7_outputs(5087) <= a and not b;
    layer7_outputs(5088) <= not a;
    layer7_outputs(5089) <= 1'b0;
    layer7_outputs(5090) <= not (a or b);
    layer7_outputs(5091) <= not b;
    layer7_outputs(5092) <= a;
    layer7_outputs(5093) <= not (a xor b);
    layer7_outputs(5094) <= not b;
    layer7_outputs(5095) <= a;
    layer7_outputs(5096) <= not a;
    layer7_outputs(5097) <= a;
    layer7_outputs(5098) <= not (a and b);
    layer7_outputs(5099) <= not b or a;
    layer7_outputs(5100) <= a or b;
    layer7_outputs(5101) <= a xor b;
    layer7_outputs(5102) <= a;
    layer7_outputs(5103) <= a xor b;
    layer7_outputs(5104) <= not (a xor b);
    layer7_outputs(5105) <= 1'b1;
    layer7_outputs(5106) <= not a;
    layer7_outputs(5107) <= b;
    layer7_outputs(5108) <= b;
    layer7_outputs(5109) <= b;
    layer7_outputs(5110) <= b;
    layer7_outputs(5111) <= b;
    layer7_outputs(5112) <= b and not a;
    layer7_outputs(5113) <= not b;
    layer7_outputs(5114) <= not a;
    layer7_outputs(5115) <= not (a xor b);
    layer7_outputs(5116) <= not a;
    layer7_outputs(5117) <= not (a and b);
    layer7_outputs(5118) <= not (a xor b);
    layer7_outputs(5119) <= not (a and b);
    layer7_outputs(5120) <= b and not a;
    layer7_outputs(5121) <= b;
    layer7_outputs(5122) <= b and not a;
    layer7_outputs(5123) <= 1'b1;
    layer7_outputs(5124) <= b and not a;
    layer7_outputs(5125) <= not a;
    layer7_outputs(5126) <= a and not b;
    layer7_outputs(5127) <= not (a or b);
    layer7_outputs(5128) <= not a;
    layer7_outputs(5129) <= not (a xor b);
    layer7_outputs(5130) <= b and not a;
    layer7_outputs(5131) <= not b;
    layer7_outputs(5132) <= not a or b;
    layer7_outputs(5133) <= not (a and b);
    layer7_outputs(5134) <= not (a xor b);
    layer7_outputs(5135) <= not a;
    layer7_outputs(5136) <= a and b;
    layer7_outputs(5137) <= not (a and b);
    layer7_outputs(5138) <= a and b;
    layer7_outputs(5139) <= a and not b;
    layer7_outputs(5140) <= not b;
    layer7_outputs(5141) <= b;
    layer7_outputs(5142) <= not (a and b);
    layer7_outputs(5143) <= not b;
    layer7_outputs(5144) <= not b or a;
    layer7_outputs(5145) <= 1'b1;
    layer7_outputs(5146) <= not b;
    layer7_outputs(5147) <= not (a or b);
    layer7_outputs(5148) <= 1'b1;
    layer7_outputs(5149) <= a xor b;
    layer7_outputs(5150) <= b;
    layer7_outputs(5151) <= a and b;
    layer7_outputs(5152) <= a and not b;
    layer7_outputs(5153) <= not a or b;
    layer7_outputs(5154) <= not (a or b);
    layer7_outputs(5155) <= a xor b;
    layer7_outputs(5156) <= not (a xor b);
    layer7_outputs(5157) <= not (a or b);
    layer7_outputs(5158) <= a;
    layer7_outputs(5159) <= a;
    layer7_outputs(5160) <= not b;
    layer7_outputs(5161) <= not (a xor b);
    layer7_outputs(5162) <= a xor b;
    layer7_outputs(5163) <= not b;
    layer7_outputs(5164) <= not a;
    layer7_outputs(5165) <= a xor b;
    layer7_outputs(5166) <= not a;
    layer7_outputs(5167) <= not a;
    layer7_outputs(5168) <= not b;
    layer7_outputs(5169) <= not b;
    layer7_outputs(5170) <= not b or a;
    layer7_outputs(5171) <= a;
    layer7_outputs(5172) <= a xor b;
    layer7_outputs(5173) <= not b;
    layer7_outputs(5174) <= b and not a;
    layer7_outputs(5175) <= b;
    layer7_outputs(5176) <= not b;
    layer7_outputs(5177) <= not b;
    layer7_outputs(5178) <= not (a or b);
    layer7_outputs(5179) <= a xor b;
    layer7_outputs(5180) <= not (a and b);
    layer7_outputs(5181) <= not b or a;
    layer7_outputs(5182) <= a;
    layer7_outputs(5183) <= not (a and b);
    layer7_outputs(5184) <= b and not a;
    layer7_outputs(5185) <= not (a and b);
    layer7_outputs(5186) <= a or b;
    layer7_outputs(5187) <= not (a and b);
    layer7_outputs(5188) <= not b;
    layer7_outputs(5189) <= a;
    layer7_outputs(5190) <= not (a or b);
    layer7_outputs(5191) <= b;
    layer7_outputs(5192) <= not b or a;
    layer7_outputs(5193) <= a xor b;
    layer7_outputs(5194) <= a or b;
    layer7_outputs(5195) <= not a or b;
    layer7_outputs(5196) <= not b;
    layer7_outputs(5197) <= a and b;
    layer7_outputs(5198) <= not a;
    layer7_outputs(5199) <= not b or a;
    layer7_outputs(5200) <= not (a or b);
    layer7_outputs(5201) <= a;
    layer7_outputs(5202) <= a;
    layer7_outputs(5203) <= b and not a;
    layer7_outputs(5204) <= not b or a;
    layer7_outputs(5205) <= a or b;
    layer7_outputs(5206) <= not b;
    layer7_outputs(5207) <= a or b;
    layer7_outputs(5208) <= b;
    layer7_outputs(5209) <= not b;
    layer7_outputs(5210) <= not (a xor b);
    layer7_outputs(5211) <= 1'b0;
    layer7_outputs(5212) <= b;
    layer7_outputs(5213) <= a and not b;
    layer7_outputs(5214) <= not a or b;
    layer7_outputs(5215) <= a and b;
    layer7_outputs(5216) <= not (a or b);
    layer7_outputs(5217) <= b;
    layer7_outputs(5218) <= a or b;
    layer7_outputs(5219) <= not b;
    layer7_outputs(5220) <= a and not b;
    layer7_outputs(5221) <= not b;
    layer7_outputs(5222) <= a xor b;
    layer7_outputs(5223) <= a and not b;
    layer7_outputs(5224) <= not b or a;
    layer7_outputs(5225) <= b;
    layer7_outputs(5226) <= a;
    layer7_outputs(5227) <= a and b;
    layer7_outputs(5228) <= not b or a;
    layer7_outputs(5229) <= not (a xor b);
    layer7_outputs(5230) <= a or b;
    layer7_outputs(5231) <= a;
    layer7_outputs(5232) <= a xor b;
    layer7_outputs(5233) <= a and b;
    layer7_outputs(5234) <= a or b;
    layer7_outputs(5235) <= not (a and b);
    layer7_outputs(5236) <= a or b;
    layer7_outputs(5237) <= not a;
    layer7_outputs(5238) <= b and not a;
    layer7_outputs(5239) <= a and b;
    layer7_outputs(5240) <= not (a and b);
    layer7_outputs(5241) <= not a or b;
    layer7_outputs(5242) <= not b;
    layer7_outputs(5243) <= not (a and b);
    layer7_outputs(5244) <= not a;
    layer7_outputs(5245) <= not (a and b);
    layer7_outputs(5246) <= not b or a;
    layer7_outputs(5247) <= a xor b;
    layer7_outputs(5248) <= b;
    layer7_outputs(5249) <= a;
    layer7_outputs(5250) <= a and b;
    layer7_outputs(5251) <= not b or a;
    layer7_outputs(5252) <= not a;
    layer7_outputs(5253) <= a xor b;
    layer7_outputs(5254) <= not a or b;
    layer7_outputs(5255) <= a;
    layer7_outputs(5256) <= not b or a;
    layer7_outputs(5257) <= a xor b;
    layer7_outputs(5258) <= not (a xor b);
    layer7_outputs(5259) <= not b;
    layer7_outputs(5260) <= not a or b;
    layer7_outputs(5261) <= not (a and b);
    layer7_outputs(5262) <= a;
    layer7_outputs(5263) <= not (a or b);
    layer7_outputs(5264) <= b;
    layer7_outputs(5265) <= b and not a;
    layer7_outputs(5266) <= a and not b;
    layer7_outputs(5267) <= not (a or b);
    layer7_outputs(5268) <= not b or a;
    layer7_outputs(5269) <= b;
    layer7_outputs(5270) <= not (a and b);
    layer7_outputs(5271) <= a;
    layer7_outputs(5272) <= a xor b;
    layer7_outputs(5273) <= not a or b;
    layer7_outputs(5274) <= a xor b;
    layer7_outputs(5275) <= a;
    layer7_outputs(5276) <= not a or b;
    layer7_outputs(5277) <= a;
    layer7_outputs(5278) <= a;
    layer7_outputs(5279) <= a and not b;
    layer7_outputs(5280) <= not b;
    layer7_outputs(5281) <= b and not a;
    layer7_outputs(5282) <= b;
    layer7_outputs(5283) <= not a;
    layer7_outputs(5284) <= 1'b0;
    layer7_outputs(5285) <= not b;
    layer7_outputs(5286) <= not (a or b);
    layer7_outputs(5287) <= a xor b;
    layer7_outputs(5288) <= not (a xor b);
    layer7_outputs(5289) <= not b or a;
    layer7_outputs(5290) <= a xor b;
    layer7_outputs(5291) <= not b;
    layer7_outputs(5292) <= not b or a;
    layer7_outputs(5293) <= a and not b;
    layer7_outputs(5294) <= a or b;
    layer7_outputs(5295) <= a;
    layer7_outputs(5296) <= not (a xor b);
    layer7_outputs(5297) <= not (a or b);
    layer7_outputs(5298) <= not (a or b);
    layer7_outputs(5299) <= a xor b;
    layer7_outputs(5300) <= not (a or b);
    layer7_outputs(5301) <= not a;
    layer7_outputs(5302) <= 1'b0;
    layer7_outputs(5303) <= a xor b;
    layer7_outputs(5304) <= a or b;
    layer7_outputs(5305) <= not (a and b);
    layer7_outputs(5306) <= not a;
    layer7_outputs(5307) <= b;
    layer7_outputs(5308) <= a and not b;
    layer7_outputs(5309) <= a and b;
    layer7_outputs(5310) <= a and b;
    layer7_outputs(5311) <= a xor b;
    layer7_outputs(5312) <= a;
    layer7_outputs(5313) <= not a;
    layer7_outputs(5314) <= a;
    layer7_outputs(5315) <= not (a and b);
    layer7_outputs(5316) <= a;
    layer7_outputs(5317) <= a or b;
    layer7_outputs(5318) <= not (a or b);
    layer7_outputs(5319) <= not a;
    layer7_outputs(5320) <= a xor b;
    layer7_outputs(5321) <= not a;
    layer7_outputs(5322) <= not (a xor b);
    layer7_outputs(5323) <= a and not b;
    layer7_outputs(5324) <= not (a and b);
    layer7_outputs(5325) <= a and b;
    layer7_outputs(5326) <= not b;
    layer7_outputs(5327) <= a and b;
    layer7_outputs(5328) <= a and not b;
    layer7_outputs(5329) <= a and not b;
    layer7_outputs(5330) <= not a;
    layer7_outputs(5331) <= a;
    layer7_outputs(5332) <= a;
    layer7_outputs(5333) <= a and not b;
    layer7_outputs(5334) <= not b or a;
    layer7_outputs(5335) <= b and not a;
    layer7_outputs(5336) <= not (a xor b);
    layer7_outputs(5337) <= b;
    layer7_outputs(5338) <= b;
    layer7_outputs(5339) <= not (a and b);
    layer7_outputs(5340) <= not b;
    layer7_outputs(5341) <= b;
    layer7_outputs(5342) <= a or b;
    layer7_outputs(5343) <= b;
    layer7_outputs(5344) <= a and not b;
    layer7_outputs(5345) <= not b;
    layer7_outputs(5346) <= a and not b;
    layer7_outputs(5347) <= a xor b;
    layer7_outputs(5348) <= a xor b;
    layer7_outputs(5349) <= not (a and b);
    layer7_outputs(5350) <= a xor b;
    layer7_outputs(5351) <= 1'b1;
    layer7_outputs(5352) <= not b or a;
    layer7_outputs(5353) <= not (a and b);
    layer7_outputs(5354) <= b;
    layer7_outputs(5355) <= not a or b;
    layer7_outputs(5356) <= not b or a;
    layer7_outputs(5357) <= not b or a;
    layer7_outputs(5358) <= not b;
    layer7_outputs(5359) <= a or b;
    layer7_outputs(5360) <= not a;
    layer7_outputs(5361) <= not a or b;
    layer7_outputs(5362) <= not b;
    layer7_outputs(5363) <= a;
    layer7_outputs(5364) <= a;
    layer7_outputs(5365) <= a and not b;
    layer7_outputs(5366) <= b;
    layer7_outputs(5367) <= not (a or b);
    layer7_outputs(5368) <= not a;
    layer7_outputs(5369) <= a;
    layer7_outputs(5370) <= a;
    layer7_outputs(5371) <= not (a xor b);
    layer7_outputs(5372) <= a and b;
    layer7_outputs(5373) <= not b;
    layer7_outputs(5374) <= not (a and b);
    layer7_outputs(5375) <= a and not b;
    layer7_outputs(5376) <= not (a xor b);
    layer7_outputs(5377) <= not b;
    layer7_outputs(5378) <= not b;
    layer7_outputs(5379) <= not (a xor b);
    layer7_outputs(5380) <= a and b;
    layer7_outputs(5381) <= b;
    layer7_outputs(5382) <= not (a or b);
    layer7_outputs(5383) <= a;
    layer7_outputs(5384) <= not (a xor b);
    layer7_outputs(5385) <= not b or a;
    layer7_outputs(5386) <= a;
    layer7_outputs(5387) <= not a;
    layer7_outputs(5388) <= b and not a;
    layer7_outputs(5389) <= a xor b;
    layer7_outputs(5390) <= not b;
    layer7_outputs(5391) <= a xor b;
    layer7_outputs(5392) <= a and b;
    layer7_outputs(5393) <= 1'b0;
    layer7_outputs(5394) <= not b or a;
    layer7_outputs(5395) <= b;
    layer7_outputs(5396) <= not b;
    layer7_outputs(5397) <= not a or b;
    layer7_outputs(5398) <= not (a and b);
    layer7_outputs(5399) <= b;
    layer7_outputs(5400) <= not (a or b);
    layer7_outputs(5401) <= a;
    layer7_outputs(5402) <= a or b;
    layer7_outputs(5403) <= a;
    layer7_outputs(5404) <= not b;
    layer7_outputs(5405) <= a;
    layer7_outputs(5406) <= not b;
    layer7_outputs(5407) <= b;
    layer7_outputs(5408) <= not (a and b);
    layer7_outputs(5409) <= a;
    layer7_outputs(5410) <= a;
    layer7_outputs(5411) <= not b;
    layer7_outputs(5412) <= not a or b;
    layer7_outputs(5413) <= not (a and b);
    layer7_outputs(5414) <= b and not a;
    layer7_outputs(5415) <= not b;
    layer7_outputs(5416) <= not a;
    layer7_outputs(5417) <= not (a or b);
    layer7_outputs(5418) <= not a or b;
    layer7_outputs(5419) <= not b;
    layer7_outputs(5420) <= b;
    layer7_outputs(5421) <= a xor b;
    layer7_outputs(5422) <= not a or b;
    layer7_outputs(5423) <= a xor b;
    layer7_outputs(5424) <= not a;
    layer7_outputs(5425) <= a xor b;
    layer7_outputs(5426) <= a xor b;
    layer7_outputs(5427) <= not (a and b);
    layer7_outputs(5428) <= not (a or b);
    layer7_outputs(5429) <= not a;
    layer7_outputs(5430) <= not a;
    layer7_outputs(5431) <= a;
    layer7_outputs(5432) <= not a;
    layer7_outputs(5433) <= b;
    layer7_outputs(5434) <= a and not b;
    layer7_outputs(5435) <= not (a xor b);
    layer7_outputs(5436) <= a xor b;
    layer7_outputs(5437) <= not b;
    layer7_outputs(5438) <= not a;
    layer7_outputs(5439) <= b and not a;
    layer7_outputs(5440) <= not (a and b);
    layer7_outputs(5441) <= not (a and b);
    layer7_outputs(5442) <= a;
    layer7_outputs(5443) <= not b;
    layer7_outputs(5444) <= a xor b;
    layer7_outputs(5445) <= a;
    layer7_outputs(5446) <= b and not a;
    layer7_outputs(5447) <= not (a xor b);
    layer7_outputs(5448) <= not (a and b);
    layer7_outputs(5449) <= a or b;
    layer7_outputs(5450) <= not a;
    layer7_outputs(5451) <= not (a or b);
    layer7_outputs(5452) <= b;
    layer7_outputs(5453) <= not a;
    layer7_outputs(5454) <= a;
    layer7_outputs(5455) <= not a or b;
    layer7_outputs(5456) <= not (a and b);
    layer7_outputs(5457) <= b and not a;
    layer7_outputs(5458) <= not b;
    layer7_outputs(5459) <= a or b;
    layer7_outputs(5460) <= a xor b;
    layer7_outputs(5461) <= a and not b;
    layer7_outputs(5462) <= not a;
    layer7_outputs(5463) <= not b;
    layer7_outputs(5464) <= a;
    layer7_outputs(5465) <= a;
    layer7_outputs(5466) <= a;
    layer7_outputs(5467) <= not (a and b);
    layer7_outputs(5468) <= not a or b;
    layer7_outputs(5469) <= a;
    layer7_outputs(5470) <= not b;
    layer7_outputs(5471) <= a and b;
    layer7_outputs(5472) <= a or b;
    layer7_outputs(5473) <= a xor b;
    layer7_outputs(5474) <= not a;
    layer7_outputs(5475) <= not (a or b);
    layer7_outputs(5476) <= not a or b;
    layer7_outputs(5477) <= a;
    layer7_outputs(5478) <= not a or b;
    layer7_outputs(5479) <= a and not b;
    layer7_outputs(5480) <= not (a xor b);
    layer7_outputs(5481) <= a;
    layer7_outputs(5482) <= a;
    layer7_outputs(5483) <= not a or b;
    layer7_outputs(5484) <= b;
    layer7_outputs(5485) <= not b;
    layer7_outputs(5486) <= a;
    layer7_outputs(5487) <= not b;
    layer7_outputs(5488) <= not a;
    layer7_outputs(5489) <= a xor b;
    layer7_outputs(5490) <= not b;
    layer7_outputs(5491) <= a and not b;
    layer7_outputs(5492) <= b and not a;
    layer7_outputs(5493) <= a and not b;
    layer7_outputs(5494) <= not a;
    layer7_outputs(5495) <= b;
    layer7_outputs(5496) <= a and not b;
    layer7_outputs(5497) <= not b;
    layer7_outputs(5498) <= not (a and b);
    layer7_outputs(5499) <= b;
    layer7_outputs(5500) <= not b or a;
    layer7_outputs(5501) <= not a or b;
    layer7_outputs(5502) <= not (a or b);
    layer7_outputs(5503) <= a;
    layer7_outputs(5504) <= b;
    layer7_outputs(5505) <= a and b;
    layer7_outputs(5506) <= a;
    layer7_outputs(5507) <= a;
    layer7_outputs(5508) <= b;
    layer7_outputs(5509) <= not (a and b);
    layer7_outputs(5510) <= not a or b;
    layer7_outputs(5511) <= a xor b;
    layer7_outputs(5512) <= not (a or b);
    layer7_outputs(5513) <= b;
    layer7_outputs(5514) <= not a;
    layer7_outputs(5515) <= not (a xor b);
    layer7_outputs(5516) <= not (a and b);
    layer7_outputs(5517) <= not b or a;
    layer7_outputs(5518) <= not a or b;
    layer7_outputs(5519) <= a and not b;
    layer7_outputs(5520) <= not a or b;
    layer7_outputs(5521) <= b;
    layer7_outputs(5522) <= a or b;
    layer7_outputs(5523) <= a;
    layer7_outputs(5524) <= not a;
    layer7_outputs(5525) <= b;
    layer7_outputs(5526) <= a xor b;
    layer7_outputs(5527) <= b;
    layer7_outputs(5528) <= not (a xor b);
    layer7_outputs(5529) <= a and b;
    layer7_outputs(5530) <= not b;
    layer7_outputs(5531) <= not b;
    layer7_outputs(5532) <= a and b;
    layer7_outputs(5533) <= a or b;
    layer7_outputs(5534) <= b;
    layer7_outputs(5535) <= a;
    layer7_outputs(5536) <= a and not b;
    layer7_outputs(5537) <= a and not b;
    layer7_outputs(5538) <= 1'b0;
    layer7_outputs(5539) <= a and not b;
    layer7_outputs(5540) <= a xor b;
    layer7_outputs(5541) <= a xor b;
    layer7_outputs(5542) <= not (a or b);
    layer7_outputs(5543) <= a or b;
    layer7_outputs(5544) <= not (a and b);
    layer7_outputs(5545) <= not b;
    layer7_outputs(5546) <= not (a or b);
    layer7_outputs(5547) <= b;
    layer7_outputs(5548) <= not b;
    layer7_outputs(5549) <= not a;
    layer7_outputs(5550) <= b;
    layer7_outputs(5551) <= not b;
    layer7_outputs(5552) <= not (a xor b);
    layer7_outputs(5553) <= not a;
    layer7_outputs(5554) <= a;
    layer7_outputs(5555) <= a;
    layer7_outputs(5556) <= a and not b;
    layer7_outputs(5557) <= not (a or b);
    layer7_outputs(5558) <= a;
    layer7_outputs(5559) <= a xor b;
    layer7_outputs(5560) <= not (a or b);
    layer7_outputs(5561) <= not b;
    layer7_outputs(5562) <= a and b;
    layer7_outputs(5563) <= not b;
    layer7_outputs(5564) <= not a or b;
    layer7_outputs(5565) <= not b;
    layer7_outputs(5566) <= not (a xor b);
    layer7_outputs(5567) <= a;
    layer7_outputs(5568) <= not b;
    layer7_outputs(5569) <= not b;
    layer7_outputs(5570) <= a or b;
    layer7_outputs(5571) <= b and not a;
    layer7_outputs(5572) <= a xor b;
    layer7_outputs(5573) <= not b;
    layer7_outputs(5574) <= b;
    layer7_outputs(5575) <= not (a and b);
    layer7_outputs(5576) <= a and not b;
    layer7_outputs(5577) <= not b;
    layer7_outputs(5578) <= b;
    layer7_outputs(5579) <= not b;
    layer7_outputs(5580) <= not (a xor b);
    layer7_outputs(5581) <= not b;
    layer7_outputs(5582) <= not (a xor b);
    layer7_outputs(5583) <= not (a xor b);
    layer7_outputs(5584) <= a xor b;
    layer7_outputs(5585) <= a and b;
    layer7_outputs(5586) <= a and b;
    layer7_outputs(5587) <= not b or a;
    layer7_outputs(5588) <= a xor b;
    layer7_outputs(5589) <= not (a or b);
    layer7_outputs(5590) <= b and not a;
    layer7_outputs(5591) <= not (a or b);
    layer7_outputs(5592) <= not b or a;
    layer7_outputs(5593) <= not a;
    layer7_outputs(5594) <= b;
    layer7_outputs(5595) <= not a;
    layer7_outputs(5596) <= not (a xor b);
    layer7_outputs(5597) <= 1'b1;
    layer7_outputs(5598) <= a xor b;
    layer7_outputs(5599) <= not (a or b);
    layer7_outputs(5600) <= b;
    layer7_outputs(5601) <= a and b;
    layer7_outputs(5602) <= a;
    layer7_outputs(5603) <= not (a and b);
    layer7_outputs(5604) <= b;
    layer7_outputs(5605) <= b;
    layer7_outputs(5606) <= a;
    layer7_outputs(5607) <= b;
    layer7_outputs(5608) <= a and not b;
    layer7_outputs(5609) <= not a;
    layer7_outputs(5610) <= a and b;
    layer7_outputs(5611) <= not (a and b);
    layer7_outputs(5612) <= b;
    layer7_outputs(5613) <= not (a xor b);
    layer7_outputs(5614) <= not a or b;
    layer7_outputs(5615) <= a and not b;
    layer7_outputs(5616) <= a;
    layer7_outputs(5617) <= a and b;
    layer7_outputs(5618) <= not (a and b);
    layer7_outputs(5619) <= not b;
    layer7_outputs(5620) <= not (a or b);
    layer7_outputs(5621) <= not (a xor b);
    layer7_outputs(5622) <= not (a xor b);
    layer7_outputs(5623) <= not (a or b);
    layer7_outputs(5624) <= 1'b1;
    layer7_outputs(5625) <= b and not a;
    layer7_outputs(5626) <= not b;
    layer7_outputs(5627) <= b;
    layer7_outputs(5628) <= a and not b;
    layer7_outputs(5629) <= not b or a;
    layer7_outputs(5630) <= not (a xor b);
    layer7_outputs(5631) <= a and not b;
    layer7_outputs(5632) <= a and b;
    layer7_outputs(5633) <= 1'b0;
    layer7_outputs(5634) <= b;
    layer7_outputs(5635) <= not b;
    layer7_outputs(5636) <= a;
    layer7_outputs(5637) <= not a;
    layer7_outputs(5638) <= not (a and b);
    layer7_outputs(5639) <= a;
    layer7_outputs(5640) <= b;
    layer7_outputs(5641) <= a;
    layer7_outputs(5642) <= not b;
    layer7_outputs(5643) <= not (a or b);
    layer7_outputs(5644) <= a;
    layer7_outputs(5645) <= b and not a;
    layer7_outputs(5646) <= a;
    layer7_outputs(5647) <= not b or a;
    layer7_outputs(5648) <= not (a xor b);
    layer7_outputs(5649) <= not a;
    layer7_outputs(5650) <= b;
    layer7_outputs(5651) <= a and b;
    layer7_outputs(5652) <= not b;
    layer7_outputs(5653) <= not a or b;
    layer7_outputs(5654) <= not a;
    layer7_outputs(5655) <= b;
    layer7_outputs(5656) <= not (a xor b);
    layer7_outputs(5657) <= a and b;
    layer7_outputs(5658) <= a;
    layer7_outputs(5659) <= b and not a;
    layer7_outputs(5660) <= not b;
    layer7_outputs(5661) <= not b;
    layer7_outputs(5662) <= a and b;
    layer7_outputs(5663) <= b and not a;
    layer7_outputs(5664) <= not b;
    layer7_outputs(5665) <= a;
    layer7_outputs(5666) <= not a;
    layer7_outputs(5667) <= a xor b;
    layer7_outputs(5668) <= not b or a;
    layer7_outputs(5669) <= not b;
    layer7_outputs(5670) <= not (a xor b);
    layer7_outputs(5671) <= not (a xor b);
    layer7_outputs(5672) <= b and not a;
    layer7_outputs(5673) <= b;
    layer7_outputs(5674) <= not a;
    layer7_outputs(5675) <= not (a xor b);
    layer7_outputs(5676) <= not b;
    layer7_outputs(5677) <= not (a xor b);
    layer7_outputs(5678) <= not b;
    layer7_outputs(5679) <= a xor b;
    layer7_outputs(5680) <= not a;
    layer7_outputs(5681) <= not a;
    layer7_outputs(5682) <= b;
    layer7_outputs(5683) <= not b;
    layer7_outputs(5684) <= not a;
    layer7_outputs(5685) <= not b;
    layer7_outputs(5686) <= not b;
    layer7_outputs(5687) <= not (a xor b);
    layer7_outputs(5688) <= not (a xor b);
    layer7_outputs(5689) <= not (a or b);
    layer7_outputs(5690) <= b;
    layer7_outputs(5691) <= not a or b;
    layer7_outputs(5692) <= a or b;
    layer7_outputs(5693) <= b;
    layer7_outputs(5694) <= a and b;
    layer7_outputs(5695) <= b;
    layer7_outputs(5696) <= a or b;
    layer7_outputs(5697) <= b;
    layer7_outputs(5698) <= not a;
    layer7_outputs(5699) <= not (a and b);
    layer7_outputs(5700) <= a;
    layer7_outputs(5701) <= b;
    layer7_outputs(5702) <= a xor b;
    layer7_outputs(5703) <= b and not a;
    layer7_outputs(5704) <= not a or b;
    layer7_outputs(5705) <= not (a xor b);
    layer7_outputs(5706) <= a and b;
    layer7_outputs(5707) <= not a;
    layer7_outputs(5708) <= a xor b;
    layer7_outputs(5709) <= b;
    layer7_outputs(5710) <= not a or b;
    layer7_outputs(5711) <= not (a xor b);
    layer7_outputs(5712) <= a xor b;
    layer7_outputs(5713) <= b;
    layer7_outputs(5714) <= not (a or b);
    layer7_outputs(5715) <= a and b;
    layer7_outputs(5716) <= a;
    layer7_outputs(5717) <= not b or a;
    layer7_outputs(5718) <= not b;
    layer7_outputs(5719) <= a and b;
    layer7_outputs(5720) <= a;
    layer7_outputs(5721) <= not (a xor b);
    layer7_outputs(5722) <= not a;
    layer7_outputs(5723) <= not (a or b);
    layer7_outputs(5724) <= not (a xor b);
    layer7_outputs(5725) <= not b or a;
    layer7_outputs(5726) <= not a or b;
    layer7_outputs(5727) <= not (a or b);
    layer7_outputs(5728) <= not b;
    layer7_outputs(5729) <= not (a xor b);
    layer7_outputs(5730) <= b and not a;
    layer7_outputs(5731) <= b;
    layer7_outputs(5732) <= not (a or b);
    layer7_outputs(5733) <= a xor b;
    layer7_outputs(5734) <= a and b;
    layer7_outputs(5735) <= a and b;
    layer7_outputs(5736) <= not (a xor b);
    layer7_outputs(5737) <= not (a xor b);
    layer7_outputs(5738) <= a xor b;
    layer7_outputs(5739) <= a and not b;
    layer7_outputs(5740) <= b and not a;
    layer7_outputs(5741) <= not b;
    layer7_outputs(5742) <= not (a xor b);
    layer7_outputs(5743) <= a and not b;
    layer7_outputs(5744) <= not (a xor b);
    layer7_outputs(5745) <= not b or a;
    layer7_outputs(5746) <= not a;
    layer7_outputs(5747) <= not (a or b);
    layer7_outputs(5748) <= a and not b;
    layer7_outputs(5749) <= not a or b;
    layer7_outputs(5750) <= not b;
    layer7_outputs(5751) <= not (a and b);
    layer7_outputs(5752) <= not (a xor b);
    layer7_outputs(5753) <= not b;
    layer7_outputs(5754) <= b;
    layer7_outputs(5755) <= not b;
    layer7_outputs(5756) <= not (a or b);
    layer7_outputs(5757) <= a xor b;
    layer7_outputs(5758) <= a;
    layer7_outputs(5759) <= not (a xor b);
    layer7_outputs(5760) <= a;
    layer7_outputs(5761) <= a and b;
    layer7_outputs(5762) <= not (a xor b);
    layer7_outputs(5763) <= not b;
    layer7_outputs(5764) <= a and not b;
    layer7_outputs(5765) <= not (a or b);
    layer7_outputs(5766) <= a;
    layer7_outputs(5767) <= a and not b;
    layer7_outputs(5768) <= a and b;
    layer7_outputs(5769) <= not b;
    layer7_outputs(5770) <= a;
    layer7_outputs(5771) <= a and b;
    layer7_outputs(5772) <= a or b;
    layer7_outputs(5773) <= a xor b;
    layer7_outputs(5774) <= not b;
    layer7_outputs(5775) <= a;
    layer7_outputs(5776) <= a xor b;
    layer7_outputs(5777) <= not (a and b);
    layer7_outputs(5778) <= not (a and b);
    layer7_outputs(5779) <= not b;
    layer7_outputs(5780) <= a;
    layer7_outputs(5781) <= not b;
    layer7_outputs(5782) <= a and not b;
    layer7_outputs(5783) <= not (a xor b);
    layer7_outputs(5784) <= not (a xor b);
    layer7_outputs(5785) <= a;
    layer7_outputs(5786) <= not (a and b);
    layer7_outputs(5787) <= a;
    layer7_outputs(5788) <= not a;
    layer7_outputs(5789) <= a xor b;
    layer7_outputs(5790) <= b;
    layer7_outputs(5791) <= not a;
    layer7_outputs(5792) <= a or b;
    layer7_outputs(5793) <= not a;
    layer7_outputs(5794) <= 1'b0;
    layer7_outputs(5795) <= not b;
    layer7_outputs(5796) <= a;
    layer7_outputs(5797) <= a xor b;
    layer7_outputs(5798) <= a;
    layer7_outputs(5799) <= not (a or b);
    layer7_outputs(5800) <= not (a xor b);
    layer7_outputs(5801) <= not b;
    layer7_outputs(5802) <= not (a or b);
    layer7_outputs(5803) <= not a;
    layer7_outputs(5804) <= not b;
    layer7_outputs(5805) <= b and not a;
    layer7_outputs(5806) <= a xor b;
    layer7_outputs(5807) <= not a;
    layer7_outputs(5808) <= not (a or b);
    layer7_outputs(5809) <= b;
    layer7_outputs(5810) <= not (a and b);
    layer7_outputs(5811) <= a and not b;
    layer7_outputs(5812) <= not b;
    layer7_outputs(5813) <= not b;
    layer7_outputs(5814) <= a or b;
    layer7_outputs(5815) <= not a;
    layer7_outputs(5816) <= b;
    layer7_outputs(5817) <= not b;
    layer7_outputs(5818) <= b and not a;
    layer7_outputs(5819) <= not a;
    layer7_outputs(5820) <= a xor b;
    layer7_outputs(5821) <= b;
    layer7_outputs(5822) <= not b;
    layer7_outputs(5823) <= not a;
    layer7_outputs(5824) <= not a or b;
    layer7_outputs(5825) <= not (a xor b);
    layer7_outputs(5826) <= b;
    layer7_outputs(5827) <= not a or b;
    layer7_outputs(5828) <= a xor b;
    layer7_outputs(5829) <= a or b;
    layer7_outputs(5830) <= not a;
    layer7_outputs(5831) <= a;
    layer7_outputs(5832) <= not b;
    layer7_outputs(5833) <= a;
    layer7_outputs(5834) <= a xor b;
    layer7_outputs(5835) <= not (a xor b);
    layer7_outputs(5836) <= b;
    layer7_outputs(5837) <= a or b;
    layer7_outputs(5838) <= not (a xor b);
    layer7_outputs(5839) <= a;
    layer7_outputs(5840) <= b and not a;
    layer7_outputs(5841) <= a and b;
    layer7_outputs(5842) <= b;
    layer7_outputs(5843) <= not b;
    layer7_outputs(5844) <= not b;
    layer7_outputs(5845) <= not (a and b);
    layer7_outputs(5846) <= not a;
    layer7_outputs(5847) <= a;
    layer7_outputs(5848) <= b;
    layer7_outputs(5849) <= a xor b;
    layer7_outputs(5850) <= b;
    layer7_outputs(5851) <= a;
    layer7_outputs(5852) <= not b;
    layer7_outputs(5853) <= not a;
    layer7_outputs(5854) <= b and not a;
    layer7_outputs(5855) <= a xor b;
    layer7_outputs(5856) <= not b;
    layer7_outputs(5857) <= a and not b;
    layer7_outputs(5858) <= not (a xor b);
    layer7_outputs(5859) <= b;
    layer7_outputs(5860) <= a;
    layer7_outputs(5861) <= not (a xor b);
    layer7_outputs(5862) <= not a;
    layer7_outputs(5863) <= not (a xor b);
    layer7_outputs(5864) <= not (a or b);
    layer7_outputs(5865) <= not a;
    layer7_outputs(5866) <= not (a or b);
    layer7_outputs(5867) <= not a;
    layer7_outputs(5868) <= a;
    layer7_outputs(5869) <= a xor b;
    layer7_outputs(5870) <= a;
    layer7_outputs(5871) <= not (a xor b);
    layer7_outputs(5872) <= not a;
    layer7_outputs(5873) <= not (a or b);
    layer7_outputs(5874) <= not a;
    layer7_outputs(5875) <= not a;
    layer7_outputs(5876) <= not (a xor b);
    layer7_outputs(5877) <= b;
    layer7_outputs(5878) <= not b;
    layer7_outputs(5879) <= a or b;
    layer7_outputs(5880) <= b;
    layer7_outputs(5881) <= b and not a;
    layer7_outputs(5882) <= a or b;
    layer7_outputs(5883) <= not a;
    layer7_outputs(5884) <= not a or b;
    layer7_outputs(5885) <= not a;
    layer7_outputs(5886) <= a xor b;
    layer7_outputs(5887) <= not (a or b);
    layer7_outputs(5888) <= a;
    layer7_outputs(5889) <= not a;
    layer7_outputs(5890) <= not b or a;
    layer7_outputs(5891) <= not a;
    layer7_outputs(5892) <= a;
    layer7_outputs(5893) <= not a;
    layer7_outputs(5894) <= b and not a;
    layer7_outputs(5895) <= not a or b;
    layer7_outputs(5896) <= b;
    layer7_outputs(5897) <= not a;
    layer7_outputs(5898) <= not (a or b);
    layer7_outputs(5899) <= a;
    layer7_outputs(5900) <= not a or b;
    layer7_outputs(5901) <= not b;
    layer7_outputs(5902) <= b;
    layer7_outputs(5903) <= b;
    layer7_outputs(5904) <= not a;
    layer7_outputs(5905) <= not b;
    layer7_outputs(5906) <= 1'b1;
    layer7_outputs(5907) <= a and b;
    layer7_outputs(5908) <= not (a xor b);
    layer7_outputs(5909) <= a xor b;
    layer7_outputs(5910) <= b and not a;
    layer7_outputs(5911) <= a;
    layer7_outputs(5912) <= a or b;
    layer7_outputs(5913) <= a or b;
    layer7_outputs(5914) <= a;
    layer7_outputs(5915) <= not a;
    layer7_outputs(5916) <= not a;
    layer7_outputs(5917) <= not b or a;
    layer7_outputs(5918) <= a or b;
    layer7_outputs(5919) <= not b;
    layer7_outputs(5920) <= a and b;
    layer7_outputs(5921) <= not b;
    layer7_outputs(5922) <= b;
    layer7_outputs(5923) <= not a;
    layer7_outputs(5924) <= not a or b;
    layer7_outputs(5925) <= a or b;
    layer7_outputs(5926) <= not (a and b);
    layer7_outputs(5927) <= not a;
    layer7_outputs(5928) <= a;
    layer7_outputs(5929) <= not (a or b);
    layer7_outputs(5930) <= not b or a;
    layer7_outputs(5931) <= a or b;
    layer7_outputs(5932) <= a and not b;
    layer7_outputs(5933) <= a and not b;
    layer7_outputs(5934) <= a or b;
    layer7_outputs(5935) <= not (a and b);
    layer7_outputs(5936) <= a xor b;
    layer7_outputs(5937) <= not b;
    layer7_outputs(5938) <= a;
    layer7_outputs(5939) <= not a;
    layer7_outputs(5940) <= not b or a;
    layer7_outputs(5941) <= not b;
    layer7_outputs(5942) <= a xor b;
    layer7_outputs(5943) <= a;
    layer7_outputs(5944) <= not (a or b);
    layer7_outputs(5945) <= b;
    layer7_outputs(5946) <= a and b;
    layer7_outputs(5947) <= a;
    layer7_outputs(5948) <= a;
    layer7_outputs(5949) <= not (a or b);
    layer7_outputs(5950) <= a;
    layer7_outputs(5951) <= not a;
    layer7_outputs(5952) <= not (a or b);
    layer7_outputs(5953) <= not (a and b);
    layer7_outputs(5954) <= b;
    layer7_outputs(5955) <= not (a xor b);
    layer7_outputs(5956) <= a;
    layer7_outputs(5957) <= not a;
    layer7_outputs(5958) <= not (a xor b);
    layer7_outputs(5959) <= a xor b;
    layer7_outputs(5960) <= a xor b;
    layer7_outputs(5961) <= not a;
    layer7_outputs(5962) <= b;
    layer7_outputs(5963) <= a and b;
    layer7_outputs(5964) <= b and not a;
    layer7_outputs(5965) <= b;
    layer7_outputs(5966) <= not (a and b);
    layer7_outputs(5967) <= not b;
    layer7_outputs(5968) <= a xor b;
    layer7_outputs(5969) <= not (a xor b);
    layer7_outputs(5970) <= not a or b;
    layer7_outputs(5971) <= not (a and b);
    layer7_outputs(5972) <= a;
    layer7_outputs(5973) <= b;
    layer7_outputs(5974) <= a or b;
    layer7_outputs(5975) <= a;
    layer7_outputs(5976) <= a and not b;
    layer7_outputs(5977) <= not (a and b);
    layer7_outputs(5978) <= a or b;
    layer7_outputs(5979) <= b;
    layer7_outputs(5980) <= a and b;
    layer7_outputs(5981) <= not b or a;
    layer7_outputs(5982) <= a;
    layer7_outputs(5983) <= not a;
    layer7_outputs(5984) <= a and not b;
    layer7_outputs(5985) <= not b;
    layer7_outputs(5986) <= not b or a;
    layer7_outputs(5987) <= not b;
    layer7_outputs(5988) <= not (a xor b);
    layer7_outputs(5989) <= not (a xor b);
    layer7_outputs(5990) <= not (a and b);
    layer7_outputs(5991) <= a xor b;
    layer7_outputs(5992) <= not b;
    layer7_outputs(5993) <= a and not b;
    layer7_outputs(5994) <= b;
    layer7_outputs(5995) <= a xor b;
    layer7_outputs(5996) <= a and not b;
    layer7_outputs(5997) <= not a;
    layer7_outputs(5998) <= a and b;
    layer7_outputs(5999) <= 1'b0;
    layer7_outputs(6000) <= a;
    layer7_outputs(6001) <= a;
    layer7_outputs(6002) <= a or b;
    layer7_outputs(6003) <= not (a xor b);
    layer7_outputs(6004) <= not b;
    layer7_outputs(6005) <= b;
    layer7_outputs(6006) <= not a or b;
    layer7_outputs(6007) <= b;
    layer7_outputs(6008) <= 1'b1;
    layer7_outputs(6009) <= b and not a;
    layer7_outputs(6010) <= not b;
    layer7_outputs(6011) <= not (a xor b);
    layer7_outputs(6012) <= not a;
    layer7_outputs(6013) <= a or b;
    layer7_outputs(6014) <= b;
    layer7_outputs(6015) <= b;
    layer7_outputs(6016) <= a;
    layer7_outputs(6017) <= b and not a;
    layer7_outputs(6018) <= not b or a;
    layer7_outputs(6019) <= a or b;
    layer7_outputs(6020) <= not (a xor b);
    layer7_outputs(6021) <= a;
    layer7_outputs(6022) <= a and not b;
    layer7_outputs(6023) <= a and not b;
    layer7_outputs(6024) <= not (a xor b);
    layer7_outputs(6025) <= not (a or b);
    layer7_outputs(6026) <= a;
    layer7_outputs(6027) <= a;
    layer7_outputs(6028) <= not b;
    layer7_outputs(6029) <= b;
    layer7_outputs(6030) <= not b;
    layer7_outputs(6031) <= a;
    layer7_outputs(6032) <= not (a xor b);
    layer7_outputs(6033) <= not (a and b);
    layer7_outputs(6034) <= a;
    layer7_outputs(6035) <= not (a xor b);
    layer7_outputs(6036) <= a;
    layer7_outputs(6037) <= a;
    layer7_outputs(6038) <= a and b;
    layer7_outputs(6039) <= not a;
    layer7_outputs(6040) <= not (a and b);
    layer7_outputs(6041) <= not a;
    layer7_outputs(6042) <= b and not a;
    layer7_outputs(6043) <= a or b;
    layer7_outputs(6044) <= not b or a;
    layer7_outputs(6045) <= 1'b0;
    layer7_outputs(6046) <= not (a xor b);
    layer7_outputs(6047) <= not (a xor b);
    layer7_outputs(6048) <= b;
    layer7_outputs(6049) <= a and not b;
    layer7_outputs(6050) <= a and b;
    layer7_outputs(6051) <= not (a or b);
    layer7_outputs(6052) <= a or b;
    layer7_outputs(6053) <= not b or a;
    layer7_outputs(6054) <= not b or a;
    layer7_outputs(6055) <= b;
    layer7_outputs(6056) <= a or b;
    layer7_outputs(6057) <= not a or b;
    layer7_outputs(6058) <= not a;
    layer7_outputs(6059) <= not (a xor b);
    layer7_outputs(6060) <= not (a xor b);
    layer7_outputs(6061) <= b;
    layer7_outputs(6062) <= not a;
    layer7_outputs(6063) <= a;
    layer7_outputs(6064) <= a xor b;
    layer7_outputs(6065) <= b and not a;
    layer7_outputs(6066) <= b and not a;
    layer7_outputs(6067) <= not (a xor b);
    layer7_outputs(6068) <= not a;
    layer7_outputs(6069) <= a xor b;
    layer7_outputs(6070) <= not a;
    layer7_outputs(6071) <= not b or a;
    layer7_outputs(6072) <= a and b;
    layer7_outputs(6073) <= b;
    layer7_outputs(6074) <= not (a or b);
    layer7_outputs(6075) <= a;
    layer7_outputs(6076) <= a and not b;
    layer7_outputs(6077) <= a or b;
    layer7_outputs(6078) <= a;
    layer7_outputs(6079) <= b;
    layer7_outputs(6080) <= a or b;
    layer7_outputs(6081) <= not b or a;
    layer7_outputs(6082) <= a;
    layer7_outputs(6083) <= a and not b;
    layer7_outputs(6084) <= a;
    layer7_outputs(6085) <= not a or b;
    layer7_outputs(6086) <= a and not b;
    layer7_outputs(6087) <= a or b;
    layer7_outputs(6088) <= not (a xor b);
    layer7_outputs(6089) <= b and not a;
    layer7_outputs(6090) <= b;
    layer7_outputs(6091) <= a and b;
    layer7_outputs(6092) <= not a;
    layer7_outputs(6093) <= a;
    layer7_outputs(6094) <= not a or b;
    layer7_outputs(6095) <= not b;
    layer7_outputs(6096) <= not (a xor b);
    layer7_outputs(6097) <= not (a or b);
    layer7_outputs(6098) <= b;
    layer7_outputs(6099) <= b and not a;
    layer7_outputs(6100) <= b;
    layer7_outputs(6101) <= not a or b;
    layer7_outputs(6102) <= not (a xor b);
    layer7_outputs(6103) <= b;
    layer7_outputs(6104) <= b;
    layer7_outputs(6105) <= not b;
    layer7_outputs(6106) <= b;
    layer7_outputs(6107) <= not b or a;
    layer7_outputs(6108) <= b;
    layer7_outputs(6109) <= b;
    layer7_outputs(6110) <= b;
    layer7_outputs(6111) <= a xor b;
    layer7_outputs(6112) <= a or b;
    layer7_outputs(6113) <= not (a or b);
    layer7_outputs(6114) <= a and b;
    layer7_outputs(6115) <= a or b;
    layer7_outputs(6116) <= not (a or b);
    layer7_outputs(6117) <= a xor b;
    layer7_outputs(6118) <= not (a or b);
    layer7_outputs(6119) <= not b;
    layer7_outputs(6120) <= not b;
    layer7_outputs(6121) <= not b or a;
    layer7_outputs(6122) <= b;
    layer7_outputs(6123) <= not b;
    layer7_outputs(6124) <= a;
    layer7_outputs(6125) <= not (a xor b);
    layer7_outputs(6126) <= b;
    layer7_outputs(6127) <= b and not a;
    layer7_outputs(6128) <= not b;
    layer7_outputs(6129) <= b and not a;
    layer7_outputs(6130) <= not b;
    layer7_outputs(6131) <= a xor b;
    layer7_outputs(6132) <= not b;
    layer7_outputs(6133) <= 1'b1;
    layer7_outputs(6134) <= not a;
    layer7_outputs(6135) <= a xor b;
    layer7_outputs(6136) <= b;
    layer7_outputs(6137) <= not a or b;
    layer7_outputs(6138) <= not (a xor b);
    layer7_outputs(6139) <= a xor b;
    layer7_outputs(6140) <= not a;
    layer7_outputs(6141) <= not b;
    layer7_outputs(6142) <= b;
    layer7_outputs(6143) <= b;
    layer7_outputs(6144) <= a;
    layer7_outputs(6145) <= b and not a;
    layer7_outputs(6146) <= not (a xor b);
    layer7_outputs(6147) <= not b;
    layer7_outputs(6148) <= a;
    layer7_outputs(6149) <= a and b;
    layer7_outputs(6150) <= a xor b;
    layer7_outputs(6151) <= not b;
    layer7_outputs(6152) <= not a or b;
    layer7_outputs(6153) <= not (a and b);
    layer7_outputs(6154) <= a and b;
    layer7_outputs(6155) <= not (a and b);
    layer7_outputs(6156) <= a;
    layer7_outputs(6157) <= not a;
    layer7_outputs(6158) <= not a;
    layer7_outputs(6159) <= not a;
    layer7_outputs(6160) <= b and not a;
    layer7_outputs(6161) <= a xor b;
    layer7_outputs(6162) <= a and b;
    layer7_outputs(6163) <= a;
    layer7_outputs(6164) <= a and not b;
    layer7_outputs(6165) <= not a;
    layer7_outputs(6166) <= not (a xor b);
    layer7_outputs(6167) <= a or b;
    layer7_outputs(6168) <= not (a and b);
    layer7_outputs(6169) <= not (a xor b);
    layer7_outputs(6170) <= a;
    layer7_outputs(6171) <= not a;
    layer7_outputs(6172) <= b;
    layer7_outputs(6173) <= not a;
    layer7_outputs(6174) <= not (a or b);
    layer7_outputs(6175) <= b;
    layer7_outputs(6176) <= not b;
    layer7_outputs(6177) <= not (a xor b);
    layer7_outputs(6178) <= b and not a;
    layer7_outputs(6179) <= not b;
    layer7_outputs(6180) <= not (a or b);
    layer7_outputs(6181) <= a;
    layer7_outputs(6182) <= a;
    layer7_outputs(6183) <= not (a and b);
    layer7_outputs(6184) <= a and b;
    layer7_outputs(6185) <= a and b;
    layer7_outputs(6186) <= b and not a;
    layer7_outputs(6187) <= b and not a;
    layer7_outputs(6188) <= b;
    layer7_outputs(6189) <= not a or b;
    layer7_outputs(6190) <= not (a xor b);
    layer7_outputs(6191) <= not (a and b);
    layer7_outputs(6192) <= a;
    layer7_outputs(6193) <= a and b;
    layer7_outputs(6194) <= a or b;
    layer7_outputs(6195) <= not a;
    layer7_outputs(6196) <= not a or b;
    layer7_outputs(6197) <= not (a or b);
    layer7_outputs(6198) <= a or b;
    layer7_outputs(6199) <= b and not a;
    layer7_outputs(6200) <= a xor b;
    layer7_outputs(6201) <= a and not b;
    layer7_outputs(6202) <= a;
    layer7_outputs(6203) <= a xor b;
    layer7_outputs(6204) <= a;
    layer7_outputs(6205) <= a and b;
    layer7_outputs(6206) <= not a;
    layer7_outputs(6207) <= a xor b;
    layer7_outputs(6208) <= a or b;
    layer7_outputs(6209) <= b;
    layer7_outputs(6210) <= a xor b;
    layer7_outputs(6211) <= not b;
    layer7_outputs(6212) <= b and not a;
    layer7_outputs(6213) <= a xor b;
    layer7_outputs(6214) <= a;
    layer7_outputs(6215) <= not (a xor b);
    layer7_outputs(6216) <= b;
    layer7_outputs(6217) <= not b;
    layer7_outputs(6218) <= b;
    layer7_outputs(6219) <= not a;
    layer7_outputs(6220) <= not b;
    layer7_outputs(6221) <= not a;
    layer7_outputs(6222) <= b and not a;
    layer7_outputs(6223) <= a or b;
    layer7_outputs(6224) <= b;
    layer7_outputs(6225) <= not b;
    layer7_outputs(6226) <= a xor b;
    layer7_outputs(6227) <= a and b;
    layer7_outputs(6228) <= a and b;
    layer7_outputs(6229) <= b;
    layer7_outputs(6230) <= not (a or b);
    layer7_outputs(6231) <= not a;
    layer7_outputs(6232) <= not a;
    layer7_outputs(6233) <= a or b;
    layer7_outputs(6234) <= not b;
    layer7_outputs(6235) <= a;
    layer7_outputs(6236) <= not b;
    layer7_outputs(6237) <= not (a or b);
    layer7_outputs(6238) <= not (a xor b);
    layer7_outputs(6239) <= not b;
    layer7_outputs(6240) <= not (a xor b);
    layer7_outputs(6241) <= b and not a;
    layer7_outputs(6242) <= not a;
    layer7_outputs(6243) <= not a;
    layer7_outputs(6244) <= not b;
    layer7_outputs(6245) <= b and not a;
    layer7_outputs(6246) <= not a;
    layer7_outputs(6247) <= a;
    layer7_outputs(6248) <= not b or a;
    layer7_outputs(6249) <= a;
    layer7_outputs(6250) <= not (a and b);
    layer7_outputs(6251) <= a;
    layer7_outputs(6252) <= a;
    layer7_outputs(6253) <= not (a and b);
    layer7_outputs(6254) <= b;
    layer7_outputs(6255) <= a;
    layer7_outputs(6256) <= a or b;
    layer7_outputs(6257) <= a and not b;
    layer7_outputs(6258) <= a and not b;
    layer7_outputs(6259) <= not a;
    layer7_outputs(6260) <= not (a or b);
    layer7_outputs(6261) <= a and b;
    layer7_outputs(6262) <= not a;
    layer7_outputs(6263) <= not b or a;
    layer7_outputs(6264) <= not b or a;
    layer7_outputs(6265) <= a and not b;
    layer7_outputs(6266) <= b and not a;
    layer7_outputs(6267) <= not a or b;
    layer7_outputs(6268) <= not b or a;
    layer7_outputs(6269) <= not a or b;
    layer7_outputs(6270) <= not a;
    layer7_outputs(6271) <= not a;
    layer7_outputs(6272) <= 1'b0;
    layer7_outputs(6273) <= not (a or b);
    layer7_outputs(6274) <= 1'b0;
    layer7_outputs(6275) <= a;
    layer7_outputs(6276) <= a and b;
    layer7_outputs(6277) <= not b;
    layer7_outputs(6278) <= b and not a;
    layer7_outputs(6279) <= not a;
    layer7_outputs(6280) <= not a;
    layer7_outputs(6281) <= b and not a;
    layer7_outputs(6282) <= not b or a;
    layer7_outputs(6283) <= not b;
    layer7_outputs(6284) <= a xor b;
    layer7_outputs(6285) <= not (a xor b);
    layer7_outputs(6286) <= not (a xor b);
    layer7_outputs(6287) <= not b or a;
    layer7_outputs(6288) <= not b;
    layer7_outputs(6289) <= b;
    layer7_outputs(6290) <= not (a xor b);
    layer7_outputs(6291) <= not (a or b);
    layer7_outputs(6292) <= not b or a;
    layer7_outputs(6293) <= not (a and b);
    layer7_outputs(6294) <= b;
    layer7_outputs(6295) <= a or b;
    layer7_outputs(6296) <= 1'b0;
    layer7_outputs(6297) <= not (a and b);
    layer7_outputs(6298) <= not a;
    layer7_outputs(6299) <= a and b;
    layer7_outputs(6300) <= a or b;
    layer7_outputs(6301) <= not (a or b);
    layer7_outputs(6302) <= a;
    layer7_outputs(6303) <= not a;
    layer7_outputs(6304) <= not (a and b);
    layer7_outputs(6305) <= not (a xor b);
    layer7_outputs(6306) <= not a or b;
    layer7_outputs(6307) <= a and b;
    layer7_outputs(6308) <= b;
    layer7_outputs(6309) <= not a;
    layer7_outputs(6310) <= not a;
    layer7_outputs(6311) <= b;
    layer7_outputs(6312) <= not a;
    layer7_outputs(6313) <= not b;
    layer7_outputs(6314) <= not b;
    layer7_outputs(6315) <= not a;
    layer7_outputs(6316) <= b;
    layer7_outputs(6317) <= not b;
    layer7_outputs(6318) <= a;
    layer7_outputs(6319) <= b and not a;
    layer7_outputs(6320) <= b and not a;
    layer7_outputs(6321) <= not (a xor b);
    layer7_outputs(6322) <= a;
    layer7_outputs(6323) <= not (a and b);
    layer7_outputs(6324) <= not b or a;
    layer7_outputs(6325) <= not b or a;
    layer7_outputs(6326) <= a and not b;
    layer7_outputs(6327) <= not a or b;
    layer7_outputs(6328) <= not b;
    layer7_outputs(6329) <= not a;
    layer7_outputs(6330) <= b;
    layer7_outputs(6331) <= not a;
    layer7_outputs(6332) <= b and not a;
    layer7_outputs(6333) <= 1'b0;
    layer7_outputs(6334) <= a xor b;
    layer7_outputs(6335) <= a and b;
    layer7_outputs(6336) <= not (a or b);
    layer7_outputs(6337) <= a xor b;
    layer7_outputs(6338) <= a;
    layer7_outputs(6339) <= b;
    layer7_outputs(6340) <= b and not a;
    layer7_outputs(6341) <= a xor b;
    layer7_outputs(6342) <= not b;
    layer7_outputs(6343) <= b;
    layer7_outputs(6344) <= not b;
    layer7_outputs(6345) <= not (a or b);
    layer7_outputs(6346) <= b;
    layer7_outputs(6347) <= not a;
    layer7_outputs(6348) <= not a;
    layer7_outputs(6349) <= not b;
    layer7_outputs(6350) <= b;
    layer7_outputs(6351) <= not (a or b);
    layer7_outputs(6352) <= not (a xor b);
    layer7_outputs(6353) <= b;
    layer7_outputs(6354) <= not b;
    layer7_outputs(6355) <= not b;
    layer7_outputs(6356) <= a and not b;
    layer7_outputs(6357) <= b and not a;
    layer7_outputs(6358) <= not b;
    layer7_outputs(6359) <= not a or b;
    layer7_outputs(6360) <= not b or a;
    layer7_outputs(6361) <= not (a and b);
    layer7_outputs(6362) <= a and not b;
    layer7_outputs(6363) <= not b;
    layer7_outputs(6364) <= a xor b;
    layer7_outputs(6365) <= a xor b;
    layer7_outputs(6366) <= a xor b;
    layer7_outputs(6367) <= not (a xor b);
    layer7_outputs(6368) <= a;
    layer7_outputs(6369) <= not (a and b);
    layer7_outputs(6370) <= a xor b;
    layer7_outputs(6371) <= a or b;
    layer7_outputs(6372) <= a and b;
    layer7_outputs(6373) <= a;
    layer7_outputs(6374) <= not b or a;
    layer7_outputs(6375) <= a;
    layer7_outputs(6376) <= a xor b;
    layer7_outputs(6377) <= not a;
    layer7_outputs(6378) <= not (a xor b);
    layer7_outputs(6379) <= a;
    layer7_outputs(6380) <= not b;
    layer7_outputs(6381) <= b and not a;
    layer7_outputs(6382) <= a xor b;
    layer7_outputs(6383) <= a and not b;
    layer7_outputs(6384) <= not a;
    layer7_outputs(6385) <= a;
    layer7_outputs(6386) <= not (a xor b);
    layer7_outputs(6387) <= 1'b1;
    layer7_outputs(6388) <= a xor b;
    layer7_outputs(6389) <= a and not b;
    layer7_outputs(6390) <= a;
    layer7_outputs(6391) <= not a or b;
    layer7_outputs(6392) <= a;
    layer7_outputs(6393) <= b and not a;
    layer7_outputs(6394) <= not (a or b);
    layer7_outputs(6395) <= b and not a;
    layer7_outputs(6396) <= 1'b1;
    layer7_outputs(6397) <= b;
    layer7_outputs(6398) <= a xor b;
    layer7_outputs(6399) <= not b or a;
    layer7_outputs(6400) <= b;
    layer7_outputs(6401) <= not (a or b);
    layer7_outputs(6402) <= a xor b;
    layer7_outputs(6403) <= b and not a;
    layer7_outputs(6404) <= not b;
    layer7_outputs(6405) <= 1'b0;
    layer7_outputs(6406) <= not (a xor b);
    layer7_outputs(6407) <= not (a or b);
    layer7_outputs(6408) <= a or b;
    layer7_outputs(6409) <= not a;
    layer7_outputs(6410) <= not a;
    layer7_outputs(6411) <= 1'b1;
    layer7_outputs(6412) <= b;
    layer7_outputs(6413) <= not (a or b);
    layer7_outputs(6414) <= not a;
    layer7_outputs(6415) <= not a;
    layer7_outputs(6416) <= not b;
    layer7_outputs(6417) <= not (a or b);
    layer7_outputs(6418) <= not a;
    layer7_outputs(6419) <= not a;
    layer7_outputs(6420) <= not a;
    layer7_outputs(6421) <= not a;
    layer7_outputs(6422) <= a;
    layer7_outputs(6423) <= not b;
    layer7_outputs(6424) <= a;
    layer7_outputs(6425) <= not b;
    layer7_outputs(6426) <= a xor b;
    layer7_outputs(6427) <= not (a xor b);
    layer7_outputs(6428) <= a;
    layer7_outputs(6429) <= not b;
    layer7_outputs(6430) <= not a;
    layer7_outputs(6431) <= not a;
    layer7_outputs(6432) <= not b;
    layer7_outputs(6433) <= a and not b;
    layer7_outputs(6434) <= not b;
    layer7_outputs(6435) <= not b or a;
    layer7_outputs(6436) <= not (a xor b);
    layer7_outputs(6437) <= a and not b;
    layer7_outputs(6438) <= not (a and b);
    layer7_outputs(6439) <= not b or a;
    layer7_outputs(6440) <= a and b;
    layer7_outputs(6441) <= 1'b0;
    layer7_outputs(6442) <= b;
    layer7_outputs(6443) <= not (a xor b);
    layer7_outputs(6444) <= not b;
    layer7_outputs(6445) <= b and not a;
    layer7_outputs(6446) <= b;
    layer7_outputs(6447) <= b;
    layer7_outputs(6448) <= not b or a;
    layer7_outputs(6449) <= not a or b;
    layer7_outputs(6450) <= not a;
    layer7_outputs(6451) <= not (a and b);
    layer7_outputs(6452) <= a and not b;
    layer7_outputs(6453) <= not b or a;
    layer7_outputs(6454) <= not (a and b);
    layer7_outputs(6455) <= a xor b;
    layer7_outputs(6456) <= not a;
    layer7_outputs(6457) <= b;
    layer7_outputs(6458) <= b and not a;
    layer7_outputs(6459) <= a and not b;
    layer7_outputs(6460) <= not b or a;
    layer7_outputs(6461) <= a;
    layer7_outputs(6462) <= b;
    layer7_outputs(6463) <= not b;
    layer7_outputs(6464) <= not b;
    layer7_outputs(6465) <= not a;
    layer7_outputs(6466) <= not a;
    layer7_outputs(6467) <= not a or b;
    layer7_outputs(6468) <= b;
    layer7_outputs(6469) <= a and b;
    layer7_outputs(6470) <= not b or a;
    layer7_outputs(6471) <= not (a or b);
    layer7_outputs(6472) <= not (a or b);
    layer7_outputs(6473) <= not (a xor b);
    layer7_outputs(6474) <= a;
    layer7_outputs(6475) <= a and not b;
    layer7_outputs(6476) <= a and not b;
    layer7_outputs(6477) <= not b;
    layer7_outputs(6478) <= a and not b;
    layer7_outputs(6479) <= a;
    layer7_outputs(6480) <= not b;
    layer7_outputs(6481) <= not a;
    layer7_outputs(6482) <= not a;
    layer7_outputs(6483) <= not a;
    layer7_outputs(6484) <= a xor b;
    layer7_outputs(6485) <= a xor b;
    layer7_outputs(6486) <= not b;
    layer7_outputs(6487) <= a and not b;
    layer7_outputs(6488) <= 1'b0;
    layer7_outputs(6489) <= 1'b1;
    layer7_outputs(6490) <= not b or a;
    layer7_outputs(6491) <= not (a xor b);
    layer7_outputs(6492) <= not a;
    layer7_outputs(6493) <= not a;
    layer7_outputs(6494) <= a;
    layer7_outputs(6495) <= b and not a;
    layer7_outputs(6496) <= b;
    layer7_outputs(6497) <= not a;
    layer7_outputs(6498) <= a and not b;
    layer7_outputs(6499) <= a or b;
    layer7_outputs(6500) <= a xor b;
    layer7_outputs(6501) <= not a;
    layer7_outputs(6502) <= not a or b;
    layer7_outputs(6503) <= a and b;
    layer7_outputs(6504) <= a and b;
    layer7_outputs(6505) <= a and not b;
    layer7_outputs(6506) <= not b;
    layer7_outputs(6507) <= not (a or b);
    layer7_outputs(6508) <= not (a or b);
    layer7_outputs(6509) <= b;
    layer7_outputs(6510) <= not (a and b);
    layer7_outputs(6511) <= a and b;
    layer7_outputs(6512) <= a and not b;
    layer7_outputs(6513) <= not a;
    layer7_outputs(6514) <= not a;
    layer7_outputs(6515) <= b and not a;
    layer7_outputs(6516) <= not a;
    layer7_outputs(6517) <= not b or a;
    layer7_outputs(6518) <= not (a and b);
    layer7_outputs(6519) <= not a or b;
    layer7_outputs(6520) <= not b or a;
    layer7_outputs(6521) <= a and not b;
    layer7_outputs(6522) <= not a;
    layer7_outputs(6523) <= a and b;
    layer7_outputs(6524) <= not (a and b);
    layer7_outputs(6525) <= a;
    layer7_outputs(6526) <= not (a xor b);
    layer7_outputs(6527) <= a;
    layer7_outputs(6528) <= not (a or b);
    layer7_outputs(6529) <= not b;
    layer7_outputs(6530) <= not a;
    layer7_outputs(6531) <= not (a or b);
    layer7_outputs(6532) <= not b;
    layer7_outputs(6533) <= a and b;
    layer7_outputs(6534) <= a or b;
    layer7_outputs(6535) <= not a;
    layer7_outputs(6536) <= not a;
    layer7_outputs(6537) <= a;
    layer7_outputs(6538) <= not b;
    layer7_outputs(6539) <= not (a and b);
    layer7_outputs(6540) <= not (a and b);
    layer7_outputs(6541) <= a and not b;
    layer7_outputs(6542) <= not a;
    layer7_outputs(6543) <= not a;
    layer7_outputs(6544) <= not a or b;
    layer7_outputs(6545) <= a xor b;
    layer7_outputs(6546) <= not (a xor b);
    layer7_outputs(6547) <= not b;
    layer7_outputs(6548) <= b and not a;
    layer7_outputs(6549) <= a and not b;
    layer7_outputs(6550) <= not a;
    layer7_outputs(6551) <= not b;
    layer7_outputs(6552) <= not (a and b);
    layer7_outputs(6553) <= a and not b;
    layer7_outputs(6554) <= not b;
    layer7_outputs(6555) <= b;
    layer7_outputs(6556) <= 1'b0;
    layer7_outputs(6557) <= b;
    layer7_outputs(6558) <= b;
    layer7_outputs(6559) <= not b;
    layer7_outputs(6560) <= not (a and b);
    layer7_outputs(6561) <= not b;
    layer7_outputs(6562) <= b and not a;
    layer7_outputs(6563) <= 1'b1;
    layer7_outputs(6564) <= not b;
    layer7_outputs(6565) <= b and not a;
    layer7_outputs(6566) <= a;
    layer7_outputs(6567) <= not (a or b);
    layer7_outputs(6568) <= not (a xor b);
    layer7_outputs(6569) <= not (a and b);
    layer7_outputs(6570) <= b;
    layer7_outputs(6571) <= b;
    layer7_outputs(6572) <= a and not b;
    layer7_outputs(6573) <= not a or b;
    layer7_outputs(6574) <= not (a xor b);
    layer7_outputs(6575) <= not a or b;
    layer7_outputs(6576) <= not b or a;
    layer7_outputs(6577) <= not b;
    layer7_outputs(6578) <= not b;
    layer7_outputs(6579) <= not b;
    layer7_outputs(6580) <= not (a xor b);
    layer7_outputs(6581) <= not a or b;
    layer7_outputs(6582) <= 1'b0;
    layer7_outputs(6583) <= not b;
    layer7_outputs(6584) <= a and b;
    layer7_outputs(6585) <= not (a and b);
    layer7_outputs(6586) <= a;
    layer7_outputs(6587) <= a;
    layer7_outputs(6588) <= not b;
    layer7_outputs(6589) <= a and not b;
    layer7_outputs(6590) <= a and b;
    layer7_outputs(6591) <= a and not b;
    layer7_outputs(6592) <= not (a and b);
    layer7_outputs(6593) <= b;
    layer7_outputs(6594) <= not b or a;
    layer7_outputs(6595) <= not b;
    layer7_outputs(6596) <= a xor b;
    layer7_outputs(6597) <= a and not b;
    layer7_outputs(6598) <= a and b;
    layer7_outputs(6599) <= not (a and b);
    layer7_outputs(6600) <= not b or a;
    layer7_outputs(6601) <= 1'b0;
    layer7_outputs(6602) <= not (a xor b);
    layer7_outputs(6603) <= not a or b;
    layer7_outputs(6604) <= not b or a;
    layer7_outputs(6605) <= b;
    layer7_outputs(6606) <= not a;
    layer7_outputs(6607) <= not b;
    layer7_outputs(6608) <= not (a xor b);
    layer7_outputs(6609) <= b;
    layer7_outputs(6610) <= not b;
    layer7_outputs(6611) <= not a or b;
    layer7_outputs(6612) <= not b or a;
    layer7_outputs(6613) <= not (a and b);
    layer7_outputs(6614) <= not b or a;
    layer7_outputs(6615) <= not a or b;
    layer7_outputs(6616) <= not (a and b);
    layer7_outputs(6617) <= b;
    layer7_outputs(6618) <= not a;
    layer7_outputs(6619) <= not b or a;
    layer7_outputs(6620) <= b and not a;
    layer7_outputs(6621) <= not (a xor b);
    layer7_outputs(6622) <= not b;
    layer7_outputs(6623) <= not a or b;
    layer7_outputs(6624) <= a and b;
    layer7_outputs(6625) <= b;
    layer7_outputs(6626) <= a;
    layer7_outputs(6627) <= not (a xor b);
    layer7_outputs(6628) <= b and not a;
    layer7_outputs(6629) <= b;
    layer7_outputs(6630) <= a or b;
    layer7_outputs(6631) <= a;
    layer7_outputs(6632) <= not a;
    layer7_outputs(6633) <= 1'b1;
    layer7_outputs(6634) <= not a or b;
    layer7_outputs(6635) <= not a;
    layer7_outputs(6636) <= not b;
    layer7_outputs(6637) <= not b;
    layer7_outputs(6638) <= 1'b0;
    layer7_outputs(6639) <= not (a and b);
    layer7_outputs(6640) <= not a;
    layer7_outputs(6641) <= not a;
    layer7_outputs(6642) <= not b;
    layer7_outputs(6643) <= not (a xor b);
    layer7_outputs(6644) <= not (a xor b);
    layer7_outputs(6645) <= b and not a;
    layer7_outputs(6646) <= not a;
    layer7_outputs(6647) <= b;
    layer7_outputs(6648) <= not b or a;
    layer7_outputs(6649) <= b and not a;
    layer7_outputs(6650) <= a;
    layer7_outputs(6651) <= b;
    layer7_outputs(6652) <= a;
    layer7_outputs(6653) <= b;
    layer7_outputs(6654) <= a xor b;
    layer7_outputs(6655) <= not a;
    layer7_outputs(6656) <= b and not a;
    layer7_outputs(6657) <= a;
    layer7_outputs(6658) <= b;
    layer7_outputs(6659) <= not b;
    layer7_outputs(6660) <= a and not b;
    layer7_outputs(6661) <= a or b;
    layer7_outputs(6662) <= not b or a;
    layer7_outputs(6663) <= not b or a;
    layer7_outputs(6664) <= not (a or b);
    layer7_outputs(6665) <= 1'b1;
    layer7_outputs(6666) <= b;
    layer7_outputs(6667) <= a xor b;
    layer7_outputs(6668) <= a;
    layer7_outputs(6669) <= not (a xor b);
    layer7_outputs(6670) <= not b;
    layer7_outputs(6671) <= a;
    layer7_outputs(6672) <= not b;
    layer7_outputs(6673) <= b;
    layer7_outputs(6674) <= a and b;
    layer7_outputs(6675) <= a or b;
    layer7_outputs(6676) <= not b;
    layer7_outputs(6677) <= not (a xor b);
    layer7_outputs(6678) <= a and not b;
    layer7_outputs(6679) <= not b;
    layer7_outputs(6680) <= a or b;
    layer7_outputs(6681) <= b and not a;
    layer7_outputs(6682) <= not b;
    layer7_outputs(6683) <= a;
    layer7_outputs(6684) <= a;
    layer7_outputs(6685) <= a or b;
    layer7_outputs(6686) <= b and not a;
    layer7_outputs(6687) <= b;
    layer7_outputs(6688) <= not a;
    layer7_outputs(6689) <= a or b;
    layer7_outputs(6690) <= a;
    layer7_outputs(6691) <= not a;
    layer7_outputs(6692) <= b;
    layer7_outputs(6693) <= not b;
    layer7_outputs(6694) <= not a or b;
    layer7_outputs(6695) <= a xor b;
    layer7_outputs(6696) <= not b;
    layer7_outputs(6697) <= not a;
    layer7_outputs(6698) <= not (a xor b);
    layer7_outputs(6699) <= not (a or b);
    layer7_outputs(6700) <= a xor b;
    layer7_outputs(6701) <= not b;
    layer7_outputs(6702) <= a;
    layer7_outputs(6703) <= a xor b;
    layer7_outputs(6704) <= not b or a;
    layer7_outputs(6705) <= not a;
    layer7_outputs(6706) <= not b or a;
    layer7_outputs(6707) <= b;
    layer7_outputs(6708) <= b;
    layer7_outputs(6709) <= a xor b;
    layer7_outputs(6710) <= a and not b;
    layer7_outputs(6711) <= b;
    layer7_outputs(6712) <= a xor b;
    layer7_outputs(6713) <= a xor b;
    layer7_outputs(6714) <= a or b;
    layer7_outputs(6715) <= not (a and b);
    layer7_outputs(6716) <= not a;
    layer7_outputs(6717) <= not (a or b);
    layer7_outputs(6718) <= b;
    layer7_outputs(6719) <= b;
    layer7_outputs(6720) <= b;
    layer7_outputs(6721) <= not (a xor b);
    layer7_outputs(6722) <= not b;
    layer7_outputs(6723) <= b and not a;
    layer7_outputs(6724) <= a or b;
    layer7_outputs(6725) <= not a or b;
    layer7_outputs(6726) <= a;
    layer7_outputs(6727) <= b and not a;
    layer7_outputs(6728) <= not b or a;
    layer7_outputs(6729) <= not (a and b);
    layer7_outputs(6730) <= b;
    layer7_outputs(6731) <= a or b;
    layer7_outputs(6732) <= not b or a;
    layer7_outputs(6733) <= a;
    layer7_outputs(6734) <= b;
    layer7_outputs(6735) <= not (a or b);
    layer7_outputs(6736) <= a or b;
    layer7_outputs(6737) <= not (a xor b);
    layer7_outputs(6738) <= a or b;
    layer7_outputs(6739) <= not b or a;
    layer7_outputs(6740) <= a and b;
    layer7_outputs(6741) <= a;
    layer7_outputs(6742) <= not (a xor b);
    layer7_outputs(6743) <= not (a xor b);
    layer7_outputs(6744) <= a;
    layer7_outputs(6745) <= not a or b;
    layer7_outputs(6746) <= not b or a;
    layer7_outputs(6747) <= a xor b;
    layer7_outputs(6748) <= a and b;
    layer7_outputs(6749) <= 1'b1;
    layer7_outputs(6750) <= not (a xor b);
    layer7_outputs(6751) <= not a or b;
    layer7_outputs(6752) <= not a;
    layer7_outputs(6753) <= b;
    layer7_outputs(6754) <= not (a xor b);
    layer7_outputs(6755) <= b;
    layer7_outputs(6756) <= b and not a;
    layer7_outputs(6757) <= not a;
    layer7_outputs(6758) <= not a;
    layer7_outputs(6759) <= a;
    layer7_outputs(6760) <= b;
    layer7_outputs(6761) <= a and b;
    layer7_outputs(6762) <= not a;
    layer7_outputs(6763) <= a;
    layer7_outputs(6764) <= a xor b;
    layer7_outputs(6765) <= not a or b;
    layer7_outputs(6766) <= not b;
    layer7_outputs(6767) <= a;
    layer7_outputs(6768) <= a;
    layer7_outputs(6769) <= a and b;
    layer7_outputs(6770) <= a and not b;
    layer7_outputs(6771) <= b;
    layer7_outputs(6772) <= not b;
    layer7_outputs(6773) <= not b;
    layer7_outputs(6774) <= not a;
    layer7_outputs(6775) <= a xor b;
    layer7_outputs(6776) <= a and not b;
    layer7_outputs(6777) <= not a or b;
    layer7_outputs(6778) <= b and not a;
    layer7_outputs(6779) <= a;
    layer7_outputs(6780) <= a;
    layer7_outputs(6781) <= 1'b0;
    layer7_outputs(6782) <= not (a xor b);
    layer7_outputs(6783) <= not (a and b);
    layer7_outputs(6784) <= not a or b;
    layer7_outputs(6785) <= not (a xor b);
    layer7_outputs(6786) <= not (a or b);
    layer7_outputs(6787) <= b;
    layer7_outputs(6788) <= not (a or b);
    layer7_outputs(6789) <= not b;
    layer7_outputs(6790) <= a xor b;
    layer7_outputs(6791) <= not a;
    layer7_outputs(6792) <= not b;
    layer7_outputs(6793) <= a;
    layer7_outputs(6794) <= not (a xor b);
    layer7_outputs(6795) <= not a;
    layer7_outputs(6796) <= not (a and b);
    layer7_outputs(6797) <= not (a or b);
    layer7_outputs(6798) <= a;
    layer7_outputs(6799) <= a or b;
    layer7_outputs(6800) <= not b;
    layer7_outputs(6801) <= not (a xor b);
    layer7_outputs(6802) <= a;
    layer7_outputs(6803) <= not a;
    layer7_outputs(6804) <= not a or b;
    layer7_outputs(6805) <= not b or a;
    layer7_outputs(6806) <= not b;
    layer7_outputs(6807) <= not a or b;
    layer7_outputs(6808) <= a xor b;
    layer7_outputs(6809) <= a xor b;
    layer7_outputs(6810) <= b;
    layer7_outputs(6811) <= not (a or b);
    layer7_outputs(6812) <= a and b;
    layer7_outputs(6813) <= not (a xor b);
    layer7_outputs(6814) <= a and not b;
    layer7_outputs(6815) <= not (a xor b);
    layer7_outputs(6816) <= a and b;
    layer7_outputs(6817) <= not b;
    layer7_outputs(6818) <= not a;
    layer7_outputs(6819) <= not a or b;
    layer7_outputs(6820) <= a;
    layer7_outputs(6821) <= b;
    layer7_outputs(6822) <= a;
    layer7_outputs(6823) <= a;
    layer7_outputs(6824) <= not (a xor b);
    layer7_outputs(6825) <= not (a or b);
    layer7_outputs(6826) <= not a;
    layer7_outputs(6827) <= not (a or b);
    layer7_outputs(6828) <= a or b;
    layer7_outputs(6829) <= not a or b;
    layer7_outputs(6830) <= b and not a;
    layer7_outputs(6831) <= b and not a;
    layer7_outputs(6832) <= not (a xor b);
    layer7_outputs(6833) <= not a;
    layer7_outputs(6834) <= not a;
    layer7_outputs(6835) <= a and b;
    layer7_outputs(6836) <= a and not b;
    layer7_outputs(6837) <= 1'b1;
    layer7_outputs(6838) <= not (a and b);
    layer7_outputs(6839) <= a;
    layer7_outputs(6840) <= a and b;
    layer7_outputs(6841) <= not a;
    layer7_outputs(6842) <= not b;
    layer7_outputs(6843) <= not b;
    layer7_outputs(6844) <= b and not a;
    layer7_outputs(6845) <= not a;
    layer7_outputs(6846) <= not b;
    layer7_outputs(6847) <= not (a or b);
    layer7_outputs(6848) <= not a;
    layer7_outputs(6849) <= b;
    layer7_outputs(6850) <= a;
    layer7_outputs(6851) <= a or b;
    layer7_outputs(6852) <= a or b;
    layer7_outputs(6853) <= not a;
    layer7_outputs(6854) <= a;
    layer7_outputs(6855) <= a;
    layer7_outputs(6856) <= not b;
    layer7_outputs(6857) <= not a;
    layer7_outputs(6858) <= not a or b;
    layer7_outputs(6859) <= not (a xor b);
    layer7_outputs(6860) <= not a;
    layer7_outputs(6861) <= not b or a;
    layer7_outputs(6862) <= not (a xor b);
    layer7_outputs(6863) <= a and b;
    layer7_outputs(6864) <= a;
    layer7_outputs(6865) <= a;
    layer7_outputs(6866) <= b;
    layer7_outputs(6867) <= a xor b;
    layer7_outputs(6868) <= a and not b;
    layer7_outputs(6869) <= a xor b;
    layer7_outputs(6870) <= a or b;
    layer7_outputs(6871) <= a and b;
    layer7_outputs(6872) <= not a or b;
    layer7_outputs(6873) <= not a;
    layer7_outputs(6874) <= not (a or b);
    layer7_outputs(6875) <= a and not b;
    layer7_outputs(6876) <= not a;
    layer7_outputs(6877) <= not a;
    layer7_outputs(6878) <= b;
    layer7_outputs(6879) <= a and not b;
    layer7_outputs(6880) <= b;
    layer7_outputs(6881) <= a or b;
    layer7_outputs(6882) <= a or b;
    layer7_outputs(6883) <= not b or a;
    layer7_outputs(6884) <= a or b;
    layer7_outputs(6885) <= b;
    layer7_outputs(6886) <= b;
    layer7_outputs(6887) <= not (a and b);
    layer7_outputs(6888) <= not (a or b);
    layer7_outputs(6889) <= b;
    layer7_outputs(6890) <= not (a xor b);
    layer7_outputs(6891) <= not a;
    layer7_outputs(6892) <= not (a xor b);
    layer7_outputs(6893) <= a xor b;
    layer7_outputs(6894) <= not a;
    layer7_outputs(6895) <= b;
    layer7_outputs(6896) <= not b or a;
    layer7_outputs(6897) <= not a;
    layer7_outputs(6898) <= not b;
    layer7_outputs(6899) <= 1'b1;
    layer7_outputs(6900) <= a and b;
    layer7_outputs(6901) <= not b;
    layer7_outputs(6902) <= not a or b;
    layer7_outputs(6903) <= b;
    layer7_outputs(6904) <= b;
    layer7_outputs(6905) <= a and b;
    layer7_outputs(6906) <= not (a xor b);
    layer7_outputs(6907) <= a;
    layer7_outputs(6908) <= a and b;
    layer7_outputs(6909) <= a and b;
    layer7_outputs(6910) <= a or b;
    layer7_outputs(6911) <= not b;
    layer7_outputs(6912) <= not (a or b);
    layer7_outputs(6913) <= a xor b;
    layer7_outputs(6914) <= a and not b;
    layer7_outputs(6915) <= not a;
    layer7_outputs(6916) <= not (a and b);
    layer7_outputs(6917) <= not b;
    layer7_outputs(6918) <= a xor b;
    layer7_outputs(6919) <= not b;
    layer7_outputs(6920) <= not (a and b);
    layer7_outputs(6921) <= a and not b;
    layer7_outputs(6922) <= not b;
    layer7_outputs(6923) <= a or b;
    layer7_outputs(6924) <= not a or b;
    layer7_outputs(6925) <= b;
    layer7_outputs(6926) <= b;
    layer7_outputs(6927) <= 1'b1;
    layer7_outputs(6928) <= b;
    layer7_outputs(6929) <= not a;
    layer7_outputs(6930) <= not (a xor b);
    layer7_outputs(6931) <= not b or a;
    layer7_outputs(6932) <= a;
    layer7_outputs(6933) <= b;
    layer7_outputs(6934) <= a;
    layer7_outputs(6935) <= not b;
    layer7_outputs(6936) <= not b;
    layer7_outputs(6937) <= a;
    layer7_outputs(6938) <= b;
    layer7_outputs(6939) <= not a or b;
    layer7_outputs(6940) <= not b;
    layer7_outputs(6941) <= not b;
    layer7_outputs(6942) <= a xor b;
    layer7_outputs(6943) <= not a;
    layer7_outputs(6944) <= not b;
    layer7_outputs(6945) <= 1'b0;
    layer7_outputs(6946) <= a xor b;
    layer7_outputs(6947) <= a;
    layer7_outputs(6948) <= not a;
    layer7_outputs(6949) <= not a or b;
    layer7_outputs(6950) <= a and b;
    layer7_outputs(6951) <= not b;
    layer7_outputs(6952) <= 1'b1;
    layer7_outputs(6953) <= not a or b;
    layer7_outputs(6954) <= a and not b;
    layer7_outputs(6955) <= a and not b;
    layer7_outputs(6956) <= not (a and b);
    layer7_outputs(6957) <= b and not a;
    layer7_outputs(6958) <= 1'b0;
    layer7_outputs(6959) <= b;
    layer7_outputs(6960) <= 1'b1;
    layer7_outputs(6961) <= not a or b;
    layer7_outputs(6962) <= not (a or b);
    layer7_outputs(6963) <= not (a and b);
    layer7_outputs(6964) <= a;
    layer7_outputs(6965) <= not a;
    layer7_outputs(6966) <= a xor b;
    layer7_outputs(6967) <= a;
    layer7_outputs(6968) <= a;
    layer7_outputs(6969) <= not a;
    layer7_outputs(6970) <= b and not a;
    layer7_outputs(6971) <= not (a or b);
    layer7_outputs(6972) <= not b or a;
    layer7_outputs(6973) <= not (a xor b);
    layer7_outputs(6974) <= not b;
    layer7_outputs(6975) <= not (a xor b);
    layer7_outputs(6976) <= b and not a;
    layer7_outputs(6977) <= not a;
    layer7_outputs(6978) <= a xor b;
    layer7_outputs(6979) <= b;
    layer7_outputs(6980) <= not b or a;
    layer7_outputs(6981) <= b;
    layer7_outputs(6982) <= a xor b;
    layer7_outputs(6983) <= a xor b;
    layer7_outputs(6984) <= 1'b0;
    layer7_outputs(6985) <= not a or b;
    layer7_outputs(6986) <= b and not a;
    layer7_outputs(6987) <= not a;
    layer7_outputs(6988) <= a xor b;
    layer7_outputs(6989) <= not (a xor b);
    layer7_outputs(6990) <= not a;
    layer7_outputs(6991) <= 1'b0;
    layer7_outputs(6992) <= not b or a;
    layer7_outputs(6993) <= not a;
    layer7_outputs(6994) <= 1'b0;
    layer7_outputs(6995) <= a;
    layer7_outputs(6996) <= not b;
    layer7_outputs(6997) <= 1'b0;
    layer7_outputs(6998) <= b and not a;
    layer7_outputs(6999) <= b and not a;
    layer7_outputs(7000) <= not (a or b);
    layer7_outputs(7001) <= not (a and b);
    layer7_outputs(7002) <= a and not b;
    layer7_outputs(7003) <= not b;
    layer7_outputs(7004) <= a;
    layer7_outputs(7005) <= not b;
    layer7_outputs(7006) <= not a or b;
    layer7_outputs(7007) <= not b or a;
    layer7_outputs(7008) <= not b or a;
    layer7_outputs(7009) <= not a or b;
    layer7_outputs(7010) <= not a;
    layer7_outputs(7011) <= a or b;
    layer7_outputs(7012) <= a xor b;
    layer7_outputs(7013) <= not a or b;
    layer7_outputs(7014) <= a;
    layer7_outputs(7015) <= a and b;
    layer7_outputs(7016) <= not (a xor b);
    layer7_outputs(7017) <= a and b;
    layer7_outputs(7018) <= b and not a;
    layer7_outputs(7019) <= a and not b;
    layer7_outputs(7020) <= b;
    layer7_outputs(7021) <= not (a and b);
    layer7_outputs(7022) <= not a;
    layer7_outputs(7023) <= b and not a;
    layer7_outputs(7024) <= a and not b;
    layer7_outputs(7025) <= b;
    layer7_outputs(7026) <= not (a xor b);
    layer7_outputs(7027) <= not b;
    layer7_outputs(7028) <= not (a xor b);
    layer7_outputs(7029) <= not b;
    layer7_outputs(7030) <= not a;
    layer7_outputs(7031) <= not (a xor b);
    layer7_outputs(7032) <= not b or a;
    layer7_outputs(7033) <= not a;
    layer7_outputs(7034) <= not (a xor b);
    layer7_outputs(7035) <= not a or b;
    layer7_outputs(7036) <= not b or a;
    layer7_outputs(7037) <= not b;
    layer7_outputs(7038) <= a or b;
    layer7_outputs(7039) <= not (a xor b);
    layer7_outputs(7040) <= not (a or b);
    layer7_outputs(7041) <= a and not b;
    layer7_outputs(7042) <= not (a xor b);
    layer7_outputs(7043) <= b and not a;
    layer7_outputs(7044) <= a;
    layer7_outputs(7045) <= not (a xor b);
    layer7_outputs(7046) <= b;
    layer7_outputs(7047) <= not (a xor b);
    layer7_outputs(7048) <= not a or b;
    layer7_outputs(7049) <= b;
    layer7_outputs(7050) <= not (a and b);
    layer7_outputs(7051) <= a and b;
    layer7_outputs(7052) <= not b or a;
    layer7_outputs(7053) <= not (a or b);
    layer7_outputs(7054) <= a;
    layer7_outputs(7055) <= not a or b;
    layer7_outputs(7056) <= b;
    layer7_outputs(7057) <= not a;
    layer7_outputs(7058) <= not (a xor b);
    layer7_outputs(7059) <= a and b;
    layer7_outputs(7060) <= 1'b0;
    layer7_outputs(7061) <= b and not a;
    layer7_outputs(7062) <= b;
    layer7_outputs(7063) <= a;
    layer7_outputs(7064) <= a;
    layer7_outputs(7065) <= not b;
    layer7_outputs(7066) <= not b or a;
    layer7_outputs(7067) <= not a;
    layer7_outputs(7068) <= not (a or b);
    layer7_outputs(7069) <= a xor b;
    layer7_outputs(7070) <= 1'b0;
    layer7_outputs(7071) <= b and not a;
    layer7_outputs(7072) <= not (a xor b);
    layer7_outputs(7073) <= not (a xor b);
    layer7_outputs(7074) <= not a;
    layer7_outputs(7075) <= not (a xor b);
    layer7_outputs(7076) <= not b;
    layer7_outputs(7077) <= not b;
    layer7_outputs(7078) <= a;
    layer7_outputs(7079) <= a and b;
    layer7_outputs(7080) <= a and b;
    layer7_outputs(7081) <= not b or a;
    layer7_outputs(7082) <= not (a or b);
    layer7_outputs(7083) <= not (a and b);
    layer7_outputs(7084) <= a;
    layer7_outputs(7085) <= b and not a;
    layer7_outputs(7086) <= a or b;
    layer7_outputs(7087) <= a and b;
    layer7_outputs(7088) <= a;
    layer7_outputs(7089) <= b and not a;
    layer7_outputs(7090) <= not a;
    layer7_outputs(7091) <= not a;
    layer7_outputs(7092) <= not (a or b);
    layer7_outputs(7093) <= a;
    layer7_outputs(7094) <= not a;
    layer7_outputs(7095) <= not b;
    layer7_outputs(7096) <= a;
    layer7_outputs(7097) <= not (a or b);
    layer7_outputs(7098) <= not (a and b);
    layer7_outputs(7099) <= a xor b;
    layer7_outputs(7100) <= a or b;
    layer7_outputs(7101) <= a xor b;
    layer7_outputs(7102) <= not (a or b);
    layer7_outputs(7103) <= b;
    layer7_outputs(7104) <= not (a and b);
    layer7_outputs(7105) <= not a;
    layer7_outputs(7106) <= not a or b;
    layer7_outputs(7107) <= a and b;
    layer7_outputs(7108) <= not a;
    layer7_outputs(7109) <= not a;
    layer7_outputs(7110) <= not b;
    layer7_outputs(7111) <= 1'b0;
    layer7_outputs(7112) <= not a;
    layer7_outputs(7113) <= b;
    layer7_outputs(7114) <= not a or b;
    layer7_outputs(7115) <= not (a and b);
    layer7_outputs(7116) <= not a or b;
    layer7_outputs(7117) <= not a or b;
    layer7_outputs(7118) <= not b or a;
    layer7_outputs(7119) <= not a or b;
    layer7_outputs(7120) <= not a;
    layer7_outputs(7121) <= not a or b;
    layer7_outputs(7122) <= not (a xor b);
    layer7_outputs(7123) <= a and b;
    layer7_outputs(7124) <= not (a or b);
    layer7_outputs(7125) <= not (a xor b);
    layer7_outputs(7126) <= b;
    layer7_outputs(7127) <= a and not b;
    layer7_outputs(7128) <= not b;
    layer7_outputs(7129) <= a;
    layer7_outputs(7130) <= not (a or b);
    layer7_outputs(7131) <= not b;
    layer7_outputs(7132) <= not a;
    layer7_outputs(7133) <= b;
    layer7_outputs(7134) <= a xor b;
    layer7_outputs(7135) <= a;
    layer7_outputs(7136) <= a and not b;
    layer7_outputs(7137) <= not b or a;
    layer7_outputs(7138) <= not (a xor b);
    layer7_outputs(7139) <= not a;
    layer7_outputs(7140) <= not (a and b);
    layer7_outputs(7141) <= not a;
    layer7_outputs(7142) <= b;
    layer7_outputs(7143) <= not a;
    layer7_outputs(7144) <= b and not a;
    layer7_outputs(7145) <= b;
    layer7_outputs(7146) <= a xor b;
    layer7_outputs(7147) <= a;
    layer7_outputs(7148) <= b;
    layer7_outputs(7149) <= not a;
    layer7_outputs(7150) <= a xor b;
    layer7_outputs(7151) <= a xor b;
    layer7_outputs(7152) <= not b;
    layer7_outputs(7153) <= not b;
    layer7_outputs(7154) <= not a;
    layer7_outputs(7155) <= 1'b1;
    layer7_outputs(7156) <= 1'b0;
    layer7_outputs(7157) <= a xor b;
    layer7_outputs(7158) <= a;
    layer7_outputs(7159) <= a and not b;
    layer7_outputs(7160) <= a;
    layer7_outputs(7161) <= not (a xor b);
    layer7_outputs(7162) <= a and not b;
    layer7_outputs(7163) <= a or b;
    layer7_outputs(7164) <= a and not b;
    layer7_outputs(7165) <= a;
    layer7_outputs(7166) <= not a or b;
    layer7_outputs(7167) <= not a;
    layer7_outputs(7168) <= not (a xor b);
    layer7_outputs(7169) <= b;
    layer7_outputs(7170) <= b;
    layer7_outputs(7171) <= not a or b;
    layer7_outputs(7172) <= b;
    layer7_outputs(7173) <= a or b;
    layer7_outputs(7174) <= not a;
    layer7_outputs(7175) <= a xor b;
    layer7_outputs(7176) <= not b;
    layer7_outputs(7177) <= not b or a;
    layer7_outputs(7178) <= a xor b;
    layer7_outputs(7179) <= a and not b;
    layer7_outputs(7180) <= a;
    layer7_outputs(7181) <= not (a and b);
    layer7_outputs(7182) <= not (a xor b);
    layer7_outputs(7183) <= not (a xor b);
    layer7_outputs(7184) <= a;
    layer7_outputs(7185) <= not (a or b);
    layer7_outputs(7186) <= b and not a;
    layer7_outputs(7187) <= not a;
    layer7_outputs(7188) <= not (a xor b);
    layer7_outputs(7189) <= a and not b;
    layer7_outputs(7190) <= not b;
    layer7_outputs(7191) <= not b or a;
    layer7_outputs(7192) <= not (a xor b);
    layer7_outputs(7193) <= a or b;
    layer7_outputs(7194) <= not (a xor b);
    layer7_outputs(7195) <= a;
    layer7_outputs(7196) <= not (a xor b);
    layer7_outputs(7197) <= not b;
    layer7_outputs(7198) <= not (a or b);
    layer7_outputs(7199) <= not b;
    layer7_outputs(7200) <= not (a and b);
    layer7_outputs(7201) <= not b;
    layer7_outputs(7202) <= not b;
    layer7_outputs(7203) <= not a;
    layer7_outputs(7204) <= b and not a;
    layer7_outputs(7205) <= not (a and b);
    layer7_outputs(7206) <= a xor b;
    layer7_outputs(7207) <= a;
    layer7_outputs(7208) <= a and b;
    layer7_outputs(7209) <= not a or b;
    layer7_outputs(7210) <= a or b;
    layer7_outputs(7211) <= 1'b0;
    layer7_outputs(7212) <= not a or b;
    layer7_outputs(7213) <= not a;
    layer7_outputs(7214) <= a;
    layer7_outputs(7215) <= a xor b;
    layer7_outputs(7216) <= b and not a;
    layer7_outputs(7217) <= not (a or b);
    layer7_outputs(7218) <= not (a or b);
    layer7_outputs(7219) <= not b;
    layer7_outputs(7220) <= not a;
    layer7_outputs(7221) <= b;
    layer7_outputs(7222) <= b and not a;
    layer7_outputs(7223) <= a;
    layer7_outputs(7224) <= not a or b;
    layer7_outputs(7225) <= not b;
    layer7_outputs(7226) <= a;
    layer7_outputs(7227) <= not (a xor b);
    layer7_outputs(7228) <= b;
    layer7_outputs(7229) <= not a or b;
    layer7_outputs(7230) <= not (a or b);
    layer7_outputs(7231) <= b and not a;
    layer7_outputs(7232) <= a;
    layer7_outputs(7233) <= b and not a;
    layer7_outputs(7234) <= a;
    layer7_outputs(7235) <= not a;
    layer7_outputs(7236) <= b;
    layer7_outputs(7237) <= b;
    layer7_outputs(7238) <= not a;
    layer7_outputs(7239) <= a xor b;
    layer7_outputs(7240) <= a xor b;
    layer7_outputs(7241) <= not (a and b);
    layer7_outputs(7242) <= a xor b;
    layer7_outputs(7243) <= b;
    layer7_outputs(7244) <= not (a xor b);
    layer7_outputs(7245) <= a;
    layer7_outputs(7246) <= a or b;
    layer7_outputs(7247) <= a or b;
    layer7_outputs(7248) <= not a;
    layer7_outputs(7249) <= a xor b;
    layer7_outputs(7250) <= not b;
    layer7_outputs(7251) <= b;
    layer7_outputs(7252) <= not (a and b);
    layer7_outputs(7253) <= not a;
    layer7_outputs(7254) <= a xor b;
    layer7_outputs(7255) <= b;
    layer7_outputs(7256) <= 1'b0;
    layer7_outputs(7257) <= a;
    layer7_outputs(7258) <= 1'b0;
    layer7_outputs(7259) <= a or b;
    layer7_outputs(7260) <= not (a or b);
    layer7_outputs(7261) <= a;
    layer7_outputs(7262) <= a xor b;
    layer7_outputs(7263) <= a;
    layer7_outputs(7264) <= a and b;
    layer7_outputs(7265) <= not (a xor b);
    layer7_outputs(7266) <= a;
    layer7_outputs(7267) <= not (a or b);
    layer7_outputs(7268) <= b;
    layer7_outputs(7269) <= not (a xor b);
    layer7_outputs(7270) <= not a;
    layer7_outputs(7271) <= not b;
    layer7_outputs(7272) <= not b;
    layer7_outputs(7273) <= not (a xor b);
    layer7_outputs(7274) <= b;
    layer7_outputs(7275) <= not b;
    layer7_outputs(7276) <= b;
    layer7_outputs(7277) <= not (a or b);
    layer7_outputs(7278) <= not (a or b);
    layer7_outputs(7279) <= not a;
    layer7_outputs(7280) <= b and not a;
    layer7_outputs(7281) <= b and not a;
    layer7_outputs(7282) <= not b;
    layer7_outputs(7283) <= a or b;
    layer7_outputs(7284) <= not a;
    layer7_outputs(7285) <= a or b;
    layer7_outputs(7286) <= b and not a;
    layer7_outputs(7287) <= a;
    layer7_outputs(7288) <= b and not a;
    layer7_outputs(7289) <= not b;
    layer7_outputs(7290) <= not b;
    layer7_outputs(7291) <= b;
    layer7_outputs(7292) <= a xor b;
    layer7_outputs(7293) <= a and not b;
    layer7_outputs(7294) <= not (a and b);
    layer7_outputs(7295) <= b;
    layer7_outputs(7296) <= not (a xor b);
    layer7_outputs(7297) <= not b;
    layer7_outputs(7298) <= not (a xor b);
    layer7_outputs(7299) <= a;
    layer7_outputs(7300) <= not b or a;
    layer7_outputs(7301) <= b;
    layer7_outputs(7302) <= not b;
    layer7_outputs(7303) <= not (a or b);
    layer7_outputs(7304) <= a and not b;
    layer7_outputs(7305) <= a xor b;
    layer7_outputs(7306) <= not (a xor b);
    layer7_outputs(7307) <= a;
    layer7_outputs(7308) <= not b;
    layer7_outputs(7309) <= not b;
    layer7_outputs(7310) <= not b or a;
    layer7_outputs(7311) <= not b;
    layer7_outputs(7312) <= b and not a;
    layer7_outputs(7313) <= b and not a;
    layer7_outputs(7314) <= a xor b;
    layer7_outputs(7315) <= not (a xor b);
    layer7_outputs(7316) <= not a;
    layer7_outputs(7317) <= not a or b;
    layer7_outputs(7318) <= a xor b;
    layer7_outputs(7319) <= 1'b1;
    layer7_outputs(7320) <= not (a or b);
    layer7_outputs(7321) <= a xor b;
    layer7_outputs(7322) <= a and not b;
    layer7_outputs(7323) <= not a;
    layer7_outputs(7324) <= not (a or b);
    layer7_outputs(7325) <= not a or b;
    layer7_outputs(7326) <= a xor b;
    layer7_outputs(7327) <= a and not b;
    layer7_outputs(7328) <= not a;
    layer7_outputs(7329) <= a or b;
    layer7_outputs(7330) <= b;
    layer7_outputs(7331) <= a and not b;
    layer7_outputs(7332) <= b;
    layer7_outputs(7333) <= a;
    layer7_outputs(7334) <= not a or b;
    layer7_outputs(7335) <= b;
    layer7_outputs(7336) <= b;
    layer7_outputs(7337) <= not (a xor b);
    layer7_outputs(7338) <= a xor b;
    layer7_outputs(7339) <= not b;
    layer7_outputs(7340) <= not (a xor b);
    layer7_outputs(7341) <= not (a xor b);
    layer7_outputs(7342) <= not (a xor b);
    layer7_outputs(7343) <= not b;
    layer7_outputs(7344) <= a xor b;
    layer7_outputs(7345) <= not (a xor b);
    layer7_outputs(7346) <= a and b;
    layer7_outputs(7347) <= b and not a;
    layer7_outputs(7348) <= not b;
    layer7_outputs(7349) <= a;
    layer7_outputs(7350) <= b;
    layer7_outputs(7351) <= a xor b;
    layer7_outputs(7352) <= a or b;
    layer7_outputs(7353) <= b;
    layer7_outputs(7354) <= b;
    layer7_outputs(7355) <= not b;
    layer7_outputs(7356) <= not b;
    layer7_outputs(7357) <= b;
    layer7_outputs(7358) <= b;
    layer7_outputs(7359) <= not b;
    layer7_outputs(7360) <= not b;
    layer7_outputs(7361) <= a or b;
    layer7_outputs(7362) <= a or b;
    layer7_outputs(7363) <= not a;
    layer7_outputs(7364) <= not (a xor b);
    layer7_outputs(7365) <= b;
    layer7_outputs(7366) <= not a;
    layer7_outputs(7367) <= not a;
    layer7_outputs(7368) <= not a or b;
    layer7_outputs(7369) <= not (a xor b);
    layer7_outputs(7370) <= a xor b;
    layer7_outputs(7371) <= not b or a;
    layer7_outputs(7372) <= not b or a;
    layer7_outputs(7373) <= not a;
    layer7_outputs(7374) <= a;
    layer7_outputs(7375) <= a and b;
    layer7_outputs(7376) <= b and not a;
    layer7_outputs(7377) <= a;
    layer7_outputs(7378) <= a;
    layer7_outputs(7379) <= not b;
    layer7_outputs(7380) <= a and b;
    layer7_outputs(7381) <= not a;
    layer7_outputs(7382) <= not b;
    layer7_outputs(7383) <= not b;
    layer7_outputs(7384) <= a and b;
    layer7_outputs(7385) <= a or b;
    layer7_outputs(7386) <= b;
    layer7_outputs(7387) <= b;
    layer7_outputs(7388) <= not a or b;
    layer7_outputs(7389) <= b;
    layer7_outputs(7390) <= a;
    layer7_outputs(7391) <= a;
    layer7_outputs(7392) <= b and not a;
    layer7_outputs(7393) <= a and not b;
    layer7_outputs(7394) <= b and not a;
    layer7_outputs(7395) <= not b or a;
    layer7_outputs(7396) <= not a or b;
    layer7_outputs(7397) <= not (a xor b);
    layer7_outputs(7398) <= not b;
    layer7_outputs(7399) <= a xor b;
    layer7_outputs(7400) <= 1'b1;
    layer7_outputs(7401) <= not (a xor b);
    layer7_outputs(7402) <= not (a or b);
    layer7_outputs(7403) <= a;
    layer7_outputs(7404) <= b;
    layer7_outputs(7405) <= b;
    layer7_outputs(7406) <= a xor b;
    layer7_outputs(7407) <= b and not a;
    layer7_outputs(7408) <= not (a or b);
    layer7_outputs(7409) <= not (a and b);
    layer7_outputs(7410) <= not b;
    layer7_outputs(7411) <= a and not b;
    layer7_outputs(7412) <= a xor b;
    layer7_outputs(7413) <= not (a xor b);
    layer7_outputs(7414) <= not b or a;
    layer7_outputs(7415) <= a xor b;
    layer7_outputs(7416) <= a and not b;
    layer7_outputs(7417) <= a xor b;
    layer7_outputs(7418) <= a and b;
    layer7_outputs(7419) <= not a;
    layer7_outputs(7420) <= not a or b;
    layer7_outputs(7421) <= a;
    layer7_outputs(7422) <= a and b;
    layer7_outputs(7423) <= not (a xor b);
    layer7_outputs(7424) <= not a;
    layer7_outputs(7425) <= a or b;
    layer7_outputs(7426) <= a xor b;
    layer7_outputs(7427) <= a;
    layer7_outputs(7428) <= not (a or b);
    layer7_outputs(7429) <= not a;
    layer7_outputs(7430) <= a or b;
    layer7_outputs(7431) <= not b or a;
    layer7_outputs(7432) <= not b or a;
    layer7_outputs(7433) <= not b or a;
    layer7_outputs(7434) <= b;
    layer7_outputs(7435) <= not a;
    layer7_outputs(7436) <= a xor b;
    layer7_outputs(7437) <= not b or a;
    layer7_outputs(7438) <= not (a or b);
    layer7_outputs(7439) <= b;
    layer7_outputs(7440) <= b;
    layer7_outputs(7441) <= not (a and b);
    layer7_outputs(7442) <= a;
    layer7_outputs(7443) <= a xor b;
    layer7_outputs(7444) <= a xor b;
    layer7_outputs(7445) <= a xor b;
    layer7_outputs(7446) <= a;
    layer7_outputs(7447) <= not a or b;
    layer7_outputs(7448) <= not b;
    layer7_outputs(7449) <= b;
    layer7_outputs(7450) <= not (a xor b);
    layer7_outputs(7451) <= a and b;
    layer7_outputs(7452) <= not b or a;
    layer7_outputs(7453) <= not b;
    layer7_outputs(7454) <= not a;
    layer7_outputs(7455) <= a and not b;
    layer7_outputs(7456) <= not b;
    layer7_outputs(7457) <= a xor b;
    layer7_outputs(7458) <= not (a or b);
    layer7_outputs(7459) <= a and not b;
    layer7_outputs(7460) <= a;
    layer7_outputs(7461) <= not a or b;
    layer7_outputs(7462) <= b;
    layer7_outputs(7463) <= b and not a;
    layer7_outputs(7464) <= not b;
    layer7_outputs(7465) <= a;
    layer7_outputs(7466) <= a xor b;
    layer7_outputs(7467) <= not a or b;
    layer7_outputs(7468) <= a xor b;
    layer7_outputs(7469) <= 1'b1;
    layer7_outputs(7470) <= not b;
    layer7_outputs(7471) <= not b;
    layer7_outputs(7472) <= not a or b;
    layer7_outputs(7473) <= not (a and b);
    layer7_outputs(7474) <= b;
    layer7_outputs(7475) <= 1'b1;
    layer7_outputs(7476) <= a;
    layer7_outputs(7477) <= a and not b;
    layer7_outputs(7478) <= not a;
    layer7_outputs(7479) <= b and not a;
    layer7_outputs(7480) <= b;
    layer7_outputs(7481) <= not a or b;
    layer7_outputs(7482) <= not a;
    layer7_outputs(7483) <= not a;
    layer7_outputs(7484) <= not b or a;
    layer7_outputs(7485) <= a and b;
    layer7_outputs(7486) <= not (a or b);
    layer7_outputs(7487) <= not b or a;
    layer7_outputs(7488) <= b;
    layer7_outputs(7489) <= b;
    layer7_outputs(7490) <= b;
    layer7_outputs(7491) <= b and not a;
    layer7_outputs(7492) <= not b;
    layer7_outputs(7493) <= a;
    layer7_outputs(7494) <= a;
    layer7_outputs(7495) <= a xor b;
    layer7_outputs(7496) <= not b;
    layer7_outputs(7497) <= not a;
    layer7_outputs(7498) <= a;
    layer7_outputs(7499) <= b;
    layer7_outputs(7500) <= a and not b;
    layer7_outputs(7501) <= not b or a;
    layer7_outputs(7502) <= not (a and b);
    layer7_outputs(7503) <= not (a xor b);
    layer7_outputs(7504) <= a or b;
    layer7_outputs(7505) <= not (a xor b);
    layer7_outputs(7506) <= b and not a;
    layer7_outputs(7507) <= a;
    layer7_outputs(7508) <= not a;
    layer7_outputs(7509) <= not a;
    layer7_outputs(7510) <= not a or b;
    layer7_outputs(7511) <= not (a xor b);
    layer7_outputs(7512) <= a and b;
    layer7_outputs(7513) <= not (a xor b);
    layer7_outputs(7514) <= a xor b;
    layer7_outputs(7515) <= a xor b;
    layer7_outputs(7516) <= b;
    layer7_outputs(7517) <= b;
    layer7_outputs(7518) <= b and not a;
    layer7_outputs(7519) <= b and not a;
    layer7_outputs(7520) <= b and not a;
    layer7_outputs(7521) <= b;
    layer7_outputs(7522) <= not a;
    layer7_outputs(7523) <= not a;
    layer7_outputs(7524) <= not (a xor b);
    layer7_outputs(7525) <= not a;
    layer7_outputs(7526) <= not (a or b);
    layer7_outputs(7527) <= not (a xor b);
    layer7_outputs(7528) <= a;
    layer7_outputs(7529) <= a;
    layer7_outputs(7530) <= not (a and b);
    layer7_outputs(7531) <= not (a xor b);
    layer7_outputs(7532) <= not (a xor b);
    layer7_outputs(7533) <= not a or b;
    layer7_outputs(7534) <= b;
    layer7_outputs(7535) <= a;
    layer7_outputs(7536) <= b;
    layer7_outputs(7537) <= not (a xor b);
    layer7_outputs(7538) <= a;
    layer7_outputs(7539) <= a xor b;
    layer7_outputs(7540) <= a and b;
    layer7_outputs(7541) <= not a;
    layer7_outputs(7542) <= a;
    layer7_outputs(7543) <= not a or b;
    layer7_outputs(7544) <= b;
    layer7_outputs(7545) <= a;
    layer7_outputs(7546) <= b and not a;
    layer7_outputs(7547) <= not b;
    layer7_outputs(7548) <= a and b;
    layer7_outputs(7549) <= a xor b;
    layer7_outputs(7550) <= a xor b;
    layer7_outputs(7551) <= a and b;
    layer7_outputs(7552) <= not (a or b);
    layer7_outputs(7553) <= a;
    layer7_outputs(7554) <= b;
    layer7_outputs(7555) <= a xor b;
    layer7_outputs(7556) <= b;
    layer7_outputs(7557) <= b;
    layer7_outputs(7558) <= not a;
    layer7_outputs(7559) <= b;
    layer7_outputs(7560) <= a and not b;
    layer7_outputs(7561) <= not a;
    layer7_outputs(7562) <= not a;
    layer7_outputs(7563) <= not b;
    layer7_outputs(7564) <= b;
    layer7_outputs(7565) <= b;
    layer7_outputs(7566) <= not a;
    layer7_outputs(7567) <= a;
    layer7_outputs(7568) <= b and not a;
    layer7_outputs(7569) <= not b or a;
    layer7_outputs(7570) <= b;
    layer7_outputs(7571) <= not b;
    layer7_outputs(7572) <= not (a xor b);
    layer7_outputs(7573) <= not a;
    layer7_outputs(7574) <= a and b;
    layer7_outputs(7575) <= not b or a;
    layer7_outputs(7576) <= a and not b;
    layer7_outputs(7577) <= a and b;
    layer7_outputs(7578) <= not (a and b);
    layer7_outputs(7579) <= not b or a;
    layer7_outputs(7580) <= not a;
    layer7_outputs(7581) <= b;
    layer7_outputs(7582) <= not a;
    layer7_outputs(7583) <= not (a xor b);
    layer7_outputs(7584) <= not b;
    layer7_outputs(7585) <= 1'b0;
    layer7_outputs(7586) <= a xor b;
    layer7_outputs(7587) <= 1'b1;
    layer7_outputs(7588) <= not a;
    layer7_outputs(7589) <= 1'b1;
    layer7_outputs(7590) <= not (a or b);
    layer7_outputs(7591) <= a or b;
    layer7_outputs(7592) <= not b;
    layer7_outputs(7593) <= b;
    layer7_outputs(7594) <= 1'b0;
    layer7_outputs(7595) <= not b;
    layer7_outputs(7596) <= not (a xor b);
    layer7_outputs(7597) <= a;
    layer7_outputs(7598) <= not (a and b);
    layer7_outputs(7599) <= b;
    layer7_outputs(7600) <= a and b;
    layer7_outputs(7601) <= a xor b;
    layer7_outputs(7602) <= not (a xor b);
    layer7_outputs(7603) <= a;
    layer7_outputs(7604) <= not a;
    layer7_outputs(7605) <= a or b;
    layer7_outputs(7606) <= not (a and b);
    layer7_outputs(7607) <= a or b;
    layer7_outputs(7608) <= not (a xor b);
    layer7_outputs(7609) <= b;
    layer7_outputs(7610) <= b and not a;
    layer7_outputs(7611) <= not a;
    layer7_outputs(7612) <= a and b;
    layer7_outputs(7613) <= b and not a;
    layer7_outputs(7614) <= not (a xor b);
    layer7_outputs(7615) <= not b;
    layer7_outputs(7616) <= not b or a;
    layer7_outputs(7617) <= b;
    layer7_outputs(7618) <= b and not a;
    layer7_outputs(7619) <= not a;
    layer7_outputs(7620) <= not a;
    layer7_outputs(7621) <= not a;
    layer7_outputs(7622) <= a;
    layer7_outputs(7623) <= a and b;
    layer7_outputs(7624) <= not a;
    layer7_outputs(7625) <= b;
    layer7_outputs(7626) <= a xor b;
    layer7_outputs(7627) <= not a or b;
    layer7_outputs(7628) <= a and b;
    layer7_outputs(7629) <= a;
    layer7_outputs(7630) <= a xor b;
    layer7_outputs(7631) <= not b;
    layer7_outputs(7632) <= b;
    layer7_outputs(7633) <= 1'b1;
    layer7_outputs(7634) <= not b or a;
    layer7_outputs(7635) <= a and b;
    layer7_outputs(7636) <= not a;
    layer7_outputs(7637) <= a and not b;
    layer7_outputs(7638) <= b;
    layer7_outputs(7639) <= not (a or b);
    layer7_outputs(7640) <= 1'b0;
    layer7_outputs(7641) <= b;
    layer7_outputs(7642) <= b;
    layer7_outputs(7643) <= not b;
    layer7_outputs(7644) <= not (a and b);
    layer7_outputs(7645) <= not a or b;
    layer7_outputs(7646) <= not a;
    layer7_outputs(7647) <= not (a xor b);
    layer7_outputs(7648) <= not b;
    layer7_outputs(7649) <= a xor b;
    layer7_outputs(7650) <= not a or b;
    layer7_outputs(7651) <= b;
    layer7_outputs(7652) <= a xor b;
    layer7_outputs(7653) <= not b or a;
    layer7_outputs(7654) <= not b;
    layer7_outputs(7655) <= a;
    layer7_outputs(7656) <= not (a or b);
    layer7_outputs(7657) <= b;
    layer7_outputs(7658) <= a or b;
    layer7_outputs(7659) <= not (a xor b);
    layer7_outputs(7660) <= not (a xor b);
    layer7_outputs(7661) <= not a or b;
    layer7_outputs(7662) <= not a;
    layer7_outputs(7663) <= a and not b;
    layer7_outputs(7664) <= not (a xor b);
    layer7_outputs(7665) <= not b;
    layer7_outputs(7666) <= a and b;
    layer7_outputs(7667) <= a or b;
    layer7_outputs(7668) <= not a or b;
    layer7_outputs(7669) <= not a;
    layer7_outputs(7670) <= a;
    layer7_outputs(7671) <= b;
    layer7_outputs(7672) <= not (a and b);
    layer7_outputs(7673) <= a or b;
    layer7_outputs(7674) <= not b;
    layer7_outputs(7675) <= not b or a;
    layer7_outputs(7676) <= a xor b;
    layer7_outputs(7677) <= not (a and b);
    layer7_outputs(7678) <= b and not a;
    layer7_outputs(7679) <= not (a and b);
    layer7_outputs(7680) <= not a or b;
    layer7_outputs(7681) <= a xor b;
    layer7_outputs(7682) <= not a;
    layer7_outputs(7683) <= not (a xor b);
    layer7_outputs(7684) <= b;
    layer7_outputs(7685) <= a;
    layer7_outputs(7686) <= not a;
    layer7_outputs(7687) <= not a;
    layer7_outputs(7688) <= not b;
    layer7_outputs(7689) <= a or b;
    layer7_outputs(7690) <= not (a or b);
    layer7_outputs(7691) <= not a;
    layer7_outputs(7692) <= not a;
    layer7_outputs(7693) <= a xor b;
    layer7_outputs(7694) <= a and not b;
    layer7_outputs(7695) <= not (a and b);
    layer7_outputs(7696) <= not (a and b);
    layer7_outputs(7697) <= not (a xor b);
    layer7_outputs(7698) <= not (a xor b);
    layer7_outputs(7699) <= not (a or b);
    layer7_outputs(7700) <= not b or a;
    layer7_outputs(7701) <= a xor b;
    layer7_outputs(7702) <= not b or a;
    layer7_outputs(7703) <= not a;
    layer7_outputs(7704) <= b;
    layer7_outputs(7705) <= not (a and b);
    layer7_outputs(7706) <= b and not a;
    layer7_outputs(7707) <= a and b;
    layer7_outputs(7708) <= not a;
    layer7_outputs(7709) <= not b;
    layer7_outputs(7710) <= not a;
    layer7_outputs(7711) <= not b;
    layer7_outputs(7712) <= a xor b;
    layer7_outputs(7713) <= not (a xor b);
    layer7_outputs(7714) <= not b;
    layer7_outputs(7715) <= not (a xor b);
    layer7_outputs(7716) <= a xor b;
    layer7_outputs(7717) <= 1'b1;
    layer7_outputs(7718) <= not b or a;
    layer7_outputs(7719) <= a and b;
    layer7_outputs(7720) <= not (a or b);
    layer7_outputs(7721) <= a xor b;
    layer7_outputs(7722) <= b;
    layer7_outputs(7723) <= b;
    layer7_outputs(7724) <= not (a xor b);
    layer7_outputs(7725) <= 1'b0;
    layer7_outputs(7726) <= not (a xor b);
    layer7_outputs(7727) <= not (a and b);
    layer7_outputs(7728) <= a;
    layer7_outputs(7729) <= not a;
    layer7_outputs(7730) <= not b or a;
    layer7_outputs(7731) <= a xor b;
    layer7_outputs(7732) <= b and not a;
    layer7_outputs(7733) <= b;
    layer7_outputs(7734) <= not b;
    layer7_outputs(7735) <= not b or a;
    layer7_outputs(7736) <= b and not a;
    layer7_outputs(7737) <= b;
    layer7_outputs(7738) <= b;
    layer7_outputs(7739) <= not a or b;
    layer7_outputs(7740) <= 1'b1;
    layer7_outputs(7741) <= not (a xor b);
    layer7_outputs(7742) <= not a;
    layer7_outputs(7743) <= b;
    layer7_outputs(7744) <= a;
    layer7_outputs(7745) <= b;
    layer7_outputs(7746) <= not b;
    layer7_outputs(7747) <= a and b;
    layer7_outputs(7748) <= a;
    layer7_outputs(7749) <= a xor b;
    layer7_outputs(7750) <= not (a xor b);
    layer7_outputs(7751) <= a and not b;
    layer7_outputs(7752) <= not a;
    layer7_outputs(7753) <= not a;
    layer7_outputs(7754) <= not b;
    layer7_outputs(7755) <= a;
    layer7_outputs(7756) <= not a;
    layer7_outputs(7757) <= b;
    layer7_outputs(7758) <= not a;
    layer7_outputs(7759) <= not a;
    layer7_outputs(7760) <= a xor b;
    layer7_outputs(7761) <= not (a or b);
    layer7_outputs(7762) <= not (a xor b);
    layer7_outputs(7763) <= a xor b;
    layer7_outputs(7764) <= not a or b;
    layer7_outputs(7765) <= not b;
    layer7_outputs(7766) <= not (a xor b);
    layer7_outputs(7767) <= not (a or b);
    layer7_outputs(7768) <= a;
    layer7_outputs(7769) <= a or b;
    layer7_outputs(7770) <= not a or b;
    layer7_outputs(7771) <= a;
    layer7_outputs(7772) <= not (a and b);
    layer7_outputs(7773) <= not a;
    layer7_outputs(7774) <= b;
    layer7_outputs(7775) <= b;
    layer7_outputs(7776) <= not a;
    layer7_outputs(7777) <= not a;
    layer7_outputs(7778) <= 1'b0;
    layer7_outputs(7779) <= a xor b;
    layer7_outputs(7780) <= b;
    layer7_outputs(7781) <= b;
    layer7_outputs(7782) <= a xor b;
    layer7_outputs(7783) <= a or b;
    layer7_outputs(7784) <= b;
    layer7_outputs(7785) <= not a or b;
    layer7_outputs(7786) <= not a;
    layer7_outputs(7787) <= b;
    layer7_outputs(7788) <= not a;
    layer7_outputs(7789) <= b;
    layer7_outputs(7790) <= b;
    layer7_outputs(7791) <= not b;
    layer7_outputs(7792) <= b;
    layer7_outputs(7793) <= b;
    layer7_outputs(7794) <= a;
    layer7_outputs(7795) <= not (a or b);
    layer7_outputs(7796) <= not b;
    layer7_outputs(7797) <= not (a and b);
    layer7_outputs(7798) <= a;
    layer7_outputs(7799) <= not (a and b);
    layer7_outputs(7800) <= not b;
    layer7_outputs(7801) <= not a;
    layer7_outputs(7802) <= a;
    layer7_outputs(7803) <= not b or a;
    layer7_outputs(7804) <= b and not a;
    layer7_outputs(7805) <= a xor b;
    layer7_outputs(7806) <= b;
    layer7_outputs(7807) <= not b or a;
    layer7_outputs(7808) <= a and not b;
    layer7_outputs(7809) <= a or b;
    layer7_outputs(7810) <= not (a or b);
    layer7_outputs(7811) <= b;
    layer7_outputs(7812) <= a and not b;
    layer7_outputs(7813) <= not b;
    layer7_outputs(7814) <= not (a and b);
    layer7_outputs(7815) <= not a;
    layer7_outputs(7816) <= not a or b;
    layer7_outputs(7817) <= b;
    layer7_outputs(7818) <= b;
    layer7_outputs(7819) <= not (a xor b);
    layer7_outputs(7820) <= not (a and b);
    layer7_outputs(7821) <= a;
    layer7_outputs(7822) <= b;
    layer7_outputs(7823) <= not (a and b);
    layer7_outputs(7824) <= b;
    layer7_outputs(7825) <= not a or b;
    layer7_outputs(7826) <= b;
    layer7_outputs(7827) <= not a or b;
    layer7_outputs(7828) <= not b;
    layer7_outputs(7829) <= a;
    layer7_outputs(7830) <= b and not a;
    layer7_outputs(7831) <= a and not b;
    layer7_outputs(7832) <= not (a xor b);
    layer7_outputs(7833) <= not (a xor b);
    layer7_outputs(7834) <= a and b;
    layer7_outputs(7835) <= a xor b;
    layer7_outputs(7836) <= not (a or b);
    layer7_outputs(7837) <= not (a or b);
    layer7_outputs(7838) <= a and not b;
    layer7_outputs(7839) <= a xor b;
    layer7_outputs(7840) <= not a;
    layer7_outputs(7841) <= b;
    layer7_outputs(7842) <= not (a or b);
    layer7_outputs(7843) <= not b;
    layer7_outputs(7844) <= not a or b;
    layer7_outputs(7845) <= b;
    layer7_outputs(7846) <= a and b;
    layer7_outputs(7847) <= not a;
    layer7_outputs(7848) <= not (a xor b);
    layer7_outputs(7849) <= not (a and b);
    layer7_outputs(7850) <= not b;
    layer7_outputs(7851) <= not b;
    layer7_outputs(7852) <= not b or a;
    layer7_outputs(7853) <= a;
    layer7_outputs(7854) <= not (a and b);
    layer7_outputs(7855) <= b;
    layer7_outputs(7856) <= not a;
    layer7_outputs(7857) <= a;
    layer7_outputs(7858) <= not b or a;
    layer7_outputs(7859) <= not (a and b);
    layer7_outputs(7860) <= a and b;
    layer7_outputs(7861) <= not a;
    layer7_outputs(7862) <= 1'b1;
    layer7_outputs(7863) <= a xor b;
    layer7_outputs(7864) <= a and not b;
    layer7_outputs(7865) <= a and not b;
    layer7_outputs(7866) <= a and b;
    layer7_outputs(7867) <= not (a xor b);
    layer7_outputs(7868) <= a and not b;
    layer7_outputs(7869) <= not (a and b);
    layer7_outputs(7870) <= a;
    layer7_outputs(7871) <= not b;
    layer7_outputs(7872) <= a;
    layer7_outputs(7873) <= not b or a;
    layer7_outputs(7874) <= not a or b;
    layer7_outputs(7875) <= not b;
    layer7_outputs(7876) <= a;
    layer7_outputs(7877) <= b;
    layer7_outputs(7878) <= not (a or b);
    layer7_outputs(7879) <= not (a and b);
    layer7_outputs(7880) <= not (a xor b);
    layer7_outputs(7881) <= a xor b;
    layer7_outputs(7882) <= a xor b;
    layer7_outputs(7883) <= b and not a;
    layer7_outputs(7884) <= not (a xor b);
    layer7_outputs(7885) <= not (a and b);
    layer7_outputs(7886) <= b;
    layer7_outputs(7887) <= not a;
    layer7_outputs(7888) <= b and not a;
    layer7_outputs(7889) <= not a;
    layer7_outputs(7890) <= not (a and b);
    layer7_outputs(7891) <= b;
    layer7_outputs(7892) <= not b;
    layer7_outputs(7893) <= b;
    layer7_outputs(7894) <= b and not a;
    layer7_outputs(7895) <= not (a xor b);
    layer7_outputs(7896) <= b;
    layer7_outputs(7897) <= a and b;
    layer7_outputs(7898) <= b and not a;
    layer7_outputs(7899) <= a and not b;
    layer7_outputs(7900) <= b;
    layer7_outputs(7901) <= not (a xor b);
    layer7_outputs(7902) <= b and not a;
    layer7_outputs(7903) <= b;
    layer7_outputs(7904) <= not b;
    layer7_outputs(7905) <= not (a xor b);
    layer7_outputs(7906) <= not (a xor b);
    layer7_outputs(7907) <= a;
    layer7_outputs(7908) <= not b or a;
    layer7_outputs(7909) <= a;
    layer7_outputs(7910) <= b and not a;
    layer7_outputs(7911) <= a and not b;
    layer7_outputs(7912) <= not a;
    layer7_outputs(7913) <= not (a xor b);
    layer7_outputs(7914) <= a and b;
    layer7_outputs(7915) <= a xor b;
    layer7_outputs(7916) <= 1'b1;
    layer7_outputs(7917) <= a or b;
    layer7_outputs(7918) <= not (a xor b);
    layer7_outputs(7919) <= b;
    layer7_outputs(7920) <= not b;
    layer7_outputs(7921) <= b;
    layer7_outputs(7922) <= not b or a;
    layer7_outputs(7923) <= a;
    layer7_outputs(7924) <= b;
    layer7_outputs(7925) <= a or b;
    layer7_outputs(7926) <= 1'b1;
    layer7_outputs(7927) <= not a;
    layer7_outputs(7928) <= 1'b1;
    layer7_outputs(7929) <= a and b;
    layer7_outputs(7930) <= a xor b;
    layer7_outputs(7931) <= not (a xor b);
    layer7_outputs(7932) <= b;
    layer7_outputs(7933) <= b;
    layer7_outputs(7934) <= a;
    layer7_outputs(7935) <= a;
    layer7_outputs(7936) <= a xor b;
    layer7_outputs(7937) <= b;
    layer7_outputs(7938) <= a and not b;
    layer7_outputs(7939) <= a and not b;
    layer7_outputs(7940) <= a xor b;
    layer7_outputs(7941) <= not b;
    layer7_outputs(7942) <= not b;
    layer7_outputs(7943) <= 1'b0;
    layer7_outputs(7944) <= a;
    layer7_outputs(7945) <= b;
    layer7_outputs(7946) <= b;
    layer7_outputs(7947) <= not a;
    layer7_outputs(7948) <= a or b;
    layer7_outputs(7949) <= not a or b;
    layer7_outputs(7950) <= b and not a;
    layer7_outputs(7951) <= a;
    layer7_outputs(7952) <= a;
    layer7_outputs(7953) <= not (a xor b);
    layer7_outputs(7954) <= a and b;
    layer7_outputs(7955) <= not b;
    layer7_outputs(7956) <= a and not b;
    layer7_outputs(7957) <= a xor b;
    layer7_outputs(7958) <= a and not b;
    layer7_outputs(7959) <= not a;
    layer7_outputs(7960) <= not b;
    layer7_outputs(7961) <= not b or a;
    layer7_outputs(7962) <= not b or a;
    layer7_outputs(7963) <= a;
    layer7_outputs(7964) <= not (a xor b);
    layer7_outputs(7965) <= not b;
    layer7_outputs(7966) <= b and not a;
    layer7_outputs(7967) <= b;
    layer7_outputs(7968) <= a and not b;
    layer7_outputs(7969) <= a;
    layer7_outputs(7970) <= a;
    layer7_outputs(7971) <= not a or b;
    layer7_outputs(7972) <= b;
    layer7_outputs(7973) <= not b;
    layer7_outputs(7974) <= a xor b;
    layer7_outputs(7975) <= a and b;
    layer7_outputs(7976) <= a and b;
    layer7_outputs(7977) <= b and not a;
    layer7_outputs(7978) <= not (a and b);
    layer7_outputs(7979) <= not (a xor b);
    layer7_outputs(7980) <= b;
    layer7_outputs(7981) <= not b;
    layer7_outputs(7982) <= a;
    layer7_outputs(7983) <= a;
    layer7_outputs(7984) <= a and b;
    layer7_outputs(7985) <= not (a xor b);
    layer7_outputs(7986) <= 1'b0;
    layer7_outputs(7987) <= not (a and b);
    layer7_outputs(7988) <= not a;
    layer7_outputs(7989) <= b;
    layer7_outputs(7990) <= not b;
    layer7_outputs(7991) <= a and not b;
    layer7_outputs(7992) <= b and not a;
    layer7_outputs(7993) <= a xor b;
    layer7_outputs(7994) <= not (a xor b);
    layer7_outputs(7995) <= not b or a;
    layer7_outputs(7996) <= not a;
    layer7_outputs(7997) <= not b or a;
    layer7_outputs(7998) <= not a;
    layer7_outputs(7999) <= a xor b;
    layer7_outputs(8000) <= not b;
    layer7_outputs(8001) <= a and not b;
    layer7_outputs(8002) <= not (a xor b);
    layer7_outputs(8003) <= b;
    layer7_outputs(8004) <= not b or a;
    layer7_outputs(8005) <= a or b;
    layer7_outputs(8006) <= a;
    layer7_outputs(8007) <= not a or b;
    layer7_outputs(8008) <= not b;
    layer7_outputs(8009) <= b;
    layer7_outputs(8010) <= not (a and b);
    layer7_outputs(8011) <= not (a xor b);
    layer7_outputs(8012) <= b;
    layer7_outputs(8013) <= not a;
    layer7_outputs(8014) <= a or b;
    layer7_outputs(8015) <= not (a and b);
    layer7_outputs(8016) <= not a or b;
    layer7_outputs(8017) <= not b;
    layer7_outputs(8018) <= not b;
    layer7_outputs(8019) <= not b;
    layer7_outputs(8020) <= a and not b;
    layer7_outputs(8021) <= not b;
    layer7_outputs(8022) <= not b;
    layer7_outputs(8023) <= not b;
    layer7_outputs(8024) <= a and b;
    layer7_outputs(8025) <= not a;
    layer7_outputs(8026) <= a and not b;
    layer7_outputs(8027) <= not (a xor b);
    layer7_outputs(8028) <= a and b;
    layer7_outputs(8029) <= a;
    layer7_outputs(8030) <= a;
    layer7_outputs(8031) <= a and not b;
    layer7_outputs(8032) <= b and not a;
    layer7_outputs(8033) <= not (a or b);
    layer7_outputs(8034) <= not (a and b);
    layer7_outputs(8035) <= not (a xor b);
    layer7_outputs(8036) <= b;
    layer7_outputs(8037) <= not a or b;
    layer7_outputs(8038) <= not (a or b);
    layer7_outputs(8039) <= a or b;
    layer7_outputs(8040) <= a xor b;
    layer7_outputs(8041) <= a;
    layer7_outputs(8042) <= a or b;
    layer7_outputs(8043) <= not (a xor b);
    layer7_outputs(8044) <= not (a xor b);
    layer7_outputs(8045) <= a;
    layer7_outputs(8046) <= not b;
    layer7_outputs(8047) <= b and not a;
    layer7_outputs(8048) <= a or b;
    layer7_outputs(8049) <= not b;
    layer7_outputs(8050) <= not a or b;
    layer7_outputs(8051) <= not a;
    layer7_outputs(8052) <= not b or a;
    layer7_outputs(8053) <= not (a and b);
    layer7_outputs(8054) <= a xor b;
    layer7_outputs(8055) <= not a;
    layer7_outputs(8056) <= b;
    layer7_outputs(8057) <= not b;
    layer7_outputs(8058) <= not a or b;
    layer7_outputs(8059) <= b;
    layer7_outputs(8060) <= not a or b;
    layer7_outputs(8061) <= a;
    layer7_outputs(8062) <= a xor b;
    layer7_outputs(8063) <= a or b;
    layer7_outputs(8064) <= not b or a;
    layer7_outputs(8065) <= not b;
    layer7_outputs(8066) <= not (a or b);
    layer7_outputs(8067) <= a;
    layer7_outputs(8068) <= not a;
    layer7_outputs(8069) <= a or b;
    layer7_outputs(8070) <= a and b;
    layer7_outputs(8071) <= not (a xor b);
    layer7_outputs(8072) <= not b;
    layer7_outputs(8073) <= not b;
    layer7_outputs(8074) <= b;
    layer7_outputs(8075) <= not (a xor b);
    layer7_outputs(8076) <= a;
    layer7_outputs(8077) <= a and b;
    layer7_outputs(8078) <= not a;
    layer7_outputs(8079) <= not b;
    layer7_outputs(8080) <= a and not b;
    layer7_outputs(8081) <= not a;
    layer7_outputs(8082) <= not (a xor b);
    layer7_outputs(8083) <= not a;
    layer7_outputs(8084) <= b;
    layer7_outputs(8085) <= a and not b;
    layer7_outputs(8086) <= b;
    layer7_outputs(8087) <= not a;
    layer7_outputs(8088) <= not (a and b);
    layer7_outputs(8089) <= a and b;
    layer7_outputs(8090) <= b;
    layer7_outputs(8091) <= not a or b;
    layer7_outputs(8092) <= not (a and b);
    layer7_outputs(8093) <= not b or a;
    layer7_outputs(8094) <= b;
    layer7_outputs(8095) <= a and b;
    layer7_outputs(8096) <= a;
    layer7_outputs(8097) <= a;
    layer7_outputs(8098) <= b;
    layer7_outputs(8099) <= not (a and b);
    layer7_outputs(8100) <= b;
    layer7_outputs(8101) <= a xor b;
    layer7_outputs(8102) <= not a;
    layer7_outputs(8103) <= not (a and b);
    layer7_outputs(8104) <= not a;
    layer7_outputs(8105) <= not b;
    layer7_outputs(8106) <= a xor b;
    layer7_outputs(8107) <= 1'b0;
    layer7_outputs(8108) <= b and not a;
    layer7_outputs(8109) <= 1'b0;
    layer7_outputs(8110) <= not (a or b);
    layer7_outputs(8111) <= not a or b;
    layer7_outputs(8112) <= not a;
    layer7_outputs(8113) <= not (a and b);
    layer7_outputs(8114) <= not (a and b);
    layer7_outputs(8115) <= a;
    layer7_outputs(8116) <= not b;
    layer7_outputs(8117) <= a;
    layer7_outputs(8118) <= not (a and b);
    layer7_outputs(8119) <= not a;
    layer7_outputs(8120) <= not (a xor b);
    layer7_outputs(8121) <= b and not a;
    layer7_outputs(8122) <= a and b;
    layer7_outputs(8123) <= not a;
    layer7_outputs(8124) <= not (a or b);
    layer7_outputs(8125) <= 1'b0;
    layer7_outputs(8126) <= b and not a;
    layer7_outputs(8127) <= b and not a;
    layer7_outputs(8128) <= not b;
    layer7_outputs(8129) <= a;
    layer7_outputs(8130) <= b;
    layer7_outputs(8131) <= a xor b;
    layer7_outputs(8132) <= not (a and b);
    layer7_outputs(8133) <= a xor b;
    layer7_outputs(8134) <= not b;
    layer7_outputs(8135) <= a;
    layer7_outputs(8136) <= a;
    layer7_outputs(8137) <= not b or a;
    layer7_outputs(8138) <= a xor b;
    layer7_outputs(8139) <= a and not b;
    layer7_outputs(8140) <= a;
    layer7_outputs(8141) <= a and not b;
    layer7_outputs(8142) <= a or b;
    layer7_outputs(8143) <= not (a xor b);
    layer7_outputs(8144) <= not a;
    layer7_outputs(8145) <= not b;
    layer7_outputs(8146) <= a xor b;
    layer7_outputs(8147) <= b and not a;
    layer7_outputs(8148) <= not b or a;
    layer7_outputs(8149) <= b;
    layer7_outputs(8150) <= not b;
    layer7_outputs(8151) <= not (a xor b);
    layer7_outputs(8152) <= not a;
    layer7_outputs(8153) <= not (a and b);
    layer7_outputs(8154) <= not (a xor b);
    layer7_outputs(8155) <= not b or a;
    layer7_outputs(8156) <= a xor b;
    layer7_outputs(8157) <= a or b;
    layer7_outputs(8158) <= not (a or b);
    layer7_outputs(8159) <= not b;
    layer7_outputs(8160) <= a;
    layer7_outputs(8161) <= a or b;
    layer7_outputs(8162) <= a xor b;
    layer7_outputs(8163) <= not b;
    layer7_outputs(8164) <= not b or a;
    layer7_outputs(8165) <= not a;
    layer7_outputs(8166) <= a or b;
    layer7_outputs(8167) <= not (a or b);
    layer7_outputs(8168) <= not (a and b);
    layer7_outputs(8169) <= a and b;
    layer7_outputs(8170) <= b and not a;
    layer7_outputs(8171) <= a;
    layer7_outputs(8172) <= b;
    layer7_outputs(8173) <= a xor b;
    layer7_outputs(8174) <= a;
    layer7_outputs(8175) <= a xor b;
    layer7_outputs(8176) <= b;
    layer7_outputs(8177) <= a;
    layer7_outputs(8178) <= a and b;
    layer7_outputs(8179) <= a and b;
    layer7_outputs(8180) <= a;
    layer7_outputs(8181) <= not (a and b);
    layer7_outputs(8182) <= not (a xor b);
    layer7_outputs(8183) <= b;
    layer7_outputs(8184) <= a xor b;
    layer7_outputs(8185) <= not (a and b);
    layer7_outputs(8186) <= not (a and b);
    layer7_outputs(8187) <= not b;
    layer7_outputs(8188) <= not a;
    layer7_outputs(8189) <= a and not b;
    layer7_outputs(8190) <= a or b;
    layer7_outputs(8191) <= not (a xor b);
    layer7_outputs(8192) <= not (a or b);
    layer7_outputs(8193) <= b;
    layer7_outputs(8194) <= not a;
    layer7_outputs(8195) <= not a or b;
    layer7_outputs(8196) <= not a;
    layer7_outputs(8197) <= a;
    layer7_outputs(8198) <= a;
    layer7_outputs(8199) <= a and b;
    layer7_outputs(8200) <= not b;
    layer7_outputs(8201) <= not (a xor b);
    layer7_outputs(8202) <= a or b;
    layer7_outputs(8203) <= b;
    layer7_outputs(8204) <= a and not b;
    layer7_outputs(8205) <= a;
    layer7_outputs(8206) <= b and not a;
    layer7_outputs(8207) <= not b;
    layer7_outputs(8208) <= a xor b;
    layer7_outputs(8209) <= a xor b;
    layer7_outputs(8210) <= not a;
    layer7_outputs(8211) <= not b or a;
    layer7_outputs(8212) <= not b or a;
    layer7_outputs(8213) <= b;
    layer7_outputs(8214) <= not a;
    layer7_outputs(8215) <= not b or a;
    layer7_outputs(8216) <= a or b;
    layer7_outputs(8217) <= not a;
    layer7_outputs(8218) <= b and not a;
    layer7_outputs(8219) <= a or b;
    layer7_outputs(8220) <= a;
    layer7_outputs(8221) <= a;
    layer7_outputs(8222) <= not (a xor b);
    layer7_outputs(8223) <= a xor b;
    layer7_outputs(8224) <= b and not a;
    layer7_outputs(8225) <= not b;
    layer7_outputs(8226) <= not b;
    layer7_outputs(8227) <= a;
    layer7_outputs(8228) <= not (a xor b);
    layer7_outputs(8229) <= b;
    layer7_outputs(8230) <= not (a xor b);
    layer7_outputs(8231) <= a xor b;
    layer7_outputs(8232) <= not b;
    layer7_outputs(8233) <= not (a xor b);
    layer7_outputs(8234) <= not (a xor b);
    layer7_outputs(8235) <= b;
    layer7_outputs(8236) <= not a;
    layer7_outputs(8237) <= b;
    layer7_outputs(8238) <= b;
    layer7_outputs(8239) <= not b;
    layer7_outputs(8240) <= b;
    layer7_outputs(8241) <= not b or a;
    layer7_outputs(8242) <= a xor b;
    layer7_outputs(8243) <= a xor b;
    layer7_outputs(8244) <= b;
    layer7_outputs(8245) <= b;
    layer7_outputs(8246) <= 1'b1;
    layer7_outputs(8247) <= 1'b1;
    layer7_outputs(8248) <= a;
    layer7_outputs(8249) <= not (a xor b);
    layer7_outputs(8250) <= b;
    layer7_outputs(8251) <= not (a xor b);
    layer7_outputs(8252) <= not (a xor b);
    layer7_outputs(8253) <= b and not a;
    layer7_outputs(8254) <= b;
    layer7_outputs(8255) <= not b;
    layer7_outputs(8256) <= not b;
    layer7_outputs(8257) <= not (a xor b);
    layer7_outputs(8258) <= not (a and b);
    layer7_outputs(8259) <= b;
    layer7_outputs(8260) <= not a or b;
    layer7_outputs(8261) <= not a;
    layer7_outputs(8262) <= b;
    layer7_outputs(8263) <= a;
    layer7_outputs(8264) <= not (a xor b);
    layer7_outputs(8265) <= not (a and b);
    layer7_outputs(8266) <= not (a or b);
    layer7_outputs(8267) <= a and b;
    layer7_outputs(8268) <= not (a and b);
    layer7_outputs(8269) <= a;
    layer7_outputs(8270) <= not a;
    layer7_outputs(8271) <= a;
    layer7_outputs(8272) <= a xor b;
    layer7_outputs(8273) <= a xor b;
    layer7_outputs(8274) <= not (a xor b);
    layer7_outputs(8275) <= 1'b0;
    layer7_outputs(8276) <= not b;
    layer7_outputs(8277) <= a;
    layer7_outputs(8278) <= not (a xor b);
    layer7_outputs(8279) <= a;
    layer7_outputs(8280) <= b;
    layer7_outputs(8281) <= b and not a;
    layer7_outputs(8282) <= b;
    layer7_outputs(8283) <= not b;
    layer7_outputs(8284) <= not (a or b);
    layer7_outputs(8285) <= b;
    layer7_outputs(8286) <= not a or b;
    layer7_outputs(8287) <= not (a and b);
    layer7_outputs(8288) <= a and b;
    layer7_outputs(8289) <= a;
    layer7_outputs(8290) <= not b or a;
    layer7_outputs(8291) <= not b;
    layer7_outputs(8292) <= not a;
    layer7_outputs(8293) <= a;
    layer7_outputs(8294) <= not a;
    layer7_outputs(8295) <= not a;
    layer7_outputs(8296) <= a or b;
    layer7_outputs(8297) <= 1'b0;
    layer7_outputs(8298) <= not (a and b);
    layer7_outputs(8299) <= not (a and b);
    layer7_outputs(8300) <= b;
    layer7_outputs(8301) <= not (a xor b);
    layer7_outputs(8302) <= a and not b;
    layer7_outputs(8303) <= b;
    layer7_outputs(8304) <= a xor b;
    layer7_outputs(8305) <= a;
    layer7_outputs(8306) <= not b;
    layer7_outputs(8307) <= not (a xor b);
    layer7_outputs(8308) <= not a;
    layer7_outputs(8309) <= a xor b;
    layer7_outputs(8310) <= a and b;
    layer7_outputs(8311) <= not b;
    layer7_outputs(8312) <= a;
    layer7_outputs(8313) <= a xor b;
    layer7_outputs(8314) <= a;
    layer7_outputs(8315) <= not a or b;
    layer7_outputs(8316) <= b;
    layer7_outputs(8317) <= not a;
    layer7_outputs(8318) <= not a;
    layer7_outputs(8319) <= not b;
    layer7_outputs(8320) <= a and not b;
    layer7_outputs(8321) <= a and not b;
    layer7_outputs(8322) <= b;
    layer7_outputs(8323) <= a xor b;
    layer7_outputs(8324) <= a and b;
    layer7_outputs(8325) <= not b or a;
    layer7_outputs(8326) <= b;
    layer7_outputs(8327) <= not (a and b);
    layer7_outputs(8328) <= a xor b;
    layer7_outputs(8329) <= not b;
    layer7_outputs(8330) <= not (a xor b);
    layer7_outputs(8331) <= not a or b;
    layer7_outputs(8332) <= b and not a;
    layer7_outputs(8333) <= not (a and b);
    layer7_outputs(8334) <= not (a and b);
    layer7_outputs(8335) <= not b;
    layer7_outputs(8336) <= not b;
    layer7_outputs(8337) <= not (a or b);
    layer7_outputs(8338) <= a;
    layer7_outputs(8339) <= not a;
    layer7_outputs(8340) <= not a;
    layer7_outputs(8341) <= not b or a;
    layer7_outputs(8342) <= not a;
    layer7_outputs(8343) <= a or b;
    layer7_outputs(8344) <= b and not a;
    layer7_outputs(8345) <= a;
    layer7_outputs(8346) <= not a;
    layer7_outputs(8347) <= a and not b;
    layer7_outputs(8348) <= not b;
    layer7_outputs(8349) <= not b;
    layer7_outputs(8350) <= not (a xor b);
    layer7_outputs(8351) <= a xor b;
    layer7_outputs(8352) <= not a;
    layer7_outputs(8353) <= b and not a;
    layer7_outputs(8354) <= a;
    layer7_outputs(8355) <= not b;
    layer7_outputs(8356) <= b;
    layer7_outputs(8357) <= not (a or b);
    layer7_outputs(8358) <= not a or b;
    layer7_outputs(8359) <= not b or a;
    layer7_outputs(8360) <= not a;
    layer7_outputs(8361) <= a;
    layer7_outputs(8362) <= a;
    layer7_outputs(8363) <= a;
    layer7_outputs(8364) <= a and not b;
    layer7_outputs(8365) <= a or b;
    layer7_outputs(8366) <= not (a and b);
    layer7_outputs(8367) <= b;
    layer7_outputs(8368) <= not b;
    layer7_outputs(8369) <= a;
    layer7_outputs(8370) <= 1'b0;
    layer7_outputs(8371) <= a xor b;
    layer7_outputs(8372) <= a;
    layer7_outputs(8373) <= a xor b;
    layer7_outputs(8374) <= not a;
    layer7_outputs(8375) <= b;
    layer7_outputs(8376) <= a;
    layer7_outputs(8377) <= b and not a;
    layer7_outputs(8378) <= not (a xor b);
    layer7_outputs(8379) <= not (a and b);
    layer7_outputs(8380) <= not b;
    layer7_outputs(8381) <= not b;
    layer7_outputs(8382) <= b and not a;
    layer7_outputs(8383) <= not b;
    layer7_outputs(8384) <= b and not a;
    layer7_outputs(8385) <= b;
    layer7_outputs(8386) <= a and b;
    layer7_outputs(8387) <= not b or a;
    layer7_outputs(8388) <= a and not b;
    layer7_outputs(8389) <= not a;
    layer7_outputs(8390) <= b and not a;
    layer7_outputs(8391) <= not a or b;
    layer7_outputs(8392) <= not (a or b);
    layer7_outputs(8393) <= not (a and b);
    layer7_outputs(8394) <= not a;
    layer7_outputs(8395) <= b and not a;
    layer7_outputs(8396) <= a and not b;
    layer7_outputs(8397) <= a and not b;
    layer7_outputs(8398) <= 1'b1;
    layer7_outputs(8399) <= b and not a;
    layer7_outputs(8400) <= not b;
    layer7_outputs(8401) <= not (a and b);
    layer7_outputs(8402) <= not b;
    layer7_outputs(8403) <= b;
    layer7_outputs(8404) <= not b;
    layer7_outputs(8405) <= not a;
    layer7_outputs(8406) <= b;
    layer7_outputs(8407) <= 1'b0;
    layer7_outputs(8408) <= a;
    layer7_outputs(8409) <= not (a or b);
    layer7_outputs(8410) <= not a;
    layer7_outputs(8411) <= b and not a;
    layer7_outputs(8412) <= not b or a;
    layer7_outputs(8413) <= not (a xor b);
    layer7_outputs(8414) <= b;
    layer7_outputs(8415) <= not (a or b);
    layer7_outputs(8416) <= not (a xor b);
    layer7_outputs(8417) <= b;
    layer7_outputs(8418) <= not a;
    layer7_outputs(8419) <= not a;
    layer7_outputs(8420) <= b;
    layer7_outputs(8421) <= a and not b;
    layer7_outputs(8422) <= not b;
    layer7_outputs(8423) <= b;
    layer7_outputs(8424) <= not a;
    layer7_outputs(8425) <= a xor b;
    layer7_outputs(8426) <= not (a xor b);
    layer7_outputs(8427) <= not (a xor b);
    layer7_outputs(8428) <= a;
    layer7_outputs(8429) <= not (a or b);
    layer7_outputs(8430) <= b;
    layer7_outputs(8431) <= a xor b;
    layer7_outputs(8432) <= a;
    layer7_outputs(8433) <= a and b;
    layer7_outputs(8434) <= a and not b;
    layer7_outputs(8435) <= not a;
    layer7_outputs(8436) <= not a;
    layer7_outputs(8437) <= a and b;
    layer7_outputs(8438) <= not a;
    layer7_outputs(8439) <= not b;
    layer7_outputs(8440) <= not b;
    layer7_outputs(8441) <= not (a or b);
    layer7_outputs(8442) <= 1'b1;
    layer7_outputs(8443) <= not (a xor b);
    layer7_outputs(8444) <= 1'b1;
    layer7_outputs(8445) <= 1'b1;
    layer7_outputs(8446) <= b;
    layer7_outputs(8447) <= b and not a;
    layer7_outputs(8448) <= not b;
    layer7_outputs(8449) <= a or b;
    layer7_outputs(8450) <= not b;
    layer7_outputs(8451) <= not (a xor b);
    layer7_outputs(8452) <= b;
    layer7_outputs(8453) <= a or b;
    layer7_outputs(8454) <= not (a xor b);
    layer7_outputs(8455) <= not b;
    layer7_outputs(8456) <= not (a xor b);
    layer7_outputs(8457) <= not b;
    layer7_outputs(8458) <= not a;
    layer7_outputs(8459) <= a;
    layer7_outputs(8460) <= not a;
    layer7_outputs(8461) <= b;
    layer7_outputs(8462) <= b and not a;
    layer7_outputs(8463) <= a or b;
    layer7_outputs(8464) <= a;
    layer7_outputs(8465) <= not a;
    layer7_outputs(8466) <= not (a or b);
    layer7_outputs(8467) <= not b;
    layer7_outputs(8468) <= a and b;
    layer7_outputs(8469) <= a xor b;
    layer7_outputs(8470) <= a;
    layer7_outputs(8471) <= a or b;
    layer7_outputs(8472) <= not (a xor b);
    layer7_outputs(8473) <= b and not a;
    layer7_outputs(8474) <= not a;
    layer7_outputs(8475) <= a and not b;
    layer7_outputs(8476) <= not a;
    layer7_outputs(8477) <= not (a and b);
    layer7_outputs(8478) <= not (a xor b);
    layer7_outputs(8479) <= not a;
    layer7_outputs(8480) <= b;
    layer7_outputs(8481) <= not a;
    layer7_outputs(8482) <= not (a xor b);
    layer7_outputs(8483) <= not (a xor b);
    layer7_outputs(8484) <= not (a xor b);
    layer7_outputs(8485) <= a or b;
    layer7_outputs(8486) <= a xor b;
    layer7_outputs(8487) <= not a;
    layer7_outputs(8488) <= b;
    layer7_outputs(8489) <= not b or a;
    layer7_outputs(8490) <= not a or b;
    layer7_outputs(8491) <= b and not a;
    layer7_outputs(8492) <= a xor b;
    layer7_outputs(8493) <= 1'b1;
    layer7_outputs(8494) <= a or b;
    layer7_outputs(8495) <= a and b;
    layer7_outputs(8496) <= not a or b;
    layer7_outputs(8497) <= not (a xor b);
    layer7_outputs(8498) <= not b or a;
    layer7_outputs(8499) <= not b;
    layer7_outputs(8500) <= not a;
    layer7_outputs(8501) <= a;
    layer7_outputs(8502) <= a xor b;
    layer7_outputs(8503) <= a;
    layer7_outputs(8504) <= not (a and b);
    layer7_outputs(8505) <= not a;
    layer7_outputs(8506) <= not a;
    layer7_outputs(8507) <= not (a and b);
    layer7_outputs(8508) <= not b or a;
    layer7_outputs(8509) <= a;
    layer7_outputs(8510) <= b and not a;
    layer7_outputs(8511) <= a;
    layer7_outputs(8512) <= not (a xor b);
    layer7_outputs(8513) <= not a;
    layer7_outputs(8514) <= not (a or b);
    layer7_outputs(8515) <= not a;
    layer7_outputs(8516) <= not (a or b);
    layer7_outputs(8517) <= not (a xor b);
    layer7_outputs(8518) <= not b;
    layer7_outputs(8519) <= b;
    layer7_outputs(8520) <= not b;
    layer7_outputs(8521) <= not b;
    layer7_outputs(8522) <= not a;
    layer7_outputs(8523) <= b;
    layer7_outputs(8524) <= not a or b;
    layer7_outputs(8525) <= not (a xor b);
    layer7_outputs(8526) <= not (a xor b);
    layer7_outputs(8527) <= not b;
    layer7_outputs(8528) <= not b;
    layer7_outputs(8529) <= not a;
    layer7_outputs(8530) <= a;
    layer7_outputs(8531) <= a and b;
    layer7_outputs(8532) <= a xor b;
    layer7_outputs(8533) <= a and b;
    layer7_outputs(8534) <= a and not b;
    layer7_outputs(8535) <= a xor b;
    layer7_outputs(8536) <= a and b;
    layer7_outputs(8537) <= not b;
    layer7_outputs(8538) <= a;
    layer7_outputs(8539) <= a xor b;
    layer7_outputs(8540) <= not (a or b);
    layer7_outputs(8541) <= not (a or b);
    layer7_outputs(8542) <= not a;
    layer7_outputs(8543) <= not (a and b);
    layer7_outputs(8544) <= a xor b;
    layer7_outputs(8545) <= not (a or b);
    layer7_outputs(8546) <= a;
    layer7_outputs(8547) <= not (a and b);
    layer7_outputs(8548) <= not b or a;
    layer7_outputs(8549) <= b and not a;
    layer7_outputs(8550) <= a and b;
    layer7_outputs(8551) <= not a;
    layer7_outputs(8552) <= not b;
    layer7_outputs(8553) <= not a or b;
    layer7_outputs(8554) <= a and b;
    layer7_outputs(8555) <= not b or a;
    layer7_outputs(8556) <= not a or b;
    layer7_outputs(8557) <= not a;
    layer7_outputs(8558) <= not b;
    layer7_outputs(8559) <= 1'b1;
    layer7_outputs(8560) <= a;
    layer7_outputs(8561) <= b;
    layer7_outputs(8562) <= not b or a;
    layer7_outputs(8563) <= not a;
    layer7_outputs(8564) <= not b or a;
    layer7_outputs(8565) <= a xor b;
    layer7_outputs(8566) <= b;
    layer7_outputs(8567) <= not b or a;
    layer7_outputs(8568) <= not a or b;
    layer7_outputs(8569) <= not a;
    layer7_outputs(8570) <= a xor b;
    layer7_outputs(8571) <= not b;
    layer7_outputs(8572) <= b;
    layer7_outputs(8573) <= b;
    layer7_outputs(8574) <= not (a or b);
    layer7_outputs(8575) <= b;
    layer7_outputs(8576) <= not (a xor b);
    layer7_outputs(8577) <= a or b;
    layer7_outputs(8578) <= not b;
    layer7_outputs(8579) <= not (a or b);
    layer7_outputs(8580) <= not b or a;
    layer7_outputs(8581) <= not (a xor b);
    layer7_outputs(8582) <= a or b;
    layer7_outputs(8583) <= a or b;
    layer7_outputs(8584) <= not b or a;
    layer7_outputs(8585) <= a and not b;
    layer7_outputs(8586) <= not a or b;
    layer7_outputs(8587) <= not b;
    layer7_outputs(8588) <= not (a xor b);
    layer7_outputs(8589) <= b;
    layer7_outputs(8590) <= b and not a;
    layer7_outputs(8591) <= not (a xor b);
    layer7_outputs(8592) <= b;
    layer7_outputs(8593) <= b;
    layer7_outputs(8594) <= a;
    layer7_outputs(8595) <= 1'b1;
    layer7_outputs(8596) <= not b;
    layer7_outputs(8597) <= not a;
    layer7_outputs(8598) <= not (a or b);
    layer7_outputs(8599) <= not (a or b);
    layer7_outputs(8600) <= not a;
    layer7_outputs(8601) <= not a;
    layer7_outputs(8602) <= not b;
    layer7_outputs(8603) <= a xor b;
    layer7_outputs(8604) <= not (a and b);
    layer7_outputs(8605) <= not a;
    layer7_outputs(8606) <= a;
    layer7_outputs(8607) <= not (a and b);
    layer7_outputs(8608) <= b;
    layer7_outputs(8609) <= a or b;
    layer7_outputs(8610) <= not (a xor b);
    layer7_outputs(8611) <= b;
    layer7_outputs(8612) <= a xor b;
    layer7_outputs(8613) <= b;
    layer7_outputs(8614) <= not b;
    layer7_outputs(8615) <= a;
    layer7_outputs(8616) <= not a;
    layer7_outputs(8617) <= not a;
    layer7_outputs(8618) <= not a;
    layer7_outputs(8619) <= not b;
    layer7_outputs(8620) <= not b or a;
    layer7_outputs(8621) <= not a or b;
    layer7_outputs(8622) <= not (a xor b);
    layer7_outputs(8623) <= not (a and b);
    layer7_outputs(8624) <= b and not a;
    layer7_outputs(8625) <= a xor b;
    layer7_outputs(8626) <= not a or b;
    layer7_outputs(8627) <= a xor b;
    layer7_outputs(8628) <= not b;
    layer7_outputs(8629) <= not (a and b);
    layer7_outputs(8630) <= a xor b;
    layer7_outputs(8631) <= not b;
    layer7_outputs(8632) <= not b;
    layer7_outputs(8633) <= b;
    layer7_outputs(8634) <= a xor b;
    layer7_outputs(8635) <= a;
    layer7_outputs(8636) <= b;
    layer7_outputs(8637) <= not b;
    layer7_outputs(8638) <= not (a and b);
    layer7_outputs(8639) <= a and not b;
    layer7_outputs(8640) <= a and b;
    layer7_outputs(8641) <= a or b;
    layer7_outputs(8642) <= a and b;
    layer7_outputs(8643) <= not a;
    layer7_outputs(8644) <= not (a xor b);
    layer7_outputs(8645) <= not (a and b);
    layer7_outputs(8646) <= b;
    layer7_outputs(8647) <= not b or a;
    layer7_outputs(8648) <= a or b;
    layer7_outputs(8649) <= a and b;
    layer7_outputs(8650) <= b and not a;
    layer7_outputs(8651) <= b;
    layer7_outputs(8652) <= not (a xor b);
    layer7_outputs(8653) <= b;
    layer7_outputs(8654) <= 1'b0;
    layer7_outputs(8655) <= not b;
    layer7_outputs(8656) <= not a;
    layer7_outputs(8657) <= a xor b;
    layer7_outputs(8658) <= not b;
    layer7_outputs(8659) <= a;
    layer7_outputs(8660) <= not a;
    layer7_outputs(8661) <= b;
    layer7_outputs(8662) <= not b;
    layer7_outputs(8663) <= not b;
    layer7_outputs(8664) <= b;
    layer7_outputs(8665) <= b;
    layer7_outputs(8666) <= not (a or b);
    layer7_outputs(8667) <= not b;
    layer7_outputs(8668) <= a and b;
    layer7_outputs(8669) <= not a;
    layer7_outputs(8670) <= b and not a;
    layer7_outputs(8671) <= not a;
    layer7_outputs(8672) <= a;
    layer7_outputs(8673) <= not b;
    layer7_outputs(8674) <= a;
    layer7_outputs(8675) <= a or b;
    layer7_outputs(8676) <= b;
    layer7_outputs(8677) <= not (a xor b);
    layer7_outputs(8678) <= not b;
    layer7_outputs(8679) <= not b or a;
    layer7_outputs(8680) <= b and not a;
    layer7_outputs(8681) <= not a;
    layer7_outputs(8682) <= not a or b;
    layer7_outputs(8683) <= b and not a;
    layer7_outputs(8684) <= a or b;
    layer7_outputs(8685) <= a;
    layer7_outputs(8686) <= not a or b;
    layer7_outputs(8687) <= not a or b;
    layer7_outputs(8688) <= a or b;
    layer7_outputs(8689) <= b;
    layer7_outputs(8690) <= a or b;
    layer7_outputs(8691) <= 1'b0;
    layer7_outputs(8692) <= a or b;
    layer7_outputs(8693) <= not a;
    layer7_outputs(8694) <= not (a xor b);
    layer7_outputs(8695) <= not a or b;
    layer7_outputs(8696) <= b;
    layer7_outputs(8697) <= not a or b;
    layer7_outputs(8698) <= not a or b;
    layer7_outputs(8699) <= b;
    layer7_outputs(8700) <= not b;
    layer7_outputs(8701) <= a;
    layer7_outputs(8702) <= not b or a;
    layer7_outputs(8703) <= a;
    layer7_outputs(8704) <= not a or b;
    layer7_outputs(8705) <= a xor b;
    layer7_outputs(8706) <= not a or b;
    layer7_outputs(8707) <= not (a and b);
    layer7_outputs(8708) <= a xor b;
    layer7_outputs(8709) <= b;
    layer7_outputs(8710) <= not b or a;
    layer7_outputs(8711) <= not (a or b);
    layer7_outputs(8712) <= not b;
    layer7_outputs(8713) <= a and b;
    layer7_outputs(8714) <= not b;
    layer7_outputs(8715) <= not (a and b);
    layer7_outputs(8716) <= not (a xor b);
    layer7_outputs(8717) <= not (a xor b);
    layer7_outputs(8718) <= a xor b;
    layer7_outputs(8719) <= not b;
    layer7_outputs(8720) <= not (a or b);
    layer7_outputs(8721) <= not (a and b);
    layer7_outputs(8722) <= not b or a;
    layer7_outputs(8723) <= not a;
    layer7_outputs(8724) <= not b or a;
    layer7_outputs(8725) <= not (a xor b);
    layer7_outputs(8726) <= a xor b;
    layer7_outputs(8727) <= a or b;
    layer7_outputs(8728) <= a;
    layer7_outputs(8729) <= not (a xor b);
    layer7_outputs(8730) <= a and not b;
    layer7_outputs(8731) <= b;
    layer7_outputs(8732) <= not (a or b);
    layer7_outputs(8733) <= a;
    layer7_outputs(8734) <= not a;
    layer7_outputs(8735) <= not a or b;
    layer7_outputs(8736) <= not (a xor b);
    layer7_outputs(8737) <= b;
    layer7_outputs(8738) <= not b;
    layer7_outputs(8739) <= not (a or b);
    layer7_outputs(8740) <= b;
    layer7_outputs(8741) <= a;
    layer7_outputs(8742) <= not b;
    layer7_outputs(8743) <= b;
    layer7_outputs(8744) <= not (a or b);
    layer7_outputs(8745) <= a and b;
    layer7_outputs(8746) <= a and b;
    layer7_outputs(8747) <= not (a and b);
    layer7_outputs(8748) <= a and b;
    layer7_outputs(8749) <= b;
    layer7_outputs(8750) <= a and not b;
    layer7_outputs(8751) <= not a;
    layer7_outputs(8752) <= b;
    layer7_outputs(8753) <= b;
    layer7_outputs(8754) <= a;
    layer7_outputs(8755) <= not (a xor b);
    layer7_outputs(8756) <= not (a and b);
    layer7_outputs(8757) <= not (a and b);
    layer7_outputs(8758) <= a or b;
    layer7_outputs(8759) <= a xor b;
    layer7_outputs(8760) <= a;
    layer7_outputs(8761) <= a;
    layer7_outputs(8762) <= b;
    layer7_outputs(8763) <= not (a and b);
    layer7_outputs(8764) <= a;
    layer7_outputs(8765) <= a;
    layer7_outputs(8766) <= a;
    layer7_outputs(8767) <= b and not a;
    layer7_outputs(8768) <= not a;
    layer7_outputs(8769) <= not (a or b);
    layer7_outputs(8770) <= b and not a;
    layer7_outputs(8771) <= a xor b;
    layer7_outputs(8772) <= a;
    layer7_outputs(8773) <= not b or a;
    layer7_outputs(8774) <= a xor b;
    layer7_outputs(8775) <= not (a and b);
    layer7_outputs(8776) <= a;
    layer7_outputs(8777) <= b;
    layer7_outputs(8778) <= not b;
    layer7_outputs(8779) <= not (a and b);
    layer7_outputs(8780) <= not (a and b);
    layer7_outputs(8781) <= not (a or b);
    layer7_outputs(8782) <= a;
    layer7_outputs(8783) <= a;
    layer7_outputs(8784) <= b;
    layer7_outputs(8785) <= not (a xor b);
    layer7_outputs(8786) <= not b or a;
    layer7_outputs(8787) <= 1'b0;
    layer7_outputs(8788) <= a;
    layer7_outputs(8789) <= a xor b;
    layer7_outputs(8790) <= not a or b;
    layer7_outputs(8791) <= not b;
    layer7_outputs(8792) <= a;
    layer7_outputs(8793) <= b;
    layer7_outputs(8794) <= not b or a;
    layer7_outputs(8795) <= 1'b1;
    layer7_outputs(8796) <= not a;
    layer7_outputs(8797) <= not (a xor b);
    layer7_outputs(8798) <= b and not a;
    layer7_outputs(8799) <= not (a or b);
    layer7_outputs(8800) <= a and not b;
    layer7_outputs(8801) <= b and not a;
    layer7_outputs(8802) <= not a;
    layer7_outputs(8803) <= not a;
    layer7_outputs(8804) <= not a;
    layer7_outputs(8805) <= not a;
    layer7_outputs(8806) <= b;
    layer7_outputs(8807) <= a;
    layer7_outputs(8808) <= not b or a;
    layer7_outputs(8809) <= b;
    layer7_outputs(8810) <= not (a and b);
    layer7_outputs(8811) <= not b;
    layer7_outputs(8812) <= not b;
    layer7_outputs(8813) <= not a;
    layer7_outputs(8814) <= not b or a;
    layer7_outputs(8815) <= a xor b;
    layer7_outputs(8816) <= a;
    layer7_outputs(8817) <= not b;
    layer7_outputs(8818) <= not b or a;
    layer7_outputs(8819) <= not (a and b);
    layer7_outputs(8820) <= not (a or b);
    layer7_outputs(8821) <= not b or a;
    layer7_outputs(8822) <= not b;
    layer7_outputs(8823) <= not b;
    layer7_outputs(8824) <= b and not a;
    layer7_outputs(8825) <= a;
    layer7_outputs(8826) <= not (a xor b);
    layer7_outputs(8827) <= not b;
    layer7_outputs(8828) <= a xor b;
    layer7_outputs(8829) <= not b;
    layer7_outputs(8830) <= a xor b;
    layer7_outputs(8831) <= not a;
    layer7_outputs(8832) <= a or b;
    layer7_outputs(8833) <= a or b;
    layer7_outputs(8834) <= not b or a;
    layer7_outputs(8835) <= a xor b;
    layer7_outputs(8836) <= not a or b;
    layer7_outputs(8837) <= not (a and b);
    layer7_outputs(8838) <= not b or a;
    layer7_outputs(8839) <= b and not a;
    layer7_outputs(8840) <= not b or a;
    layer7_outputs(8841) <= b and not a;
    layer7_outputs(8842) <= a and b;
    layer7_outputs(8843) <= not b;
    layer7_outputs(8844) <= not (a xor b);
    layer7_outputs(8845) <= not b;
    layer7_outputs(8846) <= a and not b;
    layer7_outputs(8847) <= not a;
    layer7_outputs(8848) <= not b or a;
    layer7_outputs(8849) <= not (a and b);
    layer7_outputs(8850) <= a xor b;
    layer7_outputs(8851) <= b and not a;
    layer7_outputs(8852) <= a xor b;
    layer7_outputs(8853) <= a;
    layer7_outputs(8854) <= b;
    layer7_outputs(8855) <= a;
    layer7_outputs(8856) <= not a;
    layer7_outputs(8857) <= a and b;
    layer7_outputs(8858) <= 1'b0;
    layer7_outputs(8859) <= b;
    layer7_outputs(8860) <= not (a and b);
    layer7_outputs(8861) <= a xor b;
    layer7_outputs(8862) <= not a;
    layer7_outputs(8863) <= a;
    layer7_outputs(8864) <= a;
    layer7_outputs(8865) <= a;
    layer7_outputs(8866) <= not a;
    layer7_outputs(8867) <= a;
    layer7_outputs(8868) <= b;
    layer7_outputs(8869) <= a;
    layer7_outputs(8870) <= b and not a;
    layer7_outputs(8871) <= not (a or b);
    layer7_outputs(8872) <= not a or b;
    layer7_outputs(8873) <= not (a xor b);
    layer7_outputs(8874) <= a;
    layer7_outputs(8875) <= not b or a;
    layer7_outputs(8876) <= a and not b;
    layer7_outputs(8877) <= not b or a;
    layer7_outputs(8878) <= not b;
    layer7_outputs(8879) <= b;
    layer7_outputs(8880) <= b;
    layer7_outputs(8881) <= a;
    layer7_outputs(8882) <= not b;
    layer7_outputs(8883) <= a and not b;
    layer7_outputs(8884) <= b;
    layer7_outputs(8885) <= not (a or b);
    layer7_outputs(8886) <= not (a or b);
    layer7_outputs(8887) <= not (a or b);
    layer7_outputs(8888) <= a;
    layer7_outputs(8889) <= a and b;
    layer7_outputs(8890) <= a;
    layer7_outputs(8891) <= not a;
    layer7_outputs(8892) <= a;
    layer7_outputs(8893) <= not b;
    layer7_outputs(8894) <= not a;
    layer7_outputs(8895) <= a or b;
    layer7_outputs(8896) <= not (a xor b);
    layer7_outputs(8897) <= b;
    layer7_outputs(8898) <= a and b;
    layer7_outputs(8899) <= a or b;
    layer7_outputs(8900) <= not (a xor b);
    layer7_outputs(8901) <= b;
    layer7_outputs(8902) <= not b;
    layer7_outputs(8903) <= a or b;
    layer7_outputs(8904) <= b and not a;
    layer7_outputs(8905) <= a or b;
    layer7_outputs(8906) <= a and not b;
    layer7_outputs(8907) <= not (a xor b);
    layer7_outputs(8908) <= not b;
    layer7_outputs(8909) <= not a;
    layer7_outputs(8910) <= not a;
    layer7_outputs(8911) <= a and b;
    layer7_outputs(8912) <= a;
    layer7_outputs(8913) <= not b or a;
    layer7_outputs(8914) <= a;
    layer7_outputs(8915) <= a xor b;
    layer7_outputs(8916) <= a;
    layer7_outputs(8917) <= not (a and b);
    layer7_outputs(8918) <= not a;
    layer7_outputs(8919) <= a;
    layer7_outputs(8920) <= not (a xor b);
    layer7_outputs(8921) <= a;
    layer7_outputs(8922) <= not a;
    layer7_outputs(8923) <= not (a and b);
    layer7_outputs(8924) <= not (a and b);
    layer7_outputs(8925) <= not (a and b);
    layer7_outputs(8926) <= a and not b;
    layer7_outputs(8927) <= not (a xor b);
    layer7_outputs(8928) <= not b;
    layer7_outputs(8929) <= a xor b;
    layer7_outputs(8930) <= not (a or b);
    layer7_outputs(8931) <= b;
    layer7_outputs(8932) <= a;
    layer7_outputs(8933) <= not a;
    layer7_outputs(8934) <= a or b;
    layer7_outputs(8935) <= a and b;
    layer7_outputs(8936) <= b;
    layer7_outputs(8937) <= a and b;
    layer7_outputs(8938) <= a and not b;
    layer7_outputs(8939) <= not b;
    layer7_outputs(8940) <= a and not b;
    layer7_outputs(8941) <= not (a and b);
    layer7_outputs(8942) <= not (a xor b);
    layer7_outputs(8943) <= not a;
    layer7_outputs(8944) <= b;
    layer7_outputs(8945) <= not a;
    layer7_outputs(8946) <= a and not b;
    layer7_outputs(8947) <= a;
    layer7_outputs(8948) <= a;
    layer7_outputs(8949) <= not b;
    layer7_outputs(8950) <= b;
    layer7_outputs(8951) <= not (a xor b);
    layer7_outputs(8952) <= not a or b;
    layer7_outputs(8953) <= not b;
    layer7_outputs(8954) <= a and b;
    layer7_outputs(8955) <= not (a xor b);
    layer7_outputs(8956) <= not b;
    layer7_outputs(8957) <= b and not a;
    layer7_outputs(8958) <= a;
    layer7_outputs(8959) <= b;
    layer7_outputs(8960) <= a and not b;
    layer7_outputs(8961) <= not (a and b);
    layer7_outputs(8962) <= a and not b;
    layer7_outputs(8963) <= not a;
    layer7_outputs(8964) <= not (a xor b);
    layer7_outputs(8965) <= a;
    layer7_outputs(8966) <= not (a xor b);
    layer7_outputs(8967) <= a and b;
    layer7_outputs(8968) <= a and not b;
    layer7_outputs(8969) <= b and not a;
    layer7_outputs(8970) <= b;
    layer7_outputs(8971) <= not (a xor b);
    layer7_outputs(8972) <= a;
    layer7_outputs(8973) <= a;
    layer7_outputs(8974) <= not a;
    layer7_outputs(8975) <= not b or a;
    layer7_outputs(8976) <= not a;
    layer7_outputs(8977) <= a;
    layer7_outputs(8978) <= not (a xor b);
    layer7_outputs(8979) <= a;
    layer7_outputs(8980) <= a;
    layer7_outputs(8981) <= not (a or b);
    layer7_outputs(8982) <= not (a xor b);
    layer7_outputs(8983) <= not (a xor b);
    layer7_outputs(8984) <= a and b;
    layer7_outputs(8985) <= not (a xor b);
    layer7_outputs(8986) <= not (a or b);
    layer7_outputs(8987) <= not (a or b);
    layer7_outputs(8988) <= b and not a;
    layer7_outputs(8989) <= not b or a;
    layer7_outputs(8990) <= not a or b;
    layer7_outputs(8991) <= a;
    layer7_outputs(8992) <= not (a xor b);
    layer7_outputs(8993) <= a;
    layer7_outputs(8994) <= not a or b;
    layer7_outputs(8995) <= a xor b;
    layer7_outputs(8996) <= a xor b;
    layer7_outputs(8997) <= a xor b;
    layer7_outputs(8998) <= not (a or b);
    layer7_outputs(8999) <= a or b;
    layer7_outputs(9000) <= a and not b;
    layer7_outputs(9001) <= a or b;
    layer7_outputs(9002) <= a or b;
    layer7_outputs(9003) <= not b;
    layer7_outputs(9004) <= b;
    layer7_outputs(9005) <= not a or b;
    layer7_outputs(9006) <= a;
    layer7_outputs(9007) <= a;
    layer7_outputs(9008) <= a xor b;
    layer7_outputs(9009) <= a xor b;
    layer7_outputs(9010) <= not b or a;
    layer7_outputs(9011) <= b;
    layer7_outputs(9012) <= not (a and b);
    layer7_outputs(9013) <= not (a and b);
    layer7_outputs(9014) <= a or b;
    layer7_outputs(9015) <= b;
    layer7_outputs(9016) <= b;
    layer7_outputs(9017) <= not b;
    layer7_outputs(9018) <= 1'b1;
    layer7_outputs(9019) <= not (a or b);
    layer7_outputs(9020) <= not (a and b);
    layer7_outputs(9021) <= not b;
    layer7_outputs(9022) <= not (a or b);
    layer7_outputs(9023) <= not (a xor b);
    layer7_outputs(9024) <= b and not a;
    layer7_outputs(9025) <= a xor b;
    layer7_outputs(9026) <= not b or a;
    layer7_outputs(9027) <= not a;
    layer7_outputs(9028) <= not a or b;
    layer7_outputs(9029) <= a and b;
    layer7_outputs(9030) <= a xor b;
    layer7_outputs(9031) <= not (a or b);
    layer7_outputs(9032) <= not b or a;
    layer7_outputs(9033) <= a xor b;
    layer7_outputs(9034) <= b and not a;
    layer7_outputs(9035) <= a;
    layer7_outputs(9036) <= a;
    layer7_outputs(9037) <= not (a xor b);
    layer7_outputs(9038) <= not (a xor b);
    layer7_outputs(9039) <= a and not b;
    layer7_outputs(9040) <= b;
    layer7_outputs(9041) <= not (a xor b);
    layer7_outputs(9042) <= not (a and b);
    layer7_outputs(9043) <= a;
    layer7_outputs(9044) <= a;
    layer7_outputs(9045) <= a xor b;
    layer7_outputs(9046) <= not a;
    layer7_outputs(9047) <= not (a xor b);
    layer7_outputs(9048) <= not a or b;
    layer7_outputs(9049) <= a xor b;
    layer7_outputs(9050) <= a and not b;
    layer7_outputs(9051) <= a;
    layer7_outputs(9052) <= b and not a;
    layer7_outputs(9053) <= not a or b;
    layer7_outputs(9054) <= a and not b;
    layer7_outputs(9055) <= not (a xor b);
    layer7_outputs(9056) <= b;
    layer7_outputs(9057) <= not a;
    layer7_outputs(9058) <= a and b;
    layer7_outputs(9059) <= not (a and b);
    layer7_outputs(9060) <= 1'b0;
    layer7_outputs(9061) <= not b;
    layer7_outputs(9062) <= 1'b0;
    layer7_outputs(9063) <= a or b;
    layer7_outputs(9064) <= not b;
    layer7_outputs(9065) <= not (a xor b);
    layer7_outputs(9066) <= not a;
    layer7_outputs(9067) <= a;
    layer7_outputs(9068) <= b and not a;
    layer7_outputs(9069) <= a;
    layer7_outputs(9070) <= b;
    layer7_outputs(9071) <= a xor b;
    layer7_outputs(9072) <= not b;
    layer7_outputs(9073) <= not (a xor b);
    layer7_outputs(9074) <= not b;
    layer7_outputs(9075) <= not (a xor b);
    layer7_outputs(9076) <= b;
    layer7_outputs(9077) <= not b;
    layer7_outputs(9078) <= not b;
    layer7_outputs(9079) <= a;
    layer7_outputs(9080) <= not b or a;
    layer7_outputs(9081) <= not b or a;
    layer7_outputs(9082) <= not a;
    layer7_outputs(9083) <= a and b;
    layer7_outputs(9084) <= not a;
    layer7_outputs(9085) <= 1'b1;
    layer7_outputs(9086) <= not a;
    layer7_outputs(9087) <= a;
    layer7_outputs(9088) <= b;
    layer7_outputs(9089) <= a and b;
    layer7_outputs(9090) <= not b;
    layer7_outputs(9091) <= not a;
    layer7_outputs(9092) <= not (a and b);
    layer7_outputs(9093) <= not b;
    layer7_outputs(9094) <= a;
    layer7_outputs(9095) <= b;
    layer7_outputs(9096) <= 1'b1;
    layer7_outputs(9097) <= b;
    layer7_outputs(9098) <= not a;
    layer7_outputs(9099) <= not (a or b);
    layer7_outputs(9100) <= a and b;
    layer7_outputs(9101) <= a;
    layer7_outputs(9102) <= a;
    layer7_outputs(9103) <= not b;
    layer7_outputs(9104) <= not b;
    layer7_outputs(9105) <= a and not b;
    layer7_outputs(9106) <= a;
    layer7_outputs(9107) <= a;
    layer7_outputs(9108) <= not a;
    layer7_outputs(9109) <= not (a and b);
    layer7_outputs(9110) <= not a;
    layer7_outputs(9111) <= a or b;
    layer7_outputs(9112) <= not (a xor b);
    layer7_outputs(9113) <= not b;
    layer7_outputs(9114) <= a;
    layer7_outputs(9115) <= a;
    layer7_outputs(9116) <= not a or b;
    layer7_outputs(9117) <= not (a and b);
    layer7_outputs(9118) <= a and b;
    layer7_outputs(9119) <= not (a xor b);
    layer7_outputs(9120) <= a and b;
    layer7_outputs(9121) <= not a;
    layer7_outputs(9122) <= not a or b;
    layer7_outputs(9123) <= not (a xor b);
    layer7_outputs(9124) <= a xor b;
    layer7_outputs(9125) <= 1'b0;
    layer7_outputs(9126) <= a and not b;
    layer7_outputs(9127) <= not a;
    layer7_outputs(9128) <= not a;
    layer7_outputs(9129) <= a or b;
    layer7_outputs(9130) <= not a;
    layer7_outputs(9131) <= not b;
    layer7_outputs(9132) <= a and not b;
    layer7_outputs(9133) <= not (a and b);
    layer7_outputs(9134) <= a xor b;
    layer7_outputs(9135) <= a or b;
    layer7_outputs(9136) <= a or b;
    layer7_outputs(9137) <= not b;
    layer7_outputs(9138) <= not b or a;
    layer7_outputs(9139) <= a;
    layer7_outputs(9140) <= b;
    layer7_outputs(9141) <= not (a xor b);
    layer7_outputs(9142) <= a or b;
    layer7_outputs(9143) <= a;
    layer7_outputs(9144) <= not a;
    layer7_outputs(9145) <= a or b;
    layer7_outputs(9146) <= not a;
    layer7_outputs(9147) <= a or b;
    layer7_outputs(9148) <= not a;
    layer7_outputs(9149) <= b;
    layer7_outputs(9150) <= a xor b;
    layer7_outputs(9151) <= not (a and b);
    layer7_outputs(9152) <= not (a and b);
    layer7_outputs(9153) <= a;
    layer7_outputs(9154) <= not b or a;
    layer7_outputs(9155) <= a;
    layer7_outputs(9156) <= b and not a;
    layer7_outputs(9157) <= b;
    layer7_outputs(9158) <= not a or b;
    layer7_outputs(9159) <= 1'b1;
    layer7_outputs(9160) <= a or b;
    layer7_outputs(9161) <= not (a or b);
    layer7_outputs(9162) <= a xor b;
    layer7_outputs(9163) <= a and not b;
    layer7_outputs(9164) <= not (a xor b);
    layer7_outputs(9165) <= not b or a;
    layer7_outputs(9166) <= not b;
    layer7_outputs(9167) <= a;
    layer7_outputs(9168) <= b;
    layer7_outputs(9169) <= a;
    layer7_outputs(9170) <= a;
    layer7_outputs(9171) <= 1'b0;
    layer7_outputs(9172) <= b;
    layer7_outputs(9173) <= not (a xor b);
    layer7_outputs(9174) <= not b;
    layer7_outputs(9175) <= a or b;
    layer7_outputs(9176) <= not b;
    layer7_outputs(9177) <= not b or a;
    layer7_outputs(9178) <= not a or b;
    layer7_outputs(9179) <= not (a xor b);
    layer7_outputs(9180) <= a and b;
    layer7_outputs(9181) <= not b or a;
    layer7_outputs(9182) <= not b;
    layer7_outputs(9183) <= a;
    layer7_outputs(9184) <= a or b;
    layer7_outputs(9185) <= not a;
    layer7_outputs(9186) <= not b or a;
    layer7_outputs(9187) <= a;
    layer7_outputs(9188) <= not (a and b);
    layer7_outputs(9189) <= a xor b;
    layer7_outputs(9190) <= not a or b;
    layer7_outputs(9191) <= not a or b;
    layer7_outputs(9192) <= a or b;
    layer7_outputs(9193) <= not (a xor b);
    layer7_outputs(9194) <= a and not b;
    layer7_outputs(9195) <= not a or b;
    layer7_outputs(9196) <= 1'b1;
    layer7_outputs(9197) <= not (a or b);
    layer7_outputs(9198) <= not a or b;
    layer7_outputs(9199) <= not (a xor b);
    layer7_outputs(9200) <= not b or a;
    layer7_outputs(9201) <= not a;
    layer7_outputs(9202) <= not (a xor b);
    layer7_outputs(9203) <= a and not b;
    layer7_outputs(9204) <= b;
    layer7_outputs(9205) <= not (a xor b);
    layer7_outputs(9206) <= not b;
    layer7_outputs(9207) <= b;
    layer7_outputs(9208) <= not a or b;
    layer7_outputs(9209) <= a and b;
    layer7_outputs(9210) <= not (a and b);
    layer7_outputs(9211) <= a and not b;
    layer7_outputs(9212) <= b;
    layer7_outputs(9213) <= not b;
    layer7_outputs(9214) <= not (a and b);
    layer7_outputs(9215) <= not (a xor b);
    layer7_outputs(9216) <= a xor b;
    layer7_outputs(9217) <= b;
    layer7_outputs(9218) <= not b;
    layer7_outputs(9219) <= not b;
    layer7_outputs(9220) <= not (a xor b);
    layer7_outputs(9221) <= not a;
    layer7_outputs(9222) <= a and not b;
    layer7_outputs(9223) <= not b;
    layer7_outputs(9224) <= a or b;
    layer7_outputs(9225) <= a and not b;
    layer7_outputs(9226) <= not b;
    layer7_outputs(9227) <= not a or b;
    layer7_outputs(9228) <= not (a xor b);
    layer7_outputs(9229) <= not a;
    layer7_outputs(9230) <= a xor b;
    layer7_outputs(9231) <= not a;
    layer7_outputs(9232) <= a xor b;
    layer7_outputs(9233) <= b and not a;
    layer7_outputs(9234) <= not a;
    layer7_outputs(9235) <= not a;
    layer7_outputs(9236) <= b;
    layer7_outputs(9237) <= a and not b;
    layer7_outputs(9238) <= a;
    layer7_outputs(9239) <= not a;
    layer7_outputs(9240) <= not b;
    layer7_outputs(9241) <= a xor b;
    layer7_outputs(9242) <= b;
    layer7_outputs(9243) <= not b;
    layer7_outputs(9244) <= not b or a;
    layer7_outputs(9245) <= b;
    layer7_outputs(9246) <= not (a and b);
    layer7_outputs(9247) <= a xor b;
    layer7_outputs(9248) <= a;
    layer7_outputs(9249) <= not a or b;
    layer7_outputs(9250) <= a xor b;
    layer7_outputs(9251) <= a and not b;
    layer7_outputs(9252) <= b;
    layer7_outputs(9253) <= a and b;
    layer7_outputs(9254) <= a;
    layer7_outputs(9255) <= not b;
    layer7_outputs(9256) <= not (a xor b);
    layer7_outputs(9257) <= b;
    layer7_outputs(9258) <= not b;
    layer7_outputs(9259) <= not a;
    layer7_outputs(9260) <= b;
    layer7_outputs(9261) <= a;
    layer7_outputs(9262) <= a and b;
    layer7_outputs(9263) <= a;
    layer7_outputs(9264) <= not a or b;
    layer7_outputs(9265) <= not b;
    layer7_outputs(9266) <= b;
    layer7_outputs(9267) <= a and not b;
    layer7_outputs(9268) <= b and not a;
    layer7_outputs(9269) <= a and not b;
    layer7_outputs(9270) <= not b;
    layer7_outputs(9271) <= a;
    layer7_outputs(9272) <= a xor b;
    layer7_outputs(9273) <= b;
    layer7_outputs(9274) <= not a;
    layer7_outputs(9275) <= not b;
    layer7_outputs(9276) <= not (a and b);
    layer7_outputs(9277) <= not a;
    layer7_outputs(9278) <= b and not a;
    layer7_outputs(9279) <= not a or b;
    layer7_outputs(9280) <= not (a xor b);
    layer7_outputs(9281) <= not a or b;
    layer7_outputs(9282) <= b;
    layer7_outputs(9283) <= 1'b1;
    layer7_outputs(9284) <= a;
    layer7_outputs(9285) <= a;
    layer7_outputs(9286) <= a xor b;
    layer7_outputs(9287) <= a;
    layer7_outputs(9288) <= not (a and b);
    layer7_outputs(9289) <= a and b;
    layer7_outputs(9290) <= 1'b0;
    layer7_outputs(9291) <= b;
    layer7_outputs(9292) <= not (a and b);
    layer7_outputs(9293) <= not a;
    layer7_outputs(9294) <= b;
    layer7_outputs(9295) <= a and b;
    layer7_outputs(9296) <= not a or b;
    layer7_outputs(9297) <= b;
    layer7_outputs(9298) <= not (a xor b);
    layer7_outputs(9299) <= not (a or b);
    layer7_outputs(9300) <= a xor b;
    layer7_outputs(9301) <= b and not a;
    layer7_outputs(9302) <= not b or a;
    layer7_outputs(9303) <= not b;
    layer7_outputs(9304) <= not b;
    layer7_outputs(9305) <= a xor b;
    layer7_outputs(9306) <= a and not b;
    layer7_outputs(9307) <= not b;
    layer7_outputs(9308) <= a or b;
    layer7_outputs(9309) <= not a;
    layer7_outputs(9310) <= a xor b;
    layer7_outputs(9311) <= a xor b;
    layer7_outputs(9312) <= b;
    layer7_outputs(9313) <= a and not b;
    layer7_outputs(9314) <= not (a or b);
    layer7_outputs(9315) <= not (a xor b);
    layer7_outputs(9316) <= a;
    layer7_outputs(9317) <= a and b;
    layer7_outputs(9318) <= a and b;
    layer7_outputs(9319) <= not b;
    layer7_outputs(9320) <= b;
    layer7_outputs(9321) <= b;
    layer7_outputs(9322) <= a and b;
    layer7_outputs(9323) <= not b;
    layer7_outputs(9324) <= a and b;
    layer7_outputs(9325) <= a;
    layer7_outputs(9326) <= not (a and b);
    layer7_outputs(9327) <= not b;
    layer7_outputs(9328) <= a;
    layer7_outputs(9329) <= not a or b;
    layer7_outputs(9330) <= b;
    layer7_outputs(9331) <= not a or b;
    layer7_outputs(9332) <= not a;
    layer7_outputs(9333) <= a and b;
    layer7_outputs(9334) <= a xor b;
    layer7_outputs(9335) <= a or b;
    layer7_outputs(9336) <= not b or a;
    layer7_outputs(9337) <= b;
    layer7_outputs(9338) <= a and not b;
    layer7_outputs(9339) <= a;
    layer7_outputs(9340) <= a xor b;
    layer7_outputs(9341) <= a xor b;
    layer7_outputs(9342) <= a;
    layer7_outputs(9343) <= not a or b;
    layer7_outputs(9344) <= not a;
    layer7_outputs(9345) <= a and b;
    layer7_outputs(9346) <= not a;
    layer7_outputs(9347) <= not a or b;
    layer7_outputs(9348) <= a and b;
    layer7_outputs(9349) <= a xor b;
    layer7_outputs(9350) <= not (a xor b);
    layer7_outputs(9351) <= a or b;
    layer7_outputs(9352) <= not (a or b);
    layer7_outputs(9353) <= a;
    layer7_outputs(9354) <= a xor b;
    layer7_outputs(9355) <= not a;
    layer7_outputs(9356) <= not a;
    layer7_outputs(9357) <= not (a or b);
    layer7_outputs(9358) <= a;
    layer7_outputs(9359) <= a xor b;
    layer7_outputs(9360) <= a or b;
    layer7_outputs(9361) <= not (a xor b);
    layer7_outputs(9362) <= a;
    layer7_outputs(9363) <= a and b;
    layer7_outputs(9364) <= not (a xor b);
    layer7_outputs(9365) <= not a;
    layer7_outputs(9366) <= b and not a;
    layer7_outputs(9367) <= a and not b;
    layer7_outputs(9368) <= a and b;
    layer7_outputs(9369) <= not b;
    layer7_outputs(9370) <= a;
    layer7_outputs(9371) <= not a;
    layer7_outputs(9372) <= a xor b;
    layer7_outputs(9373) <= 1'b1;
    layer7_outputs(9374) <= a;
    layer7_outputs(9375) <= a or b;
    layer7_outputs(9376) <= 1'b0;
    layer7_outputs(9377) <= a or b;
    layer7_outputs(9378) <= a or b;
    layer7_outputs(9379) <= a xor b;
    layer7_outputs(9380) <= not a;
    layer7_outputs(9381) <= not (a and b);
    layer7_outputs(9382) <= a xor b;
    layer7_outputs(9383) <= 1'b1;
    layer7_outputs(9384) <= not a;
    layer7_outputs(9385) <= a;
    layer7_outputs(9386) <= not b;
    layer7_outputs(9387) <= 1'b1;
    layer7_outputs(9388) <= b;
    layer7_outputs(9389) <= not (a xor b);
    layer7_outputs(9390) <= a and b;
    layer7_outputs(9391) <= a or b;
    layer7_outputs(9392) <= b and not a;
    layer7_outputs(9393) <= a;
    layer7_outputs(9394) <= not a;
    layer7_outputs(9395) <= a;
    layer7_outputs(9396) <= not b;
    layer7_outputs(9397) <= not a;
    layer7_outputs(9398) <= a and b;
    layer7_outputs(9399) <= not b;
    layer7_outputs(9400) <= b;
    layer7_outputs(9401) <= b;
    layer7_outputs(9402) <= not (a and b);
    layer7_outputs(9403) <= a xor b;
    layer7_outputs(9404) <= not (a and b);
    layer7_outputs(9405) <= not (a xor b);
    layer7_outputs(9406) <= a xor b;
    layer7_outputs(9407) <= b;
    layer7_outputs(9408) <= not (a and b);
    layer7_outputs(9409) <= b;
    layer7_outputs(9410) <= not b;
    layer7_outputs(9411) <= b;
    layer7_outputs(9412) <= a xor b;
    layer7_outputs(9413) <= b;
    layer7_outputs(9414) <= not a or b;
    layer7_outputs(9415) <= a and b;
    layer7_outputs(9416) <= not a or b;
    layer7_outputs(9417) <= not a;
    layer7_outputs(9418) <= not b;
    layer7_outputs(9419) <= not b;
    layer7_outputs(9420) <= not (a xor b);
    layer7_outputs(9421) <= not a;
    layer7_outputs(9422) <= not b;
    layer7_outputs(9423) <= not b;
    layer7_outputs(9424) <= a and not b;
    layer7_outputs(9425) <= a;
    layer7_outputs(9426) <= not b;
    layer7_outputs(9427) <= a and b;
    layer7_outputs(9428) <= b;
    layer7_outputs(9429) <= a xor b;
    layer7_outputs(9430) <= 1'b1;
    layer7_outputs(9431) <= a and not b;
    layer7_outputs(9432) <= not b;
    layer7_outputs(9433) <= b;
    layer7_outputs(9434) <= b and not a;
    layer7_outputs(9435) <= a;
    layer7_outputs(9436) <= not a or b;
    layer7_outputs(9437) <= a xor b;
    layer7_outputs(9438) <= not a;
    layer7_outputs(9439) <= not (a or b);
    layer7_outputs(9440) <= 1'b0;
    layer7_outputs(9441) <= a;
    layer7_outputs(9442) <= b and not a;
    layer7_outputs(9443) <= not b;
    layer7_outputs(9444) <= b and not a;
    layer7_outputs(9445) <= a xor b;
    layer7_outputs(9446) <= a;
    layer7_outputs(9447) <= a and not b;
    layer7_outputs(9448) <= not b;
    layer7_outputs(9449) <= not (a xor b);
    layer7_outputs(9450) <= not (a or b);
    layer7_outputs(9451) <= b;
    layer7_outputs(9452) <= not a;
    layer7_outputs(9453) <= b;
    layer7_outputs(9454) <= b;
    layer7_outputs(9455) <= not b;
    layer7_outputs(9456) <= not (a and b);
    layer7_outputs(9457) <= a and not b;
    layer7_outputs(9458) <= not a;
    layer7_outputs(9459) <= not (a and b);
    layer7_outputs(9460) <= a or b;
    layer7_outputs(9461) <= not b;
    layer7_outputs(9462) <= not a;
    layer7_outputs(9463) <= a;
    layer7_outputs(9464) <= not (a and b);
    layer7_outputs(9465) <= not a;
    layer7_outputs(9466) <= not a;
    layer7_outputs(9467) <= not (a and b);
    layer7_outputs(9468) <= a;
    layer7_outputs(9469) <= a;
    layer7_outputs(9470) <= b;
    layer7_outputs(9471) <= not a or b;
    layer7_outputs(9472) <= a or b;
    layer7_outputs(9473) <= b and not a;
    layer7_outputs(9474) <= a or b;
    layer7_outputs(9475) <= a or b;
    layer7_outputs(9476) <= not (a and b);
    layer7_outputs(9477) <= a;
    layer7_outputs(9478) <= a xor b;
    layer7_outputs(9479) <= not b;
    layer7_outputs(9480) <= 1'b1;
    layer7_outputs(9481) <= not (a and b);
    layer7_outputs(9482) <= a and b;
    layer7_outputs(9483) <= a;
    layer7_outputs(9484) <= not b;
    layer7_outputs(9485) <= b and not a;
    layer7_outputs(9486) <= a;
    layer7_outputs(9487) <= b and not a;
    layer7_outputs(9488) <= b;
    layer7_outputs(9489) <= not a;
    layer7_outputs(9490) <= not (a and b);
    layer7_outputs(9491) <= not b;
    layer7_outputs(9492) <= b;
    layer7_outputs(9493) <= not a;
    layer7_outputs(9494) <= b;
    layer7_outputs(9495) <= a;
    layer7_outputs(9496) <= a;
    layer7_outputs(9497) <= not a or b;
    layer7_outputs(9498) <= a and not b;
    layer7_outputs(9499) <= b;
    layer7_outputs(9500) <= not a or b;
    layer7_outputs(9501) <= not (a xor b);
    layer7_outputs(9502) <= 1'b1;
    layer7_outputs(9503) <= a;
    layer7_outputs(9504) <= b;
    layer7_outputs(9505) <= not a or b;
    layer7_outputs(9506) <= not (a or b);
    layer7_outputs(9507) <= a;
    layer7_outputs(9508) <= not a;
    layer7_outputs(9509) <= not (a or b);
    layer7_outputs(9510) <= not a or b;
    layer7_outputs(9511) <= not b;
    layer7_outputs(9512) <= not (a and b);
    layer7_outputs(9513) <= b;
    layer7_outputs(9514) <= not a;
    layer7_outputs(9515) <= not (a xor b);
    layer7_outputs(9516) <= a;
    layer7_outputs(9517) <= b;
    layer7_outputs(9518) <= not (a and b);
    layer7_outputs(9519) <= a;
    layer7_outputs(9520) <= b;
    layer7_outputs(9521) <= a;
    layer7_outputs(9522) <= 1'b0;
    layer7_outputs(9523) <= b;
    layer7_outputs(9524) <= a xor b;
    layer7_outputs(9525) <= not (a or b);
    layer7_outputs(9526) <= a xor b;
    layer7_outputs(9527) <= a;
    layer7_outputs(9528) <= not (a xor b);
    layer7_outputs(9529) <= a xor b;
    layer7_outputs(9530) <= not (a and b);
    layer7_outputs(9531) <= a and not b;
    layer7_outputs(9532) <= a and not b;
    layer7_outputs(9533) <= b;
    layer7_outputs(9534) <= a;
    layer7_outputs(9535) <= b;
    layer7_outputs(9536) <= b;
    layer7_outputs(9537) <= a and b;
    layer7_outputs(9538) <= a and b;
    layer7_outputs(9539) <= a or b;
    layer7_outputs(9540) <= not a;
    layer7_outputs(9541) <= a xor b;
    layer7_outputs(9542) <= not b;
    layer7_outputs(9543) <= not a or b;
    layer7_outputs(9544) <= b;
    layer7_outputs(9545) <= a or b;
    layer7_outputs(9546) <= a;
    layer7_outputs(9547) <= b;
    layer7_outputs(9548) <= not a;
    layer7_outputs(9549) <= a and b;
    layer7_outputs(9550) <= a;
    layer7_outputs(9551) <= b;
    layer7_outputs(9552) <= not (a xor b);
    layer7_outputs(9553) <= a;
    layer7_outputs(9554) <= not a;
    layer7_outputs(9555) <= not a;
    layer7_outputs(9556) <= a and not b;
    layer7_outputs(9557) <= not b;
    layer7_outputs(9558) <= not b;
    layer7_outputs(9559) <= not (a xor b);
    layer7_outputs(9560) <= not (a or b);
    layer7_outputs(9561) <= not a or b;
    layer7_outputs(9562) <= not a or b;
    layer7_outputs(9563) <= not a;
    layer7_outputs(9564) <= not (a and b);
    layer7_outputs(9565) <= 1'b0;
    layer7_outputs(9566) <= a and not b;
    layer7_outputs(9567) <= a xor b;
    layer7_outputs(9568) <= not b;
    layer7_outputs(9569) <= not (a and b);
    layer7_outputs(9570) <= not (a xor b);
    layer7_outputs(9571) <= a and not b;
    layer7_outputs(9572) <= not a;
    layer7_outputs(9573) <= a;
    layer7_outputs(9574) <= not a or b;
    layer7_outputs(9575) <= a and not b;
    layer7_outputs(9576) <= a xor b;
    layer7_outputs(9577) <= not (a and b);
    layer7_outputs(9578) <= not b;
    layer7_outputs(9579) <= not (a xor b);
    layer7_outputs(9580) <= not a;
    layer7_outputs(9581) <= b;
    layer7_outputs(9582) <= a xor b;
    layer7_outputs(9583) <= not a;
    layer7_outputs(9584) <= b;
    layer7_outputs(9585) <= not b or a;
    layer7_outputs(9586) <= a or b;
    layer7_outputs(9587) <= not a;
    layer7_outputs(9588) <= b;
    layer7_outputs(9589) <= not b or a;
    layer7_outputs(9590) <= a and not b;
    layer7_outputs(9591) <= not a;
    layer7_outputs(9592) <= a or b;
    layer7_outputs(9593) <= not b;
    layer7_outputs(9594) <= a xor b;
    layer7_outputs(9595) <= a xor b;
    layer7_outputs(9596) <= a or b;
    layer7_outputs(9597) <= a xor b;
    layer7_outputs(9598) <= b;
    layer7_outputs(9599) <= not (a or b);
    layer7_outputs(9600) <= not (a or b);
    layer7_outputs(9601) <= b;
    layer7_outputs(9602) <= not b;
    layer7_outputs(9603) <= not a;
    layer7_outputs(9604) <= not b;
    layer7_outputs(9605) <= a xor b;
    layer7_outputs(9606) <= a or b;
    layer7_outputs(9607) <= not b or a;
    layer7_outputs(9608) <= not (a xor b);
    layer7_outputs(9609) <= not a;
    layer7_outputs(9610) <= a or b;
    layer7_outputs(9611) <= b and not a;
    layer7_outputs(9612) <= not (a or b);
    layer7_outputs(9613) <= not (a and b);
    layer7_outputs(9614) <= a and not b;
    layer7_outputs(9615) <= not (a xor b);
    layer7_outputs(9616) <= a xor b;
    layer7_outputs(9617) <= a or b;
    layer7_outputs(9618) <= a xor b;
    layer7_outputs(9619) <= a and b;
    layer7_outputs(9620) <= a;
    layer7_outputs(9621) <= a and b;
    layer7_outputs(9622) <= 1'b1;
    layer7_outputs(9623) <= a;
    layer7_outputs(9624) <= not (a or b);
    layer7_outputs(9625) <= a;
    layer7_outputs(9626) <= b;
    layer7_outputs(9627) <= b;
    layer7_outputs(9628) <= not (a and b);
    layer7_outputs(9629) <= b;
    layer7_outputs(9630) <= a;
    layer7_outputs(9631) <= not b or a;
    layer7_outputs(9632) <= not b;
    layer7_outputs(9633) <= b;
    layer7_outputs(9634) <= a;
    layer7_outputs(9635) <= a and b;
    layer7_outputs(9636) <= not (a or b);
    layer7_outputs(9637) <= a and not b;
    layer7_outputs(9638) <= a;
    layer7_outputs(9639) <= 1'b1;
    layer7_outputs(9640) <= b;
    layer7_outputs(9641) <= a;
    layer7_outputs(9642) <= b;
    layer7_outputs(9643) <= a xor b;
    layer7_outputs(9644) <= 1'b1;
    layer7_outputs(9645) <= b and not a;
    layer7_outputs(9646) <= a or b;
    layer7_outputs(9647) <= a xor b;
    layer7_outputs(9648) <= b;
    layer7_outputs(9649) <= not a;
    layer7_outputs(9650) <= b;
    layer7_outputs(9651) <= a xor b;
    layer7_outputs(9652) <= 1'b0;
    layer7_outputs(9653) <= b;
    layer7_outputs(9654) <= a xor b;
    layer7_outputs(9655) <= b and not a;
    layer7_outputs(9656) <= b;
    layer7_outputs(9657) <= a;
    layer7_outputs(9658) <= not a;
    layer7_outputs(9659) <= not (a xor b);
    layer7_outputs(9660) <= a;
    layer7_outputs(9661) <= a;
    layer7_outputs(9662) <= a and b;
    layer7_outputs(9663) <= a;
    layer7_outputs(9664) <= b;
    layer7_outputs(9665) <= not (a xor b);
    layer7_outputs(9666) <= not b or a;
    layer7_outputs(9667) <= not a;
    layer7_outputs(9668) <= not a or b;
    layer7_outputs(9669) <= not b;
    layer7_outputs(9670) <= not a or b;
    layer7_outputs(9671) <= not b or a;
    layer7_outputs(9672) <= b and not a;
    layer7_outputs(9673) <= not a;
    layer7_outputs(9674) <= a xor b;
    layer7_outputs(9675) <= a xor b;
    layer7_outputs(9676) <= b;
    layer7_outputs(9677) <= not a;
    layer7_outputs(9678) <= not a;
    layer7_outputs(9679) <= not (a and b);
    layer7_outputs(9680) <= b;
    layer7_outputs(9681) <= not b or a;
    layer7_outputs(9682) <= a;
    layer7_outputs(9683) <= not b;
    layer7_outputs(9684) <= not (a or b);
    layer7_outputs(9685) <= not a;
    layer7_outputs(9686) <= b;
    layer7_outputs(9687) <= a xor b;
    layer7_outputs(9688) <= not a;
    layer7_outputs(9689) <= not a or b;
    layer7_outputs(9690) <= not a or b;
    layer7_outputs(9691) <= a and not b;
    layer7_outputs(9692) <= not a;
    layer7_outputs(9693) <= b;
    layer7_outputs(9694) <= a;
    layer7_outputs(9695) <= not a;
    layer7_outputs(9696) <= not (a and b);
    layer7_outputs(9697) <= a and not b;
    layer7_outputs(9698) <= not (a and b);
    layer7_outputs(9699) <= a and not b;
    layer7_outputs(9700) <= not (a xor b);
    layer7_outputs(9701) <= not b;
    layer7_outputs(9702) <= a and not b;
    layer7_outputs(9703) <= a and b;
    layer7_outputs(9704) <= not (a and b);
    layer7_outputs(9705) <= not a;
    layer7_outputs(9706) <= not b;
    layer7_outputs(9707) <= b and not a;
    layer7_outputs(9708) <= a xor b;
    layer7_outputs(9709) <= not b;
    layer7_outputs(9710) <= a and not b;
    layer7_outputs(9711) <= not (a or b);
    layer7_outputs(9712) <= not b;
    layer7_outputs(9713) <= not (a xor b);
    layer7_outputs(9714) <= a xor b;
    layer7_outputs(9715) <= not b;
    layer7_outputs(9716) <= a and b;
    layer7_outputs(9717) <= 1'b0;
    layer7_outputs(9718) <= b and not a;
    layer7_outputs(9719) <= not a;
    layer7_outputs(9720) <= not a;
    layer7_outputs(9721) <= not (a or b);
    layer7_outputs(9722) <= a;
    layer7_outputs(9723) <= not b or a;
    layer7_outputs(9724) <= 1'b0;
    layer7_outputs(9725) <= not a;
    layer7_outputs(9726) <= a or b;
    layer7_outputs(9727) <= a xor b;
    layer7_outputs(9728) <= not (a or b);
    layer7_outputs(9729) <= not a or b;
    layer7_outputs(9730) <= a xor b;
    layer7_outputs(9731) <= a or b;
    layer7_outputs(9732) <= a;
    layer7_outputs(9733) <= 1'b1;
    layer7_outputs(9734) <= a xor b;
    layer7_outputs(9735) <= not (a xor b);
    layer7_outputs(9736) <= not a or b;
    layer7_outputs(9737) <= not b or a;
    layer7_outputs(9738) <= a or b;
    layer7_outputs(9739) <= a xor b;
    layer7_outputs(9740) <= b;
    layer7_outputs(9741) <= not a;
    layer7_outputs(9742) <= a xor b;
    layer7_outputs(9743) <= a or b;
    layer7_outputs(9744) <= not (a or b);
    layer7_outputs(9745) <= a xor b;
    layer7_outputs(9746) <= not a or b;
    layer7_outputs(9747) <= not b;
    layer7_outputs(9748) <= not (a xor b);
    layer7_outputs(9749) <= a;
    layer7_outputs(9750) <= a;
    layer7_outputs(9751) <= b;
    layer7_outputs(9752) <= not a;
    layer7_outputs(9753) <= 1'b1;
    layer7_outputs(9754) <= 1'b0;
    layer7_outputs(9755) <= not b;
    layer7_outputs(9756) <= not a;
    layer7_outputs(9757) <= not (a xor b);
    layer7_outputs(9758) <= a;
    layer7_outputs(9759) <= a and not b;
    layer7_outputs(9760) <= not b;
    layer7_outputs(9761) <= not b;
    layer7_outputs(9762) <= not b;
    layer7_outputs(9763) <= not a;
    layer7_outputs(9764) <= a and not b;
    layer7_outputs(9765) <= b;
    layer7_outputs(9766) <= not (a xor b);
    layer7_outputs(9767) <= not a;
    layer7_outputs(9768) <= not b or a;
    layer7_outputs(9769) <= not b;
    layer7_outputs(9770) <= not b or a;
    layer7_outputs(9771) <= not (a and b);
    layer7_outputs(9772) <= a xor b;
    layer7_outputs(9773) <= not (a xor b);
    layer7_outputs(9774) <= not (a and b);
    layer7_outputs(9775) <= not b;
    layer7_outputs(9776) <= a xor b;
    layer7_outputs(9777) <= not b;
    layer7_outputs(9778) <= a and not b;
    layer7_outputs(9779) <= not a or b;
    layer7_outputs(9780) <= b;
    layer7_outputs(9781) <= b;
    layer7_outputs(9782) <= a;
    layer7_outputs(9783) <= b;
    layer7_outputs(9784) <= 1'b1;
    layer7_outputs(9785) <= a;
    layer7_outputs(9786) <= not a;
    layer7_outputs(9787) <= a;
    layer7_outputs(9788) <= a and b;
    layer7_outputs(9789) <= 1'b1;
    layer7_outputs(9790) <= a;
    layer7_outputs(9791) <= b;
    layer7_outputs(9792) <= b;
    layer7_outputs(9793) <= a and not b;
    layer7_outputs(9794) <= not (a or b);
    layer7_outputs(9795) <= a and b;
    layer7_outputs(9796) <= a;
    layer7_outputs(9797) <= not a or b;
    layer7_outputs(9798) <= b;
    layer7_outputs(9799) <= a xor b;
    layer7_outputs(9800) <= a or b;
    layer7_outputs(9801) <= a;
    layer7_outputs(9802) <= a and not b;
    layer7_outputs(9803) <= b;
    layer7_outputs(9804) <= not b or a;
    layer7_outputs(9805) <= b;
    layer7_outputs(9806) <= b and not a;
    layer7_outputs(9807) <= a;
    layer7_outputs(9808) <= a or b;
    layer7_outputs(9809) <= not b or a;
    layer7_outputs(9810) <= not b;
    layer7_outputs(9811) <= not a;
    layer7_outputs(9812) <= not b;
    layer7_outputs(9813) <= not (a or b);
    layer7_outputs(9814) <= a and b;
    layer7_outputs(9815) <= not a;
    layer7_outputs(9816) <= b and not a;
    layer7_outputs(9817) <= not (a or b);
    layer7_outputs(9818) <= not a or b;
    layer7_outputs(9819) <= b;
    layer7_outputs(9820) <= not a;
    layer7_outputs(9821) <= not b;
    layer7_outputs(9822) <= a xor b;
    layer7_outputs(9823) <= not a;
    layer7_outputs(9824) <= 1'b0;
    layer7_outputs(9825) <= a and b;
    layer7_outputs(9826) <= not a;
    layer7_outputs(9827) <= a xor b;
    layer7_outputs(9828) <= a and not b;
    layer7_outputs(9829) <= not a or b;
    layer7_outputs(9830) <= a and not b;
    layer7_outputs(9831) <= not (a xor b);
    layer7_outputs(9832) <= a and not b;
    layer7_outputs(9833) <= not a;
    layer7_outputs(9834) <= a and b;
    layer7_outputs(9835) <= a;
    layer7_outputs(9836) <= b and not a;
    layer7_outputs(9837) <= not (a or b);
    layer7_outputs(9838) <= a;
    layer7_outputs(9839) <= not b or a;
    layer7_outputs(9840) <= not (a or b);
    layer7_outputs(9841) <= not b or a;
    layer7_outputs(9842) <= b;
    layer7_outputs(9843) <= not (a or b);
    layer7_outputs(9844) <= not a;
    layer7_outputs(9845) <= not (a xor b);
    layer7_outputs(9846) <= not (a xor b);
    layer7_outputs(9847) <= not b;
    layer7_outputs(9848) <= not (a or b);
    layer7_outputs(9849) <= a or b;
    layer7_outputs(9850) <= not a;
    layer7_outputs(9851) <= not (a and b);
    layer7_outputs(9852) <= not b;
    layer7_outputs(9853) <= b and not a;
    layer7_outputs(9854) <= b and not a;
    layer7_outputs(9855) <= a and not b;
    layer7_outputs(9856) <= not (a and b);
    layer7_outputs(9857) <= not b;
    layer7_outputs(9858) <= not a or b;
    layer7_outputs(9859) <= not a;
    layer7_outputs(9860) <= not a;
    layer7_outputs(9861) <= b;
    layer7_outputs(9862) <= a;
    layer7_outputs(9863) <= b and not a;
    layer7_outputs(9864) <= not a or b;
    layer7_outputs(9865) <= not (a xor b);
    layer7_outputs(9866) <= a;
    layer7_outputs(9867) <= a and not b;
    layer7_outputs(9868) <= b;
    layer7_outputs(9869) <= not b;
    layer7_outputs(9870) <= not b;
    layer7_outputs(9871) <= not (a or b);
    layer7_outputs(9872) <= not (a or b);
    layer7_outputs(9873) <= b;
    layer7_outputs(9874) <= a;
    layer7_outputs(9875) <= a and b;
    layer7_outputs(9876) <= a;
    layer7_outputs(9877) <= not a;
    layer7_outputs(9878) <= not b or a;
    layer7_outputs(9879) <= not b or a;
    layer7_outputs(9880) <= not (a or b);
    layer7_outputs(9881) <= not a or b;
    layer7_outputs(9882) <= a xor b;
    layer7_outputs(9883) <= b;
    layer7_outputs(9884) <= not b;
    layer7_outputs(9885) <= not a;
    layer7_outputs(9886) <= not a or b;
    layer7_outputs(9887) <= a xor b;
    layer7_outputs(9888) <= b;
    layer7_outputs(9889) <= not a;
    layer7_outputs(9890) <= a and b;
    layer7_outputs(9891) <= a xor b;
    layer7_outputs(9892) <= a and b;
    layer7_outputs(9893) <= a xor b;
    layer7_outputs(9894) <= b and not a;
    layer7_outputs(9895) <= b;
    layer7_outputs(9896) <= not (a or b);
    layer7_outputs(9897) <= not b;
    layer7_outputs(9898) <= b and not a;
    layer7_outputs(9899) <= not b;
    layer7_outputs(9900) <= not (a or b);
    layer7_outputs(9901) <= b and not a;
    layer7_outputs(9902) <= a;
    layer7_outputs(9903) <= not b or a;
    layer7_outputs(9904) <= a xor b;
    layer7_outputs(9905) <= not b;
    layer7_outputs(9906) <= a and not b;
    layer7_outputs(9907) <= not (a xor b);
    layer7_outputs(9908) <= a;
    layer7_outputs(9909) <= a and b;
    layer7_outputs(9910) <= not (a and b);
    layer7_outputs(9911) <= a xor b;
    layer7_outputs(9912) <= not b;
    layer7_outputs(9913) <= b and not a;
    layer7_outputs(9914) <= a xor b;
    layer7_outputs(9915) <= a;
    layer7_outputs(9916) <= a and not b;
    layer7_outputs(9917) <= not a or b;
    layer7_outputs(9918) <= not a;
    layer7_outputs(9919) <= a or b;
    layer7_outputs(9920) <= b;
    layer7_outputs(9921) <= b;
    layer7_outputs(9922) <= a or b;
    layer7_outputs(9923) <= b and not a;
    layer7_outputs(9924) <= b;
    layer7_outputs(9925) <= a xor b;
    layer7_outputs(9926) <= b and not a;
    layer7_outputs(9927) <= a;
    layer7_outputs(9928) <= not b;
    layer7_outputs(9929) <= a;
    layer7_outputs(9930) <= a xor b;
    layer7_outputs(9931) <= not b;
    layer7_outputs(9932) <= b;
    layer7_outputs(9933) <= not a;
    layer7_outputs(9934) <= not b;
    layer7_outputs(9935) <= not a or b;
    layer7_outputs(9936) <= not (a xor b);
    layer7_outputs(9937) <= not (a xor b);
    layer7_outputs(9938) <= a and not b;
    layer7_outputs(9939) <= a or b;
    layer7_outputs(9940) <= a;
    layer7_outputs(9941) <= not b or a;
    layer7_outputs(9942) <= a;
    layer7_outputs(9943) <= a xor b;
    layer7_outputs(9944) <= a xor b;
    layer7_outputs(9945) <= not b or a;
    layer7_outputs(9946) <= not (a and b);
    layer7_outputs(9947) <= b and not a;
    layer7_outputs(9948) <= not (a and b);
    layer7_outputs(9949) <= not b or a;
    layer7_outputs(9950) <= a xor b;
    layer7_outputs(9951) <= a;
    layer7_outputs(9952) <= not b;
    layer7_outputs(9953) <= not b;
    layer7_outputs(9954) <= not (a xor b);
    layer7_outputs(9955) <= not b;
    layer7_outputs(9956) <= a and not b;
    layer7_outputs(9957) <= a and b;
    layer7_outputs(9958) <= a;
    layer7_outputs(9959) <= 1'b0;
    layer7_outputs(9960) <= b and not a;
    layer7_outputs(9961) <= a;
    layer7_outputs(9962) <= a xor b;
    layer7_outputs(9963) <= not (a and b);
    layer7_outputs(9964) <= not (a and b);
    layer7_outputs(9965) <= a and b;
    layer7_outputs(9966) <= a and b;
    layer7_outputs(9967) <= not (a xor b);
    layer7_outputs(9968) <= 1'b0;
    layer7_outputs(9969) <= not b;
    layer7_outputs(9970) <= not (a or b);
    layer7_outputs(9971) <= not a;
    layer7_outputs(9972) <= not (a or b);
    layer7_outputs(9973) <= not a;
    layer7_outputs(9974) <= b;
    layer7_outputs(9975) <= a xor b;
    layer7_outputs(9976) <= a and not b;
    layer7_outputs(9977) <= a xor b;
    layer7_outputs(9978) <= a or b;
    layer7_outputs(9979) <= a and b;
    layer7_outputs(9980) <= a;
    layer7_outputs(9981) <= a and not b;
    layer7_outputs(9982) <= b;
    layer7_outputs(9983) <= b;
    layer7_outputs(9984) <= not (a xor b);
    layer7_outputs(9985) <= not a;
    layer7_outputs(9986) <= a xor b;
    layer7_outputs(9987) <= not b or a;
    layer7_outputs(9988) <= not (a xor b);
    layer7_outputs(9989) <= not b;
    layer7_outputs(9990) <= b;
    layer7_outputs(9991) <= a;
    layer7_outputs(9992) <= b;
    layer7_outputs(9993) <= b;
    layer7_outputs(9994) <= not b or a;
    layer7_outputs(9995) <= a and b;
    layer7_outputs(9996) <= b;
    layer7_outputs(9997) <= a and b;
    layer7_outputs(9998) <= a;
    layer7_outputs(9999) <= not b;
    layer7_outputs(10000) <= not b;
    layer7_outputs(10001) <= b;
    layer7_outputs(10002) <= a xor b;
    layer7_outputs(10003) <= not (a xor b);
    layer7_outputs(10004) <= a;
    layer7_outputs(10005) <= a or b;
    layer7_outputs(10006) <= a;
    layer7_outputs(10007) <= a and b;
    layer7_outputs(10008) <= a and not b;
    layer7_outputs(10009) <= a or b;
    layer7_outputs(10010) <= not b;
    layer7_outputs(10011) <= not a or b;
    layer7_outputs(10012) <= a;
    layer7_outputs(10013) <= not b or a;
    layer7_outputs(10014) <= a;
    layer7_outputs(10015) <= a and not b;
    layer7_outputs(10016) <= not a;
    layer7_outputs(10017) <= a;
    layer7_outputs(10018) <= b and not a;
    layer7_outputs(10019) <= not a;
    layer7_outputs(10020) <= a or b;
    layer7_outputs(10021) <= not a;
    layer7_outputs(10022) <= not (a xor b);
    layer7_outputs(10023) <= not b;
    layer7_outputs(10024) <= b;
    layer7_outputs(10025) <= a and b;
    layer7_outputs(10026) <= not a;
    layer7_outputs(10027) <= a xor b;
    layer7_outputs(10028) <= not a;
    layer7_outputs(10029) <= a;
    layer7_outputs(10030) <= not b;
    layer7_outputs(10031) <= not b;
    layer7_outputs(10032) <= not (a or b);
    layer7_outputs(10033) <= a and not b;
    layer7_outputs(10034) <= a xor b;
    layer7_outputs(10035) <= b and not a;
    layer7_outputs(10036) <= a;
    layer7_outputs(10037) <= a;
    layer7_outputs(10038) <= a xor b;
    layer7_outputs(10039) <= not b;
    layer7_outputs(10040) <= not b;
    layer7_outputs(10041) <= b;
    layer7_outputs(10042) <= a and not b;
    layer7_outputs(10043) <= a and not b;
    layer7_outputs(10044) <= not a;
    layer7_outputs(10045) <= not (a or b);
    layer7_outputs(10046) <= b;
    layer7_outputs(10047) <= a or b;
    layer7_outputs(10048) <= not (a xor b);
    layer7_outputs(10049) <= not (a or b);
    layer7_outputs(10050) <= not (a xor b);
    layer7_outputs(10051) <= b;
    layer7_outputs(10052) <= not (a or b);
    layer7_outputs(10053) <= b;
    layer7_outputs(10054) <= b;
    layer7_outputs(10055) <= not b;
    layer7_outputs(10056) <= not a or b;
    layer7_outputs(10057) <= not (a xor b);
    layer7_outputs(10058) <= a;
    layer7_outputs(10059) <= b;
    layer7_outputs(10060) <= a xor b;
    layer7_outputs(10061) <= not b;
    layer7_outputs(10062) <= not (a or b);
    layer7_outputs(10063) <= not (a and b);
    layer7_outputs(10064) <= 1'b1;
    layer7_outputs(10065) <= b and not a;
    layer7_outputs(10066) <= b;
    layer7_outputs(10067) <= a or b;
    layer7_outputs(10068) <= a xor b;
    layer7_outputs(10069) <= not a or b;
    layer7_outputs(10070) <= not b;
    layer7_outputs(10071) <= not (a xor b);
    layer7_outputs(10072) <= not b;
    layer7_outputs(10073) <= b and not a;
    layer7_outputs(10074) <= a or b;
    layer7_outputs(10075) <= a or b;
    layer7_outputs(10076) <= b;
    layer7_outputs(10077) <= a or b;
    layer7_outputs(10078) <= b;
    layer7_outputs(10079) <= not a;
    layer7_outputs(10080) <= not a;
    layer7_outputs(10081) <= b and not a;
    layer7_outputs(10082) <= a;
    layer7_outputs(10083) <= a and not b;
    layer7_outputs(10084) <= not b;
    layer7_outputs(10085) <= a and b;
    layer7_outputs(10086) <= not b or a;
    layer7_outputs(10087) <= a xor b;
    layer7_outputs(10088) <= b;
    layer7_outputs(10089) <= not (a xor b);
    layer7_outputs(10090) <= b;
    layer7_outputs(10091) <= a and b;
    layer7_outputs(10092) <= a and not b;
    layer7_outputs(10093) <= not a;
    layer7_outputs(10094) <= not b or a;
    layer7_outputs(10095) <= a or b;
    layer7_outputs(10096) <= a;
    layer7_outputs(10097) <= not (a and b);
    layer7_outputs(10098) <= a and b;
    layer7_outputs(10099) <= a and not b;
    layer7_outputs(10100) <= not (a or b);
    layer7_outputs(10101) <= not b;
    layer7_outputs(10102) <= a;
    layer7_outputs(10103) <= 1'b1;
    layer7_outputs(10104) <= not b;
    layer7_outputs(10105) <= not (a xor b);
    layer7_outputs(10106) <= not b;
    layer7_outputs(10107) <= a and not b;
    layer7_outputs(10108) <= not a or b;
    layer7_outputs(10109) <= b and not a;
    layer7_outputs(10110) <= a xor b;
    layer7_outputs(10111) <= a and b;
    layer7_outputs(10112) <= not a or b;
    layer7_outputs(10113) <= not b;
    layer7_outputs(10114) <= not a or b;
    layer7_outputs(10115) <= b and not a;
    layer7_outputs(10116) <= not a;
    layer7_outputs(10117) <= not b;
    layer7_outputs(10118) <= b;
    layer7_outputs(10119) <= a or b;
    layer7_outputs(10120) <= not b;
    layer7_outputs(10121) <= b and not a;
    layer7_outputs(10122) <= not (a xor b);
    layer7_outputs(10123) <= a;
    layer7_outputs(10124) <= not a or b;
    layer7_outputs(10125) <= b and not a;
    layer7_outputs(10126) <= not b or a;
    layer7_outputs(10127) <= not a or b;
    layer7_outputs(10128) <= 1'b1;
    layer7_outputs(10129) <= a;
    layer7_outputs(10130) <= not a or b;
    layer7_outputs(10131) <= not a;
    layer7_outputs(10132) <= a xor b;
    layer7_outputs(10133) <= b;
    layer7_outputs(10134) <= not a;
    layer7_outputs(10135) <= b;
    layer7_outputs(10136) <= a xor b;
    layer7_outputs(10137) <= a or b;
    layer7_outputs(10138) <= a xor b;
    layer7_outputs(10139) <= not b;
    layer7_outputs(10140) <= a;
    layer7_outputs(10141) <= not (a and b);
    layer7_outputs(10142) <= a xor b;
    layer7_outputs(10143) <= not b;
    layer7_outputs(10144) <= a or b;
    layer7_outputs(10145) <= a and b;
    layer7_outputs(10146) <= not b;
    layer7_outputs(10147) <= not b;
    layer7_outputs(10148) <= not b or a;
    layer7_outputs(10149) <= not a or b;
    layer7_outputs(10150) <= a xor b;
    layer7_outputs(10151) <= b;
    layer7_outputs(10152) <= a;
    layer7_outputs(10153) <= not (a xor b);
    layer7_outputs(10154) <= not a or b;
    layer7_outputs(10155) <= not (a xor b);
    layer7_outputs(10156) <= a and not b;
    layer7_outputs(10157) <= not a;
    layer7_outputs(10158) <= a;
    layer7_outputs(10159) <= a;
    layer7_outputs(10160) <= b;
    layer7_outputs(10161) <= a or b;
    layer7_outputs(10162) <= not b;
    layer7_outputs(10163) <= a xor b;
    layer7_outputs(10164) <= a;
    layer7_outputs(10165) <= b;
    layer7_outputs(10166) <= a;
    layer7_outputs(10167) <= b and not a;
    layer7_outputs(10168) <= b;
    layer7_outputs(10169) <= not (a xor b);
    layer7_outputs(10170) <= not a or b;
    layer7_outputs(10171) <= b and not a;
    layer7_outputs(10172) <= a;
    layer7_outputs(10173) <= a;
    layer7_outputs(10174) <= b;
    layer7_outputs(10175) <= not a;
    layer7_outputs(10176) <= not a;
    layer7_outputs(10177) <= a or b;
    layer7_outputs(10178) <= not b;
    layer7_outputs(10179) <= b;
    layer7_outputs(10180) <= b;
    layer7_outputs(10181) <= not a;
    layer7_outputs(10182) <= not (a xor b);
    layer7_outputs(10183) <= not b;
    layer7_outputs(10184) <= not b;
    layer7_outputs(10185) <= a and b;
    layer7_outputs(10186) <= not (a xor b);
    layer7_outputs(10187) <= not (a and b);
    layer7_outputs(10188) <= not (a and b);
    layer7_outputs(10189) <= not a;
    layer7_outputs(10190) <= not a;
    layer7_outputs(10191) <= 1'b0;
    layer7_outputs(10192) <= b and not a;
    layer7_outputs(10193) <= not a;
    layer7_outputs(10194) <= b;
    layer7_outputs(10195) <= b and not a;
    layer7_outputs(10196) <= a xor b;
    layer7_outputs(10197) <= b;
    layer7_outputs(10198) <= not a or b;
    layer7_outputs(10199) <= not (a xor b);
    layer7_outputs(10200) <= a;
    layer7_outputs(10201) <= not (a and b);
    layer7_outputs(10202) <= a xor b;
    layer7_outputs(10203) <= a and not b;
    layer7_outputs(10204) <= not (a and b);
    layer7_outputs(10205) <= not a or b;
    layer7_outputs(10206) <= not a;
    layer7_outputs(10207) <= not (a xor b);
    layer7_outputs(10208) <= not a or b;
    layer7_outputs(10209) <= b;
    layer7_outputs(10210) <= a;
    layer7_outputs(10211) <= not b;
    layer7_outputs(10212) <= a or b;
    layer7_outputs(10213) <= not b;
    layer7_outputs(10214) <= not (a or b);
    layer7_outputs(10215) <= not (a or b);
    layer7_outputs(10216) <= not a;
    layer7_outputs(10217) <= not b;
    layer7_outputs(10218) <= not b or a;
    layer7_outputs(10219) <= a;
    layer7_outputs(10220) <= b;
    layer7_outputs(10221) <= not b or a;
    layer7_outputs(10222) <= not b or a;
    layer7_outputs(10223) <= b;
    layer7_outputs(10224) <= 1'b1;
    layer7_outputs(10225) <= not a;
    layer7_outputs(10226) <= not (a xor b);
    layer7_outputs(10227) <= not (a and b);
    layer7_outputs(10228) <= not (a or b);
    layer7_outputs(10229) <= not b;
    layer7_outputs(10230) <= not a;
    layer7_outputs(10231) <= not a or b;
    layer7_outputs(10232) <= a;
    layer7_outputs(10233) <= a xor b;
    layer7_outputs(10234) <= 1'b1;
    layer7_outputs(10235) <= a xor b;
    layer7_outputs(10236) <= 1'b0;
    layer7_outputs(10237) <= not a or b;
    layer7_outputs(10238) <= not a;
    layer7_outputs(10239) <= b;
    layer8_outputs(0) <= a or b;
    layer8_outputs(1) <= b;
    layer8_outputs(2) <= not b;
    layer8_outputs(3) <= not (a or b);
    layer8_outputs(4) <= b;
    layer8_outputs(5) <= a or b;
    layer8_outputs(6) <= not (a xor b);
    layer8_outputs(7) <= not a or b;
    layer8_outputs(8) <= b and not a;
    layer8_outputs(9) <= a;
    layer8_outputs(10) <= not (a or b);
    layer8_outputs(11) <= not (a xor b);
    layer8_outputs(12) <= not a or b;
    layer8_outputs(13) <= a;
    layer8_outputs(14) <= not a or b;
    layer8_outputs(15) <= not b;
    layer8_outputs(16) <= a;
    layer8_outputs(17) <= not b;
    layer8_outputs(18) <= a;
    layer8_outputs(19) <= a and b;
    layer8_outputs(20) <= 1'b0;
    layer8_outputs(21) <= a;
    layer8_outputs(22) <= a;
    layer8_outputs(23) <= a;
    layer8_outputs(24) <= not (a xor b);
    layer8_outputs(25) <= a;
    layer8_outputs(26) <= b and not a;
    layer8_outputs(27) <= a;
    layer8_outputs(28) <= not (a and b);
    layer8_outputs(29) <= not (a xor b);
    layer8_outputs(30) <= b and not a;
    layer8_outputs(31) <= not a;
    layer8_outputs(32) <= not a;
    layer8_outputs(33) <= a or b;
    layer8_outputs(34) <= not b;
    layer8_outputs(35) <= a xor b;
    layer8_outputs(36) <= not b;
    layer8_outputs(37) <= not b;
    layer8_outputs(38) <= a and not b;
    layer8_outputs(39) <= not b;
    layer8_outputs(40) <= not a;
    layer8_outputs(41) <= a or b;
    layer8_outputs(42) <= a;
    layer8_outputs(43) <= not (a xor b);
    layer8_outputs(44) <= not a or b;
    layer8_outputs(45) <= not b;
    layer8_outputs(46) <= not b;
    layer8_outputs(47) <= b and not a;
    layer8_outputs(48) <= a xor b;
    layer8_outputs(49) <= a xor b;
    layer8_outputs(50) <= not a;
    layer8_outputs(51) <= not (a or b);
    layer8_outputs(52) <= a and b;
    layer8_outputs(53) <= b and not a;
    layer8_outputs(54) <= a;
    layer8_outputs(55) <= not (a and b);
    layer8_outputs(56) <= not b;
    layer8_outputs(57) <= b;
    layer8_outputs(58) <= a;
    layer8_outputs(59) <= not (a and b);
    layer8_outputs(60) <= b;
    layer8_outputs(61) <= a and not b;
    layer8_outputs(62) <= a xor b;
    layer8_outputs(63) <= a or b;
    layer8_outputs(64) <= not a or b;
    layer8_outputs(65) <= not b;
    layer8_outputs(66) <= b;
    layer8_outputs(67) <= not (a and b);
    layer8_outputs(68) <= b;
    layer8_outputs(69) <= a xor b;
    layer8_outputs(70) <= a;
    layer8_outputs(71) <= b;
    layer8_outputs(72) <= not a or b;
    layer8_outputs(73) <= a;
    layer8_outputs(74) <= a;
    layer8_outputs(75) <= not a;
    layer8_outputs(76) <= not b;
    layer8_outputs(77) <= 1'b0;
    layer8_outputs(78) <= a xor b;
    layer8_outputs(79) <= not (a xor b);
    layer8_outputs(80) <= a xor b;
    layer8_outputs(81) <= not b;
    layer8_outputs(82) <= not b;
    layer8_outputs(83) <= not a or b;
    layer8_outputs(84) <= b;
    layer8_outputs(85) <= a xor b;
    layer8_outputs(86) <= not b;
    layer8_outputs(87) <= not (a xor b);
    layer8_outputs(88) <= not a;
    layer8_outputs(89) <= b;
    layer8_outputs(90) <= a xor b;
    layer8_outputs(91) <= not b or a;
    layer8_outputs(92) <= a and not b;
    layer8_outputs(93) <= a xor b;
    layer8_outputs(94) <= a xor b;
    layer8_outputs(95) <= not a or b;
    layer8_outputs(96) <= a xor b;
    layer8_outputs(97) <= not (a and b);
    layer8_outputs(98) <= a and not b;
    layer8_outputs(99) <= a;
    layer8_outputs(100) <= a or b;
    layer8_outputs(101) <= not (a xor b);
    layer8_outputs(102) <= not b;
    layer8_outputs(103) <= b;
    layer8_outputs(104) <= not b;
    layer8_outputs(105) <= not (a xor b);
    layer8_outputs(106) <= b and not a;
    layer8_outputs(107) <= a xor b;
    layer8_outputs(108) <= a and b;
    layer8_outputs(109) <= not (a or b);
    layer8_outputs(110) <= not (a or b);
    layer8_outputs(111) <= a and not b;
    layer8_outputs(112) <= not (a or b);
    layer8_outputs(113) <= not (a and b);
    layer8_outputs(114) <= not a;
    layer8_outputs(115) <= a;
    layer8_outputs(116) <= a or b;
    layer8_outputs(117) <= not (a xor b);
    layer8_outputs(118) <= not (a xor b);
    layer8_outputs(119) <= not (a and b);
    layer8_outputs(120) <= a and not b;
    layer8_outputs(121) <= not b;
    layer8_outputs(122) <= not a;
    layer8_outputs(123) <= a and b;
    layer8_outputs(124) <= not (a xor b);
    layer8_outputs(125) <= a or b;
    layer8_outputs(126) <= b;
    layer8_outputs(127) <= not b;
    layer8_outputs(128) <= a or b;
    layer8_outputs(129) <= b;
    layer8_outputs(130) <= a and not b;
    layer8_outputs(131) <= a;
    layer8_outputs(132) <= a or b;
    layer8_outputs(133) <= not b or a;
    layer8_outputs(134) <= b and not a;
    layer8_outputs(135) <= not b;
    layer8_outputs(136) <= b;
    layer8_outputs(137) <= not a or b;
    layer8_outputs(138) <= not b;
    layer8_outputs(139) <= not (a xor b);
    layer8_outputs(140) <= not b;
    layer8_outputs(141) <= not a;
    layer8_outputs(142) <= a;
    layer8_outputs(143) <= b;
    layer8_outputs(144) <= b;
    layer8_outputs(145) <= a or b;
    layer8_outputs(146) <= a or b;
    layer8_outputs(147) <= not (a xor b);
    layer8_outputs(148) <= a;
    layer8_outputs(149) <= a;
    layer8_outputs(150) <= not (a xor b);
    layer8_outputs(151) <= b;
    layer8_outputs(152) <= b;
    layer8_outputs(153) <= not a or b;
    layer8_outputs(154) <= not a;
    layer8_outputs(155) <= not a;
    layer8_outputs(156) <= not a;
    layer8_outputs(157) <= not b or a;
    layer8_outputs(158) <= not b;
    layer8_outputs(159) <= a and not b;
    layer8_outputs(160) <= not (a and b);
    layer8_outputs(161) <= b;
    layer8_outputs(162) <= b and not a;
    layer8_outputs(163) <= b and not a;
    layer8_outputs(164) <= a and b;
    layer8_outputs(165) <= not (a or b);
    layer8_outputs(166) <= a or b;
    layer8_outputs(167) <= not (a xor b);
    layer8_outputs(168) <= a or b;
    layer8_outputs(169) <= a xor b;
    layer8_outputs(170) <= a and b;
    layer8_outputs(171) <= a or b;
    layer8_outputs(172) <= not b;
    layer8_outputs(173) <= not (a xor b);
    layer8_outputs(174) <= a;
    layer8_outputs(175) <= a xor b;
    layer8_outputs(176) <= not (a xor b);
    layer8_outputs(177) <= not b or a;
    layer8_outputs(178) <= a and b;
    layer8_outputs(179) <= not (a xor b);
    layer8_outputs(180) <= not b;
    layer8_outputs(181) <= not (a or b);
    layer8_outputs(182) <= not b or a;
    layer8_outputs(183) <= not (a xor b);
    layer8_outputs(184) <= a or b;
    layer8_outputs(185) <= a xor b;
    layer8_outputs(186) <= 1'b0;
    layer8_outputs(187) <= a and b;
    layer8_outputs(188) <= not a;
    layer8_outputs(189) <= not (a xor b);
    layer8_outputs(190) <= a and b;
    layer8_outputs(191) <= a;
    layer8_outputs(192) <= a xor b;
    layer8_outputs(193) <= b;
    layer8_outputs(194) <= not b;
    layer8_outputs(195) <= not a;
    layer8_outputs(196) <= not (a xor b);
    layer8_outputs(197) <= not (a and b);
    layer8_outputs(198) <= a and not b;
    layer8_outputs(199) <= not a;
    layer8_outputs(200) <= a and not b;
    layer8_outputs(201) <= b and not a;
    layer8_outputs(202) <= not a or b;
    layer8_outputs(203) <= not b;
    layer8_outputs(204) <= b;
    layer8_outputs(205) <= not (a or b);
    layer8_outputs(206) <= a and b;
    layer8_outputs(207) <= not (a or b);
    layer8_outputs(208) <= not b;
    layer8_outputs(209) <= not (a or b);
    layer8_outputs(210) <= a or b;
    layer8_outputs(211) <= a and b;
    layer8_outputs(212) <= a or b;
    layer8_outputs(213) <= not b;
    layer8_outputs(214) <= b;
    layer8_outputs(215) <= b and not a;
    layer8_outputs(216) <= not b;
    layer8_outputs(217) <= not a;
    layer8_outputs(218) <= not b;
    layer8_outputs(219) <= b;
    layer8_outputs(220) <= not a or b;
    layer8_outputs(221) <= b and not a;
    layer8_outputs(222) <= not (a xor b);
    layer8_outputs(223) <= a;
    layer8_outputs(224) <= b;
    layer8_outputs(225) <= not a;
    layer8_outputs(226) <= a xor b;
    layer8_outputs(227) <= a;
    layer8_outputs(228) <= b;
    layer8_outputs(229) <= not (a or b);
    layer8_outputs(230) <= a xor b;
    layer8_outputs(231) <= a or b;
    layer8_outputs(232) <= b;
    layer8_outputs(233) <= a;
    layer8_outputs(234) <= not (a xor b);
    layer8_outputs(235) <= b and not a;
    layer8_outputs(236) <= 1'b1;
    layer8_outputs(237) <= not a;
    layer8_outputs(238) <= a or b;
    layer8_outputs(239) <= not a or b;
    layer8_outputs(240) <= b;
    layer8_outputs(241) <= a;
    layer8_outputs(242) <= not b;
    layer8_outputs(243) <= a;
    layer8_outputs(244) <= a xor b;
    layer8_outputs(245) <= not (a xor b);
    layer8_outputs(246) <= not (a and b);
    layer8_outputs(247) <= not (a xor b);
    layer8_outputs(248) <= not (a xor b);
    layer8_outputs(249) <= a xor b;
    layer8_outputs(250) <= b and not a;
    layer8_outputs(251) <= not (a xor b);
    layer8_outputs(252) <= a xor b;
    layer8_outputs(253) <= not (a xor b);
    layer8_outputs(254) <= not a;
    layer8_outputs(255) <= not a;
    layer8_outputs(256) <= not a;
    layer8_outputs(257) <= not b or a;
    layer8_outputs(258) <= not (a xor b);
    layer8_outputs(259) <= not b or a;
    layer8_outputs(260) <= not (a and b);
    layer8_outputs(261) <= not a or b;
    layer8_outputs(262) <= not (a or b);
    layer8_outputs(263) <= a and not b;
    layer8_outputs(264) <= a xor b;
    layer8_outputs(265) <= not a or b;
    layer8_outputs(266) <= not b or a;
    layer8_outputs(267) <= b;
    layer8_outputs(268) <= not b;
    layer8_outputs(269) <= a xor b;
    layer8_outputs(270) <= a xor b;
    layer8_outputs(271) <= not (a or b);
    layer8_outputs(272) <= not b;
    layer8_outputs(273) <= not (a and b);
    layer8_outputs(274) <= a;
    layer8_outputs(275) <= not (a and b);
    layer8_outputs(276) <= a;
    layer8_outputs(277) <= not a or b;
    layer8_outputs(278) <= not (a xor b);
    layer8_outputs(279) <= 1'b1;
    layer8_outputs(280) <= not (a xor b);
    layer8_outputs(281) <= not b or a;
    layer8_outputs(282) <= not b;
    layer8_outputs(283) <= not a or b;
    layer8_outputs(284) <= not (a or b);
    layer8_outputs(285) <= b;
    layer8_outputs(286) <= a or b;
    layer8_outputs(287) <= a xor b;
    layer8_outputs(288) <= not a;
    layer8_outputs(289) <= not a;
    layer8_outputs(290) <= not b;
    layer8_outputs(291) <= not (a xor b);
    layer8_outputs(292) <= not (a and b);
    layer8_outputs(293) <= not a or b;
    layer8_outputs(294) <= not (a or b);
    layer8_outputs(295) <= not b;
    layer8_outputs(296) <= not (a xor b);
    layer8_outputs(297) <= not a;
    layer8_outputs(298) <= not (a or b);
    layer8_outputs(299) <= a xor b;
    layer8_outputs(300) <= a and not b;
    layer8_outputs(301) <= a;
    layer8_outputs(302) <= a;
    layer8_outputs(303) <= b;
    layer8_outputs(304) <= not a;
    layer8_outputs(305) <= not (a xor b);
    layer8_outputs(306) <= a;
    layer8_outputs(307) <= a;
    layer8_outputs(308) <= not b;
    layer8_outputs(309) <= not b;
    layer8_outputs(310) <= a and not b;
    layer8_outputs(311) <= not a;
    layer8_outputs(312) <= not a;
    layer8_outputs(313) <= not b;
    layer8_outputs(314) <= a and b;
    layer8_outputs(315) <= not b or a;
    layer8_outputs(316) <= not (a or b);
    layer8_outputs(317) <= a xor b;
    layer8_outputs(318) <= not (a xor b);
    layer8_outputs(319) <= a and not b;
    layer8_outputs(320) <= a and not b;
    layer8_outputs(321) <= a or b;
    layer8_outputs(322) <= not b;
    layer8_outputs(323) <= a;
    layer8_outputs(324) <= not a;
    layer8_outputs(325) <= not (a or b);
    layer8_outputs(326) <= a xor b;
    layer8_outputs(327) <= a and b;
    layer8_outputs(328) <= not b;
    layer8_outputs(329) <= a and not b;
    layer8_outputs(330) <= not (a xor b);
    layer8_outputs(331) <= not (a and b);
    layer8_outputs(332) <= b;
    layer8_outputs(333) <= a xor b;
    layer8_outputs(334) <= not (a xor b);
    layer8_outputs(335) <= a;
    layer8_outputs(336) <= b;
    layer8_outputs(337) <= a;
    layer8_outputs(338) <= not (a and b);
    layer8_outputs(339) <= a;
    layer8_outputs(340) <= not b;
    layer8_outputs(341) <= b and not a;
    layer8_outputs(342) <= not (a xor b);
    layer8_outputs(343) <= b;
    layer8_outputs(344) <= a xor b;
    layer8_outputs(345) <= not (a xor b);
    layer8_outputs(346) <= a;
    layer8_outputs(347) <= a;
    layer8_outputs(348) <= a;
    layer8_outputs(349) <= not b;
    layer8_outputs(350) <= a;
    layer8_outputs(351) <= a xor b;
    layer8_outputs(352) <= a and not b;
    layer8_outputs(353) <= not a;
    layer8_outputs(354) <= a and not b;
    layer8_outputs(355) <= a;
    layer8_outputs(356) <= not (a xor b);
    layer8_outputs(357) <= a;
    layer8_outputs(358) <= not b;
    layer8_outputs(359) <= not a;
    layer8_outputs(360) <= b;
    layer8_outputs(361) <= b;
    layer8_outputs(362) <= a;
    layer8_outputs(363) <= a and not b;
    layer8_outputs(364) <= a xor b;
    layer8_outputs(365) <= b;
    layer8_outputs(366) <= not b;
    layer8_outputs(367) <= b;
    layer8_outputs(368) <= a and not b;
    layer8_outputs(369) <= not (a xor b);
    layer8_outputs(370) <= not a;
    layer8_outputs(371) <= a;
    layer8_outputs(372) <= not (a xor b);
    layer8_outputs(373) <= a or b;
    layer8_outputs(374) <= not (a and b);
    layer8_outputs(375) <= not a or b;
    layer8_outputs(376) <= not a;
    layer8_outputs(377) <= not b or a;
    layer8_outputs(378) <= b;
    layer8_outputs(379) <= b;
    layer8_outputs(380) <= b;
    layer8_outputs(381) <= b and not a;
    layer8_outputs(382) <= a and not b;
    layer8_outputs(383) <= not a;
    layer8_outputs(384) <= not (a and b);
    layer8_outputs(385) <= a or b;
    layer8_outputs(386) <= not a or b;
    layer8_outputs(387) <= not a;
    layer8_outputs(388) <= not a;
    layer8_outputs(389) <= not a;
    layer8_outputs(390) <= not b;
    layer8_outputs(391) <= b;
    layer8_outputs(392) <= not (a xor b);
    layer8_outputs(393) <= not b;
    layer8_outputs(394) <= a xor b;
    layer8_outputs(395) <= a;
    layer8_outputs(396) <= not a or b;
    layer8_outputs(397) <= not (a or b);
    layer8_outputs(398) <= not (a or b);
    layer8_outputs(399) <= a and not b;
    layer8_outputs(400) <= not (a xor b);
    layer8_outputs(401) <= not b;
    layer8_outputs(402) <= not (a xor b);
    layer8_outputs(403) <= a;
    layer8_outputs(404) <= not b or a;
    layer8_outputs(405) <= not (a or b);
    layer8_outputs(406) <= not (a and b);
    layer8_outputs(407) <= a xor b;
    layer8_outputs(408) <= a xor b;
    layer8_outputs(409) <= not (a xor b);
    layer8_outputs(410) <= a or b;
    layer8_outputs(411) <= b;
    layer8_outputs(412) <= not (a xor b);
    layer8_outputs(413) <= not (a and b);
    layer8_outputs(414) <= a xor b;
    layer8_outputs(415) <= a and b;
    layer8_outputs(416) <= not (a xor b);
    layer8_outputs(417) <= not a;
    layer8_outputs(418) <= not a or b;
    layer8_outputs(419) <= not b;
    layer8_outputs(420) <= not a;
    layer8_outputs(421) <= not a;
    layer8_outputs(422) <= not a or b;
    layer8_outputs(423) <= b and not a;
    layer8_outputs(424) <= a;
    layer8_outputs(425) <= not (a xor b);
    layer8_outputs(426) <= b;
    layer8_outputs(427) <= a and not b;
    layer8_outputs(428) <= not (a and b);
    layer8_outputs(429) <= a and not b;
    layer8_outputs(430) <= not (a or b);
    layer8_outputs(431) <= not a;
    layer8_outputs(432) <= b;
    layer8_outputs(433) <= not b or a;
    layer8_outputs(434) <= not b;
    layer8_outputs(435) <= not (a and b);
    layer8_outputs(436) <= a;
    layer8_outputs(437) <= a and b;
    layer8_outputs(438) <= not a or b;
    layer8_outputs(439) <= a xor b;
    layer8_outputs(440) <= b;
    layer8_outputs(441) <= a and not b;
    layer8_outputs(442) <= b;
    layer8_outputs(443) <= a and b;
    layer8_outputs(444) <= not (a xor b);
    layer8_outputs(445) <= b;
    layer8_outputs(446) <= not (a or b);
    layer8_outputs(447) <= a;
    layer8_outputs(448) <= not b or a;
    layer8_outputs(449) <= not (a xor b);
    layer8_outputs(450) <= a xor b;
    layer8_outputs(451) <= not b;
    layer8_outputs(452) <= not (a xor b);
    layer8_outputs(453) <= a or b;
    layer8_outputs(454) <= a and not b;
    layer8_outputs(455) <= a;
    layer8_outputs(456) <= not (a or b);
    layer8_outputs(457) <= not a or b;
    layer8_outputs(458) <= a xor b;
    layer8_outputs(459) <= b and not a;
    layer8_outputs(460) <= a xor b;
    layer8_outputs(461) <= a or b;
    layer8_outputs(462) <= b and not a;
    layer8_outputs(463) <= not (a xor b);
    layer8_outputs(464) <= not (a xor b);
    layer8_outputs(465) <= a or b;
    layer8_outputs(466) <= a;
    layer8_outputs(467) <= not a or b;
    layer8_outputs(468) <= not b;
    layer8_outputs(469) <= not (a or b);
    layer8_outputs(470) <= a and not b;
    layer8_outputs(471) <= not (a xor b);
    layer8_outputs(472) <= b;
    layer8_outputs(473) <= not (a xor b);
    layer8_outputs(474) <= not a;
    layer8_outputs(475) <= not a;
    layer8_outputs(476) <= a;
    layer8_outputs(477) <= a xor b;
    layer8_outputs(478) <= not (a xor b);
    layer8_outputs(479) <= a or b;
    layer8_outputs(480) <= not a;
    layer8_outputs(481) <= not (a and b);
    layer8_outputs(482) <= a;
    layer8_outputs(483) <= a xor b;
    layer8_outputs(484) <= not (a xor b);
    layer8_outputs(485) <= a xor b;
    layer8_outputs(486) <= not (a and b);
    layer8_outputs(487) <= not a;
    layer8_outputs(488) <= not (a xor b);
    layer8_outputs(489) <= a and b;
    layer8_outputs(490) <= a xor b;
    layer8_outputs(491) <= not b;
    layer8_outputs(492) <= not (a or b);
    layer8_outputs(493) <= a or b;
    layer8_outputs(494) <= b;
    layer8_outputs(495) <= a;
    layer8_outputs(496) <= not a;
    layer8_outputs(497) <= a xor b;
    layer8_outputs(498) <= a xor b;
    layer8_outputs(499) <= not (a and b);
    layer8_outputs(500) <= not (a xor b);
    layer8_outputs(501) <= b;
    layer8_outputs(502) <= not (a xor b);
    layer8_outputs(503) <= not a;
    layer8_outputs(504) <= not (a and b);
    layer8_outputs(505) <= not (a xor b);
    layer8_outputs(506) <= not b;
    layer8_outputs(507) <= not (a and b);
    layer8_outputs(508) <= not (a or b);
    layer8_outputs(509) <= not (a or b);
    layer8_outputs(510) <= not a;
    layer8_outputs(511) <= not (a xor b);
    layer8_outputs(512) <= b;
    layer8_outputs(513) <= a and not b;
    layer8_outputs(514) <= b;
    layer8_outputs(515) <= b and not a;
    layer8_outputs(516) <= not b;
    layer8_outputs(517) <= a xor b;
    layer8_outputs(518) <= b and not a;
    layer8_outputs(519) <= a xor b;
    layer8_outputs(520) <= not (a xor b);
    layer8_outputs(521) <= not a or b;
    layer8_outputs(522) <= a xor b;
    layer8_outputs(523) <= not b;
    layer8_outputs(524) <= b;
    layer8_outputs(525) <= a and not b;
    layer8_outputs(526) <= a;
    layer8_outputs(527) <= b and not a;
    layer8_outputs(528) <= not a or b;
    layer8_outputs(529) <= b and not a;
    layer8_outputs(530) <= not a;
    layer8_outputs(531) <= b and not a;
    layer8_outputs(532) <= b;
    layer8_outputs(533) <= not (a and b);
    layer8_outputs(534) <= not b;
    layer8_outputs(535) <= not a or b;
    layer8_outputs(536) <= not a;
    layer8_outputs(537) <= not (a xor b);
    layer8_outputs(538) <= not (a xor b);
    layer8_outputs(539) <= a;
    layer8_outputs(540) <= not (a or b);
    layer8_outputs(541) <= not (a xor b);
    layer8_outputs(542) <= not a;
    layer8_outputs(543) <= b;
    layer8_outputs(544) <= not b;
    layer8_outputs(545) <= a;
    layer8_outputs(546) <= a and not b;
    layer8_outputs(547) <= not a or b;
    layer8_outputs(548) <= not b;
    layer8_outputs(549) <= not (a xor b);
    layer8_outputs(550) <= not a or b;
    layer8_outputs(551) <= not a or b;
    layer8_outputs(552) <= a;
    layer8_outputs(553) <= not a or b;
    layer8_outputs(554) <= a xor b;
    layer8_outputs(555) <= b;
    layer8_outputs(556) <= a;
    layer8_outputs(557) <= not (a or b);
    layer8_outputs(558) <= not a;
    layer8_outputs(559) <= not (a xor b);
    layer8_outputs(560) <= not a or b;
    layer8_outputs(561) <= not (a xor b);
    layer8_outputs(562) <= not b or a;
    layer8_outputs(563) <= a and b;
    layer8_outputs(564) <= b;
    layer8_outputs(565) <= not (a and b);
    layer8_outputs(566) <= not b or a;
    layer8_outputs(567) <= a;
    layer8_outputs(568) <= not b;
    layer8_outputs(569) <= not a;
    layer8_outputs(570) <= not (a and b);
    layer8_outputs(571) <= not a;
    layer8_outputs(572) <= a;
    layer8_outputs(573) <= not (a or b);
    layer8_outputs(574) <= b;
    layer8_outputs(575) <= a xor b;
    layer8_outputs(576) <= b;
    layer8_outputs(577) <= not b;
    layer8_outputs(578) <= not a;
    layer8_outputs(579) <= a xor b;
    layer8_outputs(580) <= not b;
    layer8_outputs(581) <= a and not b;
    layer8_outputs(582) <= a or b;
    layer8_outputs(583) <= not a;
    layer8_outputs(584) <= a xor b;
    layer8_outputs(585) <= not (a or b);
    layer8_outputs(586) <= not a;
    layer8_outputs(587) <= not b or a;
    layer8_outputs(588) <= not (a or b);
    layer8_outputs(589) <= a;
    layer8_outputs(590) <= not a or b;
    layer8_outputs(591) <= a;
    layer8_outputs(592) <= a and not b;
    layer8_outputs(593) <= b;
    layer8_outputs(594) <= not (a and b);
    layer8_outputs(595) <= b;
    layer8_outputs(596) <= a and b;
    layer8_outputs(597) <= b and not a;
    layer8_outputs(598) <= a;
    layer8_outputs(599) <= a xor b;
    layer8_outputs(600) <= not (a xor b);
    layer8_outputs(601) <= not b or a;
    layer8_outputs(602) <= 1'b0;
    layer8_outputs(603) <= not a;
    layer8_outputs(604) <= not (a xor b);
    layer8_outputs(605) <= a;
    layer8_outputs(606) <= not (a and b);
    layer8_outputs(607) <= not b;
    layer8_outputs(608) <= a or b;
    layer8_outputs(609) <= a xor b;
    layer8_outputs(610) <= not b;
    layer8_outputs(611) <= not (a xor b);
    layer8_outputs(612) <= a or b;
    layer8_outputs(613) <= not a or b;
    layer8_outputs(614) <= b;
    layer8_outputs(615) <= not (a xor b);
    layer8_outputs(616) <= a or b;
    layer8_outputs(617) <= not (a or b);
    layer8_outputs(618) <= not b;
    layer8_outputs(619) <= not (a and b);
    layer8_outputs(620) <= a xor b;
    layer8_outputs(621) <= not (a xor b);
    layer8_outputs(622) <= not b;
    layer8_outputs(623) <= not a or b;
    layer8_outputs(624) <= not a;
    layer8_outputs(625) <= b;
    layer8_outputs(626) <= a and b;
    layer8_outputs(627) <= not a;
    layer8_outputs(628) <= a xor b;
    layer8_outputs(629) <= b and not a;
    layer8_outputs(630) <= a and b;
    layer8_outputs(631) <= not (a xor b);
    layer8_outputs(632) <= a;
    layer8_outputs(633) <= not a;
    layer8_outputs(634) <= b and not a;
    layer8_outputs(635) <= b;
    layer8_outputs(636) <= a xor b;
    layer8_outputs(637) <= a xor b;
    layer8_outputs(638) <= not b or a;
    layer8_outputs(639) <= a or b;
    layer8_outputs(640) <= b;
    layer8_outputs(641) <= b;
    layer8_outputs(642) <= not a or b;
    layer8_outputs(643) <= a or b;
    layer8_outputs(644) <= a;
    layer8_outputs(645) <= not (a xor b);
    layer8_outputs(646) <= b;
    layer8_outputs(647) <= b and not a;
    layer8_outputs(648) <= not a;
    layer8_outputs(649) <= not b;
    layer8_outputs(650) <= not (a xor b);
    layer8_outputs(651) <= not a;
    layer8_outputs(652) <= b;
    layer8_outputs(653) <= b and not a;
    layer8_outputs(654) <= not a;
    layer8_outputs(655) <= b;
    layer8_outputs(656) <= b and not a;
    layer8_outputs(657) <= b;
    layer8_outputs(658) <= 1'b0;
    layer8_outputs(659) <= not (a xor b);
    layer8_outputs(660) <= a and b;
    layer8_outputs(661) <= not a;
    layer8_outputs(662) <= b;
    layer8_outputs(663) <= not b or a;
    layer8_outputs(664) <= a;
    layer8_outputs(665) <= a and not b;
    layer8_outputs(666) <= not a;
    layer8_outputs(667) <= a or b;
    layer8_outputs(668) <= not (a xor b);
    layer8_outputs(669) <= b;
    layer8_outputs(670) <= not (a xor b);
    layer8_outputs(671) <= b;
    layer8_outputs(672) <= b;
    layer8_outputs(673) <= b;
    layer8_outputs(674) <= a xor b;
    layer8_outputs(675) <= b;
    layer8_outputs(676) <= not a or b;
    layer8_outputs(677) <= a;
    layer8_outputs(678) <= a;
    layer8_outputs(679) <= not a;
    layer8_outputs(680) <= not (a xor b);
    layer8_outputs(681) <= not b;
    layer8_outputs(682) <= b;
    layer8_outputs(683) <= not b;
    layer8_outputs(684) <= not a;
    layer8_outputs(685) <= a and b;
    layer8_outputs(686) <= b;
    layer8_outputs(687) <= not (a and b);
    layer8_outputs(688) <= a and not b;
    layer8_outputs(689) <= b;
    layer8_outputs(690) <= not b;
    layer8_outputs(691) <= b and not a;
    layer8_outputs(692) <= not a;
    layer8_outputs(693) <= not (a xor b);
    layer8_outputs(694) <= a and b;
    layer8_outputs(695) <= a and not b;
    layer8_outputs(696) <= not b;
    layer8_outputs(697) <= not (a or b);
    layer8_outputs(698) <= a;
    layer8_outputs(699) <= not a;
    layer8_outputs(700) <= a and b;
    layer8_outputs(701) <= b;
    layer8_outputs(702) <= not (a and b);
    layer8_outputs(703) <= not a;
    layer8_outputs(704) <= b and not a;
    layer8_outputs(705) <= a;
    layer8_outputs(706) <= not (a and b);
    layer8_outputs(707) <= a xor b;
    layer8_outputs(708) <= a xor b;
    layer8_outputs(709) <= not a;
    layer8_outputs(710) <= b and not a;
    layer8_outputs(711) <= a xor b;
    layer8_outputs(712) <= a;
    layer8_outputs(713) <= not a;
    layer8_outputs(714) <= not a;
    layer8_outputs(715) <= a xor b;
    layer8_outputs(716) <= b;
    layer8_outputs(717) <= not (a xor b);
    layer8_outputs(718) <= not (a xor b);
    layer8_outputs(719) <= b;
    layer8_outputs(720) <= a and not b;
    layer8_outputs(721) <= not b;
    layer8_outputs(722) <= a;
    layer8_outputs(723) <= not a;
    layer8_outputs(724) <= 1'b1;
    layer8_outputs(725) <= not (a xor b);
    layer8_outputs(726) <= not b;
    layer8_outputs(727) <= not (a xor b);
    layer8_outputs(728) <= not b or a;
    layer8_outputs(729) <= not (a xor b);
    layer8_outputs(730) <= a xor b;
    layer8_outputs(731) <= not a;
    layer8_outputs(732) <= a;
    layer8_outputs(733) <= not b or a;
    layer8_outputs(734) <= not a;
    layer8_outputs(735) <= a xor b;
    layer8_outputs(736) <= not (a or b);
    layer8_outputs(737) <= a and not b;
    layer8_outputs(738) <= b;
    layer8_outputs(739) <= not b;
    layer8_outputs(740) <= b;
    layer8_outputs(741) <= a xor b;
    layer8_outputs(742) <= not a;
    layer8_outputs(743) <= a;
    layer8_outputs(744) <= not b;
    layer8_outputs(745) <= b;
    layer8_outputs(746) <= not (a or b);
    layer8_outputs(747) <= b;
    layer8_outputs(748) <= b;
    layer8_outputs(749) <= a;
    layer8_outputs(750) <= a or b;
    layer8_outputs(751) <= a and not b;
    layer8_outputs(752) <= a and not b;
    layer8_outputs(753) <= not a;
    layer8_outputs(754) <= a xor b;
    layer8_outputs(755) <= not b;
    layer8_outputs(756) <= not a;
    layer8_outputs(757) <= not b;
    layer8_outputs(758) <= not b;
    layer8_outputs(759) <= not b;
    layer8_outputs(760) <= not a or b;
    layer8_outputs(761) <= a xor b;
    layer8_outputs(762) <= not (a xor b);
    layer8_outputs(763) <= a;
    layer8_outputs(764) <= b;
    layer8_outputs(765) <= not a;
    layer8_outputs(766) <= b and not a;
    layer8_outputs(767) <= not a;
    layer8_outputs(768) <= b and not a;
    layer8_outputs(769) <= not b;
    layer8_outputs(770) <= not (a or b);
    layer8_outputs(771) <= not b;
    layer8_outputs(772) <= 1'b0;
    layer8_outputs(773) <= not (a xor b);
    layer8_outputs(774) <= a and b;
    layer8_outputs(775) <= not b;
    layer8_outputs(776) <= a xor b;
    layer8_outputs(777) <= a xor b;
    layer8_outputs(778) <= not a;
    layer8_outputs(779) <= b and not a;
    layer8_outputs(780) <= not (a and b);
    layer8_outputs(781) <= not (a xor b);
    layer8_outputs(782) <= a xor b;
    layer8_outputs(783) <= b;
    layer8_outputs(784) <= not a or b;
    layer8_outputs(785) <= a xor b;
    layer8_outputs(786) <= b;
    layer8_outputs(787) <= not b;
    layer8_outputs(788) <= b;
    layer8_outputs(789) <= a xor b;
    layer8_outputs(790) <= not (a and b);
    layer8_outputs(791) <= not (a or b);
    layer8_outputs(792) <= not (a or b);
    layer8_outputs(793) <= a xor b;
    layer8_outputs(794) <= a;
    layer8_outputs(795) <= not b;
    layer8_outputs(796) <= b;
    layer8_outputs(797) <= a and b;
    layer8_outputs(798) <= a and not b;
    layer8_outputs(799) <= not a;
    layer8_outputs(800) <= a and b;
    layer8_outputs(801) <= not (a or b);
    layer8_outputs(802) <= a;
    layer8_outputs(803) <= not b;
    layer8_outputs(804) <= b and not a;
    layer8_outputs(805) <= not a;
    layer8_outputs(806) <= a;
    layer8_outputs(807) <= a xor b;
    layer8_outputs(808) <= not (a or b);
    layer8_outputs(809) <= not (a xor b);
    layer8_outputs(810) <= b;
    layer8_outputs(811) <= a and b;
    layer8_outputs(812) <= not a;
    layer8_outputs(813) <= a and b;
    layer8_outputs(814) <= not (a xor b);
    layer8_outputs(815) <= not b or a;
    layer8_outputs(816) <= a;
    layer8_outputs(817) <= b;
    layer8_outputs(818) <= a;
    layer8_outputs(819) <= not (a xor b);
    layer8_outputs(820) <= not b;
    layer8_outputs(821) <= b;
    layer8_outputs(822) <= not b or a;
    layer8_outputs(823) <= not b;
    layer8_outputs(824) <= b;
    layer8_outputs(825) <= a;
    layer8_outputs(826) <= not b;
    layer8_outputs(827) <= b;
    layer8_outputs(828) <= not b or a;
    layer8_outputs(829) <= not (a xor b);
    layer8_outputs(830) <= not a or b;
    layer8_outputs(831) <= a xor b;
    layer8_outputs(832) <= not b;
    layer8_outputs(833) <= not b;
    layer8_outputs(834) <= not (a xor b);
    layer8_outputs(835) <= a and b;
    layer8_outputs(836) <= a and b;
    layer8_outputs(837) <= a xor b;
    layer8_outputs(838) <= a;
    layer8_outputs(839) <= b;
    layer8_outputs(840) <= a and not b;
    layer8_outputs(841) <= a xor b;
    layer8_outputs(842) <= a xor b;
    layer8_outputs(843) <= not a;
    layer8_outputs(844) <= not (a xor b);
    layer8_outputs(845) <= b and not a;
    layer8_outputs(846) <= not a;
    layer8_outputs(847) <= not b;
    layer8_outputs(848) <= a;
    layer8_outputs(849) <= a and b;
    layer8_outputs(850) <= a xor b;
    layer8_outputs(851) <= not b;
    layer8_outputs(852) <= a xor b;
    layer8_outputs(853) <= a;
    layer8_outputs(854) <= a and b;
    layer8_outputs(855) <= not b or a;
    layer8_outputs(856) <= a xor b;
    layer8_outputs(857) <= a and not b;
    layer8_outputs(858) <= not a or b;
    layer8_outputs(859) <= a or b;
    layer8_outputs(860) <= not a;
    layer8_outputs(861) <= a xor b;
    layer8_outputs(862) <= a;
    layer8_outputs(863) <= not a;
    layer8_outputs(864) <= a xor b;
    layer8_outputs(865) <= not a or b;
    layer8_outputs(866) <= 1'b0;
    layer8_outputs(867) <= a;
    layer8_outputs(868) <= a and b;
    layer8_outputs(869) <= not a;
    layer8_outputs(870) <= not a;
    layer8_outputs(871) <= a or b;
    layer8_outputs(872) <= a and b;
    layer8_outputs(873) <= not (a xor b);
    layer8_outputs(874) <= a;
    layer8_outputs(875) <= a;
    layer8_outputs(876) <= not a;
    layer8_outputs(877) <= not b;
    layer8_outputs(878) <= not (a xor b);
    layer8_outputs(879) <= b;
    layer8_outputs(880) <= a xor b;
    layer8_outputs(881) <= b;
    layer8_outputs(882) <= not a;
    layer8_outputs(883) <= a;
    layer8_outputs(884) <= b;
    layer8_outputs(885) <= not a or b;
    layer8_outputs(886) <= a xor b;
    layer8_outputs(887) <= not a;
    layer8_outputs(888) <= a xor b;
    layer8_outputs(889) <= not (a or b);
    layer8_outputs(890) <= not a;
    layer8_outputs(891) <= b;
    layer8_outputs(892) <= a and not b;
    layer8_outputs(893) <= a;
    layer8_outputs(894) <= not b;
    layer8_outputs(895) <= not b;
    layer8_outputs(896) <= not (a xor b);
    layer8_outputs(897) <= a xor b;
    layer8_outputs(898) <= a and not b;
    layer8_outputs(899) <= a or b;
    layer8_outputs(900) <= b;
    layer8_outputs(901) <= a xor b;
    layer8_outputs(902) <= b;
    layer8_outputs(903) <= a and not b;
    layer8_outputs(904) <= b;
    layer8_outputs(905) <= b;
    layer8_outputs(906) <= b and not a;
    layer8_outputs(907) <= b;
    layer8_outputs(908) <= not a;
    layer8_outputs(909) <= b;
    layer8_outputs(910) <= b;
    layer8_outputs(911) <= a and not b;
    layer8_outputs(912) <= a xor b;
    layer8_outputs(913) <= a or b;
    layer8_outputs(914) <= b;
    layer8_outputs(915) <= not a;
    layer8_outputs(916) <= a;
    layer8_outputs(917) <= b;
    layer8_outputs(918) <= not b;
    layer8_outputs(919) <= not b;
    layer8_outputs(920) <= b and not a;
    layer8_outputs(921) <= not a;
    layer8_outputs(922) <= not a;
    layer8_outputs(923) <= not a or b;
    layer8_outputs(924) <= a;
    layer8_outputs(925) <= b;
    layer8_outputs(926) <= b;
    layer8_outputs(927) <= a and not b;
    layer8_outputs(928) <= not b or a;
    layer8_outputs(929) <= a and b;
    layer8_outputs(930) <= a;
    layer8_outputs(931) <= not (a xor b);
    layer8_outputs(932) <= not b;
    layer8_outputs(933) <= not (a or b);
    layer8_outputs(934) <= not (a xor b);
    layer8_outputs(935) <= a and not b;
    layer8_outputs(936) <= a;
    layer8_outputs(937) <= not a;
    layer8_outputs(938) <= a or b;
    layer8_outputs(939) <= a;
    layer8_outputs(940) <= not (a xor b);
    layer8_outputs(941) <= not a or b;
    layer8_outputs(942) <= not b;
    layer8_outputs(943) <= not (a xor b);
    layer8_outputs(944) <= not b or a;
    layer8_outputs(945) <= not b;
    layer8_outputs(946) <= a and b;
    layer8_outputs(947) <= not a;
    layer8_outputs(948) <= not b;
    layer8_outputs(949) <= not b;
    layer8_outputs(950) <= not b;
    layer8_outputs(951) <= a and b;
    layer8_outputs(952) <= a and b;
    layer8_outputs(953) <= a xor b;
    layer8_outputs(954) <= not b;
    layer8_outputs(955) <= not a or b;
    layer8_outputs(956) <= a xor b;
    layer8_outputs(957) <= not a;
    layer8_outputs(958) <= a xor b;
    layer8_outputs(959) <= a xor b;
    layer8_outputs(960) <= 1'b1;
    layer8_outputs(961) <= a and b;
    layer8_outputs(962) <= a xor b;
    layer8_outputs(963) <= b and not a;
    layer8_outputs(964) <= a or b;
    layer8_outputs(965) <= not (a and b);
    layer8_outputs(966) <= b;
    layer8_outputs(967) <= not (a xor b);
    layer8_outputs(968) <= not (a and b);
    layer8_outputs(969) <= a or b;
    layer8_outputs(970) <= a xor b;
    layer8_outputs(971) <= b;
    layer8_outputs(972) <= not b;
    layer8_outputs(973) <= not (a xor b);
    layer8_outputs(974) <= a;
    layer8_outputs(975) <= not a;
    layer8_outputs(976) <= not (a xor b);
    layer8_outputs(977) <= not b;
    layer8_outputs(978) <= a and b;
    layer8_outputs(979) <= not a or b;
    layer8_outputs(980) <= not (a xor b);
    layer8_outputs(981) <= not b;
    layer8_outputs(982) <= not b;
    layer8_outputs(983) <= a xor b;
    layer8_outputs(984) <= not b;
    layer8_outputs(985) <= a and b;
    layer8_outputs(986) <= a;
    layer8_outputs(987) <= a or b;
    layer8_outputs(988) <= not a or b;
    layer8_outputs(989) <= not a or b;
    layer8_outputs(990) <= b;
    layer8_outputs(991) <= not a;
    layer8_outputs(992) <= 1'b0;
    layer8_outputs(993) <= a xor b;
    layer8_outputs(994) <= not a;
    layer8_outputs(995) <= not (a xor b);
    layer8_outputs(996) <= not a or b;
    layer8_outputs(997) <= b and not a;
    layer8_outputs(998) <= a xor b;
    layer8_outputs(999) <= not b or a;
    layer8_outputs(1000) <= 1'b1;
    layer8_outputs(1001) <= a xor b;
    layer8_outputs(1002) <= not a;
    layer8_outputs(1003) <= b;
    layer8_outputs(1004) <= not b or a;
    layer8_outputs(1005) <= b;
    layer8_outputs(1006) <= not a;
    layer8_outputs(1007) <= not b;
    layer8_outputs(1008) <= a xor b;
    layer8_outputs(1009) <= not a;
    layer8_outputs(1010) <= not (a or b);
    layer8_outputs(1011) <= a xor b;
    layer8_outputs(1012) <= not a;
    layer8_outputs(1013) <= 1'b1;
    layer8_outputs(1014) <= not a;
    layer8_outputs(1015) <= b;
    layer8_outputs(1016) <= not (a xor b);
    layer8_outputs(1017) <= a xor b;
    layer8_outputs(1018) <= a xor b;
    layer8_outputs(1019) <= b;
    layer8_outputs(1020) <= not a or b;
    layer8_outputs(1021) <= a xor b;
    layer8_outputs(1022) <= a and not b;
    layer8_outputs(1023) <= not (a xor b);
    layer8_outputs(1024) <= b and not a;
    layer8_outputs(1025) <= a;
    layer8_outputs(1026) <= not (a and b);
    layer8_outputs(1027) <= a;
    layer8_outputs(1028) <= a or b;
    layer8_outputs(1029) <= a or b;
    layer8_outputs(1030) <= a;
    layer8_outputs(1031) <= not (a and b);
    layer8_outputs(1032) <= b;
    layer8_outputs(1033) <= b;
    layer8_outputs(1034) <= 1'b1;
    layer8_outputs(1035) <= a and b;
    layer8_outputs(1036) <= not (a xor b);
    layer8_outputs(1037) <= not a;
    layer8_outputs(1038) <= b;
    layer8_outputs(1039) <= b and not a;
    layer8_outputs(1040) <= not b;
    layer8_outputs(1041) <= not b;
    layer8_outputs(1042) <= a and b;
    layer8_outputs(1043) <= a;
    layer8_outputs(1044) <= a xor b;
    layer8_outputs(1045) <= not a or b;
    layer8_outputs(1046) <= not a;
    layer8_outputs(1047) <= a and not b;
    layer8_outputs(1048) <= b;
    layer8_outputs(1049) <= not a;
    layer8_outputs(1050) <= a;
    layer8_outputs(1051) <= a;
    layer8_outputs(1052) <= a or b;
    layer8_outputs(1053) <= not b;
    layer8_outputs(1054) <= a xor b;
    layer8_outputs(1055) <= not a;
    layer8_outputs(1056) <= a and b;
    layer8_outputs(1057) <= not (a xor b);
    layer8_outputs(1058) <= not a;
    layer8_outputs(1059) <= b;
    layer8_outputs(1060) <= a and b;
    layer8_outputs(1061) <= a and not b;
    layer8_outputs(1062) <= not a;
    layer8_outputs(1063) <= not (a xor b);
    layer8_outputs(1064) <= not (a or b);
    layer8_outputs(1065) <= a xor b;
    layer8_outputs(1066) <= not a;
    layer8_outputs(1067) <= a or b;
    layer8_outputs(1068) <= not a;
    layer8_outputs(1069) <= a xor b;
    layer8_outputs(1070) <= not (a xor b);
    layer8_outputs(1071) <= not b;
    layer8_outputs(1072) <= not a;
    layer8_outputs(1073) <= not b;
    layer8_outputs(1074) <= not b;
    layer8_outputs(1075) <= a;
    layer8_outputs(1076) <= not b;
    layer8_outputs(1077) <= a xor b;
    layer8_outputs(1078) <= a xor b;
    layer8_outputs(1079) <= a and b;
    layer8_outputs(1080) <= b and not a;
    layer8_outputs(1081) <= not a;
    layer8_outputs(1082) <= b and not a;
    layer8_outputs(1083) <= b;
    layer8_outputs(1084) <= a;
    layer8_outputs(1085) <= not a or b;
    layer8_outputs(1086) <= a xor b;
    layer8_outputs(1087) <= a;
    layer8_outputs(1088) <= a xor b;
    layer8_outputs(1089) <= b;
    layer8_outputs(1090) <= not a;
    layer8_outputs(1091) <= not a;
    layer8_outputs(1092) <= not b;
    layer8_outputs(1093) <= a;
    layer8_outputs(1094) <= not (a and b);
    layer8_outputs(1095) <= not (a xor b);
    layer8_outputs(1096) <= not (a xor b);
    layer8_outputs(1097) <= not a;
    layer8_outputs(1098) <= not b;
    layer8_outputs(1099) <= a xor b;
    layer8_outputs(1100) <= not a;
    layer8_outputs(1101) <= a xor b;
    layer8_outputs(1102) <= a and b;
    layer8_outputs(1103) <= a and b;
    layer8_outputs(1104) <= b;
    layer8_outputs(1105) <= a xor b;
    layer8_outputs(1106) <= b;
    layer8_outputs(1107) <= not a;
    layer8_outputs(1108) <= a;
    layer8_outputs(1109) <= b and not a;
    layer8_outputs(1110) <= a;
    layer8_outputs(1111) <= a xor b;
    layer8_outputs(1112) <= not a;
    layer8_outputs(1113) <= not b or a;
    layer8_outputs(1114) <= not (a or b);
    layer8_outputs(1115) <= a xor b;
    layer8_outputs(1116) <= not a or b;
    layer8_outputs(1117) <= not b or a;
    layer8_outputs(1118) <= not (a xor b);
    layer8_outputs(1119) <= b and not a;
    layer8_outputs(1120) <= a and b;
    layer8_outputs(1121) <= not a;
    layer8_outputs(1122) <= a xor b;
    layer8_outputs(1123) <= a;
    layer8_outputs(1124) <= b and not a;
    layer8_outputs(1125) <= not (a xor b);
    layer8_outputs(1126) <= a and b;
    layer8_outputs(1127) <= a and not b;
    layer8_outputs(1128) <= a and not b;
    layer8_outputs(1129) <= not b;
    layer8_outputs(1130) <= not b;
    layer8_outputs(1131) <= 1'b0;
    layer8_outputs(1132) <= not b or a;
    layer8_outputs(1133) <= not (a xor b);
    layer8_outputs(1134) <= not a;
    layer8_outputs(1135) <= not (a xor b);
    layer8_outputs(1136) <= a xor b;
    layer8_outputs(1137) <= not b;
    layer8_outputs(1138) <= 1'b1;
    layer8_outputs(1139) <= a or b;
    layer8_outputs(1140) <= not (a xor b);
    layer8_outputs(1141) <= a and not b;
    layer8_outputs(1142) <= not a or b;
    layer8_outputs(1143) <= a xor b;
    layer8_outputs(1144) <= not (a xor b);
    layer8_outputs(1145) <= not b or a;
    layer8_outputs(1146) <= not b;
    layer8_outputs(1147) <= a;
    layer8_outputs(1148) <= b;
    layer8_outputs(1149) <= b;
    layer8_outputs(1150) <= b;
    layer8_outputs(1151) <= not a;
    layer8_outputs(1152) <= a xor b;
    layer8_outputs(1153) <= a and b;
    layer8_outputs(1154) <= not (a xor b);
    layer8_outputs(1155) <= b;
    layer8_outputs(1156) <= a and not b;
    layer8_outputs(1157) <= a xor b;
    layer8_outputs(1158) <= a xor b;
    layer8_outputs(1159) <= b;
    layer8_outputs(1160) <= not b;
    layer8_outputs(1161) <= a;
    layer8_outputs(1162) <= a xor b;
    layer8_outputs(1163) <= not a;
    layer8_outputs(1164) <= a xor b;
    layer8_outputs(1165) <= not (a and b);
    layer8_outputs(1166) <= not (a and b);
    layer8_outputs(1167) <= not b;
    layer8_outputs(1168) <= a xor b;
    layer8_outputs(1169) <= not b or a;
    layer8_outputs(1170) <= not a;
    layer8_outputs(1171) <= not b;
    layer8_outputs(1172) <= b and not a;
    layer8_outputs(1173) <= not b;
    layer8_outputs(1174) <= not b;
    layer8_outputs(1175) <= not a;
    layer8_outputs(1176) <= a and b;
    layer8_outputs(1177) <= a and b;
    layer8_outputs(1178) <= a and b;
    layer8_outputs(1179) <= not (a and b);
    layer8_outputs(1180) <= not (a or b);
    layer8_outputs(1181) <= a or b;
    layer8_outputs(1182) <= not a;
    layer8_outputs(1183) <= a xor b;
    layer8_outputs(1184) <= a;
    layer8_outputs(1185) <= a xor b;
    layer8_outputs(1186) <= a and not b;
    layer8_outputs(1187) <= a and not b;
    layer8_outputs(1188) <= not a;
    layer8_outputs(1189) <= a;
    layer8_outputs(1190) <= b and not a;
    layer8_outputs(1191) <= b;
    layer8_outputs(1192) <= a xor b;
    layer8_outputs(1193) <= b;
    layer8_outputs(1194) <= not (a xor b);
    layer8_outputs(1195) <= a;
    layer8_outputs(1196) <= a;
    layer8_outputs(1197) <= a;
    layer8_outputs(1198) <= not a;
    layer8_outputs(1199) <= a and b;
    layer8_outputs(1200) <= not (a or b);
    layer8_outputs(1201) <= not b or a;
    layer8_outputs(1202) <= a and not b;
    layer8_outputs(1203) <= a;
    layer8_outputs(1204) <= not b;
    layer8_outputs(1205) <= b and not a;
    layer8_outputs(1206) <= not a;
    layer8_outputs(1207) <= not (a and b);
    layer8_outputs(1208) <= a;
    layer8_outputs(1209) <= not b;
    layer8_outputs(1210) <= a xor b;
    layer8_outputs(1211) <= a;
    layer8_outputs(1212) <= not b or a;
    layer8_outputs(1213) <= not b;
    layer8_outputs(1214) <= not a;
    layer8_outputs(1215) <= a;
    layer8_outputs(1216) <= not a;
    layer8_outputs(1217) <= not (a and b);
    layer8_outputs(1218) <= b;
    layer8_outputs(1219) <= not (a xor b);
    layer8_outputs(1220) <= not (a xor b);
    layer8_outputs(1221) <= a and not b;
    layer8_outputs(1222) <= not a;
    layer8_outputs(1223) <= a xor b;
    layer8_outputs(1224) <= not (a or b);
    layer8_outputs(1225) <= not (a xor b);
    layer8_outputs(1226) <= a and not b;
    layer8_outputs(1227) <= not (a xor b);
    layer8_outputs(1228) <= not b;
    layer8_outputs(1229) <= b and not a;
    layer8_outputs(1230) <= not (a xor b);
    layer8_outputs(1231) <= b;
    layer8_outputs(1232) <= b and not a;
    layer8_outputs(1233) <= not (a and b);
    layer8_outputs(1234) <= not a or b;
    layer8_outputs(1235) <= a;
    layer8_outputs(1236) <= b;
    layer8_outputs(1237) <= not a;
    layer8_outputs(1238) <= a;
    layer8_outputs(1239) <= not a;
    layer8_outputs(1240) <= not a;
    layer8_outputs(1241) <= not a;
    layer8_outputs(1242) <= a or b;
    layer8_outputs(1243) <= a and b;
    layer8_outputs(1244) <= b;
    layer8_outputs(1245) <= not (a xor b);
    layer8_outputs(1246) <= 1'b1;
    layer8_outputs(1247) <= not b;
    layer8_outputs(1248) <= a;
    layer8_outputs(1249) <= a or b;
    layer8_outputs(1250) <= b;
    layer8_outputs(1251) <= not a;
    layer8_outputs(1252) <= b;
    layer8_outputs(1253) <= not (a and b);
    layer8_outputs(1254) <= not b or a;
    layer8_outputs(1255) <= a xor b;
    layer8_outputs(1256) <= not a;
    layer8_outputs(1257) <= not b;
    layer8_outputs(1258) <= a;
    layer8_outputs(1259) <= a or b;
    layer8_outputs(1260) <= not a;
    layer8_outputs(1261) <= b;
    layer8_outputs(1262) <= not b;
    layer8_outputs(1263) <= a;
    layer8_outputs(1264) <= b;
    layer8_outputs(1265) <= not b or a;
    layer8_outputs(1266) <= a;
    layer8_outputs(1267) <= not a;
    layer8_outputs(1268) <= not a;
    layer8_outputs(1269) <= not a;
    layer8_outputs(1270) <= a;
    layer8_outputs(1271) <= not b;
    layer8_outputs(1272) <= not b;
    layer8_outputs(1273) <= a;
    layer8_outputs(1274) <= a;
    layer8_outputs(1275) <= b;
    layer8_outputs(1276) <= not b or a;
    layer8_outputs(1277) <= not (a xor b);
    layer8_outputs(1278) <= not (a xor b);
    layer8_outputs(1279) <= not (a or b);
    layer8_outputs(1280) <= a and b;
    layer8_outputs(1281) <= b;
    layer8_outputs(1282) <= not b;
    layer8_outputs(1283) <= b;
    layer8_outputs(1284) <= a;
    layer8_outputs(1285) <= 1'b1;
    layer8_outputs(1286) <= not a;
    layer8_outputs(1287) <= b;
    layer8_outputs(1288) <= not b or a;
    layer8_outputs(1289) <= a;
    layer8_outputs(1290) <= a;
    layer8_outputs(1291) <= a xor b;
    layer8_outputs(1292) <= b;
    layer8_outputs(1293) <= not (a xor b);
    layer8_outputs(1294) <= a;
    layer8_outputs(1295) <= not a;
    layer8_outputs(1296) <= not a;
    layer8_outputs(1297) <= a and b;
    layer8_outputs(1298) <= a;
    layer8_outputs(1299) <= not a or b;
    layer8_outputs(1300) <= a and b;
    layer8_outputs(1301) <= a xor b;
    layer8_outputs(1302) <= a xor b;
    layer8_outputs(1303) <= a;
    layer8_outputs(1304) <= a and not b;
    layer8_outputs(1305) <= a;
    layer8_outputs(1306) <= a xor b;
    layer8_outputs(1307) <= not (a or b);
    layer8_outputs(1308) <= not (a and b);
    layer8_outputs(1309) <= not a or b;
    layer8_outputs(1310) <= b;
    layer8_outputs(1311) <= not b;
    layer8_outputs(1312) <= not b;
    layer8_outputs(1313) <= a;
    layer8_outputs(1314) <= a or b;
    layer8_outputs(1315) <= 1'b0;
    layer8_outputs(1316) <= not b;
    layer8_outputs(1317) <= b;
    layer8_outputs(1318) <= not a;
    layer8_outputs(1319) <= not (a or b);
    layer8_outputs(1320) <= a;
    layer8_outputs(1321) <= a;
    layer8_outputs(1322) <= b;
    layer8_outputs(1323) <= not b;
    layer8_outputs(1324) <= not a;
    layer8_outputs(1325) <= a;
    layer8_outputs(1326) <= not (a xor b);
    layer8_outputs(1327) <= a;
    layer8_outputs(1328) <= a or b;
    layer8_outputs(1329) <= a;
    layer8_outputs(1330) <= b;
    layer8_outputs(1331) <= not (a xor b);
    layer8_outputs(1332) <= not a;
    layer8_outputs(1333) <= a;
    layer8_outputs(1334) <= not b;
    layer8_outputs(1335) <= a;
    layer8_outputs(1336) <= a and not b;
    layer8_outputs(1337) <= not (a and b);
    layer8_outputs(1338) <= b;
    layer8_outputs(1339) <= a;
    layer8_outputs(1340) <= b;
    layer8_outputs(1341) <= not a;
    layer8_outputs(1342) <= not (a and b);
    layer8_outputs(1343) <= a;
    layer8_outputs(1344) <= a;
    layer8_outputs(1345) <= not (a xor b);
    layer8_outputs(1346) <= not a;
    layer8_outputs(1347) <= a and not b;
    layer8_outputs(1348) <= a and b;
    layer8_outputs(1349) <= a xor b;
    layer8_outputs(1350) <= a;
    layer8_outputs(1351) <= not b;
    layer8_outputs(1352) <= not a;
    layer8_outputs(1353) <= not b;
    layer8_outputs(1354) <= not b;
    layer8_outputs(1355) <= a xor b;
    layer8_outputs(1356) <= a;
    layer8_outputs(1357) <= not a or b;
    layer8_outputs(1358) <= not b;
    layer8_outputs(1359) <= not (a xor b);
    layer8_outputs(1360) <= b;
    layer8_outputs(1361) <= a;
    layer8_outputs(1362) <= not (a xor b);
    layer8_outputs(1363) <= b;
    layer8_outputs(1364) <= 1'b1;
    layer8_outputs(1365) <= b;
    layer8_outputs(1366) <= a and not b;
    layer8_outputs(1367) <= not (a xor b);
    layer8_outputs(1368) <= not (a xor b);
    layer8_outputs(1369) <= not (a xor b);
    layer8_outputs(1370) <= a and b;
    layer8_outputs(1371) <= not (a xor b);
    layer8_outputs(1372) <= a xor b;
    layer8_outputs(1373) <= not (a or b);
    layer8_outputs(1374) <= a and b;
    layer8_outputs(1375) <= a and not b;
    layer8_outputs(1376) <= a;
    layer8_outputs(1377) <= a xor b;
    layer8_outputs(1378) <= not (a xor b);
    layer8_outputs(1379) <= b and not a;
    layer8_outputs(1380) <= a xor b;
    layer8_outputs(1381) <= a and not b;
    layer8_outputs(1382) <= not (a xor b);
    layer8_outputs(1383) <= b;
    layer8_outputs(1384) <= b and not a;
    layer8_outputs(1385) <= not a or b;
    layer8_outputs(1386) <= a;
    layer8_outputs(1387) <= not b;
    layer8_outputs(1388) <= a xor b;
    layer8_outputs(1389) <= a and b;
    layer8_outputs(1390) <= a;
    layer8_outputs(1391) <= not (a or b);
    layer8_outputs(1392) <= a and b;
    layer8_outputs(1393) <= a and b;
    layer8_outputs(1394) <= a;
    layer8_outputs(1395) <= b;
    layer8_outputs(1396) <= not a;
    layer8_outputs(1397) <= not b;
    layer8_outputs(1398) <= a;
    layer8_outputs(1399) <= not (a xor b);
    layer8_outputs(1400) <= not b or a;
    layer8_outputs(1401) <= a;
    layer8_outputs(1402) <= 1'b0;
    layer8_outputs(1403) <= b;
    layer8_outputs(1404) <= not b;
    layer8_outputs(1405) <= a;
    layer8_outputs(1406) <= not b or a;
    layer8_outputs(1407) <= a xor b;
    layer8_outputs(1408) <= not a;
    layer8_outputs(1409) <= not a;
    layer8_outputs(1410) <= a xor b;
    layer8_outputs(1411) <= not b;
    layer8_outputs(1412) <= not a;
    layer8_outputs(1413) <= b;
    layer8_outputs(1414) <= not (a xor b);
    layer8_outputs(1415) <= 1'b0;
    layer8_outputs(1416) <= not b or a;
    layer8_outputs(1417) <= not a or b;
    layer8_outputs(1418) <= a xor b;
    layer8_outputs(1419) <= not a;
    layer8_outputs(1420) <= not a;
    layer8_outputs(1421) <= a and not b;
    layer8_outputs(1422) <= a xor b;
    layer8_outputs(1423) <= 1'b1;
    layer8_outputs(1424) <= a;
    layer8_outputs(1425) <= not (a xor b);
    layer8_outputs(1426) <= b;
    layer8_outputs(1427) <= not (a xor b);
    layer8_outputs(1428) <= a and not b;
    layer8_outputs(1429) <= a xor b;
    layer8_outputs(1430) <= b;
    layer8_outputs(1431) <= not (a xor b);
    layer8_outputs(1432) <= a and not b;
    layer8_outputs(1433) <= not b or a;
    layer8_outputs(1434) <= a xor b;
    layer8_outputs(1435) <= not (a xor b);
    layer8_outputs(1436) <= not a or b;
    layer8_outputs(1437) <= b;
    layer8_outputs(1438) <= not (a or b);
    layer8_outputs(1439) <= b;
    layer8_outputs(1440) <= not a;
    layer8_outputs(1441) <= not b;
    layer8_outputs(1442) <= not b;
    layer8_outputs(1443) <= a and b;
    layer8_outputs(1444) <= b;
    layer8_outputs(1445) <= not a;
    layer8_outputs(1446) <= b and not a;
    layer8_outputs(1447) <= a xor b;
    layer8_outputs(1448) <= a;
    layer8_outputs(1449) <= a and not b;
    layer8_outputs(1450) <= a xor b;
    layer8_outputs(1451) <= not b;
    layer8_outputs(1452) <= not b;
    layer8_outputs(1453) <= b and not a;
    layer8_outputs(1454) <= a or b;
    layer8_outputs(1455) <= not (a xor b);
    layer8_outputs(1456) <= a xor b;
    layer8_outputs(1457) <= b;
    layer8_outputs(1458) <= a xor b;
    layer8_outputs(1459) <= not (a and b);
    layer8_outputs(1460) <= not b;
    layer8_outputs(1461) <= not (a xor b);
    layer8_outputs(1462) <= not a or b;
    layer8_outputs(1463) <= not (a xor b);
    layer8_outputs(1464) <= a;
    layer8_outputs(1465) <= not a;
    layer8_outputs(1466) <= not (a or b);
    layer8_outputs(1467) <= b;
    layer8_outputs(1468) <= b;
    layer8_outputs(1469) <= not a or b;
    layer8_outputs(1470) <= not (a and b);
    layer8_outputs(1471) <= not a or b;
    layer8_outputs(1472) <= a xor b;
    layer8_outputs(1473) <= a;
    layer8_outputs(1474) <= not b or a;
    layer8_outputs(1475) <= not (a and b);
    layer8_outputs(1476) <= not b or a;
    layer8_outputs(1477) <= 1'b0;
    layer8_outputs(1478) <= b;
    layer8_outputs(1479) <= not b or a;
    layer8_outputs(1480) <= a xor b;
    layer8_outputs(1481) <= a or b;
    layer8_outputs(1482) <= b and not a;
    layer8_outputs(1483) <= a xor b;
    layer8_outputs(1484) <= not (a and b);
    layer8_outputs(1485) <= b;
    layer8_outputs(1486) <= not b;
    layer8_outputs(1487) <= b and not a;
    layer8_outputs(1488) <= a or b;
    layer8_outputs(1489) <= a;
    layer8_outputs(1490) <= b;
    layer8_outputs(1491) <= a;
    layer8_outputs(1492) <= not b;
    layer8_outputs(1493) <= not a;
    layer8_outputs(1494) <= not a or b;
    layer8_outputs(1495) <= a xor b;
    layer8_outputs(1496) <= not a;
    layer8_outputs(1497) <= a;
    layer8_outputs(1498) <= b and not a;
    layer8_outputs(1499) <= not a;
    layer8_outputs(1500) <= not b;
    layer8_outputs(1501) <= not (a xor b);
    layer8_outputs(1502) <= not (a xor b);
    layer8_outputs(1503) <= a xor b;
    layer8_outputs(1504) <= a xor b;
    layer8_outputs(1505) <= a;
    layer8_outputs(1506) <= a xor b;
    layer8_outputs(1507) <= b;
    layer8_outputs(1508) <= a;
    layer8_outputs(1509) <= b and not a;
    layer8_outputs(1510) <= not a or b;
    layer8_outputs(1511) <= not a;
    layer8_outputs(1512) <= not (a xor b);
    layer8_outputs(1513) <= a;
    layer8_outputs(1514) <= b;
    layer8_outputs(1515) <= a;
    layer8_outputs(1516) <= not b;
    layer8_outputs(1517) <= not (a xor b);
    layer8_outputs(1518) <= b;
    layer8_outputs(1519) <= not a;
    layer8_outputs(1520) <= a xor b;
    layer8_outputs(1521) <= not a;
    layer8_outputs(1522) <= a and not b;
    layer8_outputs(1523) <= not b;
    layer8_outputs(1524) <= not (a or b);
    layer8_outputs(1525) <= not a;
    layer8_outputs(1526) <= not (a xor b);
    layer8_outputs(1527) <= not (a xor b);
    layer8_outputs(1528) <= b;
    layer8_outputs(1529) <= not a;
    layer8_outputs(1530) <= not (a or b);
    layer8_outputs(1531) <= b;
    layer8_outputs(1532) <= a xor b;
    layer8_outputs(1533) <= a or b;
    layer8_outputs(1534) <= a;
    layer8_outputs(1535) <= not b;
    layer8_outputs(1536) <= b and not a;
    layer8_outputs(1537) <= a or b;
    layer8_outputs(1538) <= a;
    layer8_outputs(1539) <= not a;
    layer8_outputs(1540) <= a and b;
    layer8_outputs(1541) <= a xor b;
    layer8_outputs(1542) <= not b;
    layer8_outputs(1543) <= a xor b;
    layer8_outputs(1544) <= b;
    layer8_outputs(1545) <= b;
    layer8_outputs(1546) <= b;
    layer8_outputs(1547) <= not (a xor b);
    layer8_outputs(1548) <= a or b;
    layer8_outputs(1549) <= not b or a;
    layer8_outputs(1550) <= a and not b;
    layer8_outputs(1551) <= a;
    layer8_outputs(1552) <= not (a or b);
    layer8_outputs(1553) <= not (a xor b);
    layer8_outputs(1554) <= not b;
    layer8_outputs(1555) <= b;
    layer8_outputs(1556) <= not a;
    layer8_outputs(1557) <= a or b;
    layer8_outputs(1558) <= not a or b;
    layer8_outputs(1559) <= a xor b;
    layer8_outputs(1560) <= b;
    layer8_outputs(1561) <= b;
    layer8_outputs(1562) <= a;
    layer8_outputs(1563) <= not a;
    layer8_outputs(1564) <= b;
    layer8_outputs(1565) <= a;
    layer8_outputs(1566) <= not a;
    layer8_outputs(1567) <= not (a and b);
    layer8_outputs(1568) <= not a or b;
    layer8_outputs(1569) <= a xor b;
    layer8_outputs(1570) <= not (a xor b);
    layer8_outputs(1571) <= b and not a;
    layer8_outputs(1572) <= b;
    layer8_outputs(1573) <= a xor b;
    layer8_outputs(1574) <= a and b;
    layer8_outputs(1575) <= b and not a;
    layer8_outputs(1576) <= a xor b;
    layer8_outputs(1577) <= b;
    layer8_outputs(1578) <= b;
    layer8_outputs(1579) <= not a;
    layer8_outputs(1580) <= not (a and b);
    layer8_outputs(1581) <= not b;
    layer8_outputs(1582) <= not a or b;
    layer8_outputs(1583) <= a;
    layer8_outputs(1584) <= not a;
    layer8_outputs(1585) <= not b;
    layer8_outputs(1586) <= not a or b;
    layer8_outputs(1587) <= b;
    layer8_outputs(1588) <= b;
    layer8_outputs(1589) <= a and not b;
    layer8_outputs(1590) <= a xor b;
    layer8_outputs(1591) <= a xor b;
    layer8_outputs(1592) <= not a;
    layer8_outputs(1593) <= not a;
    layer8_outputs(1594) <= not b;
    layer8_outputs(1595) <= not (a xor b);
    layer8_outputs(1596) <= not a;
    layer8_outputs(1597) <= a and not b;
    layer8_outputs(1598) <= not b;
    layer8_outputs(1599) <= a and not b;
    layer8_outputs(1600) <= a and not b;
    layer8_outputs(1601) <= a;
    layer8_outputs(1602) <= not b;
    layer8_outputs(1603) <= not b;
    layer8_outputs(1604) <= a xor b;
    layer8_outputs(1605) <= a;
    layer8_outputs(1606) <= not (a or b);
    layer8_outputs(1607) <= not a or b;
    layer8_outputs(1608) <= b;
    layer8_outputs(1609) <= b and not a;
    layer8_outputs(1610) <= not a or b;
    layer8_outputs(1611) <= a;
    layer8_outputs(1612) <= not (a and b);
    layer8_outputs(1613) <= not (a or b);
    layer8_outputs(1614) <= a or b;
    layer8_outputs(1615) <= not (a and b);
    layer8_outputs(1616) <= not a;
    layer8_outputs(1617) <= not a;
    layer8_outputs(1618) <= a xor b;
    layer8_outputs(1619) <= not b;
    layer8_outputs(1620) <= not a;
    layer8_outputs(1621) <= b;
    layer8_outputs(1622) <= not a or b;
    layer8_outputs(1623) <= not a;
    layer8_outputs(1624) <= not a or b;
    layer8_outputs(1625) <= not a;
    layer8_outputs(1626) <= a or b;
    layer8_outputs(1627) <= not b;
    layer8_outputs(1628) <= not b;
    layer8_outputs(1629) <= b;
    layer8_outputs(1630) <= not b;
    layer8_outputs(1631) <= not a;
    layer8_outputs(1632) <= a xor b;
    layer8_outputs(1633) <= not (a and b);
    layer8_outputs(1634) <= not (a xor b);
    layer8_outputs(1635) <= not (a and b);
    layer8_outputs(1636) <= not (a and b);
    layer8_outputs(1637) <= not (a or b);
    layer8_outputs(1638) <= not (a xor b);
    layer8_outputs(1639) <= a;
    layer8_outputs(1640) <= a;
    layer8_outputs(1641) <= a xor b;
    layer8_outputs(1642) <= not a;
    layer8_outputs(1643) <= not b;
    layer8_outputs(1644) <= a;
    layer8_outputs(1645) <= a xor b;
    layer8_outputs(1646) <= not b;
    layer8_outputs(1647) <= a or b;
    layer8_outputs(1648) <= not b;
    layer8_outputs(1649) <= a;
    layer8_outputs(1650) <= b;
    layer8_outputs(1651) <= not (a xor b);
    layer8_outputs(1652) <= not b or a;
    layer8_outputs(1653) <= a and not b;
    layer8_outputs(1654) <= a;
    layer8_outputs(1655) <= b;
    layer8_outputs(1656) <= a xor b;
    layer8_outputs(1657) <= not (a xor b);
    layer8_outputs(1658) <= not b;
    layer8_outputs(1659) <= not a;
    layer8_outputs(1660) <= a xor b;
    layer8_outputs(1661) <= not a or b;
    layer8_outputs(1662) <= a;
    layer8_outputs(1663) <= a;
    layer8_outputs(1664) <= not (a xor b);
    layer8_outputs(1665) <= a xor b;
    layer8_outputs(1666) <= a;
    layer8_outputs(1667) <= b;
    layer8_outputs(1668) <= a and not b;
    layer8_outputs(1669) <= not b or a;
    layer8_outputs(1670) <= b;
    layer8_outputs(1671) <= not a;
    layer8_outputs(1672) <= a and b;
    layer8_outputs(1673) <= a xor b;
    layer8_outputs(1674) <= not (a xor b);
    layer8_outputs(1675) <= a and not b;
    layer8_outputs(1676) <= not (a xor b);
    layer8_outputs(1677) <= not a;
    layer8_outputs(1678) <= not a;
    layer8_outputs(1679) <= 1'b0;
    layer8_outputs(1680) <= not b;
    layer8_outputs(1681) <= a xor b;
    layer8_outputs(1682) <= not b or a;
    layer8_outputs(1683) <= a;
    layer8_outputs(1684) <= b;
    layer8_outputs(1685) <= not a;
    layer8_outputs(1686) <= not a or b;
    layer8_outputs(1687) <= a xor b;
    layer8_outputs(1688) <= not b;
    layer8_outputs(1689) <= a;
    layer8_outputs(1690) <= not a;
    layer8_outputs(1691) <= b;
    layer8_outputs(1692) <= not b;
    layer8_outputs(1693) <= a and b;
    layer8_outputs(1694) <= a;
    layer8_outputs(1695) <= a;
    layer8_outputs(1696) <= not (a xor b);
    layer8_outputs(1697) <= a xor b;
    layer8_outputs(1698) <= not a;
    layer8_outputs(1699) <= not (a xor b);
    layer8_outputs(1700) <= not b;
    layer8_outputs(1701) <= a xor b;
    layer8_outputs(1702) <= b;
    layer8_outputs(1703) <= a xor b;
    layer8_outputs(1704) <= a and b;
    layer8_outputs(1705) <= not a or b;
    layer8_outputs(1706) <= a xor b;
    layer8_outputs(1707) <= not b;
    layer8_outputs(1708) <= not (a and b);
    layer8_outputs(1709) <= not b;
    layer8_outputs(1710) <= not b;
    layer8_outputs(1711) <= a and not b;
    layer8_outputs(1712) <= a or b;
    layer8_outputs(1713) <= not a;
    layer8_outputs(1714) <= a;
    layer8_outputs(1715) <= a and not b;
    layer8_outputs(1716) <= b;
    layer8_outputs(1717) <= not (a xor b);
    layer8_outputs(1718) <= not (a xor b);
    layer8_outputs(1719) <= a and b;
    layer8_outputs(1720) <= a and not b;
    layer8_outputs(1721) <= b and not a;
    layer8_outputs(1722) <= not (a or b);
    layer8_outputs(1723) <= a xor b;
    layer8_outputs(1724) <= a;
    layer8_outputs(1725) <= not b;
    layer8_outputs(1726) <= not b;
    layer8_outputs(1727) <= a;
    layer8_outputs(1728) <= b;
    layer8_outputs(1729) <= not b;
    layer8_outputs(1730) <= b;
    layer8_outputs(1731) <= not b;
    layer8_outputs(1732) <= a and not b;
    layer8_outputs(1733) <= not b;
    layer8_outputs(1734) <= not b or a;
    layer8_outputs(1735) <= not a;
    layer8_outputs(1736) <= not (a xor b);
    layer8_outputs(1737) <= a xor b;
    layer8_outputs(1738) <= b and not a;
    layer8_outputs(1739) <= a xor b;
    layer8_outputs(1740) <= b;
    layer8_outputs(1741) <= not a;
    layer8_outputs(1742) <= not (a xor b);
    layer8_outputs(1743) <= not a;
    layer8_outputs(1744) <= 1'b0;
    layer8_outputs(1745) <= a;
    layer8_outputs(1746) <= not b or a;
    layer8_outputs(1747) <= not a;
    layer8_outputs(1748) <= 1'b1;
    layer8_outputs(1749) <= a xor b;
    layer8_outputs(1750) <= a xor b;
    layer8_outputs(1751) <= a and b;
    layer8_outputs(1752) <= a and b;
    layer8_outputs(1753) <= not b;
    layer8_outputs(1754) <= not a;
    layer8_outputs(1755) <= b;
    layer8_outputs(1756) <= not a or b;
    layer8_outputs(1757) <= not a or b;
    layer8_outputs(1758) <= not (a xor b);
    layer8_outputs(1759) <= b and not a;
    layer8_outputs(1760) <= not (a xor b);
    layer8_outputs(1761) <= a and not b;
    layer8_outputs(1762) <= b;
    layer8_outputs(1763) <= a and b;
    layer8_outputs(1764) <= b;
    layer8_outputs(1765) <= b;
    layer8_outputs(1766) <= not b or a;
    layer8_outputs(1767) <= a and not b;
    layer8_outputs(1768) <= b and not a;
    layer8_outputs(1769) <= a xor b;
    layer8_outputs(1770) <= not b;
    layer8_outputs(1771) <= b;
    layer8_outputs(1772) <= not b;
    layer8_outputs(1773) <= b;
    layer8_outputs(1774) <= not (a and b);
    layer8_outputs(1775) <= b;
    layer8_outputs(1776) <= b and not a;
    layer8_outputs(1777) <= not b;
    layer8_outputs(1778) <= not a;
    layer8_outputs(1779) <= not b or a;
    layer8_outputs(1780) <= not (a and b);
    layer8_outputs(1781) <= not b;
    layer8_outputs(1782) <= not (a and b);
    layer8_outputs(1783) <= not (a or b);
    layer8_outputs(1784) <= b and not a;
    layer8_outputs(1785) <= not (a or b);
    layer8_outputs(1786) <= not b;
    layer8_outputs(1787) <= a;
    layer8_outputs(1788) <= not b or a;
    layer8_outputs(1789) <= a or b;
    layer8_outputs(1790) <= not (a or b);
    layer8_outputs(1791) <= a;
    layer8_outputs(1792) <= a;
    layer8_outputs(1793) <= not b;
    layer8_outputs(1794) <= not (a xor b);
    layer8_outputs(1795) <= not a;
    layer8_outputs(1796) <= a;
    layer8_outputs(1797) <= b;
    layer8_outputs(1798) <= b;
    layer8_outputs(1799) <= not (a xor b);
    layer8_outputs(1800) <= a xor b;
    layer8_outputs(1801) <= a;
    layer8_outputs(1802) <= not b;
    layer8_outputs(1803) <= not (a xor b);
    layer8_outputs(1804) <= not a or b;
    layer8_outputs(1805) <= a;
    layer8_outputs(1806) <= not b;
    layer8_outputs(1807) <= a xor b;
    layer8_outputs(1808) <= not (a xor b);
    layer8_outputs(1809) <= a;
    layer8_outputs(1810) <= not b;
    layer8_outputs(1811) <= b;
    layer8_outputs(1812) <= a;
    layer8_outputs(1813) <= 1'b1;
    layer8_outputs(1814) <= a;
    layer8_outputs(1815) <= a;
    layer8_outputs(1816) <= b;
    layer8_outputs(1817) <= b;
    layer8_outputs(1818) <= not a;
    layer8_outputs(1819) <= not a;
    layer8_outputs(1820) <= a or b;
    layer8_outputs(1821) <= a;
    layer8_outputs(1822) <= not (a xor b);
    layer8_outputs(1823) <= not (a xor b);
    layer8_outputs(1824) <= not a;
    layer8_outputs(1825) <= not (a xor b);
    layer8_outputs(1826) <= a;
    layer8_outputs(1827) <= not (a xor b);
    layer8_outputs(1828) <= a;
    layer8_outputs(1829) <= a;
    layer8_outputs(1830) <= a xor b;
    layer8_outputs(1831) <= not (a xor b);
    layer8_outputs(1832) <= b;
    layer8_outputs(1833) <= not (a or b);
    layer8_outputs(1834) <= a or b;
    layer8_outputs(1835) <= not (a or b);
    layer8_outputs(1836) <= not b;
    layer8_outputs(1837) <= a xor b;
    layer8_outputs(1838) <= a;
    layer8_outputs(1839) <= not b;
    layer8_outputs(1840) <= not (a or b);
    layer8_outputs(1841) <= a xor b;
    layer8_outputs(1842) <= a;
    layer8_outputs(1843) <= not (a xor b);
    layer8_outputs(1844) <= not a;
    layer8_outputs(1845) <= not b;
    layer8_outputs(1846) <= not b;
    layer8_outputs(1847) <= b and not a;
    layer8_outputs(1848) <= not a;
    layer8_outputs(1849) <= a;
    layer8_outputs(1850) <= a and b;
    layer8_outputs(1851) <= a xor b;
    layer8_outputs(1852) <= a xor b;
    layer8_outputs(1853) <= not (a or b);
    layer8_outputs(1854) <= a or b;
    layer8_outputs(1855) <= a and not b;
    layer8_outputs(1856) <= not (a and b);
    layer8_outputs(1857) <= a;
    layer8_outputs(1858) <= a or b;
    layer8_outputs(1859) <= not b;
    layer8_outputs(1860) <= b;
    layer8_outputs(1861) <= not (a xor b);
    layer8_outputs(1862) <= a;
    layer8_outputs(1863) <= not b;
    layer8_outputs(1864) <= a xor b;
    layer8_outputs(1865) <= not (a xor b);
    layer8_outputs(1866) <= b;
    layer8_outputs(1867) <= a;
    layer8_outputs(1868) <= a and b;
    layer8_outputs(1869) <= a;
    layer8_outputs(1870) <= a xor b;
    layer8_outputs(1871) <= a and not b;
    layer8_outputs(1872) <= not a or b;
    layer8_outputs(1873) <= a xor b;
    layer8_outputs(1874) <= b and not a;
    layer8_outputs(1875) <= not b;
    layer8_outputs(1876) <= not b;
    layer8_outputs(1877) <= a or b;
    layer8_outputs(1878) <= not b or a;
    layer8_outputs(1879) <= not b or a;
    layer8_outputs(1880) <= a and b;
    layer8_outputs(1881) <= not b;
    layer8_outputs(1882) <= a or b;
    layer8_outputs(1883) <= a xor b;
    layer8_outputs(1884) <= a;
    layer8_outputs(1885) <= not a;
    layer8_outputs(1886) <= a;
    layer8_outputs(1887) <= a or b;
    layer8_outputs(1888) <= a xor b;
    layer8_outputs(1889) <= not (a xor b);
    layer8_outputs(1890) <= not (a xor b);
    layer8_outputs(1891) <= a;
    layer8_outputs(1892) <= not a or b;
    layer8_outputs(1893) <= not a;
    layer8_outputs(1894) <= not a;
    layer8_outputs(1895) <= a or b;
    layer8_outputs(1896) <= not b;
    layer8_outputs(1897) <= 1'b1;
    layer8_outputs(1898) <= a and b;
    layer8_outputs(1899) <= a xor b;
    layer8_outputs(1900) <= a;
    layer8_outputs(1901) <= b;
    layer8_outputs(1902) <= a xor b;
    layer8_outputs(1903) <= a or b;
    layer8_outputs(1904) <= a and not b;
    layer8_outputs(1905) <= not a;
    layer8_outputs(1906) <= a xor b;
    layer8_outputs(1907) <= not b;
    layer8_outputs(1908) <= a and b;
    layer8_outputs(1909) <= not (a or b);
    layer8_outputs(1910) <= a xor b;
    layer8_outputs(1911) <= not a;
    layer8_outputs(1912) <= not b;
    layer8_outputs(1913) <= a and not b;
    layer8_outputs(1914) <= b;
    layer8_outputs(1915) <= a;
    layer8_outputs(1916) <= a;
    layer8_outputs(1917) <= not (a xor b);
    layer8_outputs(1918) <= not (a xor b);
    layer8_outputs(1919) <= not b;
    layer8_outputs(1920) <= not a;
    layer8_outputs(1921) <= a xor b;
    layer8_outputs(1922) <= not (a xor b);
    layer8_outputs(1923) <= not b or a;
    layer8_outputs(1924) <= b and not a;
    layer8_outputs(1925) <= a;
    layer8_outputs(1926) <= not (a or b);
    layer8_outputs(1927) <= not a;
    layer8_outputs(1928) <= a or b;
    layer8_outputs(1929) <= not (a and b);
    layer8_outputs(1930) <= not (a xor b);
    layer8_outputs(1931) <= not a or b;
    layer8_outputs(1932) <= a xor b;
    layer8_outputs(1933) <= not (a xor b);
    layer8_outputs(1934) <= a xor b;
    layer8_outputs(1935) <= b and not a;
    layer8_outputs(1936) <= not a;
    layer8_outputs(1937) <= not (a xor b);
    layer8_outputs(1938) <= not a;
    layer8_outputs(1939) <= b and not a;
    layer8_outputs(1940) <= a xor b;
    layer8_outputs(1941) <= b and not a;
    layer8_outputs(1942) <= not a;
    layer8_outputs(1943) <= b;
    layer8_outputs(1944) <= not a or b;
    layer8_outputs(1945) <= a;
    layer8_outputs(1946) <= b;
    layer8_outputs(1947) <= not b;
    layer8_outputs(1948) <= not a;
    layer8_outputs(1949) <= a;
    layer8_outputs(1950) <= 1'b1;
    layer8_outputs(1951) <= not a or b;
    layer8_outputs(1952) <= a and not b;
    layer8_outputs(1953) <= not (a or b);
    layer8_outputs(1954) <= not b;
    layer8_outputs(1955) <= a;
    layer8_outputs(1956) <= not b;
    layer8_outputs(1957) <= not (a xor b);
    layer8_outputs(1958) <= b and not a;
    layer8_outputs(1959) <= not b;
    layer8_outputs(1960) <= not a;
    layer8_outputs(1961) <= not (a or b);
    layer8_outputs(1962) <= a and not b;
    layer8_outputs(1963) <= a xor b;
    layer8_outputs(1964) <= a;
    layer8_outputs(1965) <= a;
    layer8_outputs(1966) <= not b;
    layer8_outputs(1967) <= not b;
    layer8_outputs(1968) <= not b;
    layer8_outputs(1969) <= a xor b;
    layer8_outputs(1970) <= not b;
    layer8_outputs(1971) <= a xor b;
    layer8_outputs(1972) <= a;
    layer8_outputs(1973) <= a and not b;
    layer8_outputs(1974) <= a;
    layer8_outputs(1975) <= not a or b;
    layer8_outputs(1976) <= a xor b;
    layer8_outputs(1977) <= a xor b;
    layer8_outputs(1978) <= b;
    layer8_outputs(1979) <= not a;
    layer8_outputs(1980) <= not (a xor b);
    layer8_outputs(1981) <= not b;
    layer8_outputs(1982) <= not a;
    layer8_outputs(1983) <= not (a and b);
    layer8_outputs(1984) <= not a;
    layer8_outputs(1985) <= a xor b;
    layer8_outputs(1986) <= b;
    layer8_outputs(1987) <= not (a xor b);
    layer8_outputs(1988) <= b;
    layer8_outputs(1989) <= not (a xor b);
    layer8_outputs(1990) <= not b;
    layer8_outputs(1991) <= a;
    layer8_outputs(1992) <= not (a or b);
    layer8_outputs(1993) <= a;
    layer8_outputs(1994) <= not a;
    layer8_outputs(1995) <= a and b;
    layer8_outputs(1996) <= not (a xor b);
    layer8_outputs(1997) <= not a;
    layer8_outputs(1998) <= not b or a;
    layer8_outputs(1999) <= not a;
    layer8_outputs(2000) <= a xor b;
    layer8_outputs(2001) <= not (a or b);
    layer8_outputs(2002) <= not (a and b);
    layer8_outputs(2003) <= a xor b;
    layer8_outputs(2004) <= a and b;
    layer8_outputs(2005) <= a;
    layer8_outputs(2006) <= a and b;
    layer8_outputs(2007) <= a or b;
    layer8_outputs(2008) <= a xor b;
    layer8_outputs(2009) <= not a;
    layer8_outputs(2010) <= a xor b;
    layer8_outputs(2011) <= not a;
    layer8_outputs(2012) <= a;
    layer8_outputs(2013) <= not (a xor b);
    layer8_outputs(2014) <= a xor b;
    layer8_outputs(2015) <= a and b;
    layer8_outputs(2016) <= not a;
    layer8_outputs(2017) <= a xor b;
    layer8_outputs(2018) <= not (a xor b);
    layer8_outputs(2019) <= a or b;
    layer8_outputs(2020) <= b and not a;
    layer8_outputs(2021) <= not (a xor b);
    layer8_outputs(2022) <= not (a xor b);
    layer8_outputs(2023) <= a or b;
    layer8_outputs(2024) <= a and not b;
    layer8_outputs(2025) <= b;
    layer8_outputs(2026) <= not (a xor b);
    layer8_outputs(2027) <= b;
    layer8_outputs(2028) <= not a;
    layer8_outputs(2029) <= b;
    layer8_outputs(2030) <= not a;
    layer8_outputs(2031) <= not (a and b);
    layer8_outputs(2032) <= a;
    layer8_outputs(2033) <= not (a xor b);
    layer8_outputs(2034) <= a xor b;
    layer8_outputs(2035) <= not b or a;
    layer8_outputs(2036) <= a;
    layer8_outputs(2037) <= not b;
    layer8_outputs(2038) <= not b;
    layer8_outputs(2039) <= a or b;
    layer8_outputs(2040) <= not (a xor b);
    layer8_outputs(2041) <= b;
    layer8_outputs(2042) <= not (a or b);
    layer8_outputs(2043) <= b and not a;
    layer8_outputs(2044) <= a and not b;
    layer8_outputs(2045) <= a and b;
    layer8_outputs(2046) <= not (a or b);
    layer8_outputs(2047) <= not (a xor b);
    layer8_outputs(2048) <= b;
    layer8_outputs(2049) <= not a;
    layer8_outputs(2050) <= not (a xor b);
    layer8_outputs(2051) <= not (a or b);
    layer8_outputs(2052) <= a xor b;
    layer8_outputs(2053) <= a;
    layer8_outputs(2054) <= b;
    layer8_outputs(2055) <= b;
    layer8_outputs(2056) <= a or b;
    layer8_outputs(2057) <= not a;
    layer8_outputs(2058) <= not a or b;
    layer8_outputs(2059) <= b and not a;
    layer8_outputs(2060) <= not (a xor b);
    layer8_outputs(2061) <= a;
    layer8_outputs(2062) <= a and not b;
    layer8_outputs(2063) <= not b;
    layer8_outputs(2064) <= not b;
    layer8_outputs(2065) <= not b;
    layer8_outputs(2066) <= b;
    layer8_outputs(2067) <= not b;
    layer8_outputs(2068) <= a xor b;
    layer8_outputs(2069) <= a and not b;
    layer8_outputs(2070) <= a;
    layer8_outputs(2071) <= not (a xor b);
    layer8_outputs(2072) <= b;
    layer8_outputs(2073) <= b;
    layer8_outputs(2074) <= a;
    layer8_outputs(2075) <= not (a xor b);
    layer8_outputs(2076) <= not a or b;
    layer8_outputs(2077) <= not (a or b);
    layer8_outputs(2078) <= not b;
    layer8_outputs(2079) <= not (a xor b);
    layer8_outputs(2080) <= b;
    layer8_outputs(2081) <= not b;
    layer8_outputs(2082) <= b;
    layer8_outputs(2083) <= a xor b;
    layer8_outputs(2084) <= not b;
    layer8_outputs(2085) <= not a;
    layer8_outputs(2086) <= not a;
    layer8_outputs(2087) <= b;
    layer8_outputs(2088) <= b and not a;
    layer8_outputs(2089) <= a;
    layer8_outputs(2090) <= 1'b0;
    layer8_outputs(2091) <= not b;
    layer8_outputs(2092) <= not b or a;
    layer8_outputs(2093) <= a;
    layer8_outputs(2094) <= not (a xor b);
    layer8_outputs(2095) <= b;
    layer8_outputs(2096) <= not (a or b);
    layer8_outputs(2097) <= b and not a;
    layer8_outputs(2098) <= not a;
    layer8_outputs(2099) <= a;
    layer8_outputs(2100) <= not a;
    layer8_outputs(2101) <= not b or a;
    layer8_outputs(2102) <= not (a or b);
    layer8_outputs(2103) <= not b;
    layer8_outputs(2104) <= a and b;
    layer8_outputs(2105) <= b;
    layer8_outputs(2106) <= not a;
    layer8_outputs(2107) <= a xor b;
    layer8_outputs(2108) <= not a or b;
    layer8_outputs(2109) <= b;
    layer8_outputs(2110) <= not (a xor b);
    layer8_outputs(2111) <= a;
    layer8_outputs(2112) <= a;
    layer8_outputs(2113) <= not (a xor b);
    layer8_outputs(2114) <= not a;
    layer8_outputs(2115) <= not b or a;
    layer8_outputs(2116) <= b and not a;
    layer8_outputs(2117) <= a;
    layer8_outputs(2118) <= a or b;
    layer8_outputs(2119) <= not (a xor b);
    layer8_outputs(2120) <= b;
    layer8_outputs(2121) <= not (a xor b);
    layer8_outputs(2122) <= not b or a;
    layer8_outputs(2123) <= a or b;
    layer8_outputs(2124) <= not (a xor b);
    layer8_outputs(2125) <= a;
    layer8_outputs(2126) <= b;
    layer8_outputs(2127) <= a and not b;
    layer8_outputs(2128) <= a and not b;
    layer8_outputs(2129) <= b;
    layer8_outputs(2130) <= a xor b;
    layer8_outputs(2131) <= b;
    layer8_outputs(2132) <= a;
    layer8_outputs(2133) <= not a;
    layer8_outputs(2134) <= a;
    layer8_outputs(2135) <= b;
    layer8_outputs(2136) <= not b;
    layer8_outputs(2137) <= not b;
    layer8_outputs(2138) <= a;
    layer8_outputs(2139) <= not a;
    layer8_outputs(2140) <= not (a xor b);
    layer8_outputs(2141) <= a or b;
    layer8_outputs(2142) <= not b;
    layer8_outputs(2143) <= a;
    layer8_outputs(2144) <= not b or a;
    layer8_outputs(2145) <= b;
    layer8_outputs(2146) <= a or b;
    layer8_outputs(2147) <= a;
    layer8_outputs(2148) <= b;
    layer8_outputs(2149) <= a xor b;
    layer8_outputs(2150) <= b and not a;
    layer8_outputs(2151) <= not b;
    layer8_outputs(2152) <= not a;
    layer8_outputs(2153) <= a;
    layer8_outputs(2154) <= a xor b;
    layer8_outputs(2155) <= a or b;
    layer8_outputs(2156) <= not (a xor b);
    layer8_outputs(2157) <= not b;
    layer8_outputs(2158) <= not b or a;
    layer8_outputs(2159) <= a;
    layer8_outputs(2160) <= b;
    layer8_outputs(2161) <= not a or b;
    layer8_outputs(2162) <= a or b;
    layer8_outputs(2163) <= a xor b;
    layer8_outputs(2164) <= not b;
    layer8_outputs(2165) <= a and not b;
    layer8_outputs(2166) <= b and not a;
    layer8_outputs(2167) <= a;
    layer8_outputs(2168) <= a or b;
    layer8_outputs(2169) <= a xor b;
    layer8_outputs(2170) <= a and not b;
    layer8_outputs(2171) <= not b;
    layer8_outputs(2172) <= not b;
    layer8_outputs(2173) <= a xor b;
    layer8_outputs(2174) <= not b or a;
    layer8_outputs(2175) <= not (a xor b);
    layer8_outputs(2176) <= not b;
    layer8_outputs(2177) <= not b;
    layer8_outputs(2178) <= not b;
    layer8_outputs(2179) <= a;
    layer8_outputs(2180) <= a;
    layer8_outputs(2181) <= a;
    layer8_outputs(2182) <= a;
    layer8_outputs(2183) <= not (a and b);
    layer8_outputs(2184) <= not (a or b);
    layer8_outputs(2185) <= a;
    layer8_outputs(2186) <= a or b;
    layer8_outputs(2187) <= not (a xor b);
    layer8_outputs(2188) <= not (a xor b);
    layer8_outputs(2189) <= not (a xor b);
    layer8_outputs(2190) <= b;
    layer8_outputs(2191) <= not a;
    layer8_outputs(2192) <= a and not b;
    layer8_outputs(2193) <= not a;
    layer8_outputs(2194) <= b and not a;
    layer8_outputs(2195) <= 1'b0;
    layer8_outputs(2196) <= not a;
    layer8_outputs(2197) <= a or b;
    layer8_outputs(2198) <= b;
    layer8_outputs(2199) <= not (a or b);
    layer8_outputs(2200) <= a;
    layer8_outputs(2201) <= not (a xor b);
    layer8_outputs(2202) <= a and not b;
    layer8_outputs(2203) <= a;
    layer8_outputs(2204) <= a and b;
    layer8_outputs(2205) <= a xor b;
    layer8_outputs(2206) <= a;
    layer8_outputs(2207) <= not a or b;
    layer8_outputs(2208) <= not (a or b);
    layer8_outputs(2209) <= not a or b;
    layer8_outputs(2210) <= a;
    layer8_outputs(2211) <= not a;
    layer8_outputs(2212) <= a xor b;
    layer8_outputs(2213) <= not (a or b);
    layer8_outputs(2214) <= a xor b;
    layer8_outputs(2215) <= not a;
    layer8_outputs(2216) <= not a or b;
    layer8_outputs(2217) <= a;
    layer8_outputs(2218) <= b;
    layer8_outputs(2219) <= b;
    layer8_outputs(2220) <= a xor b;
    layer8_outputs(2221) <= not b;
    layer8_outputs(2222) <= a or b;
    layer8_outputs(2223) <= not a or b;
    layer8_outputs(2224) <= b;
    layer8_outputs(2225) <= not (a xor b);
    layer8_outputs(2226) <= not a;
    layer8_outputs(2227) <= a;
    layer8_outputs(2228) <= 1'b1;
    layer8_outputs(2229) <= b;
    layer8_outputs(2230) <= not b;
    layer8_outputs(2231) <= a xor b;
    layer8_outputs(2232) <= not a or b;
    layer8_outputs(2233) <= b;
    layer8_outputs(2234) <= not (a xor b);
    layer8_outputs(2235) <= not a;
    layer8_outputs(2236) <= not a;
    layer8_outputs(2237) <= a or b;
    layer8_outputs(2238) <= not b;
    layer8_outputs(2239) <= a xor b;
    layer8_outputs(2240) <= a xor b;
    layer8_outputs(2241) <= b;
    layer8_outputs(2242) <= not b;
    layer8_outputs(2243) <= not a;
    layer8_outputs(2244) <= not a;
    layer8_outputs(2245) <= not b or a;
    layer8_outputs(2246) <= a or b;
    layer8_outputs(2247) <= a and b;
    layer8_outputs(2248) <= not b or a;
    layer8_outputs(2249) <= b;
    layer8_outputs(2250) <= not b;
    layer8_outputs(2251) <= not a;
    layer8_outputs(2252) <= b and not a;
    layer8_outputs(2253) <= not (a or b);
    layer8_outputs(2254) <= not a;
    layer8_outputs(2255) <= b;
    layer8_outputs(2256) <= b and not a;
    layer8_outputs(2257) <= b;
    layer8_outputs(2258) <= not b or a;
    layer8_outputs(2259) <= a xor b;
    layer8_outputs(2260) <= b;
    layer8_outputs(2261) <= not a or b;
    layer8_outputs(2262) <= not a;
    layer8_outputs(2263) <= b;
    layer8_outputs(2264) <= not b or a;
    layer8_outputs(2265) <= not b;
    layer8_outputs(2266) <= a xor b;
    layer8_outputs(2267) <= a and not b;
    layer8_outputs(2268) <= b;
    layer8_outputs(2269) <= a or b;
    layer8_outputs(2270) <= a;
    layer8_outputs(2271) <= a and not b;
    layer8_outputs(2272) <= b;
    layer8_outputs(2273) <= a xor b;
    layer8_outputs(2274) <= b;
    layer8_outputs(2275) <= a and not b;
    layer8_outputs(2276) <= a xor b;
    layer8_outputs(2277) <= a xor b;
    layer8_outputs(2278) <= not b;
    layer8_outputs(2279) <= b and not a;
    layer8_outputs(2280) <= not b;
    layer8_outputs(2281) <= not a;
    layer8_outputs(2282) <= not b;
    layer8_outputs(2283) <= not (a xor b);
    layer8_outputs(2284) <= a xor b;
    layer8_outputs(2285) <= not (a and b);
    layer8_outputs(2286) <= not b;
    layer8_outputs(2287) <= not a;
    layer8_outputs(2288) <= a;
    layer8_outputs(2289) <= not b or a;
    layer8_outputs(2290) <= a and not b;
    layer8_outputs(2291) <= not b;
    layer8_outputs(2292) <= not a;
    layer8_outputs(2293) <= not (a xor b);
    layer8_outputs(2294) <= a or b;
    layer8_outputs(2295) <= a xor b;
    layer8_outputs(2296) <= a or b;
    layer8_outputs(2297) <= not b;
    layer8_outputs(2298) <= not a or b;
    layer8_outputs(2299) <= b;
    layer8_outputs(2300) <= b;
    layer8_outputs(2301) <= a xor b;
    layer8_outputs(2302) <= not a;
    layer8_outputs(2303) <= not b;
    layer8_outputs(2304) <= not b;
    layer8_outputs(2305) <= not (a or b);
    layer8_outputs(2306) <= b;
    layer8_outputs(2307) <= a;
    layer8_outputs(2308) <= b and not a;
    layer8_outputs(2309) <= a;
    layer8_outputs(2310) <= not b;
    layer8_outputs(2311) <= a;
    layer8_outputs(2312) <= not b;
    layer8_outputs(2313) <= b;
    layer8_outputs(2314) <= a;
    layer8_outputs(2315) <= a;
    layer8_outputs(2316) <= a;
    layer8_outputs(2317) <= not (a or b);
    layer8_outputs(2318) <= a xor b;
    layer8_outputs(2319) <= not (a xor b);
    layer8_outputs(2320) <= not b;
    layer8_outputs(2321) <= b;
    layer8_outputs(2322) <= a;
    layer8_outputs(2323) <= b;
    layer8_outputs(2324) <= not b;
    layer8_outputs(2325) <= not a;
    layer8_outputs(2326) <= a xor b;
    layer8_outputs(2327) <= not (a and b);
    layer8_outputs(2328) <= not (a xor b);
    layer8_outputs(2329) <= not a or b;
    layer8_outputs(2330) <= not b;
    layer8_outputs(2331) <= a and b;
    layer8_outputs(2332) <= a xor b;
    layer8_outputs(2333) <= not (a xor b);
    layer8_outputs(2334) <= a;
    layer8_outputs(2335) <= not b;
    layer8_outputs(2336) <= not a;
    layer8_outputs(2337) <= not a;
    layer8_outputs(2338) <= a;
    layer8_outputs(2339) <= a xor b;
    layer8_outputs(2340) <= a or b;
    layer8_outputs(2341) <= a and not b;
    layer8_outputs(2342) <= a;
    layer8_outputs(2343) <= a and b;
    layer8_outputs(2344) <= not b;
    layer8_outputs(2345) <= a or b;
    layer8_outputs(2346) <= not b or a;
    layer8_outputs(2347) <= a;
    layer8_outputs(2348) <= not b;
    layer8_outputs(2349) <= b;
    layer8_outputs(2350) <= not (a xor b);
    layer8_outputs(2351) <= not (a xor b);
    layer8_outputs(2352) <= b;
    layer8_outputs(2353) <= not a;
    layer8_outputs(2354) <= a xor b;
    layer8_outputs(2355) <= a;
    layer8_outputs(2356) <= a xor b;
    layer8_outputs(2357) <= not (a and b);
    layer8_outputs(2358) <= not a;
    layer8_outputs(2359) <= a xor b;
    layer8_outputs(2360) <= not a or b;
    layer8_outputs(2361) <= a xor b;
    layer8_outputs(2362) <= not (a xor b);
    layer8_outputs(2363) <= not b;
    layer8_outputs(2364) <= not a or b;
    layer8_outputs(2365) <= a xor b;
    layer8_outputs(2366) <= not b;
    layer8_outputs(2367) <= b;
    layer8_outputs(2368) <= not (a xor b);
    layer8_outputs(2369) <= a xor b;
    layer8_outputs(2370) <= a or b;
    layer8_outputs(2371) <= a and not b;
    layer8_outputs(2372) <= a and b;
    layer8_outputs(2373) <= a or b;
    layer8_outputs(2374) <= not b;
    layer8_outputs(2375) <= a and b;
    layer8_outputs(2376) <= not (a xor b);
    layer8_outputs(2377) <= not a;
    layer8_outputs(2378) <= not (a xor b);
    layer8_outputs(2379) <= a and not b;
    layer8_outputs(2380) <= not a or b;
    layer8_outputs(2381) <= not (a xor b);
    layer8_outputs(2382) <= a and not b;
    layer8_outputs(2383) <= not (a xor b);
    layer8_outputs(2384) <= not (a and b);
    layer8_outputs(2385) <= not b;
    layer8_outputs(2386) <= a;
    layer8_outputs(2387) <= not a or b;
    layer8_outputs(2388) <= not a or b;
    layer8_outputs(2389) <= a and b;
    layer8_outputs(2390) <= not a;
    layer8_outputs(2391) <= a xor b;
    layer8_outputs(2392) <= not (a or b);
    layer8_outputs(2393) <= a xor b;
    layer8_outputs(2394) <= a xor b;
    layer8_outputs(2395) <= a xor b;
    layer8_outputs(2396) <= a;
    layer8_outputs(2397) <= a;
    layer8_outputs(2398) <= not b;
    layer8_outputs(2399) <= b;
    layer8_outputs(2400) <= a and not b;
    layer8_outputs(2401) <= b and not a;
    layer8_outputs(2402) <= a xor b;
    layer8_outputs(2403) <= a xor b;
    layer8_outputs(2404) <= a;
    layer8_outputs(2405) <= a or b;
    layer8_outputs(2406) <= b;
    layer8_outputs(2407) <= not a;
    layer8_outputs(2408) <= a or b;
    layer8_outputs(2409) <= a and not b;
    layer8_outputs(2410) <= a and not b;
    layer8_outputs(2411) <= not a;
    layer8_outputs(2412) <= not b;
    layer8_outputs(2413) <= not (a xor b);
    layer8_outputs(2414) <= b and not a;
    layer8_outputs(2415) <= not (a xor b);
    layer8_outputs(2416) <= a xor b;
    layer8_outputs(2417) <= not b;
    layer8_outputs(2418) <= not (a or b);
    layer8_outputs(2419) <= not b;
    layer8_outputs(2420) <= not (a and b);
    layer8_outputs(2421) <= 1'b1;
    layer8_outputs(2422) <= a xor b;
    layer8_outputs(2423) <= a;
    layer8_outputs(2424) <= a xor b;
    layer8_outputs(2425) <= a;
    layer8_outputs(2426) <= not (a xor b);
    layer8_outputs(2427) <= not a or b;
    layer8_outputs(2428) <= not a;
    layer8_outputs(2429) <= b;
    layer8_outputs(2430) <= not b;
    layer8_outputs(2431) <= a and not b;
    layer8_outputs(2432) <= not a;
    layer8_outputs(2433) <= not a;
    layer8_outputs(2434) <= not b;
    layer8_outputs(2435) <= a;
    layer8_outputs(2436) <= b;
    layer8_outputs(2437) <= a and not b;
    layer8_outputs(2438) <= not a;
    layer8_outputs(2439) <= not (a xor b);
    layer8_outputs(2440) <= not a;
    layer8_outputs(2441) <= a;
    layer8_outputs(2442) <= not (a xor b);
    layer8_outputs(2443) <= not b;
    layer8_outputs(2444) <= a xor b;
    layer8_outputs(2445) <= not b or a;
    layer8_outputs(2446) <= not a;
    layer8_outputs(2447) <= b;
    layer8_outputs(2448) <= not (a xor b);
    layer8_outputs(2449) <= not a or b;
    layer8_outputs(2450) <= not (a xor b);
    layer8_outputs(2451) <= not a or b;
    layer8_outputs(2452) <= not (a or b);
    layer8_outputs(2453) <= not a or b;
    layer8_outputs(2454) <= a;
    layer8_outputs(2455) <= not b;
    layer8_outputs(2456) <= b and not a;
    layer8_outputs(2457) <= b and not a;
    layer8_outputs(2458) <= a;
    layer8_outputs(2459) <= a xor b;
    layer8_outputs(2460) <= not (a and b);
    layer8_outputs(2461) <= a;
    layer8_outputs(2462) <= a xor b;
    layer8_outputs(2463) <= not b;
    layer8_outputs(2464) <= not (a and b);
    layer8_outputs(2465) <= not (a or b);
    layer8_outputs(2466) <= b and not a;
    layer8_outputs(2467) <= b;
    layer8_outputs(2468) <= a xor b;
    layer8_outputs(2469) <= a xor b;
    layer8_outputs(2470) <= a xor b;
    layer8_outputs(2471) <= a;
    layer8_outputs(2472) <= a;
    layer8_outputs(2473) <= not b;
    layer8_outputs(2474) <= not a;
    layer8_outputs(2475) <= a;
    layer8_outputs(2476) <= b and not a;
    layer8_outputs(2477) <= b;
    layer8_outputs(2478) <= not b;
    layer8_outputs(2479) <= not a or b;
    layer8_outputs(2480) <= a and not b;
    layer8_outputs(2481) <= b and not a;
    layer8_outputs(2482) <= not b;
    layer8_outputs(2483) <= not (a or b);
    layer8_outputs(2484) <= a xor b;
    layer8_outputs(2485) <= not (a and b);
    layer8_outputs(2486) <= not a;
    layer8_outputs(2487) <= not (a or b);
    layer8_outputs(2488) <= a;
    layer8_outputs(2489) <= a;
    layer8_outputs(2490) <= a and b;
    layer8_outputs(2491) <= not a;
    layer8_outputs(2492) <= not a;
    layer8_outputs(2493) <= a and b;
    layer8_outputs(2494) <= b and not a;
    layer8_outputs(2495) <= a xor b;
    layer8_outputs(2496) <= b;
    layer8_outputs(2497) <= a xor b;
    layer8_outputs(2498) <= not (a xor b);
    layer8_outputs(2499) <= b;
    layer8_outputs(2500) <= not (a or b);
    layer8_outputs(2501) <= not (a xor b);
    layer8_outputs(2502) <= b;
    layer8_outputs(2503) <= b;
    layer8_outputs(2504) <= not (a xor b);
    layer8_outputs(2505) <= not a or b;
    layer8_outputs(2506) <= a;
    layer8_outputs(2507) <= not (a xor b);
    layer8_outputs(2508) <= a and b;
    layer8_outputs(2509) <= a;
    layer8_outputs(2510) <= a xor b;
    layer8_outputs(2511) <= not b;
    layer8_outputs(2512) <= b;
    layer8_outputs(2513) <= b and not a;
    layer8_outputs(2514) <= b;
    layer8_outputs(2515) <= not (a xor b);
    layer8_outputs(2516) <= not b;
    layer8_outputs(2517) <= a xor b;
    layer8_outputs(2518) <= a or b;
    layer8_outputs(2519) <= b and not a;
    layer8_outputs(2520) <= b and not a;
    layer8_outputs(2521) <= a and b;
    layer8_outputs(2522) <= a or b;
    layer8_outputs(2523) <= b;
    layer8_outputs(2524) <= a;
    layer8_outputs(2525) <= not b;
    layer8_outputs(2526) <= not (a and b);
    layer8_outputs(2527) <= not (a xor b);
    layer8_outputs(2528) <= a and b;
    layer8_outputs(2529) <= a;
    layer8_outputs(2530) <= not b;
    layer8_outputs(2531) <= not a;
    layer8_outputs(2532) <= not a;
    layer8_outputs(2533) <= a xor b;
    layer8_outputs(2534) <= a or b;
    layer8_outputs(2535) <= not a;
    layer8_outputs(2536) <= not (a xor b);
    layer8_outputs(2537) <= b;
    layer8_outputs(2538) <= a or b;
    layer8_outputs(2539) <= 1'b1;
    layer8_outputs(2540) <= a and not b;
    layer8_outputs(2541) <= not a or b;
    layer8_outputs(2542) <= b;
    layer8_outputs(2543) <= not (a or b);
    layer8_outputs(2544) <= not b;
    layer8_outputs(2545) <= a xor b;
    layer8_outputs(2546) <= a;
    layer8_outputs(2547) <= a xor b;
    layer8_outputs(2548) <= a;
    layer8_outputs(2549) <= a xor b;
    layer8_outputs(2550) <= not (a and b);
    layer8_outputs(2551) <= a or b;
    layer8_outputs(2552) <= b and not a;
    layer8_outputs(2553) <= b;
    layer8_outputs(2554) <= not a;
    layer8_outputs(2555) <= a xor b;
    layer8_outputs(2556) <= not a;
    layer8_outputs(2557) <= not (a xor b);
    layer8_outputs(2558) <= b;
    layer8_outputs(2559) <= a;
    layer8_outputs(2560) <= a;
    layer8_outputs(2561) <= a and b;
    layer8_outputs(2562) <= not (a or b);
    layer8_outputs(2563) <= a xor b;
    layer8_outputs(2564) <= not a;
    layer8_outputs(2565) <= b;
    layer8_outputs(2566) <= a xor b;
    layer8_outputs(2567) <= not (a xor b);
    layer8_outputs(2568) <= a;
    layer8_outputs(2569) <= not (a xor b);
    layer8_outputs(2570) <= a and not b;
    layer8_outputs(2571) <= a and not b;
    layer8_outputs(2572) <= a xor b;
    layer8_outputs(2573) <= not b;
    layer8_outputs(2574) <= not b or a;
    layer8_outputs(2575) <= b;
    layer8_outputs(2576) <= a xor b;
    layer8_outputs(2577) <= not (a xor b);
    layer8_outputs(2578) <= a and not b;
    layer8_outputs(2579) <= not a;
    layer8_outputs(2580) <= a and b;
    layer8_outputs(2581) <= not a;
    layer8_outputs(2582) <= not (a or b);
    layer8_outputs(2583) <= not (a xor b);
    layer8_outputs(2584) <= a;
    layer8_outputs(2585) <= a and b;
    layer8_outputs(2586) <= a and b;
    layer8_outputs(2587) <= not b or a;
    layer8_outputs(2588) <= b and not a;
    layer8_outputs(2589) <= a;
    layer8_outputs(2590) <= a;
    layer8_outputs(2591) <= a and b;
    layer8_outputs(2592) <= not a;
    layer8_outputs(2593) <= a xor b;
    layer8_outputs(2594) <= not (a xor b);
    layer8_outputs(2595) <= not (a xor b);
    layer8_outputs(2596) <= not (a xor b);
    layer8_outputs(2597) <= not a;
    layer8_outputs(2598) <= a xor b;
    layer8_outputs(2599) <= a;
    layer8_outputs(2600) <= not (a xor b);
    layer8_outputs(2601) <= a;
    layer8_outputs(2602) <= a and b;
    layer8_outputs(2603) <= not b or a;
    layer8_outputs(2604) <= b;
    layer8_outputs(2605) <= not a;
    layer8_outputs(2606) <= a;
    layer8_outputs(2607) <= not (a and b);
    layer8_outputs(2608) <= a;
    layer8_outputs(2609) <= not (a xor b);
    layer8_outputs(2610) <= not b or a;
    layer8_outputs(2611) <= not b;
    layer8_outputs(2612) <= a and not b;
    layer8_outputs(2613) <= not b;
    layer8_outputs(2614) <= not (a xor b);
    layer8_outputs(2615) <= not b;
    layer8_outputs(2616) <= a;
    layer8_outputs(2617) <= not b;
    layer8_outputs(2618) <= b and not a;
    layer8_outputs(2619) <= 1'b0;
    layer8_outputs(2620) <= a xor b;
    layer8_outputs(2621) <= a;
    layer8_outputs(2622) <= not a;
    layer8_outputs(2623) <= a xor b;
    layer8_outputs(2624) <= a and b;
    layer8_outputs(2625) <= a xor b;
    layer8_outputs(2626) <= not a;
    layer8_outputs(2627) <= b and not a;
    layer8_outputs(2628) <= b;
    layer8_outputs(2629) <= b;
    layer8_outputs(2630) <= not b;
    layer8_outputs(2631) <= a;
    layer8_outputs(2632) <= not (a xor b);
    layer8_outputs(2633) <= a and not b;
    layer8_outputs(2634) <= b;
    layer8_outputs(2635) <= not b;
    layer8_outputs(2636) <= not (a xor b);
    layer8_outputs(2637) <= a and b;
    layer8_outputs(2638) <= not (a and b);
    layer8_outputs(2639) <= not (a xor b);
    layer8_outputs(2640) <= a or b;
    layer8_outputs(2641) <= not (a and b);
    layer8_outputs(2642) <= a xor b;
    layer8_outputs(2643) <= not a;
    layer8_outputs(2644) <= not a;
    layer8_outputs(2645) <= not b;
    layer8_outputs(2646) <= not b;
    layer8_outputs(2647) <= not (a xor b);
    layer8_outputs(2648) <= a;
    layer8_outputs(2649) <= not b or a;
    layer8_outputs(2650) <= a xor b;
    layer8_outputs(2651) <= not (a or b);
    layer8_outputs(2652) <= not b;
    layer8_outputs(2653) <= a;
    layer8_outputs(2654) <= a and b;
    layer8_outputs(2655) <= a xor b;
    layer8_outputs(2656) <= not a;
    layer8_outputs(2657) <= a and not b;
    layer8_outputs(2658) <= b and not a;
    layer8_outputs(2659) <= not a or b;
    layer8_outputs(2660) <= a xor b;
    layer8_outputs(2661) <= not (a and b);
    layer8_outputs(2662) <= not a;
    layer8_outputs(2663) <= not b;
    layer8_outputs(2664) <= b and not a;
    layer8_outputs(2665) <= not (a or b);
    layer8_outputs(2666) <= not b;
    layer8_outputs(2667) <= not b;
    layer8_outputs(2668) <= not a;
    layer8_outputs(2669) <= not (a and b);
    layer8_outputs(2670) <= a;
    layer8_outputs(2671) <= a xor b;
    layer8_outputs(2672) <= b;
    layer8_outputs(2673) <= a xor b;
    layer8_outputs(2674) <= not (a or b);
    layer8_outputs(2675) <= b;
    layer8_outputs(2676) <= b;
    layer8_outputs(2677) <= a and b;
    layer8_outputs(2678) <= a and not b;
    layer8_outputs(2679) <= a and b;
    layer8_outputs(2680) <= not a;
    layer8_outputs(2681) <= not (a xor b);
    layer8_outputs(2682) <= not b;
    layer8_outputs(2683) <= a xor b;
    layer8_outputs(2684) <= b;
    layer8_outputs(2685) <= not (a xor b);
    layer8_outputs(2686) <= a xor b;
    layer8_outputs(2687) <= a;
    layer8_outputs(2688) <= not a;
    layer8_outputs(2689) <= not (a xor b);
    layer8_outputs(2690) <= not a;
    layer8_outputs(2691) <= not (a xor b);
    layer8_outputs(2692) <= not a or b;
    layer8_outputs(2693) <= b;
    layer8_outputs(2694) <= not a or b;
    layer8_outputs(2695) <= a and not b;
    layer8_outputs(2696) <= not (a or b);
    layer8_outputs(2697) <= 1'b0;
    layer8_outputs(2698) <= not (a xor b);
    layer8_outputs(2699) <= not a;
    layer8_outputs(2700) <= not (a xor b);
    layer8_outputs(2701) <= not (a xor b);
    layer8_outputs(2702) <= a;
    layer8_outputs(2703) <= a and b;
    layer8_outputs(2704) <= not (a or b);
    layer8_outputs(2705) <= a;
    layer8_outputs(2706) <= not (a or b);
    layer8_outputs(2707) <= not (a or b);
    layer8_outputs(2708) <= not (a or b);
    layer8_outputs(2709) <= not (a xor b);
    layer8_outputs(2710) <= not b;
    layer8_outputs(2711) <= a;
    layer8_outputs(2712) <= not (a xor b);
    layer8_outputs(2713) <= not (a xor b);
    layer8_outputs(2714) <= not (a xor b);
    layer8_outputs(2715) <= a xor b;
    layer8_outputs(2716) <= a xor b;
    layer8_outputs(2717) <= not b;
    layer8_outputs(2718) <= a and not b;
    layer8_outputs(2719) <= a xor b;
    layer8_outputs(2720) <= b;
    layer8_outputs(2721) <= a;
    layer8_outputs(2722) <= a;
    layer8_outputs(2723) <= a;
    layer8_outputs(2724) <= a xor b;
    layer8_outputs(2725) <= a and not b;
    layer8_outputs(2726) <= not b;
    layer8_outputs(2727) <= not (a xor b);
    layer8_outputs(2728) <= not a or b;
    layer8_outputs(2729) <= not (a xor b);
    layer8_outputs(2730) <= a or b;
    layer8_outputs(2731) <= not (a xor b);
    layer8_outputs(2732) <= a;
    layer8_outputs(2733) <= not a;
    layer8_outputs(2734) <= a and b;
    layer8_outputs(2735) <= not (a and b);
    layer8_outputs(2736) <= b;
    layer8_outputs(2737) <= not b or a;
    layer8_outputs(2738) <= b;
    layer8_outputs(2739) <= b;
    layer8_outputs(2740) <= not a;
    layer8_outputs(2741) <= a and not b;
    layer8_outputs(2742) <= a;
    layer8_outputs(2743) <= not a;
    layer8_outputs(2744) <= a or b;
    layer8_outputs(2745) <= not b;
    layer8_outputs(2746) <= not b or a;
    layer8_outputs(2747) <= a xor b;
    layer8_outputs(2748) <= not b;
    layer8_outputs(2749) <= not b;
    layer8_outputs(2750) <= a xor b;
    layer8_outputs(2751) <= 1'b0;
    layer8_outputs(2752) <= b;
    layer8_outputs(2753) <= a and not b;
    layer8_outputs(2754) <= b and not a;
    layer8_outputs(2755) <= b;
    layer8_outputs(2756) <= a and not b;
    layer8_outputs(2757) <= not b;
    layer8_outputs(2758) <= a and b;
    layer8_outputs(2759) <= b;
    layer8_outputs(2760) <= a;
    layer8_outputs(2761) <= not (a xor b);
    layer8_outputs(2762) <= b and not a;
    layer8_outputs(2763) <= not (a xor b);
    layer8_outputs(2764) <= a;
    layer8_outputs(2765) <= not (a or b);
    layer8_outputs(2766) <= 1'b0;
    layer8_outputs(2767) <= not (a or b);
    layer8_outputs(2768) <= not (a and b);
    layer8_outputs(2769) <= a;
    layer8_outputs(2770) <= not (a xor b);
    layer8_outputs(2771) <= not b or a;
    layer8_outputs(2772) <= a;
    layer8_outputs(2773) <= not b or a;
    layer8_outputs(2774) <= not b;
    layer8_outputs(2775) <= not a;
    layer8_outputs(2776) <= a and b;
    layer8_outputs(2777) <= b;
    layer8_outputs(2778) <= a;
    layer8_outputs(2779) <= a and not b;
    layer8_outputs(2780) <= a;
    layer8_outputs(2781) <= a xor b;
    layer8_outputs(2782) <= not a;
    layer8_outputs(2783) <= b;
    layer8_outputs(2784) <= not (a and b);
    layer8_outputs(2785) <= b and not a;
    layer8_outputs(2786) <= not (a xor b);
    layer8_outputs(2787) <= a xor b;
    layer8_outputs(2788) <= not b;
    layer8_outputs(2789) <= not a;
    layer8_outputs(2790) <= b;
    layer8_outputs(2791) <= b and not a;
    layer8_outputs(2792) <= b;
    layer8_outputs(2793) <= not (a xor b);
    layer8_outputs(2794) <= not (a xor b);
    layer8_outputs(2795) <= not b;
    layer8_outputs(2796) <= b;
    layer8_outputs(2797) <= not (a xor b);
    layer8_outputs(2798) <= a;
    layer8_outputs(2799) <= not (a xor b);
    layer8_outputs(2800) <= not (a xor b);
    layer8_outputs(2801) <= b;
    layer8_outputs(2802) <= b and not a;
    layer8_outputs(2803) <= not a;
    layer8_outputs(2804) <= not (a or b);
    layer8_outputs(2805) <= not (a or b);
    layer8_outputs(2806) <= a and b;
    layer8_outputs(2807) <= not b;
    layer8_outputs(2808) <= not b;
    layer8_outputs(2809) <= a and b;
    layer8_outputs(2810) <= a;
    layer8_outputs(2811) <= not (a and b);
    layer8_outputs(2812) <= not (a and b);
    layer8_outputs(2813) <= a;
    layer8_outputs(2814) <= not (a xor b);
    layer8_outputs(2815) <= not b;
    layer8_outputs(2816) <= not a;
    layer8_outputs(2817) <= b;
    layer8_outputs(2818) <= b;
    layer8_outputs(2819) <= not b or a;
    layer8_outputs(2820) <= not (a xor b);
    layer8_outputs(2821) <= not b or a;
    layer8_outputs(2822) <= a and b;
    layer8_outputs(2823) <= not b;
    layer8_outputs(2824) <= b;
    layer8_outputs(2825) <= a;
    layer8_outputs(2826) <= a;
    layer8_outputs(2827) <= a xor b;
    layer8_outputs(2828) <= a and b;
    layer8_outputs(2829) <= b;
    layer8_outputs(2830) <= not b;
    layer8_outputs(2831) <= not b;
    layer8_outputs(2832) <= not a or b;
    layer8_outputs(2833) <= a;
    layer8_outputs(2834) <= not (a xor b);
    layer8_outputs(2835) <= not (a xor b);
    layer8_outputs(2836) <= not (a xor b);
    layer8_outputs(2837) <= a and b;
    layer8_outputs(2838) <= not a;
    layer8_outputs(2839) <= not b;
    layer8_outputs(2840) <= not b or a;
    layer8_outputs(2841) <= b;
    layer8_outputs(2842) <= not (a and b);
    layer8_outputs(2843) <= a xor b;
    layer8_outputs(2844) <= not (a xor b);
    layer8_outputs(2845) <= 1'b1;
    layer8_outputs(2846) <= a and b;
    layer8_outputs(2847) <= a xor b;
    layer8_outputs(2848) <= not b;
    layer8_outputs(2849) <= a;
    layer8_outputs(2850) <= b and not a;
    layer8_outputs(2851) <= b;
    layer8_outputs(2852) <= not b;
    layer8_outputs(2853) <= a;
    layer8_outputs(2854) <= not a;
    layer8_outputs(2855) <= a xor b;
    layer8_outputs(2856) <= a;
    layer8_outputs(2857) <= a and not b;
    layer8_outputs(2858) <= not a;
    layer8_outputs(2859) <= not b;
    layer8_outputs(2860) <= b;
    layer8_outputs(2861) <= not (a xor b);
    layer8_outputs(2862) <= a or b;
    layer8_outputs(2863) <= b;
    layer8_outputs(2864) <= not (a xor b);
    layer8_outputs(2865) <= a or b;
    layer8_outputs(2866) <= not b;
    layer8_outputs(2867) <= not a;
    layer8_outputs(2868) <= b and not a;
    layer8_outputs(2869) <= 1'b1;
    layer8_outputs(2870) <= not a;
    layer8_outputs(2871) <= not b;
    layer8_outputs(2872) <= a and not b;
    layer8_outputs(2873) <= not b;
    layer8_outputs(2874) <= b;
    layer8_outputs(2875) <= b;
    layer8_outputs(2876) <= not b;
    layer8_outputs(2877) <= not b;
    layer8_outputs(2878) <= not (a and b);
    layer8_outputs(2879) <= not b;
    layer8_outputs(2880) <= not (a or b);
    layer8_outputs(2881) <= a;
    layer8_outputs(2882) <= b;
    layer8_outputs(2883) <= not (a or b);
    layer8_outputs(2884) <= not b;
    layer8_outputs(2885) <= b;
    layer8_outputs(2886) <= b and not a;
    layer8_outputs(2887) <= not a;
    layer8_outputs(2888) <= b and not a;
    layer8_outputs(2889) <= not (a and b);
    layer8_outputs(2890) <= b;
    layer8_outputs(2891) <= a xor b;
    layer8_outputs(2892) <= a and not b;
    layer8_outputs(2893) <= not b;
    layer8_outputs(2894) <= a xor b;
    layer8_outputs(2895) <= not (a xor b);
    layer8_outputs(2896) <= a;
    layer8_outputs(2897) <= a and b;
    layer8_outputs(2898) <= not a;
    layer8_outputs(2899) <= a;
    layer8_outputs(2900) <= not (a xor b);
    layer8_outputs(2901) <= not (a xor b);
    layer8_outputs(2902) <= not b or a;
    layer8_outputs(2903) <= b and not a;
    layer8_outputs(2904) <= not a;
    layer8_outputs(2905) <= not a;
    layer8_outputs(2906) <= a;
    layer8_outputs(2907) <= a xor b;
    layer8_outputs(2908) <= not a or b;
    layer8_outputs(2909) <= b;
    layer8_outputs(2910) <= a xor b;
    layer8_outputs(2911) <= not b;
    layer8_outputs(2912) <= a;
    layer8_outputs(2913) <= a and b;
    layer8_outputs(2914) <= a xor b;
    layer8_outputs(2915) <= not a;
    layer8_outputs(2916) <= b;
    layer8_outputs(2917) <= not (a xor b);
    layer8_outputs(2918) <= b;
    layer8_outputs(2919) <= not b or a;
    layer8_outputs(2920) <= 1'b0;
    layer8_outputs(2921) <= a xor b;
    layer8_outputs(2922) <= b;
    layer8_outputs(2923) <= not b;
    layer8_outputs(2924) <= b;
    layer8_outputs(2925) <= not (a xor b);
    layer8_outputs(2926) <= b and not a;
    layer8_outputs(2927) <= not a;
    layer8_outputs(2928) <= not (a or b);
    layer8_outputs(2929) <= not a;
    layer8_outputs(2930) <= a;
    layer8_outputs(2931) <= not b or a;
    layer8_outputs(2932) <= a and not b;
    layer8_outputs(2933) <= not b;
    layer8_outputs(2934) <= not (a xor b);
    layer8_outputs(2935) <= 1'b0;
    layer8_outputs(2936) <= not (a and b);
    layer8_outputs(2937) <= not a;
    layer8_outputs(2938) <= a;
    layer8_outputs(2939) <= a and not b;
    layer8_outputs(2940) <= a;
    layer8_outputs(2941) <= b;
    layer8_outputs(2942) <= not b or a;
    layer8_outputs(2943) <= not (a and b);
    layer8_outputs(2944) <= a;
    layer8_outputs(2945) <= a xor b;
    layer8_outputs(2946) <= b and not a;
    layer8_outputs(2947) <= a;
    layer8_outputs(2948) <= not (a xor b);
    layer8_outputs(2949) <= a and not b;
    layer8_outputs(2950) <= not a or b;
    layer8_outputs(2951) <= not a;
    layer8_outputs(2952) <= not a;
    layer8_outputs(2953) <= not a;
    layer8_outputs(2954) <= b;
    layer8_outputs(2955) <= not (a and b);
    layer8_outputs(2956) <= a;
    layer8_outputs(2957) <= b;
    layer8_outputs(2958) <= not a;
    layer8_outputs(2959) <= not (a and b);
    layer8_outputs(2960) <= not b or a;
    layer8_outputs(2961) <= not b or a;
    layer8_outputs(2962) <= b and not a;
    layer8_outputs(2963) <= a;
    layer8_outputs(2964) <= not (a xor b);
    layer8_outputs(2965) <= not a or b;
    layer8_outputs(2966) <= not b;
    layer8_outputs(2967) <= b;
    layer8_outputs(2968) <= b and not a;
    layer8_outputs(2969) <= not b;
    layer8_outputs(2970) <= a xor b;
    layer8_outputs(2971) <= b;
    layer8_outputs(2972) <= not a;
    layer8_outputs(2973) <= b and not a;
    layer8_outputs(2974) <= not (a and b);
    layer8_outputs(2975) <= not b;
    layer8_outputs(2976) <= a or b;
    layer8_outputs(2977) <= not b;
    layer8_outputs(2978) <= not (a xor b);
    layer8_outputs(2979) <= not a;
    layer8_outputs(2980) <= not b;
    layer8_outputs(2981) <= not b or a;
    layer8_outputs(2982) <= not (a xor b);
    layer8_outputs(2983) <= not (a xor b);
    layer8_outputs(2984) <= not (a xor b);
    layer8_outputs(2985) <= b;
    layer8_outputs(2986) <= not a;
    layer8_outputs(2987) <= not a;
    layer8_outputs(2988) <= a;
    layer8_outputs(2989) <= not (a or b);
    layer8_outputs(2990) <= not a;
    layer8_outputs(2991) <= b;
    layer8_outputs(2992) <= not (a and b);
    layer8_outputs(2993) <= a xor b;
    layer8_outputs(2994) <= not b or a;
    layer8_outputs(2995) <= not a;
    layer8_outputs(2996) <= not (a xor b);
    layer8_outputs(2997) <= not a or b;
    layer8_outputs(2998) <= a xor b;
    layer8_outputs(2999) <= not a or b;
    layer8_outputs(3000) <= a or b;
    layer8_outputs(3001) <= not (a xor b);
    layer8_outputs(3002) <= a or b;
    layer8_outputs(3003) <= b and not a;
    layer8_outputs(3004) <= a and not b;
    layer8_outputs(3005) <= not b or a;
    layer8_outputs(3006) <= b and not a;
    layer8_outputs(3007) <= a xor b;
    layer8_outputs(3008) <= not (a and b);
    layer8_outputs(3009) <= not a or b;
    layer8_outputs(3010) <= not (a xor b);
    layer8_outputs(3011) <= not (a xor b);
    layer8_outputs(3012) <= not b;
    layer8_outputs(3013) <= not (a xor b);
    layer8_outputs(3014) <= not (a and b);
    layer8_outputs(3015) <= a and b;
    layer8_outputs(3016) <= a;
    layer8_outputs(3017) <= a xor b;
    layer8_outputs(3018) <= not b or a;
    layer8_outputs(3019) <= not (a xor b);
    layer8_outputs(3020) <= a xor b;
    layer8_outputs(3021) <= b;
    layer8_outputs(3022) <= not b or a;
    layer8_outputs(3023) <= b;
    layer8_outputs(3024) <= not a;
    layer8_outputs(3025) <= not (a and b);
    layer8_outputs(3026) <= 1'b1;
    layer8_outputs(3027) <= not b or a;
    layer8_outputs(3028) <= not b;
    layer8_outputs(3029) <= b;
    layer8_outputs(3030) <= not a or b;
    layer8_outputs(3031) <= not b;
    layer8_outputs(3032) <= not a or b;
    layer8_outputs(3033) <= not a;
    layer8_outputs(3034) <= b;
    layer8_outputs(3035) <= a or b;
    layer8_outputs(3036) <= not a;
    layer8_outputs(3037) <= a;
    layer8_outputs(3038) <= a xor b;
    layer8_outputs(3039) <= not (a or b);
    layer8_outputs(3040) <= not (a xor b);
    layer8_outputs(3041) <= not b;
    layer8_outputs(3042) <= not (a xor b);
    layer8_outputs(3043) <= b;
    layer8_outputs(3044) <= a or b;
    layer8_outputs(3045) <= not a or b;
    layer8_outputs(3046) <= not a;
    layer8_outputs(3047) <= b;
    layer8_outputs(3048) <= b;
    layer8_outputs(3049) <= b;
    layer8_outputs(3050) <= not (a xor b);
    layer8_outputs(3051) <= a xor b;
    layer8_outputs(3052) <= not (a and b);
    layer8_outputs(3053) <= a and not b;
    layer8_outputs(3054) <= a and not b;
    layer8_outputs(3055) <= not (a and b);
    layer8_outputs(3056) <= not (a and b);
    layer8_outputs(3057) <= a and b;
    layer8_outputs(3058) <= a;
    layer8_outputs(3059) <= a xor b;
    layer8_outputs(3060) <= a;
    layer8_outputs(3061) <= not b;
    layer8_outputs(3062) <= not b;
    layer8_outputs(3063) <= b;
    layer8_outputs(3064) <= not (a xor b);
    layer8_outputs(3065) <= not (a xor b);
    layer8_outputs(3066) <= not (a xor b);
    layer8_outputs(3067) <= not b;
    layer8_outputs(3068) <= not (a or b);
    layer8_outputs(3069) <= not (a xor b);
    layer8_outputs(3070) <= not a;
    layer8_outputs(3071) <= a and not b;
    layer8_outputs(3072) <= not a;
    layer8_outputs(3073) <= a;
    layer8_outputs(3074) <= a xor b;
    layer8_outputs(3075) <= not b;
    layer8_outputs(3076) <= a;
    layer8_outputs(3077) <= not a;
    layer8_outputs(3078) <= a;
    layer8_outputs(3079) <= a and b;
    layer8_outputs(3080) <= not b or a;
    layer8_outputs(3081) <= b and not a;
    layer8_outputs(3082) <= not (a and b);
    layer8_outputs(3083) <= not (a or b);
    layer8_outputs(3084) <= not b;
    layer8_outputs(3085) <= b;
    layer8_outputs(3086) <= a xor b;
    layer8_outputs(3087) <= b;
    layer8_outputs(3088) <= b;
    layer8_outputs(3089) <= a xor b;
    layer8_outputs(3090) <= b;
    layer8_outputs(3091) <= not b or a;
    layer8_outputs(3092) <= not a or b;
    layer8_outputs(3093) <= a;
    layer8_outputs(3094) <= a and b;
    layer8_outputs(3095) <= not b or a;
    layer8_outputs(3096) <= b;
    layer8_outputs(3097) <= b;
    layer8_outputs(3098) <= b;
    layer8_outputs(3099) <= not b or a;
    layer8_outputs(3100) <= b;
    layer8_outputs(3101) <= not b or a;
    layer8_outputs(3102) <= not a;
    layer8_outputs(3103) <= not (a xor b);
    layer8_outputs(3104) <= not a or b;
    layer8_outputs(3105) <= not (a xor b);
    layer8_outputs(3106) <= not (a xor b);
    layer8_outputs(3107) <= b;
    layer8_outputs(3108) <= a and not b;
    layer8_outputs(3109) <= a or b;
    layer8_outputs(3110) <= a and b;
    layer8_outputs(3111) <= a;
    layer8_outputs(3112) <= a and not b;
    layer8_outputs(3113) <= b and not a;
    layer8_outputs(3114) <= a or b;
    layer8_outputs(3115) <= a and b;
    layer8_outputs(3116) <= a;
    layer8_outputs(3117) <= b;
    layer8_outputs(3118) <= not (a xor b);
    layer8_outputs(3119) <= a and b;
    layer8_outputs(3120) <= b and not a;
    layer8_outputs(3121) <= not (a and b);
    layer8_outputs(3122) <= not a;
    layer8_outputs(3123) <= not (a xor b);
    layer8_outputs(3124) <= not b;
    layer8_outputs(3125) <= a xor b;
    layer8_outputs(3126) <= not a;
    layer8_outputs(3127) <= not b;
    layer8_outputs(3128) <= a or b;
    layer8_outputs(3129) <= b and not a;
    layer8_outputs(3130) <= a;
    layer8_outputs(3131) <= a;
    layer8_outputs(3132) <= a or b;
    layer8_outputs(3133) <= not b or a;
    layer8_outputs(3134) <= not (a xor b);
    layer8_outputs(3135) <= not a;
    layer8_outputs(3136) <= not b or a;
    layer8_outputs(3137) <= a;
    layer8_outputs(3138) <= not b;
    layer8_outputs(3139) <= a or b;
    layer8_outputs(3140) <= not b or a;
    layer8_outputs(3141) <= b;
    layer8_outputs(3142) <= not b or a;
    layer8_outputs(3143) <= b;
    layer8_outputs(3144) <= not b;
    layer8_outputs(3145) <= b;
    layer8_outputs(3146) <= not b;
    layer8_outputs(3147) <= b;
    layer8_outputs(3148) <= a xor b;
    layer8_outputs(3149) <= a;
    layer8_outputs(3150) <= not (a xor b);
    layer8_outputs(3151) <= not a;
    layer8_outputs(3152) <= not (a xor b);
    layer8_outputs(3153) <= not (a and b);
    layer8_outputs(3154) <= a and not b;
    layer8_outputs(3155) <= b;
    layer8_outputs(3156) <= not (a and b);
    layer8_outputs(3157) <= not (a xor b);
    layer8_outputs(3158) <= not a;
    layer8_outputs(3159) <= not a;
    layer8_outputs(3160) <= a xor b;
    layer8_outputs(3161) <= not (a and b);
    layer8_outputs(3162) <= a or b;
    layer8_outputs(3163) <= not a;
    layer8_outputs(3164) <= not a;
    layer8_outputs(3165) <= b;
    layer8_outputs(3166) <= not (a xor b);
    layer8_outputs(3167) <= b and not a;
    layer8_outputs(3168) <= not (a xor b);
    layer8_outputs(3169) <= b;
    layer8_outputs(3170) <= not b;
    layer8_outputs(3171) <= a and not b;
    layer8_outputs(3172) <= not a;
    layer8_outputs(3173) <= not (a xor b);
    layer8_outputs(3174) <= not b;
    layer8_outputs(3175) <= a and not b;
    layer8_outputs(3176) <= b and not a;
    layer8_outputs(3177) <= a and not b;
    layer8_outputs(3178) <= not (a xor b);
    layer8_outputs(3179) <= not (a and b);
    layer8_outputs(3180) <= a xor b;
    layer8_outputs(3181) <= not b;
    layer8_outputs(3182) <= not (a xor b);
    layer8_outputs(3183) <= b;
    layer8_outputs(3184) <= a;
    layer8_outputs(3185) <= b;
    layer8_outputs(3186) <= a;
    layer8_outputs(3187) <= b;
    layer8_outputs(3188) <= not (a xor b);
    layer8_outputs(3189) <= a;
    layer8_outputs(3190) <= not (a or b);
    layer8_outputs(3191) <= not (a xor b);
    layer8_outputs(3192) <= a xor b;
    layer8_outputs(3193) <= a xor b;
    layer8_outputs(3194) <= not b or a;
    layer8_outputs(3195) <= b and not a;
    layer8_outputs(3196) <= not a;
    layer8_outputs(3197) <= a;
    layer8_outputs(3198) <= a xor b;
    layer8_outputs(3199) <= not b;
    layer8_outputs(3200) <= not a;
    layer8_outputs(3201) <= not (a and b);
    layer8_outputs(3202) <= not (a and b);
    layer8_outputs(3203) <= not (a xor b);
    layer8_outputs(3204) <= not a;
    layer8_outputs(3205) <= b and not a;
    layer8_outputs(3206) <= 1'b1;
    layer8_outputs(3207) <= not a or b;
    layer8_outputs(3208) <= not (a or b);
    layer8_outputs(3209) <= a or b;
    layer8_outputs(3210) <= not (a and b);
    layer8_outputs(3211) <= a;
    layer8_outputs(3212) <= not b;
    layer8_outputs(3213) <= b;
    layer8_outputs(3214) <= a xor b;
    layer8_outputs(3215) <= not b;
    layer8_outputs(3216) <= b;
    layer8_outputs(3217) <= b;
    layer8_outputs(3218) <= a and not b;
    layer8_outputs(3219) <= not (a xor b);
    layer8_outputs(3220) <= not b;
    layer8_outputs(3221) <= not (a xor b);
    layer8_outputs(3222) <= not b;
    layer8_outputs(3223) <= a;
    layer8_outputs(3224) <= not a;
    layer8_outputs(3225) <= a;
    layer8_outputs(3226) <= not a or b;
    layer8_outputs(3227) <= not a;
    layer8_outputs(3228) <= not (a or b);
    layer8_outputs(3229) <= not b;
    layer8_outputs(3230) <= a;
    layer8_outputs(3231) <= a xor b;
    layer8_outputs(3232) <= not a or b;
    layer8_outputs(3233) <= a and not b;
    layer8_outputs(3234) <= b;
    layer8_outputs(3235) <= not a or b;
    layer8_outputs(3236) <= a and b;
    layer8_outputs(3237) <= a;
    layer8_outputs(3238) <= not (a xor b);
    layer8_outputs(3239) <= 1'b0;
    layer8_outputs(3240) <= b;
    layer8_outputs(3241) <= not (a and b);
    layer8_outputs(3242) <= a;
    layer8_outputs(3243) <= a;
    layer8_outputs(3244) <= not (a and b);
    layer8_outputs(3245) <= not (a xor b);
    layer8_outputs(3246) <= not (a xor b);
    layer8_outputs(3247) <= not b;
    layer8_outputs(3248) <= not a;
    layer8_outputs(3249) <= not b;
    layer8_outputs(3250) <= not (a or b);
    layer8_outputs(3251) <= a xor b;
    layer8_outputs(3252) <= not (a xor b);
    layer8_outputs(3253) <= b;
    layer8_outputs(3254) <= not b or a;
    layer8_outputs(3255) <= b;
    layer8_outputs(3256) <= not (a and b);
    layer8_outputs(3257) <= 1'b1;
    layer8_outputs(3258) <= not (a xor b);
    layer8_outputs(3259) <= b and not a;
    layer8_outputs(3260) <= not (a xor b);
    layer8_outputs(3261) <= not a;
    layer8_outputs(3262) <= b;
    layer8_outputs(3263) <= a or b;
    layer8_outputs(3264) <= not b or a;
    layer8_outputs(3265) <= 1'b0;
    layer8_outputs(3266) <= not b;
    layer8_outputs(3267) <= a xor b;
    layer8_outputs(3268) <= a or b;
    layer8_outputs(3269) <= a;
    layer8_outputs(3270) <= not b;
    layer8_outputs(3271) <= not b;
    layer8_outputs(3272) <= not (a xor b);
    layer8_outputs(3273) <= a xor b;
    layer8_outputs(3274) <= a and b;
    layer8_outputs(3275) <= not a;
    layer8_outputs(3276) <= not b;
    layer8_outputs(3277) <= a xor b;
    layer8_outputs(3278) <= not (a xor b);
    layer8_outputs(3279) <= 1'b0;
    layer8_outputs(3280) <= not b;
    layer8_outputs(3281) <= a;
    layer8_outputs(3282) <= b;
    layer8_outputs(3283) <= not a;
    layer8_outputs(3284) <= not (a xor b);
    layer8_outputs(3285) <= b;
    layer8_outputs(3286) <= not (a or b);
    layer8_outputs(3287) <= not (a xor b);
    layer8_outputs(3288) <= not b;
    layer8_outputs(3289) <= not (a xor b);
    layer8_outputs(3290) <= b;
    layer8_outputs(3291) <= not a;
    layer8_outputs(3292) <= not b;
    layer8_outputs(3293) <= a;
    layer8_outputs(3294) <= not (a xor b);
    layer8_outputs(3295) <= a;
    layer8_outputs(3296) <= a;
    layer8_outputs(3297) <= b;
    layer8_outputs(3298) <= a xor b;
    layer8_outputs(3299) <= not (a and b);
    layer8_outputs(3300) <= not (a xor b);
    layer8_outputs(3301) <= not (a xor b);
    layer8_outputs(3302) <= not (a xor b);
    layer8_outputs(3303) <= a or b;
    layer8_outputs(3304) <= b;
    layer8_outputs(3305) <= b;
    layer8_outputs(3306) <= a and not b;
    layer8_outputs(3307) <= not a or b;
    layer8_outputs(3308) <= b;
    layer8_outputs(3309) <= a;
    layer8_outputs(3310) <= not a;
    layer8_outputs(3311) <= a;
    layer8_outputs(3312) <= not (a xor b);
    layer8_outputs(3313) <= a xor b;
    layer8_outputs(3314) <= a or b;
    layer8_outputs(3315) <= b and not a;
    layer8_outputs(3316) <= a and not b;
    layer8_outputs(3317) <= a or b;
    layer8_outputs(3318) <= not (a xor b);
    layer8_outputs(3319) <= b;
    layer8_outputs(3320) <= a and b;
    layer8_outputs(3321) <= a;
    layer8_outputs(3322) <= a and not b;
    layer8_outputs(3323) <= a;
    layer8_outputs(3324) <= a xor b;
    layer8_outputs(3325) <= not (a or b);
    layer8_outputs(3326) <= a or b;
    layer8_outputs(3327) <= a xor b;
    layer8_outputs(3328) <= a;
    layer8_outputs(3329) <= b;
    layer8_outputs(3330) <= a;
    layer8_outputs(3331) <= not a;
    layer8_outputs(3332) <= not b or a;
    layer8_outputs(3333) <= a or b;
    layer8_outputs(3334) <= not b;
    layer8_outputs(3335) <= b;
    layer8_outputs(3336) <= not (a or b);
    layer8_outputs(3337) <= not (a xor b);
    layer8_outputs(3338) <= 1'b0;
    layer8_outputs(3339) <= 1'b1;
    layer8_outputs(3340) <= not (a or b);
    layer8_outputs(3341) <= not b;
    layer8_outputs(3342) <= not (a xor b);
    layer8_outputs(3343) <= not (a xor b);
    layer8_outputs(3344) <= not b;
    layer8_outputs(3345) <= not b or a;
    layer8_outputs(3346) <= a xor b;
    layer8_outputs(3347) <= not b;
    layer8_outputs(3348) <= not (a or b);
    layer8_outputs(3349) <= not (a xor b);
    layer8_outputs(3350) <= a xor b;
    layer8_outputs(3351) <= a;
    layer8_outputs(3352) <= not a;
    layer8_outputs(3353) <= not (a xor b);
    layer8_outputs(3354) <= b;
    layer8_outputs(3355) <= a and b;
    layer8_outputs(3356) <= 1'b0;
    layer8_outputs(3357) <= not a;
    layer8_outputs(3358) <= b;
    layer8_outputs(3359) <= a xor b;
    layer8_outputs(3360) <= a and not b;
    layer8_outputs(3361) <= not b;
    layer8_outputs(3362) <= a xor b;
    layer8_outputs(3363) <= b and not a;
    layer8_outputs(3364) <= not a;
    layer8_outputs(3365) <= not a or b;
    layer8_outputs(3366) <= not b;
    layer8_outputs(3367) <= a;
    layer8_outputs(3368) <= not (a xor b);
    layer8_outputs(3369) <= b;
    layer8_outputs(3370) <= not b or a;
    layer8_outputs(3371) <= b;
    layer8_outputs(3372) <= not a;
    layer8_outputs(3373) <= b;
    layer8_outputs(3374) <= not a;
    layer8_outputs(3375) <= not (a and b);
    layer8_outputs(3376) <= b;
    layer8_outputs(3377) <= not b;
    layer8_outputs(3378) <= a xor b;
    layer8_outputs(3379) <= not a;
    layer8_outputs(3380) <= not a or b;
    layer8_outputs(3381) <= not (a xor b);
    layer8_outputs(3382) <= not a;
    layer8_outputs(3383) <= not b or a;
    layer8_outputs(3384) <= a;
    layer8_outputs(3385) <= not a or b;
    layer8_outputs(3386) <= not (a and b);
    layer8_outputs(3387) <= a xor b;
    layer8_outputs(3388) <= a;
    layer8_outputs(3389) <= b;
    layer8_outputs(3390) <= a xor b;
    layer8_outputs(3391) <= b;
    layer8_outputs(3392) <= a xor b;
    layer8_outputs(3393) <= a or b;
    layer8_outputs(3394) <= a or b;
    layer8_outputs(3395) <= a;
    layer8_outputs(3396) <= not b;
    layer8_outputs(3397) <= a xor b;
    layer8_outputs(3398) <= a xor b;
    layer8_outputs(3399) <= not b;
    layer8_outputs(3400) <= not (a xor b);
    layer8_outputs(3401) <= not b;
    layer8_outputs(3402) <= not (a and b);
    layer8_outputs(3403) <= a and not b;
    layer8_outputs(3404) <= a;
    layer8_outputs(3405) <= a and not b;
    layer8_outputs(3406) <= not (a xor b);
    layer8_outputs(3407) <= not b;
    layer8_outputs(3408) <= not b;
    layer8_outputs(3409) <= a and b;
    layer8_outputs(3410) <= not b;
    layer8_outputs(3411) <= a and b;
    layer8_outputs(3412) <= not a or b;
    layer8_outputs(3413) <= not b;
    layer8_outputs(3414) <= not (a xor b);
    layer8_outputs(3415) <= b and not a;
    layer8_outputs(3416) <= a and not b;
    layer8_outputs(3417) <= not (a and b);
    layer8_outputs(3418) <= not (a xor b);
    layer8_outputs(3419) <= a and not b;
    layer8_outputs(3420) <= not (a and b);
    layer8_outputs(3421) <= a xor b;
    layer8_outputs(3422) <= not (a xor b);
    layer8_outputs(3423) <= b and not a;
    layer8_outputs(3424) <= not (a and b);
    layer8_outputs(3425) <= 1'b1;
    layer8_outputs(3426) <= not a;
    layer8_outputs(3427) <= a and b;
    layer8_outputs(3428) <= a or b;
    layer8_outputs(3429) <= a and not b;
    layer8_outputs(3430) <= not b;
    layer8_outputs(3431) <= a xor b;
    layer8_outputs(3432) <= a;
    layer8_outputs(3433) <= not b or a;
    layer8_outputs(3434) <= a;
    layer8_outputs(3435) <= not (a xor b);
    layer8_outputs(3436) <= not b;
    layer8_outputs(3437) <= not a;
    layer8_outputs(3438) <= b and not a;
    layer8_outputs(3439) <= not b or a;
    layer8_outputs(3440) <= not a;
    layer8_outputs(3441) <= not b or a;
    layer8_outputs(3442) <= not (a xor b);
    layer8_outputs(3443) <= a;
    layer8_outputs(3444) <= a xor b;
    layer8_outputs(3445) <= a and b;
    layer8_outputs(3446) <= not b;
    layer8_outputs(3447) <= a xor b;
    layer8_outputs(3448) <= not (a xor b);
    layer8_outputs(3449) <= a and b;
    layer8_outputs(3450) <= not (a or b);
    layer8_outputs(3451) <= not (a or b);
    layer8_outputs(3452) <= not (a xor b);
    layer8_outputs(3453) <= not b or a;
    layer8_outputs(3454) <= not a or b;
    layer8_outputs(3455) <= a;
    layer8_outputs(3456) <= b and not a;
    layer8_outputs(3457) <= a;
    layer8_outputs(3458) <= not (a and b);
    layer8_outputs(3459) <= not a;
    layer8_outputs(3460) <= a xor b;
    layer8_outputs(3461) <= a xor b;
    layer8_outputs(3462) <= not a;
    layer8_outputs(3463) <= a;
    layer8_outputs(3464) <= a or b;
    layer8_outputs(3465) <= not b;
    layer8_outputs(3466) <= not b or a;
    layer8_outputs(3467) <= a;
    layer8_outputs(3468) <= not b;
    layer8_outputs(3469) <= not (a xor b);
    layer8_outputs(3470) <= not b;
    layer8_outputs(3471) <= a and not b;
    layer8_outputs(3472) <= a;
    layer8_outputs(3473) <= a;
    layer8_outputs(3474) <= a;
    layer8_outputs(3475) <= a or b;
    layer8_outputs(3476) <= not a;
    layer8_outputs(3477) <= a xor b;
    layer8_outputs(3478) <= not (a xor b);
    layer8_outputs(3479) <= not a;
    layer8_outputs(3480) <= a or b;
    layer8_outputs(3481) <= b;
    layer8_outputs(3482) <= not a;
    layer8_outputs(3483) <= a xor b;
    layer8_outputs(3484) <= not a;
    layer8_outputs(3485) <= not (a xor b);
    layer8_outputs(3486) <= not b or a;
    layer8_outputs(3487) <= not a or b;
    layer8_outputs(3488) <= b;
    layer8_outputs(3489) <= not b;
    layer8_outputs(3490) <= a;
    layer8_outputs(3491) <= not (a xor b);
    layer8_outputs(3492) <= b;
    layer8_outputs(3493) <= b;
    layer8_outputs(3494) <= not b;
    layer8_outputs(3495) <= not a or b;
    layer8_outputs(3496) <= not a;
    layer8_outputs(3497) <= not (a or b);
    layer8_outputs(3498) <= not b;
    layer8_outputs(3499) <= not (a xor b);
    layer8_outputs(3500) <= b and not a;
    layer8_outputs(3501) <= a xor b;
    layer8_outputs(3502) <= a xor b;
    layer8_outputs(3503) <= b;
    layer8_outputs(3504) <= not a or b;
    layer8_outputs(3505) <= b and not a;
    layer8_outputs(3506) <= a xor b;
    layer8_outputs(3507) <= not (a xor b);
    layer8_outputs(3508) <= not a or b;
    layer8_outputs(3509) <= b and not a;
    layer8_outputs(3510) <= not (a and b);
    layer8_outputs(3511) <= not a or b;
    layer8_outputs(3512) <= a;
    layer8_outputs(3513) <= not a;
    layer8_outputs(3514) <= not a or b;
    layer8_outputs(3515) <= not b;
    layer8_outputs(3516) <= not b;
    layer8_outputs(3517) <= a;
    layer8_outputs(3518) <= a and not b;
    layer8_outputs(3519) <= not a or b;
    layer8_outputs(3520) <= not (a or b);
    layer8_outputs(3521) <= not b or a;
    layer8_outputs(3522) <= a;
    layer8_outputs(3523) <= b;
    layer8_outputs(3524) <= 1'b1;
    layer8_outputs(3525) <= a or b;
    layer8_outputs(3526) <= b;
    layer8_outputs(3527) <= not (a or b);
    layer8_outputs(3528) <= not a;
    layer8_outputs(3529) <= a;
    layer8_outputs(3530) <= not a;
    layer8_outputs(3531) <= a xor b;
    layer8_outputs(3532) <= not b or a;
    layer8_outputs(3533) <= not b or a;
    layer8_outputs(3534) <= a and b;
    layer8_outputs(3535) <= a xor b;
    layer8_outputs(3536) <= a;
    layer8_outputs(3537) <= a or b;
    layer8_outputs(3538) <= not a;
    layer8_outputs(3539) <= not a or b;
    layer8_outputs(3540) <= not b or a;
    layer8_outputs(3541) <= b;
    layer8_outputs(3542) <= a and b;
    layer8_outputs(3543) <= a and b;
    layer8_outputs(3544) <= not b or a;
    layer8_outputs(3545) <= not (a or b);
    layer8_outputs(3546) <= not b;
    layer8_outputs(3547) <= not (a or b);
    layer8_outputs(3548) <= not a;
    layer8_outputs(3549) <= a and not b;
    layer8_outputs(3550) <= not a;
    layer8_outputs(3551) <= a;
    layer8_outputs(3552) <= a;
    layer8_outputs(3553) <= not b;
    layer8_outputs(3554) <= not a;
    layer8_outputs(3555) <= a;
    layer8_outputs(3556) <= a xor b;
    layer8_outputs(3557) <= not (a xor b);
    layer8_outputs(3558) <= b;
    layer8_outputs(3559) <= not a;
    layer8_outputs(3560) <= b;
    layer8_outputs(3561) <= b;
    layer8_outputs(3562) <= a xor b;
    layer8_outputs(3563) <= a or b;
    layer8_outputs(3564) <= a and not b;
    layer8_outputs(3565) <= a;
    layer8_outputs(3566) <= not b or a;
    layer8_outputs(3567) <= not b;
    layer8_outputs(3568) <= not b;
    layer8_outputs(3569) <= not (a and b);
    layer8_outputs(3570) <= not (a and b);
    layer8_outputs(3571) <= b and not a;
    layer8_outputs(3572) <= a;
    layer8_outputs(3573) <= b;
    layer8_outputs(3574) <= a and not b;
    layer8_outputs(3575) <= a and b;
    layer8_outputs(3576) <= a xor b;
    layer8_outputs(3577) <= b and not a;
    layer8_outputs(3578) <= not a or b;
    layer8_outputs(3579) <= a;
    layer8_outputs(3580) <= not a or b;
    layer8_outputs(3581) <= a;
    layer8_outputs(3582) <= not (a xor b);
    layer8_outputs(3583) <= not a;
    layer8_outputs(3584) <= not a or b;
    layer8_outputs(3585) <= a;
    layer8_outputs(3586) <= not b or a;
    layer8_outputs(3587) <= a and b;
    layer8_outputs(3588) <= a;
    layer8_outputs(3589) <= a;
    layer8_outputs(3590) <= a xor b;
    layer8_outputs(3591) <= b;
    layer8_outputs(3592) <= a and not b;
    layer8_outputs(3593) <= a;
    layer8_outputs(3594) <= not b;
    layer8_outputs(3595) <= a xor b;
    layer8_outputs(3596) <= b;
    layer8_outputs(3597) <= not (a xor b);
    layer8_outputs(3598) <= a xor b;
    layer8_outputs(3599) <= not (a xor b);
    layer8_outputs(3600) <= b and not a;
    layer8_outputs(3601) <= a;
    layer8_outputs(3602) <= not (a xor b);
    layer8_outputs(3603) <= a xor b;
    layer8_outputs(3604) <= b and not a;
    layer8_outputs(3605) <= not a;
    layer8_outputs(3606) <= not a;
    layer8_outputs(3607) <= a or b;
    layer8_outputs(3608) <= a or b;
    layer8_outputs(3609) <= a or b;
    layer8_outputs(3610) <= b and not a;
    layer8_outputs(3611) <= not a or b;
    layer8_outputs(3612) <= not (a xor b);
    layer8_outputs(3613) <= not (a or b);
    layer8_outputs(3614) <= not b;
    layer8_outputs(3615) <= not (a xor b);
    layer8_outputs(3616) <= not b or a;
    layer8_outputs(3617) <= a and not b;
    layer8_outputs(3618) <= a xor b;
    layer8_outputs(3619) <= not (a xor b);
    layer8_outputs(3620) <= not (a xor b);
    layer8_outputs(3621) <= not a;
    layer8_outputs(3622) <= not b;
    layer8_outputs(3623) <= not b;
    layer8_outputs(3624) <= not (a xor b);
    layer8_outputs(3625) <= not (a xor b);
    layer8_outputs(3626) <= b;
    layer8_outputs(3627) <= a;
    layer8_outputs(3628) <= a and b;
    layer8_outputs(3629) <= not (a and b);
    layer8_outputs(3630) <= not a;
    layer8_outputs(3631) <= not b;
    layer8_outputs(3632) <= a;
    layer8_outputs(3633) <= not a;
    layer8_outputs(3634) <= a;
    layer8_outputs(3635) <= a xor b;
    layer8_outputs(3636) <= not b;
    layer8_outputs(3637) <= not (a or b);
    layer8_outputs(3638) <= a;
    layer8_outputs(3639) <= not b;
    layer8_outputs(3640) <= b;
    layer8_outputs(3641) <= a and not b;
    layer8_outputs(3642) <= a and b;
    layer8_outputs(3643) <= a or b;
    layer8_outputs(3644) <= not b;
    layer8_outputs(3645) <= not (a xor b);
    layer8_outputs(3646) <= not a or b;
    layer8_outputs(3647) <= not b;
    layer8_outputs(3648) <= a and b;
    layer8_outputs(3649) <= not (a xor b);
    layer8_outputs(3650) <= a xor b;
    layer8_outputs(3651) <= not (a xor b);
    layer8_outputs(3652) <= not a;
    layer8_outputs(3653) <= a and b;
    layer8_outputs(3654) <= not (a and b);
    layer8_outputs(3655) <= a;
    layer8_outputs(3656) <= a;
    layer8_outputs(3657) <= a xor b;
    layer8_outputs(3658) <= 1'b0;
    layer8_outputs(3659) <= a xor b;
    layer8_outputs(3660) <= not a;
    layer8_outputs(3661) <= a xor b;
    layer8_outputs(3662) <= not b or a;
    layer8_outputs(3663) <= not b or a;
    layer8_outputs(3664) <= b;
    layer8_outputs(3665) <= b;
    layer8_outputs(3666) <= b;
    layer8_outputs(3667) <= 1'b0;
    layer8_outputs(3668) <= a and not b;
    layer8_outputs(3669) <= not b;
    layer8_outputs(3670) <= a or b;
    layer8_outputs(3671) <= not a or b;
    layer8_outputs(3672) <= b;
    layer8_outputs(3673) <= not (a or b);
    layer8_outputs(3674) <= not (a xor b);
    layer8_outputs(3675) <= a xor b;
    layer8_outputs(3676) <= a;
    layer8_outputs(3677) <= a;
    layer8_outputs(3678) <= a and b;
    layer8_outputs(3679) <= not (a and b);
    layer8_outputs(3680) <= not b or a;
    layer8_outputs(3681) <= not (a and b);
    layer8_outputs(3682) <= a and not b;
    layer8_outputs(3683) <= not (a xor b);
    layer8_outputs(3684) <= not (a xor b);
    layer8_outputs(3685) <= not (a or b);
    layer8_outputs(3686) <= not a or b;
    layer8_outputs(3687) <= not b;
    layer8_outputs(3688) <= a xor b;
    layer8_outputs(3689) <= a;
    layer8_outputs(3690) <= a xor b;
    layer8_outputs(3691) <= not b;
    layer8_outputs(3692) <= b;
    layer8_outputs(3693) <= a;
    layer8_outputs(3694) <= a;
    layer8_outputs(3695) <= a xor b;
    layer8_outputs(3696) <= not (a xor b);
    layer8_outputs(3697) <= not a or b;
    layer8_outputs(3698) <= not (a and b);
    layer8_outputs(3699) <= not b;
    layer8_outputs(3700) <= not (a xor b);
    layer8_outputs(3701) <= not b;
    layer8_outputs(3702) <= not a or b;
    layer8_outputs(3703) <= a;
    layer8_outputs(3704) <= a;
    layer8_outputs(3705) <= a;
    layer8_outputs(3706) <= a xor b;
    layer8_outputs(3707) <= b and not a;
    layer8_outputs(3708) <= a;
    layer8_outputs(3709) <= not b;
    layer8_outputs(3710) <= not a;
    layer8_outputs(3711) <= not b;
    layer8_outputs(3712) <= not (a and b);
    layer8_outputs(3713) <= not (a or b);
    layer8_outputs(3714) <= 1'b1;
    layer8_outputs(3715) <= a or b;
    layer8_outputs(3716) <= not (a xor b);
    layer8_outputs(3717) <= b;
    layer8_outputs(3718) <= b;
    layer8_outputs(3719) <= not b;
    layer8_outputs(3720) <= not b or a;
    layer8_outputs(3721) <= b;
    layer8_outputs(3722) <= a xor b;
    layer8_outputs(3723) <= not (a xor b);
    layer8_outputs(3724) <= a xor b;
    layer8_outputs(3725) <= b;
    layer8_outputs(3726) <= not a or b;
    layer8_outputs(3727) <= b;
    layer8_outputs(3728) <= not a;
    layer8_outputs(3729) <= not b;
    layer8_outputs(3730) <= a xor b;
    layer8_outputs(3731) <= b;
    layer8_outputs(3732) <= not b or a;
    layer8_outputs(3733) <= not b or a;
    layer8_outputs(3734) <= b and not a;
    layer8_outputs(3735) <= b;
    layer8_outputs(3736) <= b;
    layer8_outputs(3737) <= a xor b;
    layer8_outputs(3738) <= a;
    layer8_outputs(3739) <= a;
    layer8_outputs(3740) <= not (a xor b);
    layer8_outputs(3741) <= not (a xor b);
    layer8_outputs(3742) <= a;
    layer8_outputs(3743) <= a and b;
    layer8_outputs(3744) <= not b;
    layer8_outputs(3745) <= a and b;
    layer8_outputs(3746) <= not (a xor b);
    layer8_outputs(3747) <= not b;
    layer8_outputs(3748) <= a;
    layer8_outputs(3749) <= not (a xor b);
    layer8_outputs(3750) <= not b;
    layer8_outputs(3751) <= not a or b;
    layer8_outputs(3752) <= 1'b1;
    layer8_outputs(3753) <= b and not a;
    layer8_outputs(3754) <= a or b;
    layer8_outputs(3755) <= not (a and b);
    layer8_outputs(3756) <= a;
    layer8_outputs(3757) <= not (a xor b);
    layer8_outputs(3758) <= b;
    layer8_outputs(3759) <= not b;
    layer8_outputs(3760) <= b;
    layer8_outputs(3761) <= not a or b;
    layer8_outputs(3762) <= a;
    layer8_outputs(3763) <= not a;
    layer8_outputs(3764) <= a and b;
    layer8_outputs(3765) <= not (a xor b);
    layer8_outputs(3766) <= a;
    layer8_outputs(3767) <= not a;
    layer8_outputs(3768) <= not b;
    layer8_outputs(3769) <= not (a xor b);
    layer8_outputs(3770) <= not b or a;
    layer8_outputs(3771) <= b and not a;
    layer8_outputs(3772) <= b;
    layer8_outputs(3773) <= not a;
    layer8_outputs(3774) <= not (a and b);
    layer8_outputs(3775) <= not b;
    layer8_outputs(3776) <= not a;
    layer8_outputs(3777) <= a;
    layer8_outputs(3778) <= b;
    layer8_outputs(3779) <= not b or a;
    layer8_outputs(3780) <= b;
    layer8_outputs(3781) <= b;
    layer8_outputs(3782) <= 1'b0;
    layer8_outputs(3783) <= not b;
    layer8_outputs(3784) <= a and not b;
    layer8_outputs(3785) <= not a;
    layer8_outputs(3786) <= not a;
    layer8_outputs(3787) <= not (a or b);
    layer8_outputs(3788) <= a xor b;
    layer8_outputs(3789) <= a xor b;
    layer8_outputs(3790) <= not b or a;
    layer8_outputs(3791) <= a and b;
    layer8_outputs(3792) <= a;
    layer8_outputs(3793) <= not a;
    layer8_outputs(3794) <= not (a and b);
    layer8_outputs(3795) <= not (a xor b);
    layer8_outputs(3796) <= not b;
    layer8_outputs(3797) <= b;
    layer8_outputs(3798) <= a xor b;
    layer8_outputs(3799) <= not b;
    layer8_outputs(3800) <= not b;
    layer8_outputs(3801) <= b;
    layer8_outputs(3802) <= a xor b;
    layer8_outputs(3803) <= b;
    layer8_outputs(3804) <= b and not a;
    layer8_outputs(3805) <= a xor b;
    layer8_outputs(3806) <= a and not b;
    layer8_outputs(3807) <= 1'b1;
    layer8_outputs(3808) <= not b;
    layer8_outputs(3809) <= not (a or b);
    layer8_outputs(3810) <= b and not a;
    layer8_outputs(3811) <= a and not b;
    layer8_outputs(3812) <= a xor b;
    layer8_outputs(3813) <= a xor b;
    layer8_outputs(3814) <= not a;
    layer8_outputs(3815) <= not b;
    layer8_outputs(3816) <= a xor b;
    layer8_outputs(3817) <= not b;
    layer8_outputs(3818) <= b;
    layer8_outputs(3819) <= not b;
    layer8_outputs(3820) <= not b;
    layer8_outputs(3821) <= a;
    layer8_outputs(3822) <= not a;
    layer8_outputs(3823) <= not (a xor b);
    layer8_outputs(3824) <= a or b;
    layer8_outputs(3825) <= not (a xor b);
    layer8_outputs(3826) <= not a;
    layer8_outputs(3827) <= a xor b;
    layer8_outputs(3828) <= not b;
    layer8_outputs(3829) <= a;
    layer8_outputs(3830) <= a xor b;
    layer8_outputs(3831) <= a xor b;
    layer8_outputs(3832) <= not (a xor b);
    layer8_outputs(3833) <= not (a or b);
    layer8_outputs(3834) <= not (a and b);
    layer8_outputs(3835) <= b and not a;
    layer8_outputs(3836) <= not (a xor b);
    layer8_outputs(3837) <= not (a or b);
    layer8_outputs(3838) <= b;
    layer8_outputs(3839) <= not b;
    layer8_outputs(3840) <= not b;
    layer8_outputs(3841) <= a xor b;
    layer8_outputs(3842) <= not (a xor b);
    layer8_outputs(3843) <= not b;
    layer8_outputs(3844) <= not b;
    layer8_outputs(3845) <= not a;
    layer8_outputs(3846) <= not a;
    layer8_outputs(3847) <= not a;
    layer8_outputs(3848) <= not a;
    layer8_outputs(3849) <= a;
    layer8_outputs(3850) <= not a;
    layer8_outputs(3851) <= not a;
    layer8_outputs(3852) <= not (a or b);
    layer8_outputs(3853) <= not a;
    layer8_outputs(3854) <= a;
    layer8_outputs(3855) <= not (a xor b);
    layer8_outputs(3856) <= a and b;
    layer8_outputs(3857) <= a xor b;
    layer8_outputs(3858) <= a xor b;
    layer8_outputs(3859) <= a and b;
    layer8_outputs(3860) <= not b;
    layer8_outputs(3861) <= a and b;
    layer8_outputs(3862) <= b;
    layer8_outputs(3863) <= not b;
    layer8_outputs(3864) <= not b;
    layer8_outputs(3865) <= a;
    layer8_outputs(3866) <= b;
    layer8_outputs(3867) <= a xor b;
    layer8_outputs(3868) <= b;
    layer8_outputs(3869) <= not (a xor b);
    layer8_outputs(3870) <= not b or a;
    layer8_outputs(3871) <= a;
    layer8_outputs(3872) <= not b;
    layer8_outputs(3873) <= not b;
    layer8_outputs(3874) <= not b;
    layer8_outputs(3875) <= not a;
    layer8_outputs(3876) <= a xor b;
    layer8_outputs(3877) <= a and b;
    layer8_outputs(3878) <= b and not a;
    layer8_outputs(3879) <= b;
    layer8_outputs(3880) <= b and not a;
    layer8_outputs(3881) <= a xor b;
    layer8_outputs(3882) <= not (a xor b);
    layer8_outputs(3883) <= b;
    layer8_outputs(3884) <= not (a xor b);
    layer8_outputs(3885) <= not (a xor b);
    layer8_outputs(3886) <= not b or a;
    layer8_outputs(3887) <= not (a and b);
    layer8_outputs(3888) <= not b or a;
    layer8_outputs(3889) <= not a or b;
    layer8_outputs(3890) <= a xor b;
    layer8_outputs(3891) <= not a;
    layer8_outputs(3892) <= not a or b;
    layer8_outputs(3893) <= not b;
    layer8_outputs(3894) <= not a;
    layer8_outputs(3895) <= not b;
    layer8_outputs(3896) <= b;
    layer8_outputs(3897) <= not b or a;
    layer8_outputs(3898) <= not (a or b);
    layer8_outputs(3899) <= not (a xor b);
    layer8_outputs(3900) <= a;
    layer8_outputs(3901) <= b;
    layer8_outputs(3902) <= a;
    layer8_outputs(3903) <= not (a xor b);
    layer8_outputs(3904) <= a;
    layer8_outputs(3905) <= not a or b;
    layer8_outputs(3906) <= not a;
    layer8_outputs(3907) <= not (a or b);
    layer8_outputs(3908) <= not b;
    layer8_outputs(3909) <= 1'b0;
    layer8_outputs(3910) <= not b;
    layer8_outputs(3911) <= a xor b;
    layer8_outputs(3912) <= not a;
    layer8_outputs(3913) <= a or b;
    layer8_outputs(3914) <= not (a and b);
    layer8_outputs(3915) <= a and b;
    layer8_outputs(3916) <= a xor b;
    layer8_outputs(3917) <= b;
    layer8_outputs(3918) <= a;
    layer8_outputs(3919) <= a and not b;
    layer8_outputs(3920) <= not b or a;
    layer8_outputs(3921) <= a xor b;
    layer8_outputs(3922) <= b and not a;
    layer8_outputs(3923) <= a and not b;
    layer8_outputs(3924) <= not a;
    layer8_outputs(3925) <= not (a and b);
    layer8_outputs(3926) <= not (a xor b);
    layer8_outputs(3927) <= a or b;
    layer8_outputs(3928) <= a or b;
    layer8_outputs(3929) <= not a;
    layer8_outputs(3930) <= a;
    layer8_outputs(3931) <= a;
    layer8_outputs(3932) <= not b;
    layer8_outputs(3933) <= not b;
    layer8_outputs(3934) <= not b;
    layer8_outputs(3935) <= a;
    layer8_outputs(3936) <= a;
    layer8_outputs(3937) <= not b;
    layer8_outputs(3938) <= not (a and b);
    layer8_outputs(3939) <= b and not a;
    layer8_outputs(3940) <= not b or a;
    layer8_outputs(3941) <= not a;
    layer8_outputs(3942) <= not (a xor b);
    layer8_outputs(3943) <= not (a and b);
    layer8_outputs(3944) <= b;
    layer8_outputs(3945) <= not (a xor b);
    layer8_outputs(3946) <= not (a xor b);
    layer8_outputs(3947) <= not (a or b);
    layer8_outputs(3948) <= not b or a;
    layer8_outputs(3949) <= not (a xor b);
    layer8_outputs(3950) <= not (a xor b);
    layer8_outputs(3951) <= a;
    layer8_outputs(3952) <= not (a xor b);
    layer8_outputs(3953) <= not b;
    layer8_outputs(3954) <= b;
    layer8_outputs(3955) <= not (a and b);
    layer8_outputs(3956) <= not b or a;
    layer8_outputs(3957) <= not a or b;
    layer8_outputs(3958) <= not b;
    layer8_outputs(3959) <= b;
    layer8_outputs(3960) <= not a;
    layer8_outputs(3961) <= b;
    layer8_outputs(3962) <= a xor b;
    layer8_outputs(3963) <= not (a xor b);
    layer8_outputs(3964) <= b and not a;
    layer8_outputs(3965) <= b;
    layer8_outputs(3966) <= not b;
    layer8_outputs(3967) <= not (a xor b);
    layer8_outputs(3968) <= not (a xor b);
    layer8_outputs(3969) <= a xor b;
    layer8_outputs(3970) <= a;
    layer8_outputs(3971) <= a or b;
    layer8_outputs(3972) <= a or b;
    layer8_outputs(3973) <= a or b;
    layer8_outputs(3974) <= a xor b;
    layer8_outputs(3975) <= a and not b;
    layer8_outputs(3976) <= b and not a;
    layer8_outputs(3977) <= b;
    layer8_outputs(3978) <= not (a xor b);
    layer8_outputs(3979) <= not a;
    layer8_outputs(3980) <= not (a and b);
    layer8_outputs(3981) <= a and b;
    layer8_outputs(3982) <= a or b;
    layer8_outputs(3983) <= not a;
    layer8_outputs(3984) <= a xor b;
    layer8_outputs(3985) <= a or b;
    layer8_outputs(3986) <= not (a and b);
    layer8_outputs(3987) <= not (a xor b);
    layer8_outputs(3988) <= not b;
    layer8_outputs(3989) <= b;
    layer8_outputs(3990) <= b;
    layer8_outputs(3991) <= a;
    layer8_outputs(3992) <= b;
    layer8_outputs(3993) <= a xor b;
    layer8_outputs(3994) <= not (a or b);
    layer8_outputs(3995) <= a;
    layer8_outputs(3996) <= not (a xor b);
    layer8_outputs(3997) <= b and not a;
    layer8_outputs(3998) <= b;
    layer8_outputs(3999) <= not b;
    layer8_outputs(4000) <= b;
    layer8_outputs(4001) <= a xor b;
    layer8_outputs(4002) <= a and not b;
    layer8_outputs(4003) <= a and b;
    layer8_outputs(4004) <= not a or b;
    layer8_outputs(4005) <= a xor b;
    layer8_outputs(4006) <= 1'b0;
    layer8_outputs(4007) <= not a;
    layer8_outputs(4008) <= not (a xor b);
    layer8_outputs(4009) <= not b or a;
    layer8_outputs(4010) <= a;
    layer8_outputs(4011) <= a and b;
    layer8_outputs(4012) <= not (a xor b);
    layer8_outputs(4013) <= not a or b;
    layer8_outputs(4014) <= not (a xor b);
    layer8_outputs(4015) <= not b;
    layer8_outputs(4016) <= not (a xor b);
    layer8_outputs(4017) <= not (a xor b);
    layer8_outputs(4018) <= a xor b;
    layer8_outputs(4019) <= a xor b;
    layer8_outputs(4020) <= a and not b;
    layer8_outputs(4021) <= not (a xor b);
    layer8_outputs(4022) <= b;
    layer8_outputs(4023) <= a;
    layer8_outputs(4024) <= not a or b;
    layer8_outputs(4025) <= b;
    layer8_outputs(4026) <= not (a xor b);
    layer8_outputs(4027) <= not (a xor b);
    layer8_outputs(4028) <= b;
    layer8_outputs(4029) <= a;
    layer8_outputs(4030) <= not a;
    layer8_outputs(4031) <= not (a and b);
    layer8_outputs(4032) <= a;
    layer8_outputs(4033) <= not (a and b);
    layer8_outputs(4034) <= not a;
    layer8_outputs(4035) <= not a;
    layer8_outputs(4036) <= not (a or b);
    layer8_outputs(4037) <= not b or a;
    layer8_outputs(4038) <= a and not b;
    layer8_outputs(4039) <= a or b;
    layer8_outputs(4040) <= b;
    layer8_outputs(4041) <= a xor b;
    layer8_outputs(4042) <= a xor b;
    layer8_outputs(4043) <= a;
    layer8_outputs(4044) <= a and b;
    layer8_outputs(4045) <= not a;
    layer8_outputs(4046) <= a or b;
    layer8_outputs(4047) <= not a;
    layer8_outputs(4048) <= not a;
    layer8_outputs(4049) <= a xor b;
    layer8_outputs(4050) <= not (a xor b);
    layer8_outputs(4051) <= not b;
    layer8_outputs(4052) <= a xor b;
    layer8_outputs(4053) <= not a;
    layer8_outputs(4054) <= not b;
    layer8_outputs(4055) <= not (a xor b);
    layer8_outputs(4056) <= a and not b;
    layer8_outputs(4057) <= a;
    layer8_outputs(4058) <= not b;
    layer8_outputs(4059) <= not b;
    layer8_outputs(4060) <= not (a xor b);
    layer8_outputs(4061) <= not a;
    layer8_outputs(4062) <= a or b;
    layer8_outputs(4063) <= a or b;
    layer8_outputs(4064) <= not (a xor b);
    layer8_outputs(4065) <= a and b;
    layer8_outputs(4066) <= not a or b;
    layer8_outputs(4067) <= a;
    layer8_outputs(4068) <= b;
    layer8_outputs(4069) <= a xor b;
    layer8_outputs(4070) <= a;
    layer8_outputs(4071) <= b;
    layer8_outputs(4072) <= not a;
    layer8_outputs(4073) <= a;
    layer8_outputs(4074) <= not a or b;
    layer8_outputs(4075) <= not b;
    layer8_outputs(4076) <= a and not b;
    layer8_outputs(4077) <= a and b;
    layer8_outputs(4078) <= a xor b;
    layer8_outputs(4079) <= a and b;
    layer8_outputs(4080) <= not (a xor b);
    layer8_outputs(4081) <= not (a xor b);
    layer8_outputs(4082) <= not (a xor b);
    layer8_outputs(4083) <= b;
    layer8_outputs(4084) <= not b;
    layer8_outputs(4085) <= not (a and b);
    layer8_outputs(4086) <= not (a xor b);
    layer8_outputs(4087) <= not b;
    layer8_outputs(4088) <= a;
    layer8_outputs(4089) <= a or b;
    layer8_outputs(4090) <= a xor b;
    layer8_outputs(4091) <= a;
    layer8_outputs(4092) <= not (a and b);
    layer8_outputs(4093) <= a;
    layer8_outputs(4094) <= b;
    layer8_outputs(4095) <= not (a or b);
    layer8_outputs(4096) <= not b;
    layer8_outputs(4097) <= b;
    layer8_outputs(4098) <= a and b;
    layer8_outputs(4099) <= a or b;
    layer8_outputs(4100) <= 1'b1;
    layer8_outputs(4101) <= not a or b;
    layer8_outputs(4102) <= a;
    layer8_outputs(4103) <= not b or a;
    layer8_outputs(4104) <= not (a xor b);
    layer8_outputs(4105) <= a;
    layer8_outputs(4106) <= not a;
    layer8_outputs(4107) <= a and not b;
    layer8_outputs(4108) <= not b;
    layer8_outputs(4109) <= not b;
    layer8_outputs(4110) <= not a;
    layer8_outputs(4111) <= not a;
    layer8_outputs(4112) <= not (a xor b);
    layer8_outputs(4113) <= not a;
    layer8_outputs(4114) <= not a;
    layer8_outputs(4115) <= not a;
    layer8_outputs(4116) <= not (a and b);
    layer8_outputs(4117) <= not b or a;
    layer8_outputs(4118) <= a xor b;
    layer8_outputs(4119) <= not a;
    layer8_outputs(4120) <= a;
    layer8_outputs(4121) <= a xor b;
    layer8_outputs(4122) <= a xor b;
    layer8_outputs(4123) <= a;
    layer8_outputs(4124) <= a and b;
    layer8_outputs(4125) <= b;
    layer8_outputs(4126) <= a and not b;
    layer8_outputs(4127) <= a xor b;
    layer8_outputs(4128) <= not b;
    layer8_outputs(4129) <= not b or a;
    layer8_outputs(4130) <= a xor b;
    layer8_outputs(4131) <= a or b;
    layer8_outputs(4132) <= not b;
    layer8_outputs(4133) <= not b;
    layer8_outputs(4134) <= not a or b;
    layer8_outputs(4135) <= a xor b;
    layer8_outputs(4136) <= a or b;
    layer8_outputs(4137) <= not b or a;
    layer8_outputs(4138) <= b and not a;
    layer8_outputs(4139) <= not b;
    layer8_outputs(4140) <= not (a and b);
    layer8_outputs(4141) <= not a;
    layer8_outputs(4142) <= b;
    layer8_outputs(4143) <= a or b;
    layer8_outputs(4144) <= not (a xor b);
    layer8_outputs(4145) <= b and not a;
    layer8_outputs(4146) <= not b;
    layer8_outputs(4147) <= b;
    layer8_outputs(4148) <= a or b;
    layer8_outputs(4149) <= not (a xor b);
    layer8_outputs(4150) <= not (a xor b);
    layer8_outputs(4151) <= a;
    layer8_outputs(4152) <= not a or b;
    layer8_outputs(4153) <= b;
    layer8_outputs(4154) <= not (a xor b);
    layer8_outputs(4155) <= not (a xor b);
    layer8_outputs(4156) <= not (a xor b);
    layer8_outputs(4157) <= a;
    layer8_outputs(4158) <= b;
    layer8_outputs(4159) <= not a;
    layer8_outputs(4160) <= not (a xor b);
    layer8_outputs(4161) <= b;
    layer8_outputs(4162) <= b and not a;
    layer8_outputs(4163) <= not b or a;
    layer8_outputs(4164) <= a xor b;
    layer8_outputs(4165) <= not (a xor b);
    layer8_outputs(4166) <= a xor b;
    layer8_outputs(4167) <= not (a xor b);
    layer8_outputs(4168) <= a and b;
    layer8_outputs(4169) <= not b;
    layer8_outputs(4170) <= a or b;
    layer8_outputs(4171) <= a or b;
    layer8_outputs(4172) <= a;
    layer8_outputs(4173) <= a and b;
    layer8_outputs(4174) <= not (a or b);
    layer8_outputs(4175) <= a;
    layer8_outputs(4176) <= not b;
    layer8_outputs(4177) <= a;
    layer8_outputs(4178) <= b;
    layer8_outputs(4179) <= not (a and b);
    layer8_outputs(4180) <= a and b;
    layer8_outputs(4181) <= a;
    layer8_outputs(4182) <= a;
    layer8_outputs(4183) <= not (a or b);
    layer8_outputs(4184) <= a and not b;
    layer8_outputs(4185) <= a xor b;
    layer8_outputs(4186) <= not a or b;
    layer8_outputs(4187) <= not b;
    layer8_outputs(4188) <= a xor b;
    layer8_outputs(4189) <= not a;
    layer8_outputs(4190) <= a and b;
    layer8_outputs(4191) <= not (a and b);
    layer8_outputs(4192) <= a and not b;
    layer8_outputs(4193) <= b and not a;
    layer8_outputs(4194) <= a;
    layer8_outputs(4195) <= not a;
    layer8_outputs(4196) <= b and not a;
    layer8_outputs(4197) <= not a;
    layer8_outputs(4198) <= not a;
    layer8_outputs(4199) <= not a;
    layer8_outputs(4200) <= b;
    layer8_outputs(4201) <= not b or a;
    layer8_outputs(4202) <= b and not a;
    layer8_outputs(4203) <= not (a or b);
    layer8_outputs(4204) <= not b or a;
    layer8_outputs(4205) <= not b;
    layer8_outputs(4206) <= 1'b1;
    layer8_outputs(4207) <= b and not a;
    layer8_outputs(4208) <= not (a and b);
    layer8_outputs(4209) <= not b;
    layer8_outputs(4210) <= not (a xor b);
    layer8_outputs(4211) <= not b;
    layer8_outputs(4212) <= not a;
    layer8_outputs(4213) <= not a;
    layer8_outputs(4214) <= not (a xor b);
    layer8_outputs(4215) <= a;
    layer8_outputs(4216) <= b;
    layer8_outputs(4217) <= a or b;
    layer8_outputs(4218) <= b and not a;
    layer8_outputs(4219) <= a;
    layer8_outputs(4220) <= a;
    layer8_outputs(4221) <= a or b;
    layer8_outputs(4222) <= a xor b;
    layer8_outputs(4223) <= not (a xor b);
    layer8_outputs(4224) <= not b;
    layer8_outputs(4225) <= a and not b;
    layer8_outputs(4226) <= not a;
    layer8_outputs(4227) <= not a or b;
    layer8_outputs(4228) <= not (a or b);
    layer8_outputs(4229) <= a and b;
    layer8_outputs(4230) <= not a or b;
    layer8_outputs(4231) <= b and not a;
    layer8_outputs(4232) <= not (a and b);
    layer8_outputs(4233) <= a and not b;
    layer8_outputs(4234) <= not (a or b);
    layer8_outputs(4235) <= not b or a;
    layer8_outputs(4236) <= not (a or b);
    layer8_outputs(4237) <= 1'b0;
    layer8_outputs(4238) <= not a;
    layer8_outputs(4239) <= a xor b;
    layer8_outputs(4240) <= a xor b;
    layer8_outputs(4241) <= a;
    layer8_outputs(4242) <= a xor b;
    layer8_outputs(4243) <= a;
    layer8_outputs(4244) <= not (a or b);
    layer8_outputs(4245) <= not (a xor b);
    layer8_outputs(4246) <= a;
    layer8_outputs(4247) <= not a;
    layer8_outputs(4248) <= not a;
    layer8_outputs(4249) <= not (a or b);
    layer8_outputs(4250) <= not b;
    layer8_outputs(4251) <= not (a or b);
    layer8_outputs(4252) <= b;
    layer8_outputs(4253) <= not (a or b);
    layer8_outputs(4254) <= a;
    layer8_outputs(4255) <= a and b;
    layer8_outputs(4256) <= not (a xor b);
    layer8_outputs(4257) <= not (a xor b);
    layer8_outputs(4258) <= not b;
    layer8_outputs(4259) <= 1'b0;
    layer8_outputs(4260) <= a and not b;
    layer8_outputs(4261) <= not (a xor b);
    layer8_outputs(4262) <= not b;
    layer8_outputs(4263) <= a xor b;
    layer8_outputs(4264) <= not b;
    layer8_outputs(4265) <= a or b;
    layer8_outputs(4266) <= b;
    layer8_outputs(4267) <= b;
    layer8_outputs(4268) <= not a;
    layer8_outputs(4269) <= not a;
    layer8_outputs(4270) <= not (a xor b);
    layer8_outputs(4271) <= a;
    layer8_outputs(4272) <= not b or a;
    layer8_outputs(4273) <= a;
    layer8_outputs(4274) <= b;
    layer8_outputs(4275) <= b and not a;
    layer8_outputs(4276) <= a;
    layer8_outputs(4277) <= a;
    layer8_outputs(4278) <= b;
    layer8_outputs(4279) <= a xor b;
    layer8_outputs(4280) <= a xor b;
    layer8_outputs(4281) <= not a or b;
    layer8_outputs(4282) <= b;
    layer8_outputs(4283) <= not b;
    layer8_outputs(4284) <= a and b;
    layer8_outputs(4285) <= not (a or b);
    layer8_outputs(4286) <= not b;
    layer8_outputs(4287) <= b;
    layer8_outputs(4288) <= a xor b;
    layer8_outputs(4289) <= not a;
    layer8_outputs(4290) <= not (a xor b);
    layer8_outputs(4291) <= not (a xor b);
    layer8_outputs(4292) <= 1'b0;
    layer8_outputs(4293) <= a;
    layer8_outputs(4294) <= not a;
    layer8_outputs(4295) <= a;
    layer8_outputs(4296) <= not (a or b);
    layer8_outputs(4297) <= a xor b;
    layer8_outputs(4298) <= a and not b;
    layer8_outputs(4299) <= b;
    layer8_outputs(4300) <= a xor b;
    layer8_outputs(4301) <= not a;
    layer8_outputs(4302) <= not b;
    layer8_outputs(4303) <= a or b;
    layer8_outputs(4304) <= not a;
    layer8_outputs(4305) <= a xor b;
    layer8_outputs(4306) <= a;
    layer8_outputs(4307) <= not b;
    layer8_outputs(4308) <= b and not a;
    layer8_outputs(4309) <= not (a and b);
    layer8_outputs(4310) <= not (a or b);
    layer8_outputs(4311) <= not (a and b);
    layer8_outputs(4312) <= b;
    layer8_outputs(4313) <= not b or a;
    layer8_outputs(4314) <= not b or a;
    layer8_outputs(4315) <= not b;
    layer8_outputs(4316) <= a;
    layer8_outputs(4317) <= not (a or b);
    layer8_outputs(4318) <= not (a and b);
    layer8_outputs(4319) <= not a or b;
    layer8_outputs(4320) <= not (a xor b);
    layer8_outputs(4321) <= a xor b;
    layer8_outputs(4322) <= a;
    layer8_outputs(4323) <= not b;
    layer8_outputs(4324) <= not (a or b);
    layer8_outputs(4325) <= not a;
    layer8_outputs(4326) <= a;
    layer8_outputs(4327) <= b;
    layer8_outputs(4328) <= not (a xor b);
    layer8_outputs(4329) <= not b;
    layer8_outputs(4330) <= a xor b;
    layer8_outputs(4331) <= 1'b1;
    layer8_outputs(4332) <= not (a and b);
    layer8_outputs(4333) <= not (a xor b);
    layer8_outputs(4334) <= not a;
    layer8_outputs(4335) <= not b;
    layer8_outputs(4336) <= a;
    layer8_outputs(4337) <= b;
    layer8_outputs(4338) <= a and b;
    layer8_outputs(4339) <= not a;
    layer8_outputs(4340) <= a and b;
    layer8_outputs(4341) <= not a;
    layer8_outputs(4342) <= not b or a;
    layer8_outputs(4343) <= not a;
    layer8_outputs(4344) <= not b or a;
    layer8_outputs(4345) <= not b;
    layer8_outputs(4346) <= not b or a;
    layer8_outputs(4347) <= a xor b;
    layer8_outputs(4348) <= 1'b0;
    layer8_outputs(4349) <= 1'b0;
    layer8_outputs(4350) <= a;
    layer8_outputs(4351) <= not (a and b);
    layer8_outputs(4352) <= b;
    layer8_outputs(4353) <= a or b;
    layer8_outputs(4354) <= a or b;
    layer8_outputs(4355) <= a;
    layer8_outputs(4356) <= not b;
    layer8_outputs(4357) <= b;
    layer8_outputs(4358) <= a xor b;
    layer8_outputs(4359) <= not a;
    layer8_outputs(4360) <= not (a xor b);
    layer8_outputs(4361) <= 1'b0;
    layer8_outputs(4362) <= not (a xor b);
    layer8_outputs(4363) <= not a;
    layer8_outputs(4364) <= not (a xor b);
    layer8_outputs(4365) <= not (a or b);
    layer8_outputs(4366) <= not a or b;
    layer8_outputs(4367) <= not (a xor b);
    layer8_outputs(4368) <= not b;
    layer8_outputs(4369) <= a or b;
    layer8_outputs(4370) <= a;
    layer8_outputs(4371) <= a or b;
    layer8_outputs(4372) <= a;
    layer8_outputs(4373) <= b and not a;
    layer8_outputs(4374) <= b;
    layer8_outputs(4375) <= not (a xor b);
    layer8_outputs(4376) <= b;
    layer8_outputs(4377) <= not (a and b);
    layer8_outputs(4378) <= not b;
    layer8_outputs(4379) <= not a;
    layer8_outputs(4380) <= b;
    layer8_outputs(4381) <= a;
    layer8_outputs(4382) <= a xor b;
    layer8_outputs(4383) <= not b or a;
    layer8_outputs(4384) <= not (a xor b);
    layer8_outputs(4385) <= not (a xor b);
    layer8_outputs(4386) <= not a;
    layer8_outputs(4387) <= not b or a;
    layer8_outputs(4388) <= not b;
    layer8_outputs(4389) <= b;
    layer8_outputs(4390) <= not a or b;
    layer8_outputs(4391) <= b;
    layer8_outputs(4392) <= not b or a;
    layer8_outputs(4393) <= not (a xor b);
    layer8_outputs(4394) <= a or b;
    layer8_outputs(4395) <= a xor b;
    layer8_outputs(4396) <= not a or b;
    layer8_outputs(4397) <= not a;
    layer8_outputs(4398) <= a xor b;
    layer8_outputs(4399) <= not (a and b);
    layer8_outputs(4400) <= a;
    layer8_outputs(4401) <= a;
    layer8_outputs(4402) <= not (a or b);
    layer8_outputs(4403) <= not a or b;
    layer8_outputs(4404) <= a;
    layer8_outputs(4405) <= a;
    layer8_outputs(4406) <= a;
    layer8_outputs(4407) <= b;
    layer8_outputs(4408) <= a and b;
    layer8_outputs(4409) <= not (a xor b);
    layer8_outputs(4410) <= b;
    layer8_outputs(4411) <= b and not a;
    layer8_outputs(4412) <= not b;
    layer8_outputs(4413) <= not a or b;
    layer8_outputs(4414) <= not (a and b);
    layer8_outputs(4415) <= not (a xor b);
    layer8_outputs(4416) <= not b;
    layer8_outputs(4417) <= not b or a;
    layer8_outputs(4418) <= not (a xor b);
    layer8_outputs(4419) <= not b;
    layer8_outputs(4420) <= not a or b;
    layer8_outputs(4421) <= not b;
    layer8_outputs(4422) <= a;
    layer8_outputs(4423) <= not b or a;
    layer8_outputs(4424) <= not b;
    layer8_outputs(4425) <= a or b;
    layer8_outputs(4426) <= not b;
    layer8_outputs(4427) <= b;
    layer8_outputs(4428) <= not (a and b);
    layer8_outputs(4429) <= a xor b;
    layer8_outputs(4430) <= a xor b;
    layer8_outputs(4431) <= 1'b1;
    layer8_outputs(4432) <= not (a and b);
    layer8_outputs(4433) <= not (a and b);
    layer8_outputs(4434) <= a xor b;
    layer8_outputs(4435) <= b;
    layer8_outputs(4436) <= not b;
    layer8_outputs(4437) <= a or b;
    layer8_outputs(4438) <= not b;
    layer8_outputs(4439) <= not b or a;
    layer8_outputs(4440) <= a and b;
    layer8_outputs(4441) <= not (a xor b);
    layer8_outputs(4442) <= not (a or b);
    layer8_outputs(4443) <= b;
    layer8_outputs(4444) <= not (a and b);
    layer8_outputs(4445) <= b;
    layer8_outputs(4446) <= not (a and b);
    layer8_outputs(4447) <= 1'b0;
    layer8_outputs(4448) <= b;
    layer8_outputs(4449) <= a xor b;
    layer8_outputs(4450) <= a xor b;
    layer8_outputs(4451) <= a xor b;
    layer8_outputs(4452) <= a or b;
    layer8_outputs(4453) <= a xor b;
    layer8_outputs(4454) <= a and not b;
    layer8_outputs(4455) <= a;
    layer8_outputs(4456) <= a and b;
    layer8_outputs(4457) <= a and not b;
    layer8_outputs(4458) <= a;
    layer8_outputs(4459) <= not b;
    layer8_outputs(4460) <= not (a xor b);
    layer8_outputs(4461) <= not (a xor b);
    layer8_outputs(4462) <= a and b;
    layer8_outputs(4463) <= not (a or b);
    layer8_outputs(4464) <= not (a xor b);
    layer8_outputs(4465) <= a;
    layer8_outputs(4466) <= a and not b;
    layer8_outputs(4467) <= not a or b;
    layer8_outputs(4468) <= a xor b;
    layer8_outputs(4469) <= not b;
    layer8_outputs(4470) <= a or b;
    layer8_outputs(4471) <= not b;
    layer8_outputs(4472) <= not b;
    layer8_outputs(4473) <= b;
    layer8_outputs(4474) <= b;
    layer8_outputs(4475) <= b;
    layer8_outputs(4476) <= not b or a;
    layer8_outputs(4477) <= b;
    layer8_outputs(4478) <= a;
    layer8_outputs(4479) <= not a;
    layer8_outputs(4480) <= not b or a;
    layer8_outputs(4481) <= 1'b0;
    layer8_outputs(4482) <= not (a and b);
    layer8_outputs(4483) <= not a or b;
    layer8_outputs(4484) <= b;
    layer8_outputs(4485) <= not (a xor b);
    layer8_outputs(4486) <= not (a xor b);
    layer8_outputs(4487) <= not a;
    layer8_outputs(4488) <= not a;
    layer8_outputs(4489) <= not (a xor b);
    layer8_outputs(4490) <= a xor b;
    layer8_outputs(4491) <= not (a or b);
    layer8_outputs(4492) <= b;
    layer8_outputs(4493) <= a;
    layer8_outputs(4494) <= a;
    layer8_outputs(4495) <= a xor b;
    layer8_outputs(4496) <= not b;
    layer8_outputs(4497) <= a xor b;
    layer8_outputs(4498) <= a;
    layer8_outputs(4499) <= a;
    layer8_outputs(4500) <= not a or b;
    layer8_outputs(4501) <= a xor b;
    layer8_outputs(4502) <= not a;
    layer8_outputs(4503) <= not b;
    layer8_outputs(4504) <= not a;
    layer8_outputs(4505) <= a xor b;
    layer8_outputs(4506) <= not (a or b);
    layer8_outputs(4507) <= a and b;
    layer8_outputs(4508) <= a xor b;
    layer8_outputs(4509) <= not a;
    layer8_outputs(4510) <= a;
    layer8_outputs(4511) <= not a;
    layer8_outputs(4512) <= a and b;
    layer8_outputs(4513) <= not b;
    layer8_outputs(4514) <= not (a xor b);
    layer8_outputs(4515) <= not (a xor b);
    layer8_outputs(4516) <= a and b;
    layer8_outputs(4517) <= a xor b;
    layer8_outputs(4518) <= b;
    layer8_outputs(4519) <= not a or b;
    layer8_outputs(4520) <= not (a or b);
    layer8_outputs(4521) <= a;
    layer8_outputs(4522) <= b and not a;
    layer8_outputs(4523) <= not b or a;
    layer8_outputs(4524) <= a;
    layer8_outputs(4525) <= not (a xor b);
    layer8_outputs(4526) <= not a or b;
    layer8_outputs(4527) <= a or b;
    layer8_outputs(4528) <= a or b;
    layer8_outputs(4529) <= a xor b;
    layer8_outputs(4530) <= a;
    layer8_outputs(4531) <= a;
    layer8_outputs(4532) <= not (a and b);
    layer8_outputs(4533) <= not (a or b);
    layer8_outputs(4534) <= a and b;
    layer8_outputs(4535) <= a;
    layer8_outputs(4536) <= not a or b;
    layer8_outputs(4537) <= b;
    layer8_outputs(4538) <= a;
    layer8_outputs(4539) <= not b;
    layer8_outputs(4540) <= not a;
    layer8_outputs(4541) <= not (a and b);
    layer8_outputs(4542) <= b;
    layer8_outputs(4543) <= not (a xor b);
    layer8_outputs(4544) <= a xor b;
    layer8_outputs(4545) <= not a;
    layer8_outputs(4546) <= not b or a;
    layer8_outputs(4547) <= not b or a;
    layer8_outputs(4548) <= a;
    layer8_outputs(4549) <= a;
    layer8_outputs(4550) <= a or b;
    layer8_outputs(4551) <= not a;
    layer8_outputs(4552) <= not (a xor b);
    layer8_outputs(4553) <= a xor b;
    layer8_outputs(4554) <= a and not b;
    layer8_outputs(4555) <= not a or b;
    layer8_outputs(4556) <= a xor b;
    layer8_outputs(4557) <= not (a xor b);
    layer8_outputs(4558) <= not (a xor b);
    layer8_outputs(4559) <= not (a xor b);
    layer8_outputs(4560) <= b;
    layer8_outputs(4561) <= not a or b;
    layer8_outputs(4562) <= a and b;
    layer8_outputs(4563) <= a and not b;
    layer8_outputs(4564) <= a or b;
    layer8_outputs(4565) <= not (a and b);
    layer8_outputs(4566) <= not (a and b);
    layer8_outputs(4567) <= not b;
    layer8_outputs(4568) <= not a;
    layer8_outputs(4569) <= not b or a;
    layer8_outputs(4570) <= b;
    layer8_outputs(4571) <= not a;
    layer8_outputs(4572) <= a or b;
    layer8_outputs(4573) <= a xor b;
    layer8_outputs(4574) <= b and not a;
    layer8_outputs(4575) <= b;
    layer8_outputs(4576) <= not a or b;
    layer8_outputs(4577) <= not (a or b);
    layer8_outputs(4578) <= a xor b;
    layer8_outputs(4579) <= not a;
    layer8_outputs(4580) <= a xor b;
    layer8_outputs(4581) <= a and not b;
    layer8_outputs(4582) <= a or b;
    layer8_outputs(4583) <= not (a and b);
    layer8_outputs(4584) <= not (a xor b);
    layer8_outputs(4585) <= b;
    layer8_outputs(4586) <= not b;
    layer8_outputs(4587) <= b;
    layer8_outputs(4588) <= a xor b;
    layer8_outputs(4589) <= not a;
    layer8_outputs(4590) <= a xor b;
    layer8_outputs(4591) <= a and b;
    layer8_outputs(4592) <= not b;
    layer8_outputs(4593) <= a and b;
    layer8_outputs(4594) <= not a;
    layer8_outputs(4595) <= a xor b;
    layer8_outputs(4596) <= not a or b;
    layer8_outputs(4597) <= a xor b;
    layer8_outputs(4598) <= not (a xor b);
    layer8_outputs(4599) <= b;
    layer8_outputs(4600) <= not (a xor b);
    layer8_outputs(4601) <= not (a or b);
    layer8_outputs(4602) <= b;
    layer8_outputs(4603) <= not (a xor b);
    layer8_outputs(4604) <= not (a and b);
    layer8_outputs(4605) <= not b;
    layer8_outputs(4606) <= not b;
    layer8_outputs(4607) <= a and b;
    layer8_outputs(4608) <= a;
    layer8_outputs(4609) <= not (a xor b);
    layer8_outputs(4610) <= b;
    layer8_outputs(4611) <= a;
    layer8_outputs(4612) <= a and not b;
    layer8_outputs(4613) <= b and not a;
    layer8_outputs(4614) <= a and not b;
    layer8_outputs(4615) <= not (a xor b);
    layer8_outputs(4616) <= a xor b;
    layer8_outputs(4617) <= a xor b;
    layer8_outputs(4618) <= not a;
    layer8_outputs(4619) <= a;
    layer8_outputs(4620) <= not b or a;
    layer8_outputs(4621) <= not a;
    layer8_outputs(4622) <= a or b;
    layer8_outputs(4623) <= a xor b;
    layer8_outputs(4624) <= a and not b;
    layer8_outputs(4625) <= not (a or b);
    layer8_outputs(4626) <= a;
    layer8_outputs(4627) <= a xor b;
    layer8_outputs(4628) <= a xor b;
    layer8_outputs(4629) <= not b;
    layer8_outputs(4630) <= not a or b;
    layer8_outputs(4631) <= b;
    layer8_outputs(4632) <= a xor b;
    layer8_outputs(4633) <= not (a xor b);
    layer8_outputs(4634) <= not a;
    layer8_outputs(4635) <= a xor b;
    layer8_outputs(4636) <= b;
    layer8_outputs(4637) <= b;
    layer8_outputs(4638) <= not a;
    layer8_outputs(4639) <= a and b;
    layer8_outputs(4640) <= not (a and b);
    layer8_outputs(4641) <= a;
    layer8_outputs(4642) <= not (a xor b);
    layer8_outputs(4643) <= not b or a;
    layer8_outputs(4644) <= not (a xor b);
    layer8_outputs(4645) <= not (a or b);
    layer8_outputs(4646) <= a or b;
    layer8_outputs(4647) <= a xor b;
    layer8_outputs(4648) <= not b or a;
    layer8_outputs(4649) <= not b or a;
    layer8_outputs(4650) <= not b or a;
    layer8_outputs(4651) <= not b;
    layer8_outputs(4652) <= a;
    layer8_outputs(4653) <= not a or b;
    layer8_outputs(4654) <= not a;
    layer8_outputs(4655) <= b;
    layer8_outputs(4656) <= b;
    layer8_outputs(4657) <= a xor b;
    layer8_outputs(4658) <= a xor b;
    layer8_outputs(4659) <= not a or b;
    layer8_outputs(4660) <= a and b;
    layer8_outputs(4661) <= b;
    layer8_outputs(4662) <= a xor b;
    layer8_outputs(4663) <= not b;
    layer8_outputs(4664) <= not a;
    layer8_outputs(4665) <= a and b;
    layer8_outputs(4666) <= a;
    layer8_outputs(4667) <= b;
    layer8_outputs(4668) <= not (a or b);
    layer8_outputs(4669) <= not b or a;
    layer8_outputs(4670) <= not a;
    layer8_outputs(4671) <= b and not a;
    layer8_outputs(4672) <= a xor b;
    layer8_outputs(4673) <= not a;
    layer8_outputs(4674) <= not (a and b);
    layer8_outputs(4675) <= a xor b;
    layer8_outputs(4676) <= b and not a;
    layer8_outputs(4677) <= not b;
    layer8_outputs(4678) <= a;
    layer8_outputs(4679) <= not (a xor b);
    layer8_outputs(4680) <= a and b;
    layer8_outputs(4681) <= not a or b;
    layer8_outputs(4682) <= not a;
    layer8_outputs(4683) <= not b;
    layer8_outputs(4684) <= a or b;
    layer8_outputs(4685) <= a;
    layer8_outputs(4686) <= not (a xor b);
    layer8_outputs(4687) <= a or b;
    layer8_outputs(4688) <= b and not a;
    layer8_outputs(4689) <= a and b;
    layer8_outputs(4690) <= a;
    layer8_outputs(4691) <= a xor b;
    layer8_outputs(4692) <= a xor b;
    layer8_outputs(4693) <= b;
    layer8_outputs(4694) <= b;
    layer8_outputs(4695) <= b and not a;
    layer8_outputs(4696) <= a;
    layer8_outputs(4697) <= not b;
    layer8_outputs(4698) <= not a or b;
    layer8_outputs(4699) <= not b;
    layer8_outputs(4700) <= a or b;
    layer8_outputs(4701) <= a and not b;
    layer8_outputs(4702) <= a xor b;
    layer8_outputs(4703) <= a;
    layer8_outputs(4704) <= a;
    layer8_outputs(4705) <= not b;
    layer8_outputs(4706) <= not (a and b);
    layer8_outputs(4707) <= a and not b;
    layer8_outputs(4708) <= not a;
    layer8_outputs(4709) <= not a;
    layer8_outputs(4710) <= b;
    layer8_outputs(4711) <= b;
    layer8_outputs(4712) <= not b;
    layer8_outputs(4713) <= b;
    layer8_outputs(4714) <= not b or a;
    layer8_outputs(4715) <= not b;
    layer8_outputs(4716) <= a and b;
    layer8_outputs(4717) <= a xor b;
    layer8_outputs(4718) <= a xor b;
    layer8_outputs(4719) <= b;
    layer8_outputs(4720) <= a or b;
    layer8_outputs(4721) <= a;
    layer8_outputs(4722) <= b;
    layer8_outputs(4723) <= b;
    layer8_outputs(4724) <= 1'b0;
    layer8_outputs(4725) <= not b;
    layer8_outputs(4726) <= not a;
    layer8_outputs(4727) <= not b;
    layer8_outputs(4728) <= not (a and b);
    layer8_outputs(4729) <= not a;
    layer8_outputs(4730) <= a and not b;
    layer8_outputs(4731) <= b and not a;
    layer8_outputs(4732) <= not b;
    layer8_outputs(4733) <= b and not a;
    layer8_outputs(4734) <= not (a and b);
    layer8_outputs(4735) <= not (a and b);
    layer8_outputs(4736) <= a;
    layer8_outputs(4737) <= not b or a;
    layer8_outputs(4738) <= not a;
    layer8_outputs(4739) <= a;
    layer8_outputs(4740) <= a xor b;
    layer8_outputs(4741) <= not (a xor b);
    layer8_outputs(4742) <= a;
    layer8_outputs(4743) <= not (a or b);
    layer8_outputs(4744) <= not a;
    layer8_outputs(4745) <= not a;
    layer8_outputs(4746) <= a;
    layer8_outputs(4747) <= a xor b;
    layer8_outputs(4748) <= b;
    layer8_outputs(4749) <= not a;
    layer8_outputs(4750) <= a xor b;
    layer8_outputs(4751) <= not (a xor b);
    layer8_outputs(4752) <= a or b;
    layer8_outputs(4753) <= not b or a;
    layer8_outputs(4754) <= not (a xor b);
    layer8_outputs(4755) <= b and not a;
    layer8_outputs(4756) <= a xor b;
    layer8_outputs(4757) <= a or b;
    layer8_outputs(4758) <= a and b;
    layer8_outputs(4759) <= not a or b;
    layer8_outputs(4760) <= b;
    layer8_outputs(4761) <= not (a or b);
    layer8_outputs(4762) <= a or b;
    layer8_outputs(4763) <= b;
    layer8_outputs(4764) <= a xor b;
    layer8_outputs(4765) <= not (a xor b);
    layer8_outputs(4766) <= a;
    layer8_outputs(4767) <= a and b;
    layer8_outputs(4768) <= not (a xor b);
    layer8_outputs(4769) <= not a;
    layer8_outputs(4770) <= a;
    layer8_outputs(4771) <= a xor b;
    layer8_outputs(4772) <= not (a xor b);
    layer8_outputs(4773) <= not b;
    layer8_outputs(4774) <= not (a xor b);
    layer8_outputs(4775) <= a xor b;
    layer8_outputs(4776) <= not a;
    layer8_outputs(4777) <= not a;
    layer8_outputs(4778) <= a and not b;
    layer8_outputs(4779) <= a xor b;
    layer8_outputs(4780) <= a or b;
    layer8_outputs(4781) <= not a;
    layer8_outputs(4782) <= a;
    layer8_outputs(4783) <= not (a xor b);
    layer8_outputs(4784) <= a and not b;
    layer8_outputs(4785) <= not (a xor b);
    layer8_outputs(4786) <= not b;
    layer8_outputs(4787) <= not b or a;
    layer8_outputs(4788) <= not (a and b);
    layer8_outputs(4789) <= a;
    layer8_outputs(4790) <= a and b;
    layer8_outputs(4791) <= not b;
    layer8_outputs(4792) <= not a;
    layer8_outputs(4793) <= a or b;
    layer8_outputs(4794) <= a xor b;
    layer8_outputs(4795) <= a;
    layer8_outputs(4796) <= not a;
    layer8_outputs(4797) <= not b;
    layer8_outputs(4798) <= b;
    layer8_outputs(4799) <= a;
    layer8_outputs(4800) <= not (a and b);
    layer8_outputs(4801) <= a xor b;
    layer8_outputs(4802) <= not (a and b);
    layer8_outputs(4803) <= not (a or b);
    layer8_outputs(4804) <= not (a or b);
    layer8_outputs(4805) <= not (a xor b);
    layer8_outputs(4806) <= not (a or b);
    layer8_outputs(4807) <= not (a and b);
    layer8_outputs(4808) <= a xor b;
    layer8_outputs(4809) <= a;
    layer8_outputs(4810) <= not a;
    layer8_outputs(4811) <= not a;
    layer8_outputs(4812) <= not a;
    layer8_outputs(4813) <= a xor b;
    layer8_outputs(4814) <= not (a xor b);
    layer8_outputs(4815) <= a;
    layer8_outputs(4816) <= a and not b;
    layer8_outputs(4817) <= a and b;
    layer8_outputs(4818) <= a;
    layer8_outputs(4819) <= not a;
    layer8_outputs(4820) <= not a or b;
    layer8_outputs(4821) <= a and b;
    layer8_outputs(4822) <= a;
    layer8_outputs(4823) <= b and not a;
    layer8_outputs(4824) <= not b;
    layer8_outputs(4825) <= a xor b;
    layer8_outputs(4826) <= b;
    layer8_outputs(4827) <= a xor b;
    layer8_outputs(4828) <= b;
    layer8_outputs(4829) <= not a;
    layer8_outputs(4830) <= not (a and b);
    layer8_outputs(4831) <= a xor b;
    layer8_outputs(4832) <= a;
    layer8_outputs(4833) <= 1'b1;
    layer8_outputs(4834) <= a xor b;
    layer8_outputs(4835) <= a xor b;
    layer8_outputs(4836) <= a and b;
    layer8_outputs(4837) <= a and b;
    layer8_outputs(4838) <= a xor b;
    layer8_outputs(4839) <= 1'b1;
    layer8_outputs(4840) <= 1'b1;
    layer8_outputs(4841) <= b;
    layer8_outputs(4842) <= b;
    layer8_outputs(4843) <= not a;
    layer8_outputs(4844) <= not b;
    layer8_outputs(4845) <= a;
    layer8_outputs(4846) <= a;
    layer8_outputs(4847) <= not b;
    layer8_outputs(4848) <= b;
    layer8_outputs(4849) <= a;
    layer8_outputs(4850) <= not (a or b);
    layer8_outputs(4851) <= not (a xor b);
    layer8_outputs(4852) <= not b;
    layer8_outputs(4853) <= a xor b;
    layer8_outputs(4854) <= a and b;
    layer8_outputs(4855) <= a and not b;
    layer8_outputs(4856) <= not (a xor b);
    layer8_outputs(4857) <= a;
    layer8_outputs(4858) <= not a;
    layer8_outputs(4859) <= not (a or b);
    layer8_outputs(4860) <= b;
    layer8_outputs(4861) <= a;
    layer8_outputs(4862) <= b;
    layer8_outputs(4863) <= a;
    layer8_outputs(4864) <= not (a or b);
    layer8_outputs(4865) <= 1'b0;
    layer8_outputs(4866) <= not (a xor b);
    layer8_outputs(4867) <= not (a and b);
    layer8_outputs(4868) <= a;
    layer8_outputs(4869) <= b and not a;
    layer8_outputs(4870) <= a or b;
    layer8_outputs(4871) <= not b;
    layer8_outputs(4872) <= a;
    layer8_outputs(4873) <= b;
    layer8_outputs(4874) <= a xor b;
    layer8_outputs(4875) <= a;
    layer8_outputs(4876) <= b;
    layer8_outputs(4877) <= not a;
    layer8_outputs(4878) <= a and not b;
    layer8_outputs(4879) <= not a;
    layer8_outputs(4880) <= a xor b;
    layer8_outputs(4881) <= not a;
    layer8_outputs(4882) <= not b;
    layer8_outputs(4883) <= b;
    layer8_outputs(4884) <= a xor b;
    layer8_outputs(4885) <= 1'b1;
    layer8_outputs(4886) <= a and b;
    layer8_outputs(4887) <= a and b;
    layer8_outputs(4888) <= not a;
    layer8_outputs(4889) <= a xor b;
    layer8_outputs(4890) <= not (a xor b);
    layer8_outputs(4891) <= a;
    layer8_outputs(4892) <= a;
    layer8_outputs(4893) <= a and not b;
    layer8_outputs(4894) <= a and b;
    layer8_outputs(4895) <= not (a xor b);
    layer8_outputs(4896) <= not b;
    layer8_outputs(4897) <= not b;
    layer8_outputs(4898) <= not (a or b);
    layer8_outputs(4899) <= a and not b;
    layer8_outputs(4900) <= a and b;
    layer8_outputs(4901) <= b and not a;
    layer8_outputs(4902) <= not (a and b);
    layer8_outputs(4903) <= b;
    layer8_outputs(4904) <= a xor b;
    layer8_outputs(4905) <= a;
    layer8_outputs(4906) <= b;
    layer8_outputs(4907) <= not a or b;
    layer8_outputs(4908) <= b;
    layer8_outputs(4909) <= a;
    layer8_outputs(4910) <= 1'b1;
    layer8_outputs(4911) <= not b;
    layer8_outputs(4912) <= not a;
    layer8_outputs(4913) <= a and b;
    layer8_outputs(4914) <= b;
    layer8_outputs(4915) <= a xor b;
    layer8_outputs(4916) <= a and not b;
    layer8_outputs(4917) <= a xor b;
    layer8_outputs(4918) <= not (a xor b);
    layer8_outputs(4919) <= not (a or b);
    layer8_outputs(4920) <= b;
    layer8_outputs(4921) <= not a or b;
    layer8_outputs(4922) <= not (a or b);
    layer8_outputs(4923) <= not b;
    layer8_outputs(4924) <= not a;
    layer8_outputs(4925) <= not (a and b);
    layer8_outputs(4926) <= not (a xor b);
    layer8_outputs(4927) <= not (a and b);
    layer8_outputs(4928) <= not b;
    layer8_outputs(4929) <= not (a and b);
    layer8_outputs(4930) <= a and not b;
    layer8_outputs(4931) <= not (a xor b);
    layer8_outputs(4932) <= b and not a;
    layer8_outputs(4933) <= not a;
    layer8_outputs(4934) <= not (a and b);
    layer8_outputs(4935) <= not b;
    layer8_outputs(4936) <= not (a or b);
    layer8_outputs(4937) <= a and not b;
    layer8_outputs(4938) <= b;
    layer8_outputs(4939) <= not (a xor b);
    layer8_outputs(4940) <= not b;
    layer8_outputs(4941) <= not (a xor b);
    layer8_outputs(4942) <= not b or a;
    layer8_outputs(4943) <= b;
    layer8_outputs(4944) <= a;
    layer8_outputs(4945) <= not a;
    layer8_outputs(4946) <= not (a or b);
    layer8_outputs(4947) <= not (a or b);
    layer8_outputs(4948) <= not (a or b);
    layer8_outputs(4949) <= not (a or b);
    layer8_outputs(4950) <= a;
    layer8_outputs(4951) <= not (a xor b);
    layer8_outputs(4952) <= not a;
    layer8_outputs(4953) <= a or b;
    layer8_outputs(4954) <= a or b;
    layer8_outputs(4955) <= not a;
    layer8_outputs(4956) <= a xor b;
    layer8_outputs(4957) <= not b;
    layer8_outputs(4958) <= a xor b;
    layer8_outputs(4959) <= not (a xor b);
    layer8_outputs(4960) <= not a;
    layer8_outputs(4961) <= a;
    layer8_outputs(4962) <= not a;
    layer8_outputs(4963) <= not b;
    layer8_outputs(4964) <= a xor b;
    layer8_outputs(4965) <= a;
    layer8_outputs(4966) <= a and not b;
    layer8_outputs(4967) <= not b or a;
    layer8_outputs(4968) <= not (a or b);
    layer8_outputs(4969) <= a and not b;
    layer8_outputs(4970) <= not (a and b);
    layer8_outputs(4971) <= not (a and b);
    layer8_outputs(4972) <= a and not b;
    layer8_outputs(4973) <= a xor b;
    layer8_outputs(4974) <= a and not b;
    layer8_outputs(4975) <= a and b;
    layer8_outputs(4976) <= a and b;
    layer8_outputs(4977) <= not (a xor b);
    layer8_outputs(4978) <= a and b;
    layer8_outputs(4979) <= not (a xor b);
    layer8_outputs(4980) <= not (a xor b);
    layer8_outputs(4981) <= b;
    layer8_outputs(4982) <= b and not a;
    layer8_outputs(4983) <= a;
    layer8_outputs(4984) <= 1'b1;
    layer8_outputs(4985) <= b;
    layer8_outputs(4986) <= a;
    layer8_outputs(4987) <= a;
    layer8_outputs(4988) <= a;
    layer8_outputs(4989) <= not (a xor b);
    layer8_outputs(4990) <= a;
    layer8_outputs(4991) <= not (a xor b);
    layer8_outputs(4992) <= not b;
    layer8_outputs(4993) <= not (a xor b);
    layer8_outputs(4994) <= a or b;
    layer8_outputs(4995) <= a;
    layer8_outputs(4996) <= not (a xor b);
    layer8_outputs(4997) <= not b;
    layer8_outputs(4998) <= a;
    layer8_outputs(4999) <= a xor b;
    layer8_outputs(5000) <= not a or b;
    layer8_outputs(5001) <= not (a xor b);
    layer8_outputs(5002) <= a xor b;
    layer8_outputs(5003) <= a and not b;
    layer8_outputs(5004) <= a and not b;
    layer8_outputs(5005) <= a xor b;
    layer8_outputs(5006) <= not b;
    layer8_outputs(5007) <= not (a and b);
    layer8_outputs(5008) <= a;
    layer8_outputs(5009) <= a xor b;
    layer8_outputs(5010) <= not (a xor b);
    layer8_outputs(5011) <= not b;
    layer8_outputs(5012) <= 1'b1;
    layer8_outputs(5013) <= a and b;
    layer8_outputs(5014) <= not (a xor b);
    layer8_outputs(5015) <= not b;
    layer8_outputs(5016) <= a;
    layer8_outputs(5017) <= not (a and b);
    layer8_outputs(5018) <= b;
    layer8_outputs(5019) <= not (a or b);
    layer8_outputs(5020) <= not (a and b);
    layer8_outputs(5021) <= a xor b;
    layer8_outputs(5022) <= not b;
    layer8_outputs(5023) <= a;
    layer8_outputs(5024) <= not (a xor b);
    layer8_outputs(5025) <= not a;
    layer8_outputs(5026) <= a and not b;
    layer8_outputs(5027) <= not b;
    layer8_outputs(5028) <= a and b;
    layer8_outputs(5029) <= not a;
    layer8_outputs(5030) <= a xor b;
    layer8_outputs(5031) <= not b or a;
    layer8_outputs(5032) <= a or b;
    layer8_outputs(5033) <= a xor b;
    layer8_outputs(5034) <= b;
    layer8_outputs(5035) <= b;
    layer8_outputs(5036) <= b and not a;
    layer8_outputs(5037) <= a;
    layer8_outputs(5038) <= a xor b;
    layer8_outputs(5039) <= a;
    layer8_outputs(5040) <= b and not a;
    layer8_outputs(5041) <= b;
    layer8_outputs(5042) <= 1'b0;
    layer8_outputs(5043) <= a;
    layer8_outputs(5044) <= 1'b1;
    layer8_outputs(5045) <= b;
    layer8_outputs(5046) <= not a;
    layer8_outputs(5047) <= not (a and b);
    layer8_outputs(5048) <= b;
    layer8_outputs(5049) <= a xor b;
    layer8_outputs(5050) <= b;
    layer8_outputs(5051) <= b;
    layer8_outputs(5052) <= a or b;
    layer8_outputs(5053) <= a;
    layer8_outputs(5054) <= not a or b;
    layer8_outputs(5055) <= b;
    layer8_outputs(5056) <= a xor b;
    layer8_outputs(5057) <= not b;
    layer8_outputs(5058) <= b;
    layer8_outputs(5059) <= b;
    layer8_outputs(5060) <= not (a or b);
    layer8_outputs(5061) <= not a;
    layer8_outputs(5062) <= b;
    layer8_outputs(5063) <= not a;
    layer8_outputs(5064) <= b and not a;
    layer8_outputs(5065) <= not b or a;
    layer8_outputs(5066) <= b and not a;
    layer8_outputs(5067) <= a or b;
    layer8_outputs(5068) <= not a;
    layer8_outputs(5069) <= a and b;
    layer8_outputs(5070) <= not b;
    layer8_outputs(5071) <= a and b;
    layer8_outputs(5072) <= a and b;
    layer8_outputs(5073) <= a or b;
    layer8_outputs(5074) <= not a;
    layer8_outputs(5075) <= not a or b;
    layer8_outputs(5076) <= a;
    layer8_outputs(5077) <= b;
    layer8_outputs(5078) <= a;
    layer8_outputs(5079) <= not (a xor b);
    layer8_outputs(5080) <= a or b;
    layer8_outputs(5081) <= not (a or b);
    layer8_outputs(5082) <= not a or b;
    layer8_outputs(5083) <= not (a xor b);
    layer8_outputs(5084) <= not (a xor b);
    layer8_outputs(5085) <= b;
    layer8_outputs(5086) <= a xor b;
    layer8_outputs(5087) <= b and not a;
    layer8_outputs(5088) <= not b or a;
    layer8_outputs(5089) <= a or b;
    layer8_outputs(5090) <= b and not a;
    layer8_outputs(5091) <= not b or a;
    layer8_outputs(5092) <= not (a xor b);
    layer8_outputs(5093) <= not a;
    layer8_outputs(5094) <= not (a and b);
    layer8_outputs(5095) <= not a;
    layer8_outputs(5096) <= a;
    layer8_outputs(5097) <= not (a and b);
    layer8_outputs(5098) <= not a;
    layer8_outputs(5099) <= not a or b;
    layer8_outputs(5100) <= a or b;
    layer8_outputs(5101) <= b;
    layer8_outputs(5102) <= not (a and b);
    layer8_outputs(5103) <= a and not b;
    layer8_outputs(5104) <= not a;
    layer8_outputs(5105) <= not b;
    layer8_outputs(5106) <= b;
    layer8_outputs(5107) <= not a;
    layer8_outputs(5108) <= not (a xor b);
    layer8_outputs(5109) <= a xor b;
    layer8_outputs(5110) <= not (a and b);
    layer8_outputs(5111) <= a;
    layer8_outputs(5112) <= not b;
    layer8_outputs(5113) <= not b;
    layer8_outputs(5114) <= a;
    layer8_outputs(5115) <= not (a xor b);
    layer8_outputs(5116) <= a xor b;
    layer8_outputs(5117) <= not (a xor b);
    layer8_outputs(5118) <= not a;
    layer8_outputs(5119) <= not (a xor b);
    layer8_outputs(5120) <= a xor b;
    layer8_outputs(5121) <= not b;
    layer8_outputs(5122) <= not a or b;
    layer8_outputs(5123) <= a or b;
    layer8_outputs(5124) <= not a;
    layer8_outputs(5125) <= a;
    layer8_outputs(5126) <= not (a or b);
    layer8_outputs(5127) <= not (a xor b);
    layer8_outputs(5128) <= not b;
    layer8_outputs(5129) <= a xor b;
    layer8_outputs(5130) <= 1'b1;
    layer8_outputs(5131) <= a and not b;
    layer8_outputs(5132) <= a xor b;
    layer8_outputs(5133) <= not a;
    layer8_outputs(5134) <= a xor b;
    layer8_outputs(5135) <= a xor b;
    layer8_outputs(5136) <= not (a xor b);
    layer8_outputs(5137) <= not a;
    layer8_outputs(5138) <= a xor b;
    layer8_outputs(5139) <= not a or b;
    layer8_outputs(5140) <= not b;
    layer8_outputs(5141) <= not b;
    layer8_outputs(5142) <= not b;
    layer8_outputs(5143) <= not (a xor b);
    layer8_outputs(5144) <= not b;
    layer8_outputs(5145) <= not (a and b);
    layer8_outputs(5146) <= not b;
    layer8_outputs(5147) <= a;
    layer8_outputs(5148) <= not (a or b);
    layer8_outputs(5149) <= not a;
    layer8_outputs(5150) <= not (a and b);
    layer8_outputs(5151) <= not (a and b);
    layer8_outputs(5152) <= a xor b;
    layer8_outputs(5153) <= b and not a;
    layer8_outputs(5154) <= not a or b;
    layer8_outputs(5155) <= not (a xor b);
    layer8_outputs(5156) <= b;
    layer8_outputs(5157) <= b and not a;
    layer8_outputs(5158) <= not a;
    layer8_outputs(5159) <= not (a xor b);
    layer8_outputs(5160) <= a;
    layer8_outputs(5161) <= not b;
    layer8_outputs(5162) <= not (a or b);
    layer8_outputs(5163) <= not b;
    layer8_outputs(5164) <= a xor b;
    layer8_outputs(5165) <= b;
    layer8_outputs(5166) <= a xor b;
    layer8_outputs(5167) <= not b or a;
    layer8_outputs(5168) <= not (a and b);
    layer8_outputs(5169) <= not b;
    layer8_outputs(5170) <= a and not b;
    layer8_outputs(5171) <= not b;
    layer8_outputs(5172) <= a xor b;
    layer8_outputs(5173) <= b;
    layer8_outputs(5174) <= not b;
    layer8_outputs(5175) <= a and b;
    layer8_outputs(5176) <= a and b;
    layer8_outputs(5177) <= not (a and b);
    layer8_outputs(5178) <= b;
    layer8_outputs(5179) <= a or b;
    layer8_outputs(5180) <= not b or a;
    layer8_outputs(5181) <= not b;
    layer8_outputs(5182) <= a or b;
    layer8_outputs(5183) <= not a;
    layer8_outputs(5184) <= b;
    layer8_outputs(5185) <= 1'b0;
    layer8_outputs(5186) <= a;
    layer8_outputs(5187) <= not (a xor b);
    layer8_outputs(5188) <= not (a xor b);
    layer8_outputs(5189) <= not a;
    layer8_outputs(5190) <= a xor b;
    layer8_outputs(5191) <= a;
    layer8_outputs(5192) <= not (a xor b);
    layer8_outputs(5193) <= b;
    layer8_outputs(5194) <= not a or b;
    layer8_outputs(5195) <= not a or b;
    layer8_outputs(5196) <= not b;
    layer8_outputs(5197) <= a and not b;
    layer8_outputs(5198) <= not (a xor b);
    layer8_outputs(5199) <= a xor b;
    layer8_outputs(5200) <= a;
    layer8_outputs(5201) <= not (a xor b);
    layer8_outputs(5202) <= b and not a;
    layer8_outputs(5203) <= b and not a;
    layer8_outputs(5204) <= not (a xor b);
    layer8_outputs(5205) <= a and b;
    layer8_outputs(5206) <= a xor b;
    layer8_outputs(5207) <= a and b;
    layer8_outputs(5208) <= 1'b0;
    layer8_outputs(5209) <= not (a and b);
    layer8_outputs(5210) <= 1'b0;
    layer8_outputs(5211) <= not (a or b);
    layer8_outputs(5212) <= not (a xor b);
    layer8_outputs(5213) <= a and b;
    layer8_outputs(5214) <= a;
    layer8_outputs(5215) <= a;
    layer8_outputs(5216) <= b and not a;
    layer8_outputs(5217) <= not a;
    layer8_outputs(5218) <= not (a or b);
    layer8_outputs(5219) <= not a;
    layer8_outputs(5220) <= b;
    layer8_outputs(5221) <= b;
    layer8_outputs(5222) <= not (a xor b);
    layer8_outputs(5223) <= not b or a;
    layer8_outputs(5224) <= a;
    layer8_outputs(5225) <= not a;
    layer8_outputs(5226) <= a xor b;
    layer8_outputs(5227) <= not (a xor b);
    layer8_outputs(5228) <= not (a and b);
    layer8_outputs(5229) <= not a;
    layer8_outputs(5230) <= a xor b;
    layer8_outputs(5231) <= a xor b;
    layer8_outputs(5232) <= a and not b;
    layer8_outputs(5233) <= b;
    layer8_outputs(5234) <= a;
    layer8_outputs(5235) <= b;
    layer8_outputs(5236) <= a;
    layer8_outputs(5237) <= a and b;
    layer8_outputs(5238) <= a xor b;
    layer8_outputs(5239) <= not b;
    layer8_outputs(5240) <= not a;
    layer8_outputs(5241) <= a or b;
    layer8_outputs(5242) <= a xor b;
    layer8_outputs(5243) <= a;
    layer8_outputs(5244) <= a;
    layer8_outputs(5245) <= a xor b;
    layer8_outputs(5246) <= a and b;
    layer8_outputs(5247) <= not (a xor b);
    layer8_outputs(5248) <= not b;
    layer8_outputs(5249) <= not b;
    layer8_outputs(5250) <= a;
    layer8_outputs(5251) <= not b;
    layer8_outputs(5252) <= a and not b;
    layer8_outputs(5253) <= a or b;
    layer8_outputs(5254) <= not a;
    layer8_outputs(5255) <= not a or b;
    layer8_outputs(5256) <= not (a xor b);
    layer8_outputs(5257) <= not (a or b);
    layer8_outputs(5258) <= a xor b;
    layer8_outputs(5259) <= not b or a;
    layer8_outputs(5260) <= a;
    layer8_outputs(5261) <= not b;
    layer8_outputs(5262) <= not b;
    layer8_outputs(5263) <= b;
    layer8_outputs(5264) <= a;
    layer8_outputs(5265) <= b;
    layer8_outputs(5266) <= not (a or b);
    layer8_outputs(5267) <= a and not b;
    layer8_outputs(5268) <= not (a or b);
    layer8_outputs(5269) <= a or b;
    layer8_outputs(5270) <= a and b;
    layer8_outputs(5271) <= a or b;
    layer8_outputs(5272) <= not a or b;
    layer8_outputs(5273) <= not (a or b);
    layer8_outputs(5274) <= a;
    layer8_outputs(5275) <= not (a xor b);
    layer8_outputs(5276) <= b and not a;
    layer8_outputs(5277) <= not a or b;
    layer8_outputs(5278) <= a or b;
    layer8_outputs(5279) <= not b;
    layer8_outputs(5280) <= b;
    layer8_outputs(5281) <= b and not a;
    layer8_outputs(5282) <= not b or a;
    layer8_outputs(5283) <= b;
    layer8_outputs(5284) <= not (a or b);
    layer8_outputs(5285) <= a and not b;
    layer8_outputs(5286) <= a;
    layer8_outputs(5287) <= a;
    layer8_outputs(5288) <= not b;
    layer8_outputs(5289) <= not a;
    layer8_outputs(5290) <= not b;
    layer8_outputs(5291) <= b;
    layer8_outputs(5292) <= a xor b;
    layer8_outputs(5293) <= not a;
    layer8_outputs(5294) <= not a;
    layer8_outputs(5295) <= not b;
    layer8_outputs(5296) <= a and not b;
    layer8_outputs(5297) <= a and not b;
    layer8_outputs(5298) <= a xor b;
    layer8_outputs(5299) <= a;
    layer8_outputs(5300) <= a;
    layer8_outputs(5301) <= not b;
    layer8_outputs(5302) <= a or b;
    layer8_outputs(5303) <= not (a or b);
    layer8_outputs(5304) <= a xor b;
    layer8_outputs(5305) <= not a;
    layer8_outputs(5306) <= a and not b;
    layer8_outputs(5307) <= b and not a;
    layer8_outputs(5308) <= a and not b;
    layer8_outputs(5309) <= b;
    layer8_outputs(5310) <= not b;
    layer8_outputs(5311) <= a;
    layer8_outputs(5312) <= not (a xor b);
    layer8_outputs(5313) <= a;
    layer8_outputs(5314) <= a;
    layer8_outputs(5315) <= not a;
    layer8_outputs(5316) <= a;
    layer8_outputs(5317) <= a xor b;
    layer8_outputs(5318) <= a and not b;
    layer8_outputs(5319) <= not b or a;
    layer8_outputs(5320) <= a and b;
    layer8_outputs(5321) <= not (a xor b);
    layer8_outputs(5322) <= a and b;
    layer8_outputs(5323) <= not (a xor b);
    layer8_outputs(5324) <= a or b;
    layer8_outputs(5325) <= a xor b;
    layer8_outputs(5326) <= not a;
    layer8_outputs(5327) <= not a;
    layer8_outputs(5328) <= not (a xor b);
    layer8_outputs(5329) <= not a or b;
    layer8_outputs(5330) <= not a;
    layer8_outputs(5331) <= a;
    layer8_outputs(5332) <= not (a xor b);
    layer8_outputs(5333) <= not b or a;
    layer8_outputs(5334) <= a xor b;
    layer8_outputs(5335) <= not a;
    layer8_outputs(5336) <= not b or a;
    layer8_outputs(5337) <= not b or a;
    layer8_outputs(5338) <= a and not b;
    layer8_outputs(5339) <= a xor b;
    layer8_outputs(5340) <= not a;
    layer8_outputs(5341) <= a;
    layer8_outputs(5342) <= not (a xor b);
    layer8_outputs(5343) <= not b;
    layer8_outputs(5344) <= not b;
    layer8_outputs(5345) <= not (a and b);
    layer8_outputs(5346) <= not b;
    layer8_outputs(5347) <= a xor b;
    layer8_outputs(5348) <= a;
    layer8_outputs(5349) <= not b;
    layer8_outputs(5350) <= not (a xor b);
    layer8_outputs(5351) <= a or b;
    layer8_outputs(5352) <= b;
    layer8_outputs(5353) <= a xor b;
    layer8_outputs(5354) <= not b;
    layer8_outputs(5355) <= a xor b;
    layer8_outputs(5356) <= a xor b;
    layer8_outputs(5357) <= not b;
    layer8_outputs(5358) <= not a;
    layer8_outputs(5359) <= b;
    layer8_outputs(5360) <= not (a xor b);
    layer8_outputs(5361) <= a and b;
    layer8_outputs(5362) <= a xor b;
    layer8_outputs(5363) <= not a;
    layer8_outputs(5364) <= not b;
    layer8_outputs(5365) <= a or b;
    layer8_outputs(5366) <= not a;
    layer8_outputs(5367) <= not b;
    layer8_outputs(5368) <= b;
    layer8_outputs(5369) <= not b;
    layer8_outputs(5370) <= a;
    layer8_outputs(5371) <= not a;
    layer8_outputs(5372) <= a and b;
    layer8_outputs(5373) <= not a or b;
    layer8_outputs(5374) <= not a;
    layer8_outputs(5375) <= a and not b;
    layer8_outputs(5376) <= not (a or b);
    layer8_outputs(5377) <= not b or a;
    layer8_outputs(5378) <= a xor b;
    layer8_outputs(5379) <= not a or b;
    layer8_outputs(5380) <= a and b;
    layer8_outputs(5381) <= a;
    layer8_outputs(5382) <= not (a xor b);
    layer8_outputs(5383) <= not (a and b);
    layer8_outputs(5384) <= not b;
    layer8_outputs(5385) <= a or b;
    layer8_outputs(5386) <= a xor b;
    layer8_outputs(5387) <= a xor b;
    layer8_outputs(5388) <= not a;
    layer8_outputs(5389) <= b;
    layer8_outputs(5390) <= not a;
    layer8_outputs(5391) <= not a;
    layer8_outputs(5392) <= not (a and b);
    layer8_outputs(5393) <= a and b;
    layer8_outputs(5394) <= a xor b;
    layer8_outputs(5395) <= a and b;
    layer8_outputs(5396) <= not a or b;
    layer8_outputs(5397) <= a;
    layer8_outputs(5398) <= not a;
    layer8_outputs(5399) <= not a;
    layer8_outputs(5400) <= b;
    layer8_outputs(5401) <= a and not b;
    layer8_outputs(5402) <= b;
    layer8_outputs(5403) <= not (a and b);
    layer8_outputs(5404) <= a or b;
    layer8_outputs(5405) <= not b or a;
    layer8_outputs(5406) <= not b;
    layer8_outputs(5407) <= a and b;
    layer8_outputs(5408) <= not a;
    layer8_outputs(5409) <= not (a xor b);
    layer8_outputs(5410) <= not a;
    layer8_outputs(5411) <= not b;
    layer8_outputs(5412) <= not b;
    layer8_outputs(5413) <= a;
    layer8_outputs(5414) <= not a;
    layer8_outputs(5415) <= a xor b;
    layer8_outputs(5416) <= not (a xor b);
    layer8_outputs(5417) <= not a;
    layer8_outputs(5418) <= a xor b;
    layer8_outputs(5419) <= a xor b;
    layer8_outputs(5420) <= not b;
    layer8_outputs(5421) <= a and not b;
    layer8_outputs(5422) <= a;
    layer8_outputs(5423) <= not b;
    layer8_outputs(5424) <= a;
    layer8_outputs(5425) <= not (a xor b);
    layer8_outputs(5426) <= not b or a;
    layer8_outputs(5427) <= b;
    layer8_outputs(5428) <= a xor b;
    layer8_outputs(5429) <= not b;
    layer8_outputs(5430) <= not (a xor b);
    layer8_outputs(5431) <= a and not b;
    layer8_outputs(5432) <= not (a or b);
    layer8_outputs(5433) <= b;
    layer8_outputs(5434) <= a;
    layer8_outputs(5435) <= not b;
    layer8_outputs(5436) <= a;
    layer8_outputs(5437) <= not (a and b);
    layer8_outputs(5438) <= not b;
    layer8_outputs(5439) <= not a;
    layer8_outputs(5440) <= a;
    layer8_outputs(5441) <= not (a and b);
    layer8_outputs(5442) <= not a;
    layer8_outputs(5443) <= not b or a;
    layer8_outputs(5444) <= not a;
    layer8_outputs(5445) <= b;
    layer8_outputs(5446) <= a or b;
    layer8_outputs(5447) <= a or b;
    layer8_outputs(5448) <= a xor b;
    layer8_outputs(5449) <= not (a or b);
    layer8_outputs(5450) <= a;
    layer8_outputs(5451) <= not a;
    layer8_outputs(5452) <= a or b;
    layer8_outputs(5453) <= b;
    layer8_outputs(5454) <= b;
    layer8_outputs(5455) <= not a;
    layer8_outputs(5456) <= not (a xor b);
    layer8_outputs(5457) <= b;
    layer8_outputs(5458) <= a xor b;
    layer8_outputs(5459) <= not a;
    layer8_outputs(5460) <= a xor b;
    layer8_outputs(5461) <= not (a or b);
    layer8_outputs(5462) <= a;
    layer8_outputs(5463) <= b and not a;
    layer8_outputs(5464) <= a and b;
    layer8_outputs(5465) <= not b;
    layer8_outputs(5466) <= not b or a;
    layer8_outputs(5467) <= a and not b;
    layer8_outputs(5468) <= not b or a;
    layer8_outputs(5469) <= not (a xor b);
    layer8_outputs(5470) <= not a;
    layer8_outputs(5471) <= not b;
    layer8_outputs(5472) <= b;
    layer8_outputs(5473) <= not b;
    layer8_outputs(5474) <= a;
    layer8_outputs(5475) <= not a;
    layer8_outputs(5476) <= not (a and b);
    layer8_outputs(5477) <= not (a xor b);
    layer8_outputs(5478) <= a xor b;
    layer8_outputs(5479) <= b;
    layer8_outputs(5480) <= a xor b;
    layer8_outputs(5481) <= a;
    layer8_outputs(5482) <= a xor b;
    layer8_outputs(5483) <= not a;
    layer8_outputs(5484) <= not b or a;
    layer8_outputs(5485) <= a and not b;
    layer8_outputs(5486) <= b and not a;
    layer8_outputs(5487) <= a;
    layer8_outputs(5488) <= not b or a;
    layer8_outputs(5489) <= a xor b;
    layer8_outputs(5490) <= a xor b;
    layer8_outputs(5491) <= not (a xor b);
    layer8_outputs(5492) <= not a or b;
    layer8_outputs(5493) <= a;
    layer8_outputs(5494) <= not b;
    layer8_outputs(5495) <= a;
    layer8_outputs(5496) <= a and b;
    layer8_outputs(5497) <= a and not b;
    layer8_outputs(5498) <= not b;
    layer8_outputs(5499) <= a and not b;
    layer8_outputs(5500) <= a and not b;
    layer8_outputs(5501) <= a xor b;
    layer8_outputs(5502) <= not (a xor b);
    layer8_outputs(5503) <= not (a or b);
    layer8_outputs(5504) <= b and not a;
    layer8_outputs(5505) <= a;
    layer8_outputs(5506) <= a and b;
    layer8_outputs(5507) <= a;
    layer8_outputs(5508) <= b;
    layer8_outputs(5509) <= not (a xor b);
    layer8_outputs(5510) <= a;
    layer8_outputs(5511) <= not a;
    layer8_outputs(5512) <= not b;
    layer8_outputs(5513) <= a xor b;
    layer8_outputs(5514) <= b;
    layer8_outputs(5515) <= not (a xor b);
    layer8_outputs(5516) <= a;
    layer8_outputs(5517) <= a and not b;
    layer8_outputs(5518) <= not b or a;
    layer8_outputs(5519) <= not a;
    layer8_outputs(5520) <= not (a or b);
    layer8_outputs(5521) <= not (a xor b);
    layer8_outputs(5522) <= b and not a;
    layer8_outputs(5523) <= not (a xor b);
    layer8_outputs(5524) <= a and not b;
    layer8_outputs(5525) <= not (a xor b);
    layer8_outputs(5526) <= not b;
    layer8_outputs(5527) <= a and b;
    layer8_outputs(5528) <= a;
    layer8_outputs(5529) <= not a;
    layer8_outputs(5530) <= not (a xor b);
    layer8_outputs(5531) <= a xor b;
    layer8_outputs(5532) <= a and not b;
    layer8_outputs(5533) <= b;
    layer8_outputs(5534) <= a and b;
    layer8_outputs(5535) <= b;
    layer8_outputs(5536) <= not (a xor b);
    layer8_outputs(5537) <= not (a xor b);
    layer8_outputs(5538) <= not (a and b);
    layer8_outputs(5539) <= a and not b;
    layer8_outputs(5540) <= a;
    layer8_outputs(5541) <= not a;
    layer8_outputs(5542) <= not a;
    layer8_outputs(5543) <= not (a or b);
    layer8_outputs(5544) <= a xor b;
    layer8_outputs(5545) <= a;
    layer8_outputs(5546) <= a and not b;
    layer8_outputs(5547) <= not b;
    layer8_outputs(5548) <= a xor b;
    layer8_outputs(5549) <= 1'b0;
    layer8_outputs(5550) <= a;
    layer8_outputs(5551) <= b;
    layer8_outputs(5552) <= not b;
    layer8_outputs(5553) <= a xor b;
    layer8_outputs(5554) <= not (a xor b);
    layer8_outputs(5555) <= not (a xor b);
    layer8_outputs(5556) <= not a or b;
    layer8_outputs(5557) <= a and b;
    layer8_outputs(5558) <= not a or b;
    layer8_outputs(5559) <= not b or a;
    layer8_outputs(5560) <= a xor b;
    layer8_outputs(5561) <= not (a or b);
    layer8_outputs(5562) <= a and b;
    layer8_outputs(5563) <= a;
    layer8_outputs(5564) <= a xor b;
    layer8_outputs(5565) <= 1'b0;
    layer8_outputs(5566) <= a;
    layer8_outputs(5567) <= not a;
    layer8_outputs(5568) <= a and not b;
    layer8_outputs(5569) <= a xor b;
    layer8_outputs(5570) <= not (a and b);
    layer8_outputs(5571) <= not b or a;
    layer8_outputs(5572) <= not a;
    layer8_outputs(5573) <= not a;
    layer8_outputs(5574) <= not (a xor b);
    layer8_outputs(5575) <= not (a xor b);
    layer8_outputs(5576) <= a xor b;
    layer8_outputs(5577) <= a xor b;
    layer8_outputs(5578) <= not a;
    layer8_outputs(5579) <= a;
    layer8_outputs(5580) <= a;
    layer8_outputs(5581) <= not a;
    layer8_outputs(5582) <= not b or a;
    layer8_outputs(5583) <= not a or b;
    layer8_outputs(5584) <= not a;
    layer8_outputs(5585) <= a and b;
    layer8_outputs(5586) <= b;
    layer8_outputs(5587) <= not (a or b);
    layer8_outputs(5588) <= not (a and b);
    layer8_outputs(5589) <= a;
    layer8_outputs(5590) <= a and b;
    layer8_outputs(5591) <= not a;
    layer8_outputs(5592) <= not (a or b);
    layer8_outputs(5593) <= b;
    layer8_outputs(5594) <= not b;
    layer8_outputs(5595) <= a;
    layer8_outputs(5596) <= a;
    layer8_outputs(5597) <= not b;
    layer8_outputs(5598) <= 1'b0;
    layer8_outputs(5599) <= a xor b;
    layer8_outputs(5600) <= a;
    layer8_outputs(5601) <= b;
    layer8_outputs(5602) <= b;
    layer8_outputs(5603) <= not b or a;
    layer8_outputs(5604) <= a and b;
    layer8_outputs(5605) <= not (a xor b);
    layer8_outputs(5606) <= not (a xor b);
    layer8_outputs(5607) <= a;
    layer8_outputs(5608) <= a or b;
    layer8_outputs(5609) <= b;
    layer8_outputs(5610) <= a and b;
    layer8_outputs(5611) <= not (a xor b);
    layer8_outputs(5612) <= a xor b;
    layer8_outputs(5613) <= not b;
    layer8_outputs(5614) <= b;
    layer8_outputs(5615) <= not a;
    layer8_outputs(5616) <= not b;
    layer8_outputs(5617) <= a;
    layer8_outputs(5618) <= not a;
    layer8_outputs(5619) <= a and not b;
    layer8_outputs(5620) <= a xor b;
    layer8_outputs(5621) <= a;
    layer8_outputs(5622) <= not b;
    layer8_outputs(5623) <= not b;
    layer8_outputs(5624) <= not a;
    layer8_outputs(5625) <= not (a or b);
    layer8_outputs(5626) <= a;
    layer8_outputs(5627) <= not (a xor b);
    layer8_outputs(5628) <= not (a and b);
    layer8_outputs(5629) <= a and not b;
    layer8_outputs(5630) <= not (a or b);
    layer8_outputs(5631) <= not b;
    layer8_outputs(5632) <= b;
    layer8_outputs(5633) <= not (a xor b);
    layer8_outputs(5634) <= not b;
    layer8_outputs(5635) <= b and not a;
    layer8_outputs(5636) <= not a;
    layer8_outputs(5637) <= a xor b;
    layer8_outputs(5638) <= not a;
    layer8_outputs(5639) <= a;
    layer8_outputs(5640) <= not a or b;
    layer8_outputs(5641) <= not (a or b);
    layer8_outputs(5642) <= not b;
    layer8_outputs(5643) <= b and not a;
    layer8_outputs(5644) <= not a;
    layer8_outputs(5645) <= a;
    layer8_outputs(5646) <= not a or b;
    layer8_outputs(5647) <= a xor b;
    layer8_outputs(5648) <= a;
    layer8_outputs(5649) <= a and b;
    layer8_outputs(5650) <= a;
    layer8_outputs(5651) <= a and not b;
    layer8_outputs(5652) <= not b;
    layer8_outputs(5653) <= b;
    layer8_outputs(5654) <= a;
    layer8_outputs(5655) <= not a;
    layer8_outputs(5656) <= a and b;
    layer8_outputs(5657) <= not (a xor b);
    layer8_outputs(5658) <= a xor b;
    layer8_outputs(5659) <= a;
    layer8_outputs(5660) <= a;
    layer8_outputs(5661) <= a;
    layer8_outputs(5662) <= a or b;
    layer8_outputs(5663) <= not (a and b);
    layer8_outputs(5664) <= b;
    layer8_outputs(5665) <= a;
    layer8_outputs(5666) <= not b;
    layer8_outputs(5667) <= a xor b;
    layer8_outputs(5668) <= a xor b;
    layer8_outputs(5669) <= a xor b;
    layer8_outputs(5670) <= b and not a;
    layer8_outputs(5671) <= b;
    layer8_outputs(5672) <= not a or b;
    layer8_outputs(5673) <= a xor b;
    layer8_outputs(5674) <= a and b;
    layer8_outputs(5675) <= not a;
    layer8_outputs(5676) <= not (a xor b);
    layer8_outputs(5677) <= not (a xor b);
    layer8_outputs(5678) <= not b;
    layer8_outputs(5679) <= a xor b;
    layer8_outputs(5680) <= not (a xor b);
    layer8_outputs(5681) <= not a;
    layer8_outputs(5682) <= not (a xor b);
    layer8_outputs(5683) <= not (a xor b);
    layer8_outputs(5684) <= not (a xor b);
    layer8_outputs(5685) <= a and not b;
    layer8_outputs(5686) <= a and not b;
    layer8_outputs(5687) <= b and not a;
    layer8_outputs(5688) <= a and b;
    layer8_outputs(5689) <= not b or a;
    layer8_outputs(5690) <= not (a or b);
    layer8_outputs(5691) <= not b;
    layer8_outputs(5692) <= not a;
    layer8_outputs(5693) <= a xor b;
    layer8_outputs(5694) <= not (a or b);
    layer8_outputs(5695) <= not (a or b);
    layer8_outputs(5696) <= b;
    layer8_outputs(5697) <= b;
    layer8_outputs(5698) <= not b;
    layer8_outputs(5699) <= b;
    layer8_outputs(5700) <= not (a xor b);
    layer8_outputs(5701) <= not (a or b);
    layer8_outputs(5702) <= not (a or b);
    layer8_outputs(5703) <= b;
    layer8_outputs(5704) <= a xor b;
    layer8_outputs(5705) <= not (a and b);
    layer8_outputs(5706) <= b and not a;
    layer8_outputs(5707) <= a xor b;
    layer8_outputs(5708) <= not a;
    layer8_outputs(5709) <= not (a or b);
    layer8_outputs(5710) <= not (a xor b);
    layer8_outputs(5711) <= a or b;
    layer8_outputs(5712) <= not (a xor b);
    layer8_outputs(5713) <= not a;
    layer8_outputs(5714) <= not a;
    layer8_outputs(5715) <= not (a and b);
    layer8_outputs(5716) <= not a;
    layer8_outputs(5717) <= a and not b;
    layer8_outputs(5718) <= not (a and b);
    layer8_outputs(5719) <= b;
    layer8_outputs(5720) <= not a;
    layer8_outputs(5721) <= a and not b;
    layer8_outputs(5722) <= not b or a;
    layer8_outputs(5723) <= a;
    layer8_outputs(5724) <= not a;
    layer8_outputs(5725) <= a xor b;
    layer8_outputs(5726) <= not (a xor b);
    layer8_outputs(5727) <= not b;
    layer8_outputs(5728) <= a and not b;
    layer8_outputs(5729) <= a;
    layer8_outputs(5730) <= not b;
    layer8_outputs(5731) <= a and not b;
    layer8_outputs(5732) <= not a;
    layer8_outputs(5733) <= not b;
    layer8_outputs(5734) <= not a or b;
    layer8_outputs(5735) <= a and b;
    layer8_outputs(5736) <= a xor b;
    layer8_outputs(5737) <= a;
    layer8_outputs(5738) <= not b;
    layer8_outputs(5739) <= a or b;
    layer8_outputs(5740) <= not a;
    layer8_outputs(5741) <= not b or a;
    layer8_outputs(5742) <= a and b;
    layer8_outputs(5743) <= not (a and b);
    layer8_outputs(5744) <= not b;
    layer8_outputs(5745) <= not a;
    layer8_outputs(5746) <= a;
    layer8_outputs(5747) <= not b;
    layer8_outputs(5748) <= not a;
    layer8_outputs(5749) <= b;
    layer8_outputs(5750) <= a;
    layer8_outputs(5751) <= not a or b;
    layer8_outputs(5752) <= b;
    layer8_outputs(5753) <= a;
    layer8_outputs(5754) <= a xor b;
    layer8_outputs(5755) <= not b;
    layer8_outputs(5756) <= a and not b;
    layer8_outputs(5757) <= a and not b;
    layer8_outputs(5758) <= a xor b;
    layer8_outputs(5759) <= b;
    layer8_outputs(5760) <= not a;
    layer8_outputs(5761) <= a;
    layer8_outputs(5762) <= not (a xor b);
    layer8_outputs(5763) <= b;
    layer8_outputs(5764) <= b;
    layer8_outputs(5765) <= not a;
    layer8_outputs(5766) <= not b;
    layer8_outputs(5767) <= a or b;
    layer8_outputs(5768) <= not b;
    layer8_outputs(5769) <= a xor b;
    layer8_outputs(5770) <= not (a xor b);
    layer8_outputs(5771) <= not (a and b);
    layer8_outputs(5772) <= a xor b;
    layer8_outputs(5773) <= not a or b;
    layer8_outputs(5774) <= not (a or b);
    layer8_outputs(5775) <= a xor b;
    layer8_outputs(5776) <= not a or b;
    layer8_outputs(5777) <= not a;
    layer8_outputs(5778) <= a;
    layer8_outputs(5779) <= not a;
    layer8_outputs(5780) <= not (a xor b);
    layer8_outputs(5781) <= b;
    layer8_outputs(5782) <= not a;
    layer8_outputs(5783) <= not (a and b);
    layer8_outputs(5784) <= b;
    layer8_outputs(5785) <= not b;
    layer8_outputs(5786) <= not b;
    layer8_outputs(5787) <= a xor b;
    layer8_outputs(5788) <= a or b;
    layer8_outputs(5789) <= b;
    layer8_outputs(5790) <= not (a or b);
    layer8_outputs(5791) <= not b;
    layer8_outputs(5792) <= a;
    layer8_outputs(5793) <= not (a and b);
    layer8_outputs(5794) <= not (a xor b);
    layer8_outputs(5795) <= a;
    layer8_outputs(5796) <= b;
    layer8_outputs(5797) <= b and not a;
    layer8_outputs(5798) <= a xor b;
    layer8_outputs(5799) <= not b or a;
    layer8_outputs(5800) <= b;
    layer8_outputs(5801) <= not (a xor b);
    layer8_outputs(5802) <= 1'b0;
    layer8_outputs(5803) <= a or b;
    layer8_outputs(5804) <= 1'b1;
    layer8_outputs(5805) <= not (a or b);
    layer8_outputs(5806) <= not (a xor b);
    layer8_outputs(5807) <= a;
    layer8_outputs(5808) <= a;
    layer8_outputs(5809) <= a and not b;
    layer8_outputs(5810) <= a xor b;
    layer8_outputs(5811) <= not (a and b);
    layer8_outputs(5812) <= b;
    layer8_outputs(5813) <= a xor b;
    layer8_outputs(5814) <= not b or a;
    layer8_outputs(5815) <= not b;
    layer8_outputs(5816) <= a and b;
    layer8_outputs(5817) <= not b;
    layer8_outputs(5818) <= a xor b;
    layer8_outputs(5819) <= not (a xor b);
    layer8_outputs(5820) <= a;
    layer8_outputs(5821) <= b;
    layer8_outputs(5822) <= a;
    layer8_outputs(5823) <= a xor b;
    layer8_outputs(5824) <= a or b;
    layer8_outputs(5825) <= b;
    layer8_outputs(5826) <= not (a xor b);
    layer8_outputs(5827) <= 1'b0;
    layer8_outputs(5828) <= not (a or b);
    layer8_outputs(5829) <= not (a xor b);
    layer8_outputs(5830) <= a and not b;
    layer8_outputs(5831) <= b;
    layer8_outputs(5832) <= a or b;
    layer8_outputs(5833) <= not b;
    layer8_outputs(5834) <= not a;
    layer8_outputs(5835) <= b and not a;
    layer8_outputs(5836) <= not b;
    layer8_outputs(5837) <= a and not b;
    layer8_outputs(5838) <= a and not b;
    layer8_outputs(5839) <= a xor b;
    layer8_outputs(5840) <= not a;
    layer8_outputs(5841) <= not (a xor b);
    layer8_outputs(5842) <= 1'b0;
    layer8_outputs(5843) <= not a;
    layer8_outputs(5844) <= not (a xor b);
    layer8_outputs(5845) <= a xor b;
    layer8_outputs(5846) <= not (a xor b);
    layer8_outputs(5847) <= not (a or b);
    layer8_outputs(5848) <= a xor b;
    layer8_outputs(5849) <= a and b;
    layer8_outputs(5850) <= not b;
    layer8_outputs(5851) <= b;
    layer8_outputs(5852) <= b;
    layer8_outputs(5853) <= b;
    layer8_outputs(5854) <= not a;
    layer8_outputs(5855) <= not (a xor b);
    layer8_outputs(5856) <= not b;
    layer8_outputs(5857) <= a and b;
    layer8_outputs(5858) <= b;
    layer8_outputs(5859) <= b and not a;
    layer8_outputs(5860) <= b and not a;
    layer8_outputs(5861) <= b and not a;
    layer8_outputs(5862) <= not (a or b);
    layer8_outputs(5863) <= b;
    layer8_outputs(5864) <= not (a xor b);
    layer8_outputs(5865) <= not b or a;
    layer8_outputs(5866) <= b;
    layer8_outputs(5867) <= a xor b;
    layer8_outputs(5868) <= not b;
    layer8_outputs(5869) <= not (a xor b);
    layer8_outputs(5870) <= 1'b1;
    layer8_outputs(5871) <= not (a xor b);
    layer8_outputs(5872) <= not b;
    layer8_outputs(5873) <= not b or a;
    layer8_outputs(5874) <= a;
    layer8_outputs(5875) <= not b or a;
    layer8_outputs(5876) <= not (a or b);
    layer8_outputs(5877) <= not a;
    layer8_outputs(5878) <= not b or a;
    layer8_outputs(5879) <= not (a xor b);
    layer8_outputs(5880) <= not (a or b);
    layer8_outputs(5881) <= not (a and b);
    layer8_outputs(5882) <= a or b;
    layer8_outputs(5883) <= not (a xor b);
    layer8_outputs(5884) <= a or b;
    layer8_outputs(5885) <= a and b;
    layer8_outputs(5886) <= not (a or b);
    layer8_outputs(5887) <= a;
    layer8_outputs(5888) <= a xor b;
    layer8_outputs(5889) <= not a or b;
    layer8_outputs(5890) <= not b;
    layer8_outputs(5891) <= a xor b;
    layer8_outputs(5892) <= a and b;
    layer8_outputs(5893) <= not (a and b);
    layer8_outputs(5894) <= not (a xor b);
    layer8_outputs(5895) <= a and b;
    layer8_outputs(5896) <= a and not b;
    layer8_outputs(5897) <= 1'b0;
    layer8_outputs(5898) <= b;
    layer8_outputs(5899) <= a;
    layer8_outputs(5900) <= a;
    layer8_outputs(5901) <= not (a xor b);
    layer8_outputs(5902) <= not b;
    layer8_outputs(5903) <= a;
    layer8_outputs(5904) <= not a;
    layer8_outputs(5905) <= not a or b;
    layer8_outputs(5906) <= a or b;
    layer8_outputs(5907) <= b and not a;
    layer8_outputs(5908) <= not b;
    layer8_outputs(5909) <= not a;
    layer8_outputs(5910) <= not b;
    layer8_outputs(5911) <= not a;
    layer8_outputs(5912) <= b;
    layer8_outputs(5913) <= a and not b;
    layer8_outputs(5914) <= b;
    layer8_outputs(5915) <= not (a or b);
    layer8_outputs(5916) <= b;
    layer8_outputs(5917) <= not a;
    layer8_outputs(5918) <= not (a or b);
    layer8_outputs(5919) <= not a;
    layer8_outputs(5920) <= a and b;
    layer8_outputs(5921) <= b and not a;
    layer8_outputs(5922) <= not (a and b);
    layer8_outputs(5923) <= b and not a;
    layer8_outputs(5924) <= not a;
    layer8_outputs(5925) <= b;
    layer8_outputs(5926) <= b and not a;
    layer8_outputs(5927) <= not (a xor b);
    layer8_outputs(5928) <= not (a xor b);
    layer8_outputs(5929) <= not a or b;
    layer8_outputs(5930) <= not b or a;
    layer8_outputs(5931) <= a;
    layer8_outputs(5932) <= not (a or b);
    layer8_outputs(5933) <= b and not a;
    layer8_outputs(5934) <= a;
    layer8_outputs(5935) <= not a;
    layer8_outputs(5936) <= a xor b;
    layer8_outputs(5937) <= a xor b;
    layer8_outputs(5938) <= a or b;
    layer8_outputs(5939) <= not (a xor b);
    layer8_outputs(5940) <= not b;
    layer8_outputs(5941) <= b and not a;
    layer8_outputs(5942) <= a xor b;
    layer8_outputs(5943) <= not a or b;
    layer8_outputs(5944) <= not (a xor b);
    layer8_outputs(5945) <= a;
    layer8_outputs(5946) <= a;
    layer8_outputs(5947) <= not a or b;
    layer8_outputs(5948) <= not a;
    layer8_outputs(5949) <= not a;
    layer8_outputs(5950) <= a or b;
    layer8_outputs(5951) <= a or b;
    layer8_outputs(5952) <= not a;
    layer8_outputs(5953) <= not a;
    layer8_outputs(5954) <= not b;
    layer8_outputs(5955) <= b and not a;
    layer8_outputs(5956) <= a;
    layer8_outputs(5957) <= b;
    layer8_outputs(5958) <= a;
    layer8_outputs(5959) <= b;
    layer8_outputs(5960) <= a;
    layer8_outputs(5961) <= not (a xor b);
    layer8_outputs(5962) <= not b;
    layer8_outputs(5963) <= not a or b;
    layer8_outputs(5964) <= a and not b;
    layer8_outputs(5965) <= a;
    layer8_outputs(5966) <= a;
    layer8_outputs(5967) <= not a;
    layer8_outputs(5968) <= a or b;
    layer8_outputs(5969) <= a xor b;
    layer8_outputs(5970) <= not b;
    layer8_outputs(5971) <= b;
    layer8_outputs(5972) <= not (a or b);
    layer8_outputs(5973) <= not a or b;
    layer8_outputs(5974) <= not a or b;
    layer8_outputs(5975) <= a;
    layer8_outputs(5976) <= not (a or b);
    layer8_outputs(5977) <= not b;
    layer8_outputs(5978) <= a or b;
    layer8_outputs(5979) <= not b;
    layer8_outputs(5980) <= not b;
    layer8_outputs(5981) <= not a;
    layer8_outputs(5982) <= not (a xor b);
    layer8_outputs(5983) <= not a;
    layer8_outputs(5984) <= b;
    layer8_outputs(5985) <= not b;
    layer8_outputs(5986) <= a xor b;
    layer8_outputs(5987) <= not a;
    layer8_outputs(5988) <= not (a and b);
    layer8_outputs(5989) <= not (a xor b);
    layer8_outputs(5990) <= not b;
    layer8_outputs(5991) <= not a;
    layer8_outputs(5992) <= a;
    layer8_outputs(5993) <= not (a xor b);
    layer8_outputs(5994) <= not (a or b);
    layer8_outputs(5995) <= not (a xor b);
    layer8_outputs(5996) <= not a or b;
    layer8_outputs(5997) <= not a;
    layer8_outputs(5998) <= b;
    layer8_outputs(5999) <= a and b;
    layer8_outputs(6000) <= a and not b;
    layer8_outputs(6001) <= a;
    layer8_outputs(6002) <= a xor b;
    layer8_outputs(6003) <= not (a xor b);
    layer8_outputs(6004) <= not (a xor b);
    layer8_outputs(6005) <= a and not b;
    layer8_outputs(6006) <= not (a xor b);
    layer8_outputs(6007) <= not b;
    layer8_outputs(6008) <= a or b;
    layer8_outputs(6009) <= not a;
    layer8_outputs(6010) <= a or b;
    layer8_outputs(6011) <= a xor b;
    layer8_outputs(6012) <= b and not a;
    layer8_outputs(6013) <= b and not a;
    layer8_outputs(6014) <= not (a and b);
    layer8_outputs(6015) <= not b;
    layer8_outputs(6016) <= a and b;
    layer8_outputs(6017) <= b;
    layer8_outputs(6018) <= not b or a;
    layer8_outputs(6019) <= b;
    layer8_outputs(6020) <= not b;
    layer8_outputs(6021) <= not b or a;
    layer8_outputs(6022) <= b and not a;
    layer8_outputs(6023) <= not b;
    layer8_outputs(6024) <= not (a xor b);
    layer8_outputs(6025) <= not a;
    layer8_outputs(6026) <= not b;
    layer8_outputs(6027) <= 1'b1;
    layer8_outputs(6028) <= a or b;
    layer8_outputs(6029) <= a xor b;
    layer8_outputs(6030) <= a xor b;
    layer8_outputs(6031) <= not (a xor b);
    layer8_outputs(6032) <= not a or b;
    layer8_outputs(6033) <= not (a xor b);
    layer8_outputs(6034) <= b;
    layer8_outputs(6035) <= a xor b;
    layer8_outputs(6036) <= not (a or b);
    layer8_outputs(6037) <= not a;
    layer8_outputs(6038) <= b;
    layer8_outputs(6039) <= not a;
    layer8_outputs(6040) <= not a;
    layer8_outputs(6041) <= a;
    layer8_outputs(6042) <= 1'b0;
    layer8_outputs(6043) <= b;
    layer8_outputs(6044) <= a and not b;
    layer8_outputs(6045) <= not (a xor b);
    layer8_outputs(6046) <= b;
    layer8_outputs(6047) <= not (a xor b);
    layer8_outputs(6048) <= not a;
    layer8_outputs(6049) <= not a;
    layer8_outputs(6050) <= a or b;
    layer8_outputs(6051) <= not b or a;
    layer8_outputs(6052) <= not b;
    layer8_outputs(6053) <= a and not b;
    layer8_outputs(6054) <= a;
    layer8_outputs(6055) <= b;
    layer8_outputs(6056) <= 1'b0;
    layer8_outputs(6057) <= not (a xor b);
    layer8_outputs(6058) <= not (a xor b);
    layer8_outputs(6059) <= a and b;
    layer8_outputs(6060) <= a xor b;
    layer8_outputs(6061) <= not a;
    layer8_outputs(6062) <= not a or b;
    layer8_outputs(6063) <= a;
    layer8_outputs(6064) <= a xor b;
    layer8_outputs(6065) <= not b or a;
    layer8_outputs(6066) <= a xor b;
    layer8_outputs(6067) <= a xor b;
    layer8_outputs(6068) <= a;
    layer8_outputs(6069) <= b;
    layer8_outputs(6070) <= not a;
    layer8_outputs(6071) <= b;
    layer8_outputs(6072) <= not b or a;
    layer8_outputs(6073) <= b;
    layer8_outputs(6074) <= a or b;
    layer8_outputs(6075) <= a and not b;
    layer8_outputs(6076) <= a;
    layer8_outputs(6077) <= not (a or b);
    layer8_outputs(6078) <= not a or b;
    layer8_outputs(6079) <= not b;
    layer8_outputs(6080) <= not b;
    layer8_outputs(6081) <= a;
    layer8_outputs(6082) <= b and not a;
    layer8_outputs(6083) <= a xor b;
    layer8_outputs(6084) <= a;
    layer8_outputs(6085) <= b;
    layer8_outputs(6086) <= a and b;
    layer8_outputs(6087) <= not a;
    layer8_outputs(6088) <= a or b;
    layer8_outputs(6089) <= a xor b;
    layer8_outputs(6090) <= not b;
    layer8_outputs(6091) <= not (a xor b);
    layer8_outputs(6092) <= not b;
    layer8_outputs(6093) <= not b;
    layer8_outputs(6094) <= a xor b;
    layer8_outputs(6095) <= a;
    layer8_outputs(6096) <= not a;
    layer8_outputs(6097) <= not (a xor b);
    layer8_outputs(6098) <= b;
    layer8_outputs(6099) <= a;
    layer8_outputs(6100) <= a xor b;
    layer8_outputs(6101) <= a xor b;
    layer8_outputs(6102) <= not a;
    layer8_outputs(6103) <= a or b;
    layer8_outputs(6104) <= a;
    layer8_outputs(6105) <= b;
    layer8_outputs(6106) <= not (a xor b);
    layer8_outputs(6107) <= b;
    layer8_outputs(6108) <= a;
    layer8_outputs(6109) <= a or b;
    layer8_outputs(6110) <= a and b;
    layer8_outputs(6111) <= b;
    layer8_outputs(6112) <= not (a and b);
    layer8_outputs(6113) <= not b;
    layer8_outputs(6114) <= b;
    layer8_outputs(6115) <= not (a and b);
    layer8_outputs(6116) <= a or b;
    layer8_outputs(6117) <= a;
    layer8_outputs(6118) <= not a or b;
    layer8_outputs(6119) <= not a;
    layer8_outputs(6120) <= a xor b;
    layer8_outputs(6121) <= b;
    layer8_outputs(6122) <= not (a xor b);
    layer8_outputs(6123) <= not b;
    layer8_outputs(6124) <= not a;
    layer8_outputs(6125) <= b and not a;
    layer8_outputs(6126) <= not (a xor b);
    layer8_outputs(6127) <= a xor b;
    layer8_outputs(6128) <= b and not a;
    layer8_outputs(6129) <= not (a and b);
    layer8_outputs(6130) <= not a;
    layer8_outputs(6131) <= b;
    layer8_outputs(6132) <= not b;
    layer8_outputs(6133) <= not b;
    layer8_outputs(6134) <= a xor b;
    layer8_outputs(6135) <= not a;
    layer8_outputs(6136) <= not (a xor b);
    layer8_outputs(6137) <= not (a xor b);
    layer8_outputs(6138) <= b;
    layer8_outputs(6139) <= a;
    layer8_outputs(6140) <= not (a or b);
    layer8_outputs(6141) <= b;
    layer8_outputs(6142) <= b;
    layer8_outputs(6143) <= not (a or b);
    layer8_outputs(6144) <= a;
    layer8_outputs(6145) <= not (a or b);
    layer8_outputs(6146) <= not b;
    layer8_outputs(6147) <= a;
    layer8_outputs(6148) <= b;
    layer8_outputs(6149) <= a;
    layer8_outputs(6150) <= b;
    layer8_outputs(6151) <= a;
    layer8_outputs(6152) <= b;
    layer8_outputs(6153) <= a xor b;
    layer8_outputs(6154) <= not b;
    layer8_outputs(6155) <= a and not b;
    layer8_outputs(6156) <= a;
    layer8_outputs(6157) <= not b;
    layer8_outputs(6158) <= b;
    layer8_outputs(6159) <= not a or b;
    layer8_outputs(6160) <= not b or a;
    layer8_outputs(6161) <= b;
    layer8_outputs(6162) <= a and not b;
    layer8_outputs(6163) <= a or b;
    layer8_outputs(6164) <= not (a xor b);
    layer8_outputs(6165) <= a xor b;
    layer8_outputs(6166) <= not (a xor b);
    layer8_outputs(6167) <= not a or b;
    layer8_outputs(6168) <= not a or b;
    layer8_outputs(6169) <= not (a xor b);
    layer8_outputs(6170) <= a xor b;
    layer8_outputs(6171) <= not (a xor b);
    layer8_outputs(6172) <= not (a and b);
    layer8_outputs(6173) <= b and not a;
    layer8_outputs(6174) <= not b or a;
    layer8_outputs(6175) <= a and b;
    layer8_outputs(6176) <= not a or b;
    layer8_outputs(6177) <= a xor b;
    layer8_outputs(6178) <= a xor b;
    layer8_outputs(6179) <= a;
    layer8_outputs(6180) <= a;
    layer8_outputs(6181) <= not (a xor b);
    layer8_outputs(6182) <= not b;
    layer8_outputs(6183) <= a;
    layer8_outputs(6184) <= not (a xor b);
    layer8_outputs(6185) <= a;
    layer8_outputs(6186) <= not (a xor b);
    layer8_outputs(6187) <= a and b;
    layer8_outputs(6188) <= not (a xor b);
    layer8_outputs(6189) <= 1'b1;
    layer8_outputs(6190) <= a;
    layer8_outputs(6191) <= not b or a;
    layer8_outputs(6192) <= b;
    layer8_outputs(6193) <= not a;
    layer8_outputs(6194) <= not (a xor b);
    layer8_outputs(6195) <= not (a or b);
    layer8_outputs(6196) <= not (a or b);
    layer8_outputs(6197) <= not b;
    layer8_outputs(6198) <= a and b;
    layer8_outputs(6199) <= a xor b;
    layer8_outputs(6200) <= a xor b;
    layer8_outputs(6201) <= b and not a;
    layer8_outputs(6202) <= not (a or b);
    layer8_outputs(6203) <= a xor b;
    layer8_outputs(6204) <= b and not a;
    layer8_outputs(6205) <= a xor b;
    layer8_outputs(6206) <= not b;
    layer8_outputs(6207) <= a;
    layer8_outputs(6208) <= not a;
    layer8_outputs(6209) <= not (a xor b);
    layer8_outputs(6210) <= a;
    layer8_outputs(6211) <= b and not a;
    layer8_outputs(6212) <= a xor b;
    layer8_outputs(6213) <= a and not b;
    layer8_outputs(6214) <= not a;
    layer8_outputs(6215) <= not (a xor b);
    layer8_outputs(6216) <= not b;
    layer8_outputs(6217) <= a xor b;
    layer8_outputs(6218) <= not (a xor b);
    layer8_outputs(6219) <= not b;
    layer8_outputs(6220) <= not a or b;
    layer8_outputs(6221) <= not (a xor b);
    layer8_outputs(6222) <= not a;
    layer8_outputs(6223) <= not b;
    layer8_outputs(6224) <= a xor b;
    layer8_outputs(6225) <= a;
    layer8_outputs(6226) <= not b or a;
    layer8_outputs(6227) <= b;
    layer8_outputs(6228) <= not (a xor b);
    layer8_outputs(6229) <= b;
    layer8_outputs(6230) <= not (a xor b);
    layer8_outputs(6231) <= not b;
    layer8_outputs(6232) <= not b or a;
    layer8_outputs(6233) <= not (a or b);
    layer8_outputs(6234) <= not (a xor b);
    layer8_outputs(6235) <= not a or b;
    layer8_outputs(6236) <= not (a xor b);
    layer8_outputs(6237) <= not b;
    layer8_outputs(6238) <= not a;
    layer8_outputs(6239) <= 1'b0;
    layer8_outputs(6240) <= not (a xor b);
    layer8_outputs(6241) <= not (a xor b);
    layer8_outputs(6242) <= not (a xor b);
    layer8_outputs(6243) <= a and not b;
    layer8_outputs(6244) <= a;
    layer8_outputs(6245) <= a and b;
    layer8_outputs(6246) <= not a;
    layer8_outputs(6247) <= not b;
    layer8_outputs(6248) <= not b;
    layer8_outputs(6249) <= not b or a;
    layer8_outputs(6250) <= a and not b;
    layer8_outputs(6251) <= not a;
    layer8_outputs(6252) <= not b or a;
    layer8_outputs(6253) <= not (a xor b);
    layer8_outputs(6254) <= 1'b1;
    layer8_outputs(6255) <= not b;
    layer8_outputs(6256) <= not (a xor b);
    layer8_outputs(6257) <= not a;
    layer8_outputs(6258) <= b;
    layer8_outputs(6259) <= not (a or b);
    layer8_outputs(6260) <= not a;
    layer8_outputs(6261) <= not (a and b);
    layer8_outputs(6262) <= a xor b;
    layer8_outputs(6263) <= a and not b;
    layer8_outputs(6264) <= not a;
    layer8_outputs(6265) <= b;
    layer8_outputs(6266) <= not a;
    layer8_outputs(6267) <= not a;
    layer8_outputs(6268) <= not b;
    layer8_outputs(6269) <= not (a xor b);
    layer8_outputs(6270) <= not b or a;
    layer8_outputs(6271) <= not (a xor b);
    layer8_outputs(6272) <= not (a xor b);
    layer8_outputs(6273) <= not (a xor b);
    layer8_outputs(6274) <= not (a or b);
    layer8_outputs(6275) <= b;
    layer8_outputs(6276) <= not a;
    layer8_outputs(6277) <= a or b;
    layer8_outputs(6278) <= b and not a;
    layer8_outputs(6279) <= not (a or b);
    layer8_outputs(6280) <= not b;
    layer8_outputs(6281) <= b;
    layer8_outputs(6282) <= a and not b;
    layer8_outputs(6283) <= a;
    layer8_outputs(6284) <= not (a xor b);
    layer8_outputs(6285) <= a;
    layer8_outputs(6286) <= not a;
    layer8_outputs(6287) <= not (a and b);
    layer8_outputs(6288) <= a xor b;
    layer8_outputs(6289) <= not (a and b);
    layer8_outputs(6290) <= a or b;
    layer8_outputs(6291) <= not a;
    layer8_outputs(6292) <= a and not b;
    layer8_outputs(6293) <= not a or b;
    layer8_outputs(6294) <= b and not a;
    layer8_outputs(6295) <= a;
    layer8_outputs(6296) <= a and b;
    layer8_outputs(6297) <= not (a xor b);
    layer8_outputs(6298) <= a xor b;
    layer8_outputs(6299) <= b;
    layer8_outputs(6300) <= not a;
    layer8_outputs(6301) <= a xor b;
    layer8_outputs(6302) <= not b;
    layer8_outputs(6303) <= not b;
    layer8_outputs(6304) <= b;
    layer8_outputs(6305) <= not b;
    layer8_outputs(6306) <= not b;
    layer8_outputs(6307) <= not b or a;
    layer8_outputs(6308) <= not b;
    layer8_outputs(6309) <= b and not a;
    layer8_outputs(6310) <= a xor b;
    layer8_outputs(6311) <= not (a xor b);
    layer8_outputs(6312) <= a or b;
    layer8_outputs(6313) <= a xor b;
    layer8_outputs(6314) <= not (a and b);
    layer8_outputs(6315) <= b;
    layer8_outputs(6316) <= not a;
    layer8_outputs(6317) <= a xor b;
    layer8_outputs(6318) <= not (a xor b);
    layer8_outputs(6319) <= b;
    layer8_outputs(6320) <= not a or b;
    layer8_outputs(6321) <= not a;
    layer8_outputs(6322) <= not (a and b);
    layer8_outputs(6323) <= a;
    layer8_outputs(6324) <= a;
    layer8_outputs(6325) <= not b;
    layer8_outputs(6326) <= a;
    layer8_outputs(6327) <= not (a xor b);
    layer8_outputs(6328) <= not a or b;
    layer8_outputs(6329) <= not a;
    layer8_outputs(6330) <= b;
    layer8_outputs(6331) <= a and b;
    layer8_outputs(6332) <= not a;
    layer8_outputs(6333) <= a and b;
    layer8_outputs(6334) <= a xor b;
    layer8_outputs(6335) <= b and not a;
    layer8_outputs(6336) <= not (a xor b);
    layer8_outputs(6337) <= a and not b;
    layer8_outputs(6338) <= not a;
    layer8_outputs(6339) <= not (a and b);
    layer8_outputs(6340) <= a;
    layer8_outputs(6341) <= not (a or b);
    layer8_outputs(6342) <= b and not a;
    layer8_outputs(6343) <= not (a xor b);
    layer8_outputs(6344) <= a xor b;
    layer8_outputs(6345) <= b;
    layer8_outputs(6346) <= a or b;
    layer8_outputs(6347) <= a;
    layer8_outputs(6348) <= not a;
    layer8_outputs(6349) <= 1'b1;
    layer8_outputs(6350) <= a and b;
    layer8_outputs(6351) <= a;
    layer8_outputs(6352) <= a xor b;
    layer8_outputs(6353) <= not a;
    layer8_outputs(6354) <= not b;
    layer8_outputs(6355) <= a and b;
    layer8_outputs(6356) <= a;
    layer8_outputs(6357) <= not (a xor b);
    layer8_outputs(6358) <= not b;
    layer8_outputs(6359) <= a xor b;
    layer8_outputs(6360) <= b and not a;
    layer8_outputs(6361) <= a;
    layer8_outputs(6362) <= b and not a;
    layer8_outputs(6363) <= not b or a;
    layer8_outputs(6364) <= a;
    layer8_outputs(6365) <= not b or a;
    layer8_outputs(6366) <= a xor b;
    layer8_outputs(6367) <= b;
    layer8_outputs(6368) <= b and not a;
    layer8_outputs(6369) <= a xor b;
    layer8_outputs(6370) <= a;
    layer8_outputs(6371) <= a and not b;
    layer8_outputs(6372) <= a and b;
    layer8_outputs(6373) <= not b;
    layer8_outputs(6374) <= a and b;
    layer8_outputs(6375) <= not b;
    layer8_outputs(6376) <= b;
    layer8_outputs(6377) <= not (a and b);
    layer8_outputs(6378) <= a;
    layer8_outputs(6379) <= a xor b;
    layer8_outputs(6380) <= a and not b;
    layer8_outputs(6381) <= not (a xor b);
    layer8_outputs(6382) <= not (a or b);
    layer8_outputs(6383) <= a;
    layer8_outputs(6384) <= not b;
    layer8_outputs(6385) <= a and b;
    layer8_outputs(6386) <= a;
    layer8_outputs(6387) <= not a;
    layer8_outputs(6388) <= not (a and b);
    layer8_outputs(6389) <= a and not b;
    layer8_outputs(6390) <= b;
    layer8_outputs(6391) <= not b;
    layer8_outputs(6392) <= b;
    layer8_outputs(6393) <= a;
    layer8_outputs(6394) <= b;
    layer8_outputs(6395) <= b;
    layer8_outputs(6396) <= a xor b;
    layer8_outputs(6397) <= not a;
    layer8_outputs(6398) <= not a or b;
    layer8_outputs(6399) <= a;
    layer8_outputs(6400) <= not (a xor b);
    layer8_outputs(6401) <= a or b;
    layer8_outputs(6402) <= not a;
    layer8_outputs(6403) <= a or b;
    layer8_outputs(6404) <= a;
    layer8_outputs(6405) <= a xor b;
    layer8_outputs(6406) <= a;
    layer8_outputs(6407) <= a xor b;
    layer8_outputs(6408) <= not a;
    layer8_outputs(6409) <= not a;
    layer8_outputs(6410) <= not a or b;
    layer8_outputs(6411) <= not (a xor b);
    layer8_outputs(6412) <= a xor b;
    layer8_outputs(6413) <= not (a xor b);
    layer8_outputs(6414) <= not b or a;
    layer8_outputs(6415) <= not a;
    layer8_outputs(6416) <= not (a and b);
    layer8_outputs(6417) <= a;
    layer8_outputs(6418) <= not b;
    layer8_outputs(6419) <= not a;
    layer8_outputs(6420) <= a;
    layer8_outputs(6421) <= b;
    layer8_outputs(6422) <= not (a xor b);
    layer8_outputs(6423) <= not (a or b);
    layer8_outputs(6424) <= a or b;
    layer8_outputs(6425) <= not b;
    layer8_outputs(6426) <= not b or a;
    layer8_outputs(6427) <= b;
    layer8_outputs(6428) <= a and not b;
    layer8_outputs(6429) <= a xor b;
    layer8_outputs(6430) <= not a;
    layer8_outputs(6431) <= not (a xor b);
    layer8_outputs(6432) <= b;
    layer8_outputs(6433) <= not b;
    layer8_outputs(6434) <= a xor b;
    layer8_outputs(6435) <= not b;
    layer8_outputs(6436) <= not (a xor b);
    layer8_outputs(6437) <= not a;
    layer8_outputs(6438) <= b;
    layer8_outputs(6439) <= a and not b;
    layer8_outputs(6440) <= a xor b;
    layer8_outputs(6441) <= not a;
    layer8_outputs(6442) <= not (a xor b);
    layer8_outputs(6443) <= a and not b;
    layer8_outputs(6444) <= b;
    layer8_outputs(6445) <= a or b;
    layer8_outputs(6446) <= not a or b;
    layer8_outputs(6447) <= not b;
    layer8_outputs(6448) <= not (a or b);
    layer8_outputs(6449) <= not b;
    layer8_outputs(6450) <= a xor b;
    layer8_outputs(6451) <= a or b;
    layer8_outputs(6452) <= a xor b;
    layer8_outputs(6453) <= not (a xor b);
    layer8_outputs(6454) <= not a;
    layer8_outputs(6455) <= b;
    layer8_outputs(6456) <= b;
    layer8_outputs(6457) <= b;
    layer8_outputs(6458) <= not a;
    layer8_outputs(6459) <= a;
    layer8_outputs(6460) <= not b or a;
    layer8_outputs(6461) <= not a;
    layer8_outputs(6462) <= b;
    layer8_outputs(6463) <= not b;
    layer8_outputs(6464) <= not a or b;
    layer8_outputs(6465) <= not (a or b);
    layer8_outputs(6466) <= not a;
    layer8_outputs(6467) <= b and not a;
    layer8_outputs(6468) <= 1'b0;
    layer8_outputs(6469) <= b;
    layer8_outputs(6470) <= not (a xor b);
    layer8_outputs(6471) <= a;
    layer8_outputs(6472) <= not a;
    layer8_outputs(6473) <= a or b;
    layer8_outputs(6474) <= a xor b;
    layer8_outputs(6475) <= a;
    layer8_outputs(6476) <= a xor b;
    layer8_outputs(6477) <= b;
    layer8_outputs(6478) <= not (a xor b);
    layer8_outputs(6479) <= not (a xor b);
    layer8_outputs(6480) <= a;
    layer8_outputs(6481) <= b;
    layer8_outputs(6482) <= a;
    layer8_outputs(6483) <= not (a xor b);
    layer8_outputs(6484) <= not (a or b);
    layer8_outputs(6485) <= a;
    layer8_outputs(6486) <= b;
    layer8_outputs(6487) <= b;
    layer8_outputs(6488) <= not a or b;
    layer8_outputs(6489) <= not a or b;
    layer8_outputs(6490) <= not a;
    layer8_outputs(6491) <= b;
    layer8_outputs(6492) <= not (a xor b);
    layer8_outputs(6493) <= not (a or b);
    layer8_outputs(6494) <= not b or a;
    layer8_outputs(6495) <= a xor b;
    layer8_outputs(6496) <= not b;
    layer8_outputs(6497) <= a;
    layer8_outputs(6498) <= not b or a;
    layer8_outputs(6499) <= not b;
    layer8_outputs(6500) <= not (a xor b);
    layer8_outputs(6501) <= b;
    layer8_outputs(6502) <= not a or b;
    layer8_outputs(6503) <= a or b;
    layer8_outputs(6504) <= a and b;
    layer8_outputs(6505) <= not b;
    layer8_outputs(6506) <= a and b;
    layer8_outputs(6507) <= not (a xor b);
    layer8_outputs(6508) <= b;
    layer8_outputs(6509) <= not a;
    layer8_outputs(6510) <= not b;
    layer8_outputs(6511) <= a and not b;
    layer8_outputs(6512) <= not (a xor b);
    layer8_outputs(6513) <= a;
    layer8_outputs(6514) <= not b;
    layer8_outputs(6515) <= b;
    layer8_outputs(6516) <= not (a xor b);
    layer8_outputs(6517) <= a and b;
    layer8_outputs(6518) <= not b;
    layer8_outputs(6519) <= not (a xor b);
    layer8_outputs(6520) <= a;
    layer8_outputs(6521) <= not a or b;
    layer8_outputs(6522) <= a;
    layer8_outputs(6523) <= a and b;
    layer8_outputs(6524) <= a and not b;
    layer8_outputs(6525) <= a;
    layer8_outputs(6526) <= a and b;
    layer8_outputs(6527) <= not (a xor b);
    layer8_outputs(6528) <= a xor b;
    layer8_outputs(6529) <= a and not b;
    layer8_outputs(6530) <= b;
    layer8_outputs(6531) <= a xor b;
    layer8_outputs(6532) <= not (a xor b);
    layer8_outputs(6533) <= b;
    layer8_outputs(6534) <= b and not a;
    layer8_outputs(6535) <= a xor b;
    layer8_outputs(6536) <= a;
    layer8_outputs(6537) <= a;
    layer8_outputs(6538) <= not (a xor b);
    layer8_outputs(6539) <= b;
    layer8_outputs(6540) <= a;
    layer8_outputs(6541) <= a xor b;
    layer8_outputs(6542) <= not (a xor b);
    layer8_outputs(6543) <= a xor b;
    layer8_outputs(6544) <= b;
    layer8_outputs(6545) <= b;
    layer8_outputs(6546) <= a;
    layer8_outputs(6547) <= not (a xor b);
    layer8_outputs(6548) <= not a;
    layer8_outputs(6549) <= not (a or b);
    layer8_outputs(6550) <= a xor b;
    layer8_outputs(6551) <= a xor b;
    layer8_outputs(6552) <= a xor b;
    layer8_outputs(6553) <= a;
    layer8_outputs(6554) <= not (a xor b);
    layer8_outputs(6555) <= not a;
    layer8_outputs(6556) <= not b;
    layer8_outputs(6557) <= a and b;
    layer8_outputs(6558) <= not b;
    layer8_outputs(6559) <= a and b;
    layer8_outputs(6560) <= not (a xor b);
    layer8_outputs(6561) <= a or b;
    layer8_outputs(6562) <= not a;
    layer8_outputs(6563) <= not (a or b);
    layer8_outputs(6564) <= not (a and b);
    layer8_outputs(6565) <= not a;
    layer8_outputs(6566) <= a and b;
    layer8_outputs(6567) <= not a or b;
    layer8_outputs(6568) <= not b;
    layer8_outputs(6569) <= a;
    layer8_outputs(6570) <= not a;
    layer8_outputs(6571) <= b;
    layer8_outputs(6572) <= a xor b;
    layer8_outputs(6573) <= not (a xor b);
    layer8_outputs(6574) <= not b or a;
    layer8_outputs(6575) <= b;
    layer8_outputs(6576) <= b;
    layer8_outputs(6577) <= b;
    layer8_outputs(6578) <= not b;
    layer8_outputs(6579) <= not (a xor b);
    layer8_outputs(6580) <= not (a xor b);
    layer8_outputs(6581) <= not (a xor b);
    layer8_outputs(6582) <= not a or b;
    layer8_outputs(6583) <= a and b;
    layer8_outputs(6584) <= a and not b;
    layer8_outputs(6585) <= not a;
    layer8_outputs(6586) <= not a;
    layer8_outputs(6587) <= not (a and b);
    layer8_outputs(6588) <= not (a and b);
    layer8_outputs(6589) <= a xor b;
    layer8_outputs(6590) <= not (a and b);
    layer8_outputs(6591) <= a;
    layer8_outputs(6592) <= a and not b;
    layer8_outputs(6593) <= not (a xor b);
    layer8_outputs(6594) <= b and not a;
    layer8_outputs(6595) <= a xor b;
    layer8_outputs(6596) <= b;
    layer8_outputs(6597) <= a xor b;
    layer8_outputs(6598) <= not (a xor b);
    layer8_outputs(6599) <= not (a and b);
    layer8_outputs(6600) <= b and not a;
    layer8_outputs(6601) <= not (a or b);
    layer8_outputs(6602) <= not a;
    layer8_outputs(6603) <= a and not b;
    layer8_outputs(6604) <= a xor b;
    layer8_outputs(6605) <= a xor b;
    layer8_outputs(6606) <= not a;
    layer8_outputs(6607) <= a or b;
    layer8_outputs(6608) <= not b;
    layer8_outputs(6609) <= a;
    layer8_outputs(6610) <= not (a and b);
    layer8_outputs(6611) <= b;
    layer8_outputs(6612) <= a;
    layer8_outputs(6613) <= not b;
    layer8_outputs(6614) <= not a or b;
    layer8_outputs(6615) <= b;
    layer8_outputs(6616) <= a;
    layer8_outputs(6617) <= not (a xor b);
    layer8_outputs(6618) <= not (a xor b);
    layer8_outputs(6619) <= not (a xor b);
    layer8_outputs(6620) <= not a;
    layer8_outputs(6621) <= b and not a;
    layer8_outputs(6622) <= a or b;
    layer8_outputs(6623) <= not (a xor b);
    layer8_outputs(6624) <= not b;
    layer8_outputs(6625) <= a;
    layer8_outputs(6626) <= b;
    layer8_outputs(6627) <= a;
    layer8_outputs(6628) <= not (a and b);
    layer8_outputs(6629) <= not b or a;
    layer8_outputs(6630) <= a xor b;
    layer8_outputs(6631) <= a or b;
    layer8_outputs(6632) <= not a;
    layer8_outputs(6633) <= not (a or b);
    layer8_outputs(6634) <= b and not a;
    layer8_outputs(6635) <= a xor b;
    layer8_outputs(6636) <= not (a xor b);
    layer8_outputs(6637) <= not b;
    layer8_outputs(6638) <= b;
    layer8_outputs(6639) <= not a;
    layer8_outputs(6640) <= a;
    layer8_outputs(6641) <= a;
    layer8_outputs(6642) <= a;
    layer8_outputs(6643) <= a and b;
    layer8_outputs(6644) <= not (a or b);
    layer8_outputs(6645) <= not b;
    layer8_outputs(6646) <= b and not a;
    layer8_outputs(6647) <= b and not a;
    layer8_outputs(6648) <= a and not b;
    layer8_outputs(6649) <= a and not b;
    layer8_outputs(6650) <= a xor b;
    layer8_outputs(6651) <= a or b;
    layer8_outputs(6652) <= a and b;
    layer8_outputs(6653) <= not (a or b);
    layer8_outputs(6654) <= not (a xor b);
    layer8_outputs(6655) <= a xor b;
    layer8_outputs(6656) <= a or b;
    layer8_outputs(6657) <= not b or a;
    layer8_outputs(6658) <= not a;
    layer8_outputs(6659) <= not (a and b);
    layer8_outputs(6660) <= a;
    layer8_outputs(6661) <= a xor b;
    layer8_outputs(6662) <= a xor b;
    layer8_outputs(6663) <= not b or a;
    layer8_outputs(6664) <= not (a or b);
    layer8_outputs(6665) <= a xor b;
    layer8_outputs(6666) <= not a or b;
    layer8_outputs(6667) <= not (a and b);
    layer8_outputs(6668) <= b and not a;
    layer8_outputs(6669) <= a;
    layer8_outputs(6670) <= a xor b;
    layer8_outputs(6671) <= b;
    layer8_outputs(6672) <= a or b;
    layer8_outputs(6673) <= not (a xor b);
    layer8_outputs(6674) <= a;
    layer8_outputs(6675) <= a xor b;
    layer8_outputs(6676) <= not (a or b);
    layer8_outputs(6677) <= not b or a;
    layer8_outputs(6678) <= b and not a;
    layer8_outputs(6679) <= not (a xor b);
    layer8_outputs(6680) <= not b or a;
    layer8_outputs(6681) <= b;
    layer8_outputs(6682) <= not b;
    layer8_outputs(6683) <= not b or a;
    layer8_outputs(6684) <= not (a xor b);
    layer8_outputs(6685) <= not a;
    layer8_outputs(6686) <= not a;
    layer8_outputs(6687) <= 1'b1;
    layer8_outputs(6688) <= not (a or b);
    layer8_outputs(6689) <= not (a or b);
    layer8_outputs(6690) <= b and not a;
    layer8_outputs(6691) <= a;
    layer8_outputs(6692) <= not (a or b);
    layer8_outputs(6693) <= not (a and b);
    layer8_outputs(6694) <= b and not a;
    layer8_outputs(6695) <= a xor b;
    layer8_outputs(6696) <= not a or b;
    layer8_outputs(6697) <= not b;
    layer8_outputs(6698) <= not a;
    layer8_outputs(6699) <= not (a xor b);
    layer8_outputs(6700) <= not a;
    layer8_outputs(6701) <= a and b;
    layer8_outputs(6702) <= not (a xor b);
    layer8_outputs(6703) <= not b;
    layer8_outputs(6704) <= not a or b;
    layer8_outputs(6705) <= a or b;
    layer8_outputs(6706) <= a and not b;
    layer8_outputs(6707) <= a;
    layer8_outputs(6708) <= not b;
    layer8_outputs(6709) <= b and not a;
    layer8_outputs(6710) <= a;
    layer8_outputs(6711) <= a or b;
    layer8_outputs(6712) <= not b;
    layer8_outputs(6713) <= not (a xor b);
    layer8_outputs(6714) <= not (a and b);
    layer8_outputs(6715) <= a and b;
    layer8_outputs(6716) <= a and b;
    layer8_outputs(6717) <= a and not b;
    layer8_outputs(6718) <= not (a and b);
    layer8_outputs(6719) <= not a or b;
    layer8_outputs(6720) <= not (a and b);
    layer8_outputs(6721) <= a xor b;
    layer8_outputs(6722) <= not (a xor b);
    layer8_outputs(6723) <= not (a and b);
    layer8_outputs(6724) <= not a;
    layer8_outputs(6725) <= not (a or b);
    layer8_outputs(6726) <= not a or b;
    layer8_outputs(6727) <= not a;
    layer8_outputs(6728) <= a and not b;
    layer8_outputs(6729) <= not b;
    layer8_outputs(6730) <= a;
    layer8_outputs(6731) <= not (a xor b);
    layer8_outputs(6732) <= not (a xor b);
    layer8_outputs(6733) <= not (a xor b);
    layer8_outputs(6734) <= b;
    layer8_outputs(6735) <= b;
    layer8_outputs(6736) <= not b;
    layer8_outputs(6737) <= not a;
    layer8_outputs(6738) <= not a;
    layer8_outputs(6739) <= not a;
    layer8_outputs(6740) <= not (a or b);
    layer8_outputs(6741) <= not b or a;
    layer8_outputs(6742) <= b;
    layer8_outputs(6743) <= not (a and b);
    layer8_outputs(6744) <= b;
    layer8_outputs(6745) <= not (a xor b);
    layer8_outputs(6746) <= not a;
    layer8_outputs(6747) <= not b or a;
    layer8_outputs(6748) <= not (a xor b);
    layer8_outputs(6749) <= not b or a;
    layer8_outputs(6750) <= a;
    layer8_outputs(6751) <= not b;
    layer8_outputs(6752) <= a;
    layer8_outputs(6753) <= a xor b;
    layer8_outputs(6754) <= not a;
    layer8_outputs(6755) <= not b or a;
    layer8_outputs(6756) <= not a;
    layer8_outputs(6757) <= not a or b;
    layer8_outputs(6758) <= a and not b;
    layer8_outputs(6759) <= not a or b;
    layer8_outputs(6760) <= b and not a;
    layer8_outputs(6761) <= not (a or b);
    layer8_outputs(6762) <= not b;
    layer8_outputs(6763) <= b;
    layer8_outputs(6764) <= not b;
    layer8_outputs(6765) <= not b;
    layer8_outputs(6766) <= a and not b;
    layer8_outputs(6767) <= not a;
    layer8_outputs(6768) <= b;
    layer8_outputs(6769) <= not a or b;
    layer8_outputs(6770) <= a and b;
    layer8_outputs(6771) <= b;
    layer8_outputs(6772) <= a or b;
    layer8_outputs(6773) <= not a or b;
    layer8_outputs(6774) <= not a;
    layer8_outputs(6775) <= not b;
    layer8_outputs(6776) <= b;
    layer8_outputs(6777) <= a;
    layer8_outputs(6778) <= a and b;
    layer8_outputs(6779) <= not b or a;
    layer8_outputs(6780) <= a;
    layer8_outputs(6781) <= a or b;
    layer8_outputs(6782) <= a;
    layer8_outputs(6783) <= not a;
    layer8_outputs(6784) <= not b;
    layer8_outputs(6785) <= not a;
    layer8_outputs(6786) <= not b;
    layer8_outputs(6787) <= not b;
    layer8_outputs(6788) <= a and b;
    layer8_outputs(6789) <= b and not a;
    layer8_outputs(6790) <= a xor b;
    layer8_outputs(6791) <= not a or b;
    layer8_outputs(6792) <= a xor b;
    layer8_outputs(6793) <= a;
    layer8_outputs(6794) <= not (a or b);
    layer8_outputs(6795) <= a xor b;
    layer8_outputs(6796) <= a and b;
    layer8_outputs(6797) <= a xor b;
    layer8_outputs(6798) <= not a;
    layer8_outputs(6799) <= a xor b;
    layer8_outputs(6800) <= a and not b;
    layer8_outputs(6801) <= b and not a;
    layer8_outputs(6802) <= b and not a;
    layer8_outputs(6803) <= a and b;
    layer8_outputs(6804) <= a;
    layer8_outputs(6805) <= a;
    layer8_outputs(6806) <= a and b;
    layer8_outputs(6807) <= a;
    layer8_outputs(6808) <= b;
    layer8_outputs(6809) <= a xor b;
    layer8_outputs(6810) <= not a;
    layer8_outputs(6811) <= a xor b;
    layer8_outputs(6812) <= not (a and b);
    layer8_outputs(6813) <= not (a or b);
    layer8_outputs(6814) <= not a;
    layer8_outputs(6815) <= b;
    layer8_outputs(6816) <= a;
    layer8_outputs(6817) <= a or b;
    layer8_outputs(6818) <= b;
    layer8_outputs(6819) <= not a;
    layer8_outputs(6820) <= not b or a;
    layer8_outputs(6821) <= not b;
    layer8_outputs(6822) <= not b;
    layer8_outputs(6823) <= not b;
    layer8_outputs(6824) <= not b or a;
    layer8_outputs(6825) <= a;
    layer8_outputs(6826) <= not (a xor b);
    layer8_outputs(6827) <= a;
    layer8_outputs(6828) <= not (a and b);
    layer8_outputs(6829) <= b;
    layer8_outputs(6830) <= a;
    layer8_outputs(6831) <= b;
    layer8_outputs(6832) <= b;
    layer8_outputs(6833) <= a xor b;
    layer8_outputs(6834) <= a xor b;
    layer8_outputs(6835) <= a and b;
    layer8_outputs(6836) <= a or b;
    layer8_outputs(6837) <= b;
    layer8_outputs(6838) <= not (a xor b);
    layer8_outputs(6839) <= not (a xor b);
    layer8_outputs(6840) <= a;
    layer8_outputs(6841) <= a xor b;
    layer8_outputs(6842) <= a or b;
    layer8_outputs(6843) <= a xor b;
    layer8_outputs(6844) <= a xor b;
    layer8_outputs(6845) <= not (a xor b);
    layer8_outputs(6846) <= not b;
    layer8_outputs(6847) <= not a;
    layer8_outputs(6848) <= not (a xor b);
    layer8_outputs(6849) <= not a;
    layer8_outputs(6850) <= not b or a;
    layer8_outputs(6851) <= b;
    layer8_outputs(6852) <= a;
    layer8_outputs(6853) <= a;
    layer8_outputs(6854) <= not b;
    layer8_outputs(6855) <= b and not a;
    layer8_outputs(6856) <= b;
    layer8_outputs(6857) <= not (a and b);
    layer8_outputs(6858) <= not a;
    layer8_outputs(6859) <= not (a or b);
    layer8_outputs(6860) <= a and b;
    layer8_outputs(6861) <= a xor b;
    layer8_outputs(6862) <= a and b;
    layer8_outputs(6863) <= a xor b;
    layer8_outputs(6864) <= a xor b;
    layer8_outputs(6865) <= not a or b;
    layer8_outputs(6866) <= a and b;
    layer8_outputs(6867) <= b;
    layer8_outputs(6868) <= a and not b;
    layer8_outputs(6869) <= b;
    layer8_outputs(6870) <= not (a xor b);
    layer8_outputs(6871) <= a;
    layer8_outputs(6872) <= not (a xor b);
    layer8_outputs(6873) <= a or b;
    layer8_outputs(6874) <= b;
    layer8_outputs(6875) <= not b;
    layer8_outputs(6876) <= b and not a;
    layer8_outputs(6877) <= not (a and b);
    layer8_outputs(6878) <= b;
    layer8_outputs(6879) <= not a;
    layer8_outputs(6880) <= a xor b;
    layer8_outputs(6881) <= not b or a;
    layer8_outputs(6882) <= not (a or b);
    layer8_outputs(6883) <= not a or b;
    layer8_outputs(6884) <= a xor b;
    layer8_outputs(6885) <= not (a xor b);
    layer8_outputs(6886) <= not b;
    layer8_outputs(6887) <= a and not b;
    layer8_outputs(6888) <= 1'b1;
    layer8_outputs(6889) <= b;
    layer8_outputs(6890) <= b and not a;
    layer8_outputs(6891) <= not a;
    layer8_outputs(6892) <= not b;
    layer8_outputs(6893) <= b;
    layer8_outputs(6894) <= not (a xor b);
    layer8_outputs(6895) <= not a;
    layer8_outputs(6896) <= not (a xor b);
    layer8_outputs(6897) <= b;
    layer8_outputs(6898) <= a and not b;
    layer8_outputs(6899) <= not b;
    layer8_outputs(6900) <= not (a and b);
    layer8_outputs(6901) <= a xor b;
    layer8_outputs(6902) <= a;
    layer8_outputs(6903) <= a;
    layer8_outputs(6904) <= 1'b0;
    layer8_outputs(6905) <= a or b;
    layer8_outputs(6906) <= not a;
    layer8_outputs(6907) <= not b;
    layer8_outputs(6908) <= b and not a;
    layer8_outputs(6909) <= b;
    layer8_outputs(6910) <= not (a xor b);
    layer8_outputs(6911) <= a xor b;
    layer8_outputs(6912) <= not a;
    layer8_outputs(6913) <= not (a xor b);
    layer8_outputs(6914) <= not (a xor b);
    layer8_outputs(6915) <= b;
    layer8_outputs(6916) <= a;
    layer8_outputs(6917) <= not b;
    layer8_outputs(6918) <= not a;
    layer8_outputs(6919) <= a;
    layer8_outputs(6920) <= a or b;
    layer8_outputs(6921) <= a xor b;
    layer8_outputs(6922) <= a xor b;
    layer8_outputs(6923) <= not a;
    layer8_outputs(6924) <= a xor b;
    layer8_outputs(6925) <= a xor b;
    layer8_outputs(6926) <= not (a xor b);
    layer8_outputs(6927) <= not (a xor b);
    layer8_outputs(6928) <= not b;
    layer8_outputs(6929) <= not a;
    layer8_outputs(6930) <= not (a xor b);
    layer8_outputs(6931) <= not (a xor b);
    layer8_outputs(6932) <= not (a xor b);
    layer8_outputs(6933) <= b and not a;
    layer8_outputs(6934) <= not a;
    layer8_outputs(6935) <= not (a xor b);
    layer8_outputs(6936) <= not b;
    layer8_outputs(6937) <= not (a xor b);
    layer8_outputs(6938) <= not (a and b);
    layer8_outputs(6939) <= a xor b;
    layer8_outputs(6940) <= a;
    layer8_outputs(6941) <= b;
    layer8_outputs(6942) <= not b or a;
    layer8_outputs(6943) <= not (a xor b);
    layer8_outputs(6944) <= a;
    layer8_outputs(6945) <= not b;
    layer8_outputs(6946) <= a or b;
    layer8_outputs(6947) <= not b;
    layer8_outputs(6948) <= not a;
    layer8_outputs(6949) <= not (a and b);
    layer8_outputs(6950) <= a xor b;
    layer8_outputs(6951) <= not (a xor b);
    layer8_outputs(6952) <= not (a or b);
    layer8_outputs(6953) <= not (a and b);
    layer8_outputs(6954) <= not (a or b);
    layer8_outputs(6955) <= b;
    layer8_outputs(6956) <= not b or a;
    layer8_outputs(6957) <= not a;
    layer8_outputs(6958) <= a and b;
    layer8_outputs(6959) <= a xor b;
    layer8_outputs(6960) <= not (a xor b);
    layer8_outputs(6961) <= not (a xor b);
    layer8_outputs(6962) <= not (a xor b);
    layer8_outputs(6963) <= not (a xor b);
    layer8_outputs(6964) <= not b;
    layer8_outputs(6965) <= not (a xor b);
    layer8_outputs(6966) <= a;
    layer8_outputs(6967) <= not a;
    layer8_outputs(6968) <= not a;
    layer8_outputs(6969) <= a or b;
    layer8_outputs(6970) <= not b;
    layer8_outputs(6971) <= not (a xor b);
    layer8_outputs(6972) <= b;
    layer8_outputs(6973) <= not a;
    layer8_outputs(6974) <= a and not b;
    layer8_outputs(6975) <= b;
    layer8_outputs(6976) <= a xor b;
    layer8_outputs(6977) <= a;
    layer8_outputs(6978) <= a;
    layer8_outputs(6979) <= not a or b;
    layer8_outputs(6980) <= not b;
    layer8_outputs(6981) <= a xor b;
    layer8_outputs(6982) <= not b;
    layer8_outputs(6983) <= b;
    layer8_outputs(6984) <= not b;
    layer8_outputs(6985) <= not a or b;
    layer8_outputs(6986) <= 1'b0;
    layer8_outputs(6987) <= not a;
    layer8_outputs(6988) <= b and not a;
    layer8_outputs(6989) <= not a;
    layer8_outputs(6990) <= b;
    layer8_outputs(6991) <= not a;
    layer8_outputs(6992) <= b;
    layer8_outputs(6993) <= b;
    layer8_outputs(6994) <= a xor b;
    layer8_outputs(6995) <= a;
    layer8_outputs(6996) <= not (a and b);
    layer8_outputs(6997) <= a;
    layer8_outputs(6998) <= not a;
    layer8_outputs(6999) <= a and not b;
    layer8_outputs(7000) <= not a or b;
    layer8_outputs(7001) <= b and not a;
    layer8_outputs(7002) <= a and not b;
    layer8_outputs(7003) <= not b or a;
    layer8_outputs(7004) <= a and not b;
    layer8_outputs(7005) <= 1'b0;
    layer8_outputs(7006) <= not (a and b);
    layer8_outputs(7007) <= not (a and b);
    layer8_outputs(7008) <= not a;
    layer8_outputs(7009) <= not a or b;
    layer8_outputs(7010) <= a;
    layer8_outputs(7011) <= not b;
    layer8_outputs(7012) <= a;
    layer8_outputs(7013) <= a xor b;
    layer8_outputs(7014) <= a;
    layer8_outputs(7015) <= b;
    layer8_outputs(7016) <= not (a xor b);
    layer8_outputs(7017) <= b;
    layer8_outputs(7018) <= not (a xor b);
    layer8_outputs(7019) <= b;
    layer8_outputs(7020) <= a xor b;
    layer8_outputs(7021) <= a xor b;
    layer8_outputs(7022) <= not a;
    layer8_outputs(7023) <= not a;
    layer8_outputs(7024) <= a;
    layer8_outputs(7025) <= not (a and b);
    layer8_outputs(7026) <= not b;
    layer8_outputs(7027) <= b and not a;
    layer8_outputs(7028) <= not b or a;
    layer8_outputs(7029) <= a;
    layer8_outputs(7030) <= a xor b;
    layer8_outputs(7031) <= a;
    layer8_outputs(7032) <= b;
    layer8_outputs(7033) <= a;
    layer8_outputs(7034) <= not (a and b);
    layer8_outputs(7035) <= not (a and b);
    layer8_outputs(7036) <= a and not b;
    layer8_outputs(7037) <= a xor b;
    layer8_outputs(7038) <= a;
    layer8_outputs(7039) <= not (a xor b);
    layer8_outputs(7040) <= 1'b0;
    layer8_outputs(7041) <= not b;
    layer8_outputs(7042) <= a and b;
    layer8_outputs(7043) <= not b;
    layer8_outputs(7044) <= a and b;
    layer8_outputs(7045) <= b;
    layer8_outputs(7046) <= a or b;
    layer8_outputs(7047) <= a;
    layer8_outputs(7048) <= not a;
    layer8_outputs(7049) <= not (a or b);
    layer8_outputs(7050) <= not a;
    layer8_outputs(7051) <= b and not a;
    layer8_outputs(7052) <= a and not b;
    layer8_outputs(7053) <= a;
    layer8_outputs(7054) <= a and b;
    layer8_outputs(7055) <= a and b;
    layer8_outputs(7056) <= not (a xor b);
    layer8_outputs(7057) <= a and not b;
    layer8_outputs(7058) <= not b or a;
    layer8_outputs(7059) <= a;
    layer8_outputs(7060) <= a;
    layer8_outputs(7061) <= a and not b;
    layer8_outputs(7062) <= a;
    layer8_outputs(7063) <= b and not a;
    layer8_outputs(7064) <= b;
    layer8_outputs(7065) <= a xor b;
    layer8_outputs(7066) <= a xor b;
    layer8_outputs(7067) <= not (a xor b);
    layer8_outputs(7068) <= a;
    layer8_outputs(7069) <= a xor b;
    layer8_outputs(7070) <= a xor b;
    layer8_outputs(7071) <= a and b;
    layer8_outputs(7072) <= not (a and b);
    layer8_outputs(7073) <= not a;
    layer8_outputs(7074) <= not b;
    layer8_outputs(7075) <= a or b;
    layer8_outputs(7076) <= not a;
    layer8_outputs(7077) <= not (a xor b);
    layer8_outputs(7078) <= not b;
    layer8_outputs(7079) <= b and not a;
    layer8_outputs(7080) <= 1'b1;
    layer8_outputs(7081) <= not (a xor b);
    layer8_outputs(7082) <= a or b;
    layer8_outputs(7083) <= not a;
    layer8_outputs(7084) <= a xor b;
    layer8_outputs(7085) <= 1'b0;
    layer8_outputs(7086) <= not (a xor b);
    layer8_outputs(7087) <= not a;
    layer8_outputs(7088) <= not (a and b);
    layer8_outputs(7089) <= not a;
    layer8_outputs(7090) <= b;
    layer8_outputs(7091) <= a xor b;
    layer8_outputs(7092) <= b and not a;
    layer8_outputs(7093) <= not b;
    layer8_outputs(7094) <= not a or b;
    layer8_outputs(7095) <= not b;
    layer8_outputs(7096) <= a and b;
    layer8_outputs(7097) <= b;
    layer8_outputs(7098) <= a and b;
    layer8_outputs(7099) <= a;
    layer8_outputs(7100) <= not a;
    layer8_outputs(7101) <= a xor b;
    layer8_outputs(7102) <= not b or a;
    layer8_outputs(7103) <= a and b;
    layer8_outputs(7104) <= not b;
    layer8_outputs(7105) <= not a;
    layer8_outputs(7106) <= not (a xor b);
    layer8_outputs(7107) <= not a;
    layer8_outputs(7108) <= a or b;
    layer8_outputs(7109) <= a or b;
    layer8_outputs(7110) <= 1'b0;
    layer8_outputs(7111) <= not (a or b);
    layer8_outputs(7112) <= a;
    layer8_outputs(7113) <= not b or a;
    layer8_outputs(7114) <= a;
    layer8_outputs(7115) <= not a or b;
    layer8_outputs(7116) <= a and not b;
    layer8_outputs(7117) <= a;
    layer8_outputs(7118) <= not a;
    layer8_outputs(7119) <= not b;
    layer8_outputs(7120) <= a;
    layer8_outputs(7121) <= not b;
    layer8_outputs(7122) <= a xor b;
    layer8_outputs(7123) <= not a;
    layer8_outputs(7124) <= not b;
    layer8_outputs(7125) <= b and not a;
    layer8_outputs(7126) <= a;
    layer8_outputs(7127) <= b;
    layer8_outputs(7128) <= not a;
    layer8_outputs(7129) <= not (a xor b);
    layer8_outputs(7130) <= b;
    layer8_outputs(7131) <= a xor b;
    layer8_outputs(7132) <= b;
    layer8_outputs(7133) <= not b;
    layer8_outputs(7134) <= not (a or b);
    layer8_outputs(7135) <= 1'b0;
    layer8_outputs(7136) <= not (a or b);
    layer8_outputs(7137) <= a xor b;
    layer8_outputs(7138) <= b;
    layer8_outputs(7139) <= not b;
    layer8_outputs(7140) <= a;
    layer8_outputs(7141) <= a;
    layer8_outputs(7142) <= a and not b;
    layer8_outputs(7143) <= not (a xor b);
    layer8_outputs(7144) <= b;
    layer8_outputs(7145) <= not (a xor b);
    layer8_outputs(7146) <= a;
    layer8_outputs(7147) <= a and b;
    layer8_outputs(7148) <= not b;
    layer8_outputs(7149) <= b and not a;
    layer8_outputs(7150) <= a xor b;
    layer8_outputs(7151) <= not a;
    layer8_outputs(7152) <= not (a xor b);
    layer8_outputs(7153) <= not (a xor b);
    layer8_outputs(7154) <= a and not b;
    layer8_outputs(7155) <= a and not b;
    layer8_outputs(7156) <= not a;
    layer8_outputs(7157) <= not a;
    layer8_outputs(7158) <= b and not a;
    layer8_outputs(7159) <= b;
    layer8_outputs(7160) <= not (a xor b);
    layer8_outputs(7161) <= not a;
    layer8_outputs(7162) <= not a;
    layer8_outputs(7163) <= not a or b;
    layer8_outputs(7164) <= a;
    layer8_outputs(7165) <= a xor b;
    layer8_outputs(7166) <= a xor b;
    layer8_outputs(7167) <= not b;
    layer8_outputs(7168) <= b;
    layer8_outputs(7169) <= not a;
    layer8_outputs(7170) <= not a;
    layer8_outputs(7171) <= a;
    layer8_outputs(7172) <= not b or a;
    layer8_outputs(7173) <= b and not a;
    layer8_outputs(7174) <= a and b;
    layer8_outputs(7175) <= a and not b;
    layer8_outputs(7176) <= not a;
    layer8_outputs(7177) <= a or b;
    layer8_outputs(7178) <= not (a xor b);
    layer8_outputs(7179) <= b;
    layer8_outputs(7180) <= a xor b;
    layer8_outputs(7181) <= not a or b;
    layer8_outputs(7182) <= not b;
    layer8_outputs(7183) <= b and not a;
    layer8_outputs(7184) <= a and not b;
    layer8_outputs(7185) <= a;
    layer8_outputs(7186) <= not a or b;
    layer8_outputs(7187) <= not b;
    layer8_outputs(7188) <= not b;
    layer8_outputs(7189) <= b;
    layer8_outputs(7190) <= not (a xor b);
    layer8_outputs(7191) <= b;
    layer8_outputs(7192) <= a xor b;
    layer8_outputs(7193) <= a and b;
    layer8_outputs(7194) <= not (a xor b);
    layer8_outputs(7195) <= not (a xor b);
    layer8_outputs(7196) <= b;
    layer8_outputs(7197) <= a xor b;
    layer8_outputs(7198) <= not b;
    layer8_outputs(7199) <= b;
    layer8_outputs(7200) <= not a;
    layer8_outputs(7201) <= a;
    layer8_outputs(7202) <= a xor b;
    layer8_outputs(7203) <= a;
    layer8_outputs(7204) <= a xor b;
    layer8_outputs(7205) <= b;
    layer8_outputs(7206) <= a;
    layer8_outputs(7207) <= a xor b;
    layer8_outputs(7208) <= a xor b;
    layer8_outputs(7209) <= not (a or b);
    layer8_outputs(7210) <= not b;
    layer8_outputs(7211) <= a xor b;
    layer8_outputs(7212) <= not b or a;
    layer8_outputs(7213) <= a xor b;
    layer8_outputs(7214) <= not (a xor b);
    layer8_outputs(7215) <= a xor b;
    layer8_outputs(7216) <= b;
    layer8_outputs(7217) <= b;
    layer8_outputs(7218) <= not a or b;
    layer8_outputs(7219) <= not (a or b);
    layer8_outputs(7220) <= not a;
    layer8_outputs(7221) <= b and not a;
    layer8_outputs(7222) <= a and b;
    layer8_outputs(7223) <= a;
    layer8_outputs(7224) <= not (a xor b);
    layer8_outputs(7225) <= a xor b;
    layer8_outputs(7226) <= not b;
    layer8_outputs(7227) <= a;
    layer8_outputs(7228) <= not (a xor b);
    layer8_outputs(7229) <= not a;
    layer8_outputs(7230) <= not (a xor b);
    layer8_outputs(7231) <= a or b;
    layer8_outputs(7232) <= not (a and b);
    layer8_outputs(7233) <= not (a and b);
    layer8_outputs(7234) <= not b or a;
    layer8_outputs(7235) <= a xor b;
    layer8_outputs(7236) <= not (a or b);
    layer8_outputs(7237) <= a or b;
    layer8_outputs(7238) <= not (a xor b);
    layer8_outputs(7239) <= a;
    layer8_outputs(7240) <= a and b;
    layer8_outputs(7241) <= b;
    layer8_outputs(7242) <= b;
    layer8_outputs(7243) <= not a;
    layer8_outputs(7244) <= not a;
    layer8_outputs(7245) <= a and b;
    layer8_outputs(7246) <= not a or b;
    layer8_outputs(7247) <= a xor b;
    layer8_outputs(7248) <= a or b;
    layer8_outputs(7249) <= not b;
    layer8_outputs(7250) <= a;
    layer8_outputs(7251) <= not b;
    layer8_outputs(7252) <= b;
    layer8_outputs(7253) <= a or b;
    layer8_outputs(7254) <= not a;
    layer8_outputs(7255) <= a or b;
    layer8_outputs(7256) <= a;
    layer8_outputs(7257) <= b and not a;
    layer8_outputs(7258) <= not (a and b);
    layer8_outputs(7259) <= not (a and b);
    layer8_outputs(7260) <= not (a xor b);
    layer8_outputs(7261) <= a or b;
    layer8_outputs(7262) <= b;
    layer8_outputs(7263) <= not b;
    layer8_outputs(7264) <= b and not a;
    layer8_outputs(7265) <= a and not b;
    layer8_outputs(7266) <= not (a xor b);
    layer8_outputs(7267) <= a xor b;
    layer8_outputs(7268) <= not b;
    layer8_outputs(7269) <= a;
    layer8_outputs(7270) <= a and b;
    layer8_outputs(7271) <= not (a xor b);
    layer8_outputs(7272) <= b;
    layer8_outputs(7273) <= not a;
    layer8_outputs(7274) <= a xor b;
    layer8_outputs(7275) <= b;
    layer8_outputs(7276) <= not b;
    layer8_outputs(7277) <= not b;
    layer8_outputs(7278) <= not (a xor b);
    layer8_outputs(7279) <= b;
    layer8_outputs(7280) <= a or b;
    layer8_outputs(7281) <= a and b;
    layer8_outputs(7282) <= a;
    layer8_outputs(7283) <= b;
    layer8_outputs(7284) <= not a or b;
    layer8_outputs(7285) <= not a or b;
    layer8_outputs(7286) <= a xor b;
    layer8_outputs(7287) <= not a;
    layer8_outputs(7288) <= a and b;
    layer8_outputs(7289) <= not b;
    layer8_outputs(7290) <= not b;
    layer8_outputs(7291) <= a xor b;
    layer8_outputs(7292) <= not (a xor b);
    layer8_outputs(7293) <= not a;
    layer8_outputs(7294) <= b;
    layer8_outputs(7295) <= not (a or b);
    layer8_outputs(7296) <= not b;
    layer8_outputs(7297) <= not (a and b);
    layer8_outputs(7298) <= a and b;
    layer8_outputs(7299) <= not a;
    layer8_outputs(7300) <= not (a xor b);
    layer8_outputs(7301) <= b;
    layer8_outputs(7302) <= not a;
    layer8_outputs(7303) <= not a;
    layer8_outputs(7304) <= a xor b;
    layer8_outputs(7305) <= a and not b;
    layer8_outputs(7306) <= not (a xor b);
    layer8_outputs(7307) <= not (a or b);
    layer8_outputs(7308) <= not (a xor b);
    layer8_outputs(7309) <= b;
    layer8_outputs(7310) <= not (a xor b);
    layer8_outputs(7311) <= not a;
    layer8_outputs(7312) <= a or b;
    layer8_outputs(7313) <= a;
    layer8_outputs(7314) <= not b;
    layer8_outputs(7315) <= a;
    layer8_outputs(7316) <= a;
    layer8_outputs(7317) <= a xor b;
    layer8_outputs(7318) <= b;
    layer8_outputs(7319) <= a and b;
    layer8_outputs(7320) <= not (a or b);
    layer8_outputs(7321) <= not (a xor b);
    layer8_outputs(7322) <= b and not a;
    layer8_outputs(7323) <= a and not b;
    layer8_outputs(7324) <= not (a xor b);
    layer8_outputs(7325) <= a;
    layer8_outputs(7326) <= b and not a;
    layer8_outputs(7327) <= a and b;
    layer8_outputs(7328) <= not a;
    layer8_outputs(7329) <= not a or b;
    layer8_outputs(7330) <= a xor b;
    layer8_outputs(7331) <= a or b;
    layer8_outputs(7332) <= not a;
    layer8_outputs(7333) <= not (a and b);
    layer8_outputs(7334) <= a or b;
    layer8_outputs(7335) <= not a;
    layer8_outputs(7336) <= a xor b;
    layer8_outputs(7337) <= b;
    layer8_outputs(7338) <= a and not b;
    layer8_outputs(7339) <= not (a and b);
    layer8_outputs(7340) <= a xor b;
    layer8_outputs(7341) <= b;
    layer8_outputs(7342) <= b;
    layer8_outputs(7343) <= not (a xor b);
    layer8_outputs(7344) <= not b;
    layer8_outputs(7345) <= not (a xor b);
    layer8_outputs(7346) <= a;
    layer8_outputs(7347) <= a and b;
    layer8_outputs(7348) <= not (a or b);
    layer8_outputs(7349) <= a xor b;
    layer8_outputs(7350) <= not b or a;
    layer8_outputs(7351) <= not (a and b);
    layer8_outputs(7352) <= a and not b;
    layer8_outputs(7353) <= not b;
    layer8_outputs(7354) <= not (a xor b);
    layer8_outputs(7355) <= b and not a;
    layer8_outputs(7356) <= a and b;
    layer8_outputs(7357) <= a xor b;
    layer8_outputs(7358) <= a or b;
    layer8_outputs(7359) <= a;
    layer8_outputs(7360) <= a and not b;
    layer8_outputs(7361) <= not (a or b);
    layer8_outputs(7362) <= a and b;
    layer8_outputs(7363) <= a or b;
    layer8_outputs(7364) <= a xor b;
    layer8_outputs(7365) <= not a or b;
    layer8_outputs(7366) <= a xor b;
    layer8_outputs(7367) <= a and b;
    layer8_outputs(7368) <= a;
    layer8_outputs(7369) <= b and not a;
    layer8_outputs(7370) <= b;
    layer8_outputs(7371) <= b and not a;
    layer8_outputs(7372) <= not a;
    layer8_outputs(7373) <= a;
    layer8_outputs(7374) <= not (a xor b);
    layer8_outputs(7375) <= a;
    layer8_outputs(7376) <= not (a xor b);
    layer8_outputs(7377) <= not (a xor b);
    layer8_outputs(7378) <= not b;
    layer8_outputs(7379) <= b;
    layer8_outputs(7380) <= b;
    layer8_outputs(7381) <= b and not a;
    layer8_outputs(7382) <= not b or a;
    layer8_outputs(7383) <= not b;
    layer8_outputs(7384) <= a or b;
    layer8_outputs(7385) <= a xor b;
    layer8_outputs(7386) <= not (a xor b);
    layer8_outputs(7387) <= b;
    layer8_outputs(7388) <= not b;
    layer8_outputs(7389) <= not b;
    layer8_outputs(7390) <= not a;
    layer8_outputs(7391) <= not (a or b);
    layer8_outputs(7392) <= not a or b;
    layer8_outputs(7393) <= a and b;
    layer8_outputs(7394) <= not (a xor b);
    layer8_outputs(7395) <= not a;
    layer8_outputs(7396) <= not b;
    layer8_outputs(7397) <= a;
    layer8_outputs(7398) <= a;
    layer8_outputs(7399) <= not b;
    layer8_outputs(7400) <= a;
    layer8_outputs(7401) <= not b;
    layer8_outputs(7402) <= b;
    layer8_outputs(7403) <= a and b;
    layer8_outputs(7404) <= b;
    layer8_outputs(7405) <= not a;
    layer8_outputs(7406) <= b;
    layer8_outputs(7407) <= not (a and b);
    layer8_outputs(7408) <= not b;
    layer8_outputs(7409) <= a;
    layer8_outputs(7410) <= b;
    layer8_outputs(7411) <= not (a xor b);
    layer8_outputs(7412) <= a and not b;
    layer8_outputs(7413) <= a xor b;
    layer8_outputs(7414) <= a or b;
    layer8_outputs(7415) <= not a;
    layer8_outputs(7416) <= not (a xor b);
    layer8_outputs(7417) <= not b or a;
    layer8_outputs(7418) <= not b;
    layer8_outputs(7419) <= b;
    layer8_outputs(7420) <= a xor b;
    layer8_outputs(7421) <= a;
    layer8_outputs(7422) <= a;
    layer8_outputs(7423) <= not (a and b);
    layer8_outputs(7424) <= a xor b;
    layer8_outputs(7425) <= not b or a;
    layer8_outputs(7426) <= not (a and b);
    layer8_outputs(7427) <= not b or a;
    layer8_outputs(7428) <= not (a xor b);
    layer8_outputs(7429) <= a and b;
    layer8_outputs(7430) <= a;
    layer8_outputs(7431) <= not (a and b);
    layer8_outputs(7432) <= not a;
    layer8_outputs(7433) <= not b;
    layer8_outputs(7434) <= not (a xor b);
    layer8_outputs(7435) <= b;
    layer8_outputs(7436) <= a and b;
    layer8_outputs(7437) <= b and not a;
    layer8_outputs(7438) <= b;
    layer8_outputs(7439) <= not (a or b);
    layer8_outputs(7440) <= b;
    layer8_outputs(7441) <= not a;
    layer8_outputs(7442) <= b and not a;
    layer8_outputs(7443) <= a xor b;
    layer8_outputs(7444) <= a and b;
    layer8_outputs(7445) <= a and b;
    layer8_outputs(7446) <= b;
    layer8_outputs(7447) <= not b;
    layer8_outputs(7448) <= a;
    layer8_outputs(7449) <= a and not b;
    layer8_outputs(7450) <= not b;
    layer8_outputs(7451) <= not (a xor b);
    layer8_outputs(7452) <= a xor b;
    layer8_outputs(7453) <= not (a xor b);
    layer8_outputs(7454) <= not b;
    layer8_outputs(7455) <= not (a or b);
    layer8_outputs(7456) <= a or b;
    layer8_outputs(7457) <= not a;
    layer8_outputs(7458) <= a xor b;
    layer8_outputs(7459) <= not (a xor b);
    layer8_outputs(7460) <= a and b;
    layer8_outputs(7461) <= not b;
    layer8_outputs(7462) <= not b;
    layer8_outputs(7463) <= b;
    layer8_outputs(7464) <= b and not a;
    layer8_outputs(7465) <= not b or a;
    layer8_outputs(7466) <= a or b;
    layer8_outputs(7467) <= not (a xor b);
    layer8_outputs(7468) <= not b or a;
    layer8_outputs(7469) <= not (a xor b);
    layer8_outputs(7470) <= a and b;
    layer8_outputs(7471) <= not a;
    layer8_outputs(7472) <= not a;
    layer8_outputs(7473) <= a;
    layer8_outputs(7474) <= not (a xor b);
    layer8_outputs(7475) <= a and not b;
    layer8_outputs(7476) <= not a or b;
    layer8_outputs(7477) <= b;
    layer8_outputs(7478) <= a;
    layer8_outputs(7479) <= b;
    layer8_outputs(7480) <= a and b;
    layer8_outputs(7481) <= a xor b;
    layer8_outputs(7482) <= a;
    layer8_outputs(7483) <= not (a xor b);
    layer8_outputs(7484) <= not b;
    layer8_outputs(7485) <= a and b;
    layer8_outputs(7486) <= b;
    layer8_outputs(7487) <= not (a xor b);
    layer8_outputs(7488) <= not a;
    layer8_outputs(7489) <= a;
    layer8_outputs(7490) <= not b;
    layer8_outputs(7491) <= a or b;
    layer8_outputs(7492) <= a or b;
    layer8_outputs(7493) <= a;
    layer8_outputs(7494) <= not b;
    layer8_outputs(7495) <= not (a or b);
    layer8_outputs(7496) <= a;
    layer8_outputs(7497) <= a;
    layer8_outputs(7498) <= not (a xor b);
    layer8_outputs(7499) <= not (a xor b);
    layer8_outputs(7500) <= a and not b;
    layer8_outputs(7501) <= a xor b;
    layer8_outputs(7502) <= a xor b;
    layer8_outputs(7503) <= a or b;
    layer8_outputs(7504) <= b;
    layer8_outputs(7505) <= not (a xor b);
    layer8_outputs(7506) <= a and b;
    layer8_outputs(7507) <= a;
    layer8_outputs(7508) <= not (a xor b);
    layer8_outputs(7509) <= b;
    layer8_outputs(7510) <= a xor b;
    layer8_outputs(7511) <= 1'b0;
    layer8_outputs(7512) <= not a or b;
    layer8_outputs(7513) <= not a;
    layer8_outputs(7514) <= not a or b;
    layer8_outputs(7515) <= not (a xor b);
    layer8_outputs(7516) <= not b or a;
    layer8_outputs(7517) <= not a or b;
    layer8_outputs(7518) <= b;
    layer8_outputs(7519) <= a or b;
    layer8_outputs(7520) <= a xor b;
    layer8_outputs(7521) <= not (a xor b);
    layer8_outputs(7522) <= a xor b;
    layer8_outputs(7523) <= not b;
    layer8_outputs(7524) <= not a or b;
    layer8_outputs(7525) <= a xor b;
    layer8_outputs(7526) <= not a;
    layer8_outputs(7527) <= b;
    layer8_outputs(7528) <= a;
    layer8_outputs(7529) <= not a;
    layer8_outputs(7530) <= a or b;
    layer8_outputs(7531) <= not a or b;
    layer8_outputs(7532) <= not b;
    layer8_outputs(7533) <= not b;
    layer8_outputs(7534) <= not b;
    layer8_outputs(7535) <= a xor b;
    layer8_outputs(7536) <= b;
    layer8_outputs(7537) <= not b;
    layer8_outputs(7538) <= not (a xor b);
    layer8_outputs(7539) <= not (a xor b);
    layer8_outputs(7540) <= not a;
    layer8_outputs(7541) <= a xor b;
    layer8_outputs(7542) <= not a;
    layer8_outputs(7543) <= a;
    layer8_outputs(7544) <= a or b;
    layer8_outputs(7545) <= a xor b;
    layer8_outputs(7546) <= b;
    layer8_outputs(7547) <= not b or a;
    layer8_outputs(7548) <= b;
    layer8_outputs(7549) <= a;
    layer8_outputs(7550) <= not b or a;
    layer8_outputs(7551) <= not a or b;
    layer8_outputs(7552) <= a;
    layer8_outputs(7553) <= not b;
    layer8_outputs(7554) <= a;
    layer8_outputs(7555) <= a xor b;
    layer8_outputs(7556) <= not (a xor b);
    layer8_outputs(7557) <= not (a xor b);
    layer8_outputs(7558) <= a xor b;
    layer8_outputs(7559) <= not (a xor b);
    layer8_outputs(7560) <= not (a xor b);
    layer8_outputs(7561) <= a xor b;
    layer8_outputs(7562) <= a xor b;
    layer8_outputs(7563) <= not b;
    layer8_outputs(7564) <= a xor b;
    layer8_outputs(7565) <= not (a or b);
    layer8_outputs(7566) <= a and b;
    layer8_outputs(7567) <= not (a xor b);
    layer8_outputs(7568) <= b;
    layer8_outputs(7569) <= a or b;
    layer8_outputs(7570) <= a or b;
    layer8_outputs(7571) <= not (a and b);
    layer8_outputs(7572) <= b;
    layer8_outputs(7573) <= b;
    layer8_outputs(7574) <= a xor b;
    layer8_outputs(7575) <= not a or b;
    layer8_outputs(7576) <= not (a xor b);
    layer8_outputs(7577) <= a or b;
    layer8_outputs(7578) <= a and b;
    layer8_outputs(7579) <= not b;
    layer8_outputs(7580) <= b;
    layer8_outputs(7581) <= 1'b0;
    layer8_outputs(7582) <= a and not b;
    layer8_outputs(7583) <= not a;
    layer8_outputs(7584) <= not a or b;
    layer8_outputs(7585) <= not b;
    layer8_outputs(7586) <= b;
    layer8_outputs(7587) <= not a;
    layer8_outputs(7588) <= not (a xor b);
    layer8_outputs(7589) <= not (a or b);
    layer8_outputs(7590) <= a;
    layer8_outputs(7591) <= a xor b;
    layer8_outputs(7592) <= b;
    layer8_outputs(7593) <= b and not a;
    layer8_outputs(7594) <= not (a and b);
    layer8_outputs(7595) <= not a;
    layer8_outputs(7596) <= a;
    layer8_outputs(7597) <= a;
    layer8_outputs(7598) <= not (a and b);
    layer8_outputs(7599) <= a;
    layer8_outputs(7600) <= not (a or b);
    layer8_outputs(7601) <= b;
    layer8_outputs(7602) <= a;
    layer8_outputs(7603) <= a;
    layer8_outputs(7604) <= a;
    layer8_outputs(7605) <= b and not a;
    layer8_outputs(7606) <= a xor b;
    layer8_outputs(7607) <= a xor b;
    layer8_outputs(7608) <= a xor b;
    layer8_outputs(7609) <= b;
    layer8_outputs(7610) <= not b;
    layer8_outputs(7611) <= not (a xor b);
    layer8_outputs(7612) <= not (a xor b);
    layer8_outputs(7613) <= b;
    layer8_outputs(7614) <= not b or a;
    layer8_outputs(7615) <= a xor b;
    layer8_outputs(7616) <= a or b;
    layer8_outputs(7617) <= a;
    layer8_outputs(7618) <= b;
    layer8_outputs(7619) <= not b or a;
    layer8_outputs(7620) <= not b or a;
    layer8_outputs(7621) <= a xor b;
    layer8_outputs(7622) <= not a or b;
    layer8_outputs(7623) <= not a;
    layer8_outputs(7624) <= a xor b;
    layer8_outputs(7625) <= not b or a;
    layer8_outputs(7626) <= a xor b;
    layer8_outputs(7627) <= not b or a;
    layer8_outputs(7628) <= b;
    layer8_outputs(7629) <= b;
    layer8_outputs(7630) <= a and b;
    layer8_outputs(7631) <= not a;
    layer8_outputs(7632) <= not (a and b);
    layer8_outputs(7633) <= b and not a;
    layer8_outputs(7634) <= a xor b;
    layer8_outputs(7635) <= a;
    layer8_outputs(7636) <= not (a and b);
    layer8_outputs(7637) <= not b;
    layer8_outputs(7638) <= not (a or b);
    layer8_outputs(7639) <= not a;
    layer8_outputs(7640) <= not a;
    layer8_outputs(7641) <= a or b;
    layer8_outputs(7642) <= b and not a;
    layer8_outputs(7643) <= a xor b;
    layer8_outputs(7644) <= b and not a;
    layer8_outputs(7645) <= a;
    layer8_outputs(7646) <= a;
    layer8_outputs(7647) <= a;
    layer8_outputs(7648) <= not a or b;
    layer8_outputs(7649) <= a and not b;
    layer8_outputs(7650) <= a;
    layer8_outputs(7651) <= not (a and b);
    layer8_outputs(7652) <= a xor b;
    layer8_outputs(7653) <= not (a and b);
    layer8_outputs(7654) <= not a or b;
    layer8_outputs(7655) <= b;
    layer8_outputs(7656) <= a xor b;
    layer8_outputs(7657) <= not (a and b);
    layer8_outputs(7658) <= b;
    layer8_outputs(7659) <= not b;
    layer8_outputs(7660) <= a and b;
    layer8_outputs(7661) <= b;
    layer8_outputs(7662) <= a;
    layer8_outputs(7663) <= a xor b;
    layer8_outputs(7664) <= a and not b;
    layer8_outputs(7665) <= not a;
    layer8_outputs(7666) <= not (a or b);
    layer8_outputs(7667) <= b and not a;
    layer8_outputs(7668) <= a xor b;
    layer8_outputs(7669) <= not a or b;
    layer8_outputs(7670) <= not (a xor b);
    layer8_outputs(7671) <= not a or b;
    layer8_outputs(7672) <= not (a and b);
    layer8_outputs(7673) <= not a;
    layer8_outputs(7674) <= not a or b;
    layer8_outputs(7675) <= a xor b;
    layer8_outputs(7676) <= a and not b;
    layer8_outputs(7677) <= not b or a;
    layer8_outputs(7678) <= 1'b1;
    layer8_outputs(7679) <= a or b;
    layer8_outputs(7680) <= b;
    layer8_outputs(7681) <= not (a xor b);
    layer8_outputs(7682) <= a;
    layer8_outputs(7683) <= a and not b;
    layer8_outputs(7684) <= a and not b;
    layer8_outputs(7685) <= not a;
    layer8_outputs(7686) <= a xor b;
    layer8_outputs(7687) <= a or b;
    layer8_outputs(7688) <= not (a xor b);
    layer8_outputs(7689) <= a xor b;
    layer8_outputs(7690) <= not a;
    layer8_outputs(7691) <= a and not b;
    layer8_outputs(7692) <= a xor b;
    layer8_outputs(7693) <= not (a and b);
    layer8_outputs(7694) <= a;
    layer8_outputs(7695) <= not (a xor b);
    layer8_outputs(7696) <= b;
    layer8_outputs(7697) <= a;
    layer8_outputs(7698) <= a and not b;
    layer8_outputs(7699) <= b;
    layer8_outputs(7700) <= not b;
    layer8_outputs(7701) <= b;
    layer8_outputs(7702) <= not (a or b);
    layer8_outputs(7703) <= not (a xor b);
    layer8_outputs(7704) <= b;
    layer8_outputs(7705) <= b;
    layer8_outputs(7706) <= not a;
    layer8_outputs(7707) <= not b;
    layer8_outputs(7708) <= not b;
    layer8_outputs(7709) <= a and not b;
    layer8_outputs(7710) <= a;
    layer8_outputs(7711) <= not b or a;
    layer8_outputs(7712) <= not (a and b);
    layer8_outputs(7713) <= not (a xor b);
    layer8_outputs(7714) <= not (a xor b);
    layer8_outputs(7715) <= not b;
    layer8_outputs(7716) <= not b or a;
    layer8_outputs(7717) <= b and not a;
    layer8_outputs(7718) <= not b;
    layer8_outputs(7719) <= b;
    layer8_outputs(7720) <= b;
    layer8_outputs(7721) <= not (a xor b);
    layer8_outputs(7722) <= not (a and b);
    layer8_outputs(7723) <= b and not a;
    layer8_outputs(7724) <= not a;
    layer8_outputs(7725) <= a xor b;
    layer8_outputs(7726) <= a;
    layer8_outputs(7727) <= not (a xor b);
    layer8_outputs(7728) <= not a or b;
    layer8_outputs(7729) <= a;
    layer8_outputs(7730) <= b;
    layer8_outputs(7731) <= a;
    layer8_outputs(7732) <= b and not a;
    layer8_outputs(7733) <= a;
    layer8_outputs(7734) <= not b;
    layer8_outputs(7735) <= b;
    layer8_outputs(7736) <= not b or a;
    layer8_outputs(7737) <= b;
    layer8_outputs(7738) <= a;
    layer8_outputs(7739) <= not a;
    layer8_outputs(7740) <= a xor b;
    layer8_outputs(7741) <= a xor b;
    layer8_outputs(7742) <= not a;
    layer8_outputs(7743) <= a and not b;
    layer8_outputs(7744) <= not b;
    layer8_outputs(7745) <= b and not a;
    layer8_outputs(7746) <= not b;
    layer8_outputs(7747) <= a xor b;
    layer8_outputs(7748) <= a;
    layer8_outputs(7749) <= a and b;
    layer8_outputs(7750) <= a and not b;
    layer8_outputs(7751) <= a xor b;
    layer8_outputs(7752) <= b and not a;
    layer8_outputs(7753) <= b;
    layer8_outputs(7754) <= not b;
    layer8_outputs(7755) <= not a or b;
    layer8_outputs(7756) <= not b or a;
    layer8_outputs(7757) <= not b;
    layer8_outputs(7758) <= not a;
    layer8_outputs(7759) <= a and b;
    layer8_outputs(7760) <= not a;
    layer8_outputs(7761) <= a xor b;
    layer8_outputs(7762) <= b;
    layer8_outputs(7763) <= not b;
    layer8_outputs(7764) <= a xor b;
    layer8_outputs(7765) <= b;
    layer8_outputs(7766) <= not (a or b);
    layer8_outputs(7767) <= not a;
    layer8_outputs(7768) <= a;
    layer8_outputs(7769) <= b and not a;
    layer8_outputs(7770) <= not a or b;
    layer8_outputs(7771) <= a and b;
    layer8_outputs(7772) <= a;
    layer8_outputs(7773) <= not (a and b);
    layer8_outputs(7774) <= a and not b;
    layer8_outputs(7775) <= not a;
    layer8_outputs(7776) <= a and b;
    layer8_outputs(7777) <= b;
    layer8_outputs(7778) <= not (a or b);
    layer8_outputs(7779) <= b;
    layer8_outputs(7780) <= b;
    layer8_outputs(7781) <= not a;
    layer8_outputs(7782) <= not b;
    layer8_outputs(7783) <= b and not a;
    layer8_outputs(7784) <= not (a xor b);
    layer8_outputs(7785) <= a;
    layer8_outputs(7786) <= a;
    layer8_outputs(7787) <= b;
    layer8_outputs(7788) <= not a;
    layer8_outputs(7789) <= a;
    layer8_outputs(7790) <= 1'b1;
    layer8_outputs(7791) <= a and b;
    layer8_outputs(7792) <= a xor b;
    layer8_outputs(7793) <= not b or a;
    layer8_outputs(7794) <= not a;
    layer8_outputs(7795) <= not a or b;
    layer8_outputs(7796) <= a xor b;
    layer8_outputs(7797) <= b;
    layer8_outputs(7798) <= not a;
    layer8_outputs(7799) <= not b;
    layer8_outputs(7800) <= not (a or b);
    layer8_outputs(7801) <= not (a xor b);
    layer8_outputs(7802) <= a and b;
    layer8_outputs(7803) <= b;
    layer8_outputs(7804) <= not (a or b);
    layer8_outputs(7805) <= not a;
    layer8_outputs(7806) <= a;
    layer8_outputs(7807) <= b;
    layer8_outputs(7808) <= b;
    layer8_outputs(7809) <= a and not b;
    layer8_outputs(7810) <= not a;
    layer8_outputs(7811) <= a;
    layer8_outputs(7812) <= a;
    layer8_outputs(7813) <= not (a and b);
    layer8_outputs(7814) <= a;
    layer8_outputs(7815) <= b;
    layer8_outputs(7816) <= b;
    layer8_outputs(7817) <= a or b;
    layer8_outputs(7818) <= b and not a;
    layer8_outputs(7819) <= not b;
    layer8_outputs(7820) <= not a or b;
    layer8_outputs(7821) <= a and b;
    layer8_outputs(7822) <= b;
    layer8_outputs(7823) <= not b;
    layer8_outputs(7824) <= a or b;
    layer8_outputs(7825) <= a and b;
    layer8_outputs(7826) <= not (a and b);
    layer8_outputs(7827) <= a and b;
    layer8_outputs(7828) <= b;
    layer8_outputs(7829) <= not a;
    layer8_outputs(7830) <= b;
    layer8_outputs(7831) <= not (a xor b);
    layer8_outputs(7832) <= a and not b;
    layer8_outputs(7833) <= not (a xor b);
    layer8_outputs(7834) <= not b;
    layer8_outputs(7835) <= not a or b;
    layer8_outputs(7836) <= a and b;
    layer8_outputs(7837) <= not (a xor b);
    layer8_outputs(7838) <= a xor b;
    layer8_outputs(7839) <= a or b;
    layer8_outputs(7840) <= not b;
    layer8_outputs(7841) <= a or b;
    layer8_outputs(7842) <= a xor b;
    layer8_outputs(7843) <= not b;
    layer8_outputs(7844) <= a or b;
    layer8_outputs(7845) <= not b;
    layer8_outputs(7846) <= a and not b;
    layer8_outputs(7847) <= not (a or b);
    layer8_outputs(7848) <= not a;
    layer8_outputs(7849) <= not a;
    layer8_outputs(7850) <= a xor b;
    layer8_outputs(7851) <= a and not b;
    layer8_outputs(7852) <= a xor b;
    layer8_outputs(7853) <= a xor b;
    layer8_outputs(7854) <= not (a xor b);
    layer8_outputs(7855) <= not a or b;
    layer8_outputs(7856) <= a and b;
    layer8_outputs(7857) <= not b;
    layer8_outputs(7858) <= not (a and b);
    layer8_outputs(7859) <= not (a or b);
    layer8_outputs(7860) <= not b;
    layer8_outputs(7861) <= 1'b0;
    layer8_outputs(7862) <= not b or a;
    layer8_outputs(7863) <= not b or a;
    layer8_outputs(7864) <= not b;
    layer8_outputs(7865) <= not a;
    layer8_outputs(7866) <= not (a or b);
    layer8_outputs(7867) <= b;
    layer8_outputs(7868) <= not (a xor b);
    layer8_outputs(7869) <= not (a and b);
    layer8_outputs(7870) <= b;
    layer8_outputs(7871) <= not a;
    layer8_outputs(7872) <= a;
    layer8_outputs(7873) <= a xor b;
    layer8_outputs(7874) <= b;
    layer8_outputs(7875) <= b;
    layer8_outputs(7876) <= a;
    layer8_outputs(7877) <= a and b;
    layer8_outputs(7878) <= a or b;
    layer8_outputs(7879) <= b;
    layer8_outputs(7880) <= not (a xor b);
    layer8_outputs(7881) <= not b;
    layer8_outputs(7882) <= not (a or b);
    layer8_outputs(7883) <= not b;
    layer8_outputs(7884) <= a xor b;
    layer8_outputs(7885) <= not a;
    layer8_outputs(7886) <= a xor b;
    layer8_outputs(7887) <= a or b;
    layer8_outputs(7888) <= a and b;
    layer8_outputs(7889) <= not (a xor b);
    layer8_outputs(7890) <= not a or b;
    layer8_outputs(7891) <= a xor b;
    layer8_outputs(7892) <= a;
    layer8_outputs(7893) <= not (a xor b);
    layer8_outputs(7894) <= a and b;
    layer8_outputs(7895) <= a;
    layer8_outputs(7896) <= a;
    layer8_outputs(7897) <= not b;
    layer8_outputs(7898) <= b and not a;
    layer8_outputs(7899) <= a and not b;
    layer8_outputs(7900) <= a;
    layer8_outputs(7901) <= not (a and b);
    layer8_outputs(7902) <= a xor b;
    layer8_outputs(7903) <= a xor b;
    layer8_outputs(7904) <= not a;
    layer8_outputs(7905) <= a and b;
    layer8_outputs(7906) <= b and not a;
    layer8_outputs(7907) <= b;
    layer8_outputs(7908) <= not (a xor b);
    layer8_outputs(7909) <= not (a and b);
    layer8_outputs(7910) <= not a;
    layer8_outputs(7911) <= not (a xor b);
    layer8_outputs(7912) <= not (a xor b);
    layer8_outputs(7913) <= not b;
    layer8_outputs(7914) <= b and not a;
    layer8_outputs(7915) <= a and b;
    layer8_outputs(7916) <= not a;
    layer8_outputs(7917) <= a xor b;
    layer8_outputs(7918) <= a;
    layer8_outputs(7919) <= not a;
    layer8_outputs(7920) <= b;
    layer8_outputs(7921) <= not (a or b);
    layer8_outputs(7922) <= a and not b;
    layer8_outputs(7923) <= not a;
    layer8_outputs(7924) <= a xor b;
    layer8_outputs(7925) <= not (a xor b);
    layer8_outputs(7926) <= not a;
    layer8_outputs(7927) <= b and not a;
    layer8_outputs(7928) <= b;
    layer8_outputs(7929) <= a or b;
    layer8_outputs(7930) <= not (a or b);
    layer8_outputs(7931) <= not b;
    layer8_outputs(7932) <= a xor b;
    layer8_outputs(7933) <= not b or a;
    layer8_outputs(7934) <= not b;
    layer8_outputs(7935) <= b;
    layer8_outputs(7936) <= not b;
    layer8_outputs(7937) <= a or b;
    layer8_outputs(7938) <= a and not b;
    layer8_outputs(7939) <= not (a or b);
    layer8_outputs(7940) <= not (a xor b);
    layer8_outputs(7941) <= not (a xor b);
    layer8_outputs(7942) <= not (a and b);
    layer8_outputs(7943) <= not a;
    layer8_outputs(7944) <= not a or b;
    layer8_outputs(7945) <= a and b;
    layer8_outputs(7946) <= a xor b;
    layer8_outputs(7947) <= a and not b;
    layer8_outputs(7948) <= a xor b;
    layer8_outputs(7949) <= not b;
    layer8_outputs(7950) <= a or b;
    layer8_outputs(7951) <= 1'b1;
    layer8_outputs(7952) <= not (a xor b);
    layer8_outputs(7953) <= not b;
    layer8_outputs(7954) <= not (a xor b);
    layer8_outputs(7955) <= a and b;
    layer8_outputs(7956) <= not a;
    layer8_outputs(7957) <= not (a and b);
    layer8_outputs(7958) <= not a;
    layer8_outputs(7959) <= not b;
    layer8_outputs(7960) <= not a or b;
    layer8_outputs(7961) <= a and b;
    layer8_outputs(7962) <= a and b;
    layer8_outputs(7963) <= not b;
    layer8_outputs(7964) <= a or b;
    layer8_outputs(7965) <= not b;
    layer8_outputs(7966) <= a;
    layer8_outputs(7967) <= b;
    layer8_outputs(7968) <= not (a xor b);
    layer8_outputs(7969) <= b;
    layer8_outputs(7970) <= not a or b;
    layer8_outputs(7971) <= a and b;
    layer8_outputs(7972) <= not (a or b);
    layer8_outputs(7973) <= not a;
    layer8_outputs(7974) <= not a or b;
    layer8_outputs(7975) <= not (a xor b);
    layer8_outputs(7976) <= not (a or b);
    layer8_outputs(7977) <= not (a xor b);
    layer8_outputs(7978) <= a;
    layer8_outputs(7979) <= not a;
    layer8_outputs(7980) <= not b;
    layer8_outputs(7981) <= a;
    layer8_outputs(7982) <= a;
    layer8_outputs(7983) <= not (a xor b);
    layer8_outputs(7984) <= not (a and b);
    layer8_outputs(7985) <= a xor b;
    layer8_outputs(7986) <= not b or a;
    layer8_outputs(7987) <= a xor b;
    layer8_outputs(7988) <= not b;
    layer8_outputs(7989) <= b;
    layer8_outputs(7990) <= not b;
    layer8_outputs(7991) <= not a;
    layer8_outputs(7992) <= a and not b;
    layer8_outputs(7993) <= a;
    layer8_outputs(7994) <= b;
    layer8_outputs(7995) <= not (a or b);
    layer8_outputs(7996) <= not (a xor b);
    layer8_outputs(7997) <= a and b;
    layer8_outputs(7998) <= not b or a;
    layer8_outputs(7999) <= not (a and b);
    layer8_outputs(8000) <= a and not b;
    layer8_outputs(8001) <= not (a xor b);
    layer8_outputs(8002) <= a and b;
    layer8_outputs(8003) <= not (a xor b);
    layer8_outputs(8004) <= not (a and b);
    layer8_outputs(8005) <= not b;
    layer8_outputs(8006) <= b;
    layer8_outputs(8007) <= not (a xor b);
    layer8_outputs(8008) <= a or b;
    layer8_outputs(8009) <= b;
    layer8_outputs(8010) <= not a;
    layer8_outputs(8011) <= a;
    layer8_outputs(8012) <= a;
    layer8_outputs(8013) <= not (a or b);
    layer8_outputs(8014) <= b;
    layer8_outputs(8015) <= b;
    layer8_outputs(8016) <= not (a xor b);
    layer8_outputs(8017) <= not b;
    layer8_outputs(8018) <= not (a and b);
    layer8_outputs(8019) <= b and not a;
    layer8_outputs(8020) <= not b or a;
    layer8_outputs(8021) <= 1'b0;
    layer8_outputs(8022) <= not (a xor b);
    layer8_outputs(8023) <= not b;
    layer8_outputs(8024) <= a xor b;
    layer8_outputs(8025) <= a xor b;
    layer8_outputs(8026) <= a and not b;
    layer8_outputs(8027) <= b;
    layer8_outputs(8028) <= a xor b;
    layer8_outputs(8029) <= not b;
    layer8_outputs(8030) <= b;
    layer8_outputs(8031) <= a;
    layer8_outputs(8032) <= a xor b;
    layer8_outputs(8033) <= a;
    layer8_outputs(8034) <= a;
    layer8_outputs(8035) <= b;
    layer8_outputs(8036) <= a;
    layer8_outputs(8037) <= not a;
    layer8_outputs(8038) <= a;
    layer8_outputs(8039) <= not (a or b);
    layer8_outputs(8040) <= not a;
    layer8_outputs(8041) <= not (a xor b);
    layer8_outputs(8042) <= not a or b;
    layer8_outputs(8043) <= not a;
    layer8_outputs(8044) <= b;
    layer8_outputs(8045) <= a;
    layer8_outputs(8046) <= not b;
    layer8_outputs(8047) <= b;
    layer8_outputs(8048) <= not (a and b);
    layer8_outputs(8049) <= a xor b;
    layer8_outputs(8050) <= a xor b;
    layer8_outputs(8051) <= a or b;
    layer8_outputs(8052) <= not (a xor b);
    layer8_outputs(8053) <= a and b;
    layer8_outputs(8054) <= not a;
    layer8_outputs(8055) <= not (a and b);
    layer8_outputs(8056) <= not a;
    layer8_outputs(8057) <= not b or a;
    layer8_outputs(8058) <= not (a or b);
    layer8_outputs(8059) <= b;
    layer8_outputs(8060) <= a xor b;
    layer8_outputs(8061) <= a and not b;
    layer8_outputs(8062) <= not (a or b);
    layer8_outputs(8063) <= b;
    layer8_outputs(8064) <= a xor b;
    layer8_outputs(8065) <= not b;
    layer8_outputs(8066) <= not b;
    layer8_outputs(8067) <= a xor b;
    layer8_outputs(8068) <= not b;
    layer8_outputs(8069) <= not b;
    layer8_outputs(8070) <= not (a xor b);
    layer8_outputs(8071) <= a;
    layer8_outputs(8072) <= b and not a;
    layer8_outputs(8073) <= not a;
    layer8_outputs(8074) <= a;
    layer8_outputs(8075) <= not b;
    layer8_outputs(8076) <= not (a xor b);
    layer8_outputs(8077) <= not (a xor b);
    layer8_outputs(8078) <= a xor b;
    layer8_outputs(8079) <= not b;
    layer8_outputs(8080) <= not (a xor b);
    layer8_outputs(8081) <= not a;
    layer8_outputs(8082) <= a and b;
    layer8_outputs(8083) <= not a;
    layer8_outputs(8084) <= a xor b;
    layer8_outputs(8085) <= b;
    layer8_outputs(8086) <= not a or b;
    layer8_outputs(8087) <= not (a xor b);
    layer8_outputs(8088) <= not b;
    layer8_outputs(8089) <= b;
    layer8_outputs(8090) <= not a or b;
    layer8_outputs(8091) <= a xor b;
    layer8_outputs(8092) <= not (a xor b);
    layer8_outputs(8093) <= not b;
    layer8_outputs(8094) <= a xor b;
    layer8_outputs(8095) <= 1'b1;
    layer8_outputs(8096) <= not b;
    layer8_outputs(8097) <= not a or b;
    layer8_outputs(8098) <= not (a and b);
    layer8_outputs(8099) <= not a;
    layer8_outputs(8100) <= not a;
    layer8_outputs(8101) <= not b;
    layer8_outputs(8102) <= not a;
    layer8_outputs(8103) <= not (a xor b);
    layer8_outputs(8104) <= not (a xor b);
    layer8_outputs(8105) <= a and not b;
    layer8_outputs(8106) <= not b or a;
    layer8_outputs(8107) <= a;
    layer8_outputs(8108) <= not (a xor b);
    layer8_outputs(8109) <= a;
    layer8_outputs(8110) <= a;
    layer8_outputs(8111) <= b;
    layer8_outputs(8112) <= not b;
    layer8_outputs(8113) <= not a;
    layer8_outputs(8114) <= b;
    layer8_outputs(8115) <= not a;
    layer8_outputs(8116) <= not a;
    layer8_outputs(8117) <= not a or b;
    layer8_outputs(8118) <= not (a xor b);
    layer8_outputs(8119) <= a or b;
    layer8_outputs(8120) <= not a;
    layer8_outputs(8121) <= b and not a;
    layer8_outputs(8122) <= not (a xor b);
    layer8_outputs(8123) <= not a;
    layer8_outputs(8124) <= a or b;
    layer8_outputs(8125) <= a xor b;
    layer8_outputs(8126) <= b;
    layer8_outputs(8127) <= not b;
    layer8_outputs(8128) <= a xor b;
    layer8_outputs(8129) <= a and b;
    layer8_outputs(8130) <= not b or a;
    layer8_outputs(8131) <= not b or a;
    layer8_outputs(8132) <= a;
    layer8_outputs(8133) <= not b or a;
    layer8_outputs(8134) <= not a;
    layer8_outputs(8135) <= not a;
    layer8_outputs(8136) <= not b or a;
    layer8_outputs(8137) <= a;
    layer8_outputs(8138) <= a and not b;
    layer8_outputs(8139) <= a or b;
    layer8_outputs(8140) <= not (a xor b);
    layer8_outputs(8141) <= not (a or b);
    layer8_outputs(8142) <= a xor b;
    layer8_outputs(8143) <= not b;
    layer8_outputs(8144) <= not a;
    layer8_outputs(8145) <= not b or a;
    layer8_outputs(8146) <= a xor b;
    layer8_outputs(8147) <= a and not b;
    layer8_outputs(8148) <= a;
    layer8_outputs(8149) <= a;
    layer8_outputs(8150) <= a and not b;
    layer8_outputs(8151) <= a or b;
    layer8_outputs(8152) <= b;
    layer8_outputs(8153) <= a xor b;
    layer8_outputs(8154) <= not b or a;
    layer8_outputs(8155) <= not b;
    layer8_outputs(8156) <= b;
    layer8_outputs(8157) <= not (a or b);
    layer8_outputs(8158) <= a and not b;
    layer8_outputs(8159) <= not (a or b);
    layer8_outputs(8160) <= a xor b;
    layer8_outputs(8161) <= a and not b;
    layer8_outputs(8162) <= not (a and b);
    layer8_outputs(8163) <= a;
    layer8_outputs(8164) <= not b or a;
    layer8_outputs(8165) <= a or b;
    layer8_outputs(8166) <= not a or b;
    layer8_outputs(8167) <= not b;
    layer8_outputs(8168) <= not b;
    layer8_outputs(8169) <= not b;
    layer8_outputs(8170) <= b and not a;
    layer8_outputs(8171) <= a and not b;
    layer8_outputs(8172) <= a;
    layer8_outputs(8173) <= a and not b;
    layer8_outputs(8174) <= a;
    layer8_outputs(8175) <= a;
    layer8_outputs(8176) <= b and not a;
    layer8_outputs(8177) <= a;
    layer8_outputs(8178) <= a;
    layer8_outputs(8179) <= a xor b;
    layer8_outputs(8180) <= not a;
    layer8_outputs(8181) <= not (a xor b);
    layer8_outputs(8182) <= a and not b;
    layer8_outputs(8183) <= a and not b;
    layer8_outputs(8184) <= not a;
    layer8_outputs(8185) <= not b;
    layer8_outputs(8186) <= not a;
    layer8_outputs(8187) <= not (a or b);
    layer8_outputs(8188) <= a xor b;
    layer8_outputs(8189) <= not (a and b);
    layer8_outputs(8190) <= a or b;
    layer8_outputs(8191) <= a xor b;
    layer8_outputs(8192) <= not (a or b);
    layer8_outputs(8193) <= b and not a;
    layer8_outputs(8194) <= b and not a;
    layer8_outputs(8195) <= b and not a;
    layer8_outputs(8196) <= a xor b;
    layer8_outputs(8197) <= not (a xor b);
    layer8_outputs(8198) <= a xor b;
    layer8_outputs(8199) <= not b;
    layer8_outputs(8200) <= not a or b;
    layer8_outputs(8201) <= a and b;
    layer8_outputs(8202) <= not (a xor b);
    layer8_outputs(8203) <= not (a xor b);
    layer8_outputs(8204) <= not (a xor b);
    layer8_outputs(8205) <= a or b;
    layer8_outputs(8206) <= a xor b;
    layer8_outputs(8207) <= b and not a;
    layer8_outputs(8208) <= not (a xor b);
    layer8_outputs(8209) <= not b or a;
    layer8_outputs(8210) <= b;
    layer8_outputs(8211) <= b;
    layer8_outputs(8212) <= b;
    layer8_outputs(8213) <= not b;
    layer8_outputs(8214) <= not b;
    layer8_outputs(8215) <= not b;
    layer8_outputs(8216) <= a and b;
    layer8_outputs(8217) <= a or b;
    layer8_outputs(8218) <= a and b;
    layer8_outputs(8219) <= not a or b;
    layer8_outputs(8220) <= not a;
    layer8_outputs(8221) <= 1'b1;
    layer8_outputs(8222) <= 1'b1;
    layer8_outputs(8223) <= not (a and b);
    layer8_outputs(8224) <= not a or b;
    layer8_outputs(8225) <= not (a xor b);
    layer8_outputs(8226) <= b and not a;
    layer8_outputs(8227) <= b;
    layer8_outputs(8228) <= a;
    layer8_outputs(8229) <= a;
    layer8_outputs(8230) <= not (a xor b);
    layer8_outputs(8231) <= a;
    layer8_outputs(8232) <= a and not b;
    layer8_outputs(8233) <= not b;
    layer8_outputs(8234) <= not a or b;
    layer8_outputs(8235) <= not a;
    layer8_outputs(8236) <= not (a xor b);
    layer8_outputs(8237) <= a and b;
    layer8_outputs(8238) <= b;
    layer8_outputs(8239) <= not b;
    layer8_outputs(8240) <= a and not b;
    layer8_outputs(8241) <= b and not a;
    layer8_outputs(8242) <= b;
    layer8_outputs(8243) <= b;
    layer8_outputs(8244) <= not b or a;
    layer8_outputs(8245) <= not (a xor b);
    layer8_outputs(8246) <= a or b;
    layer8_outputs(8247) <= b;
    layer8_outputs(8248) <= not a;
    layer8_outputs(8249) <= a;
    layer8_outputs(8250) <= not a or b;
    layer8_outputs(8251) <= not (a and b);
    layer8_outputs(8252) <= a xor b;
    layer8_outputs(8253) <= a or b;
    layer8_outputs(8254) <= not a;
    layer8_outputs(8255) <= b;
    layer8_outputs(8256) <= not (a or b);
    layer8_outputs(8257) <= a;
    layer8_outputs(8258) <= not b or a;
    layer8_outputs(8259) <= not (a or b);
    layer8_outputs(8260) <= not b;
    layer8_outputs(8261) <= a;
    layer8_outputs(8262) <= not b;
    layer8_outputs(8263) <= a and not b;
    layer8_outputs(8264) <= not a or b;
    layer8_outputs(8265) <= not a or b;
    layer8_outputs(8266) <= not a;
    layer8_outputs(8267) <= a and not b;
    layer8_outputs(8268) <= not b;
    layer8_outputs(8269) <= b;
    layer8_outputs(8270) <= not b;
    layer8_outputs(8271) <= not b or a;
    layer8_outputs(8272) <= not (a xor b);
    layer8_outputs(8273) <= not b or a;
    layer8_outputs(8274) <= not a or b;
    layer8_outputs(8275) <= not (a xor b);
    layer8_outputs(8276) <= b;
    layer8_outputs(8277) <= a xor b;
    layer8_outputs(8278) <= a and b;
    layer8_outputs(8279) <= not a or b;
    layer8_outputs(8280) <= b;
    layer8_outputs(8281) <= not (a xor b);
    layer8_outputs(8282) <= a;
    layer8_outputs(8283) <= not (a xor b);
    layer8_outputs(8284) <= not b or a;
    layer8_outputs(8285) <= not b;
    layer8_outputs(8286) <= b;
    layer8_outputs(8287) <= not (a xor b);
    layer8_outputs(8288) <= a;
    layer8_outputs(8289) <= 1'b0;
    layer8_outputs(8290) <= a;
    layer8_outputs(8291) <= not (a xor b);
    layer8_outputs(8292) <= not b or a;
    layer8_outputs(8293) <= not b;
    layer8_outputs(8294) <= not (a xor b);
    layer8_outputs(8295) <= not a;
    layer8_outputs(8296) <= not (a or b);
    layer8_outputs(8297) <= a xor b;
    layer8_outputs(8298) <= not a;
    layer8_outputs(8299) <= a and not b;
    layer8_outputs(8300) <= not a;
    layer8_outputs(8301) <= not (a xor b);
    layer8_outputs(8302) <= b;
    layer8_outputs(8303) <= a xor b;
    layer8_outputs(8304) <= not (a xor b);
    layer8_outputs(8305) <= not b;
    layer8_outputs(8306) <= a or b;
    layer8_outputs(8307) <= b and not a;
    layer8_outputs(8308) <= not b;
    layer8_outputs(8309) <= not b;
    layer8_outputs(8310) <= a;
    layer8_outputs(8311) <= not (a xor b);
    layer8_outputs(8312) <= b;
    layer8_outputs(8313) <= not b or a;
    layer8_outputs(8314) <= not (a or b);
    layer8_outputs(8315) <= b;
    layer8_outputs(8316) <= b;
    layer8_outputs(8317) <= a and b;
    layer8_outputs(8318) <= a;
    layer8_outputs(8319) <= a;
    layer8_outputs(8320) <= a xor b;
    layer8_outputs(8321) <= not (a xor b);
    layer8_outputs(8322) <= not b;
    layer8_outputs(8323) <= not (a xor b);
    layer8_outputs(8324) <= not b;
    layer8_outputs(8325) <= a and b;
    layer8_outputs(8326) <= a or b;
    layer8_outputs(8327) <= a and not b;
    layer8_outputs(8328) <= a;
    layer8_outputs(8329) <= not a;
    layer8_outputs(8330) <= not a;
    layer8_outputs(8331) <= a or b;
    layer8_outputs(8332) <= not (a or b);
    layer8_outputs(8333) <= not a or b;
    layer8_outputs(8334) <= b;
    layer8_outputs(8335) <= not b or a;
    layer8_outputs(8336) <= b;
    layer8_outputs(8337) <= b and not a;
    layer8_outputs(8338) <= a xor b;
    layer8_outputs(8339) <= not a;
    layer8_outputs(8340) <= not (a xor b);
    layer8_outputs(8341) <= not a;
    layer8_outputs(8342) <= not (a and b);
    layer8_outputs(8343) <= not b;
    layer8_outputs(8344) <= a;
    layer8_outputs(8345) <= a;
    layer8_outputs(8346) <= not (a and b);
    layer8_outputs(8347) <= a;
    layer8_outputs(8348) <= not (a or b);
    layer8_outputs(8349) <= a xor b;
    layer8_outputs(8350) <= not a or b;
    layer8_outputs(8351) <= a or b;
    layer8_outputs(8352) <= not a;
    layer8_outputs(8353) <= 1'b0;
    layer8_outputs(8354) <= not b;
    layer8_outputs(8355) <= b;
    layer8_outputs(8356) <= not b;
    layer8_outputs(8357) <= b;
    layer8_outputs(8358) <= not (a xor b);
    layer8_outputs(8359) <= b;
    layer8_outputs(8360) <= not b;
    layer8_outputs(8361) <= a;
    layer8_outputs(8362) <= b and not a;
    layer8_outputs(8363) <= a xor b;
    layer8_outputs(8364) <= not (a xor b);
    layer8_outputs(8365) <= not (a xor b);
    layer8_outputs(8366) <= not b;
    layer8_outputs(8367) <= not (a xor b);
    layer8_outputs(8368) <= b;
    layer8_outputs(8369) <= a xor b;
    layer8_outputs(8370) <= b;
    layer8_outputs(8371) <= not a or b;
    layer8_outputs(8372) <= a and not b;
    layer8_outputs(8373) <= a or b;
    layer8_outputs(8374) <= b;
    layer8_outputs(8375) <= not (a xor b);
    layer8_outputs(8376) <= not (a xor b);
    layer8_outputs(8377) <= a xor b;
    layer8_outputs(8378) <= not (a xor b);
    layer8_outputs(8379) <= not b;
    layer8_outputs(8380) <= not a;
    layer8_outputs(8381) <= not (a and b);
    layer8_outputs(8382) <= b;
    layer8_outputs(8383) <= not (a xor b);
    layer8_outputs(8384) <= not (a xor b);
    layer8_outputs(8385) <= not a;
    layer8_outputs(8386) <= b;
    layer8_outputs(8387) <= a xor b;
    layer8_outputs(8388) <= 1'b0;
    layer8_outputs(8389) <= not b or a;
    layer8_outputs(8390) <= not b;
    layer8_outputs(8391) <= not a or b;
    layer8_outputs(8392) <= b;
    layer8_outputs(8393) <= not a;
    layer8_outputs(8394) <= a or b;
    layer8_outputs(8395) <= not a;
    layer8_outputs(8396) <= a xor b;
    layer8_outputs(8397) <= not (a or b);
    layer8_outputs(8398) <= a;
    layer8_outputs(8399) <= not (a xor b);
    layer8_outputs(8400) <= not (a xor b);
    layer8_outputs(8401) <= not (a or b);
    layer8_outputs(8402) <= a xor b;
    layer8_outputs(8403) <= not (a xor b);
    layer8_outputs(8404) <= a and b;
    layer8_outputs(8405) <= b;
    layer8_outputs(8406) <= a and not b;
    layer8_outputs(8407) <= not a;
    layer8_outputs(8408) <= not (a xor b);
    layer8_outputs(8409) <= not a or b;
    layer8_outputs(8410) <= not (a xor b);
    layer8_outputs(8411) <= b and not a;
    layer8_outputs(8412) <= not (a and b);
    layer8_outputs(8413) <= b;
    layer8_outputs(8414) <= not a;
    layer8_outputs(8415) <= 1'b0;
    layer8_outputs(8416) <= b;
    layer8_outputs(8417) <= not a;
    layer8_outputs(8418) <= a;
    layer8_outputs(8419) <= not a;
    layer8_outputs(8420) <= not a;
    layer8_outputs(8421) <= not b;
    layer8_outputs(8422) <= a or b;
    layer8_outputs(8423) <= not b;
    layer8_outputs(8424) <= b;
    layer8_outputs(8425) <= b and not a;
    layer8_outputs(8426) <= b and not a;
    layer8_outputs(8427) <= b;
    layer8_outputs(8428) <= b;
    layer8_outputs(8429) <= a;
    layer8_outputs(8430) <= not a;
    layer8_outputs(8431) <= not b;
    layer8_outputs(8432) <= not (a or b);
    layer8_outputs(8433) <= not b;
    layer8_outputs(8434) <= not a;
    layer8_outputs(8435) <= not (a xor b);
    layer8_outputs(8436) <= not (a and b);
    layer8_outputs(8437) <= not b;
    layer8_outputs(8438) <= a;
    layer8_outputs(8439) <= not (a and b);
    layer8_outputs(8440) <= b and not a;
    layer8_outputs(8441) <= b;
    layer8_outputs(8442) <= not (a or b);
    layer8_outputs(8443) <= a;
    layer8_outputs(8444) <= not (a xor b);
    layer8_outputs(8445) <= not (a xor b);
    layer8_outputs(8446) <= not b;
    layer8_outputs(8447) <= a;
    layer8_outputs(8448) <= not (a or b);
    layer8_outputs(8449) <= b and not a;
    layer8_outputs(8450) <= b and not a;
    layer8_outputs(8451) <= 1'b1;
    layer8_outputs(8452) <= not (a xor b);
    layer8_outputs(8453) <= not b;
    layer8_outputs(8454) <= not (a and b);
    layer8_outputs(8455) <= not b;
    layer8_outputs(8456) <= b;
    layer8_outputs(8457) <= not a;
    layer8_outputs(8458) <= not (a and b);
    layer8_outputs(8459) <= not b;
    layer8_outputs(8460) <= b;
    layer8_outputs(8461) <= not (a or b);
    layer8_outputs(8462) <= not b;
    layer8_outputs(8463) <= 1'b1;
    layer8_outputs(8464) <= a xor b;
    layer8_outputs(8465) <= a;
    layer8_outputs(8466) <= not b or a;
    layer8_outputs(8467) <= not a or b;
    layer8_outputs(8468) <= a xor b;
    layer8_outputs(8469) <= not (a xor b);
    layer8_outputs(8470) <= not a;
    layer8_outputs(8471) <= a and b;
    layer8_outputs(8472) <= not b or a;
    layer8_outputs(8473) <= not a or b;
    layer8_outputs(8474) <= a xor b;
    layer8_outputs(8475) <= not a or b;
    layer8_outputs(8476) <= not a;
    layer8_outputs(8477) <= b and not a;
    layer8_outputs(8478) <= b and not a;
    layer8_outputs(8479) <= not (a xor b);
    layer8_outputs(8480) <= b;
    layer8_outputs(8481) <= a;
    layer8_outputs(8482) <= not a;
    layer8_outputs(8483) <= a xor b;
    layer8_outputs(8484) <= b;
    layer8_outputs(8485) <= b;
    layer8_outputs(8486) <= not (a xor b);
    layer8_outputs(8487) <= not (a or b);
    layer8_outputs(8488) <= a xor b;
    layer8_outputs(8489) <= not b;
    layer8_outputs(8490) <= a and b;
    layer8_outputs(8491) <= b;
    layer8_outputs(8492) <= b;
    layer8_outputs(8493) <= not (a or b);
    layer8_outputs(8494) <= b;
    layer8_outputs(8495) <= not a;
    layer8_outputs(8496) <= a;
    layer8_outputs(8497) <= not a or b;
    layer8_outputs(8498) <= not (a and b);
    layer8_outputs(8499) <= a or b;
    layer8_outputs(8500) <= a and b;
    layer8_outputs(8501) <= a and b;
    layer8_outputs(8502) <= not (a or b);
    layer8_outputs(8503) <= not a;
    layer8_outputs(8504) <= b;
    layer8_outputs(8505) <= not (a xor b);
    layer8_outputs(8506) <= a or b;
    layer8_outputs(8507) <= a;
    layer8_outputs(8508) <= not a;
    layer8_outputs(8509) <= not a;
    layer8_outputs(8510) <= not (a or b);
    layer8_outputs(8511) <= not (a xor b);
    layer8_outputs(8512) <= b;
    layer8_outputs(8513) <= not b;
    layer8_outputs(8514) <= b;
    layer8_outputs(8515) <= not a;
    layer8_outputs(8516) <= a;
    layer8_outputs(8517) <= 1'b0;
    layer8_outputs(8518) <= not a or b;
    layer8_outputs(8519) <= b;
    layer8_outputs(8520) <= b and not a;
    layer8_outputs(8521) <= a;
    layer8_outputs(8522) <= not (a xor b);
    layer8_outputs(8523) <= not (a and b);
    layer8_outputs(8524) <= a xor b;
    layer8_outputs(8525) <= not a;
    layer8_outputs(8526) <= a;
    layer8_outputs(8527) <= a xor b;
    layer8_outputs(8528) <= a xor b;
    layer8_outputs(8529) <= b and not a;
    layer8_outputs(8530) <= a;
    layer8_outputs(8531) <= a and b;
    layer8_outputs(8532) <= b and not a;
    layer8_outputs(8533) <= b;
    layer8_outputs(8534) <= b;
    layer8_outputs(8535) <= a xor b;
    layer8_outputs(8536) <= not a;
    layer8_outputs(8537) <= a and b;
    layer8_outputs(8538) <= a and b;
    layer8_outputs(8539) <= not a or b;
    layer8_outputs(8540) <= not b;
    layer8_outputs(8541) <= not b;
    layer8_outputs(8542) <= not (a or b);
    layer8_outputs(8543) <= not a or b;
    layer8_outputs(8544) <= a;
    layer8_outputs(8545) <= b;
    layer8_outputs(8546) <= not a;
    layer8_outputs(8547) <= not a;
    layer8_outputs(8548) <= a xor b;
    layer8_outputs(8549) <= a;
    layer8_outputs(8550) <= a;
    layer8_outputs(8551) <= not b;
    layer8_outputs(8552) <= not (a xor b);
    layer8_outputs(8553) <= 1'b0;
    layer8_outputs(8554) <= not (a and b);
    layer8_outputs(8555) <= not b or a;
    layer8_outputs(8556) <= a xor b;
    layer8_outputs(8557) <= a xor b;
    layer8_outputs(8558) <= not b;
    layer8_outputs(8559) <= a;
    layer8_outputs(8560) <= a;
    layer8_outputs(8561) <= not (a xor b);
    layer8_outputs(8562) <= not (a xor b);
    layer8_outputs(8563) <= not (a xor b);
    layer8_outputs(8564) <= 1'b1;
    layer8_outputs(8565) <= a xor b;
    layer8_outputs(8566) <= b;
    layer8_outputs(8567) <= not (a xor b);
    layer8_outputs(8568) <= a and not b;
    layer8_outputs(8569) <= b;
    layer8_outputs(8570) <= b;
    layer8_outputs(8571) <= b and not a;
    layer8_outputs(8572) <= not b;
    layer8_outputs(8573) <= not (a xor b);
    layer8_outputs(8574) <= b and not a;
    layer8_outputs(8575) <= not b;
    layer8_outputs(8576) <= not a;
    layer8_outputs(8577) <= not (a and b);
    layer8_outputs(8578) <= not (a and b);
    layer8_outputs(8579) <= a;
    layer8_outputs(8580) <= a xor b;
    layer8_outputs(8581) <= b;
    layer8_outputs(8582) <= not a or b;
    layer8_outputs(8583) <= not (a xor b);
    layer8_outputs(8584) <= b;
    layer8_outputs(8585) <= a xor b;
    layer8_outputs(8586) <= not a;
    layer8_outputs(8587) <= b and not a;
    layer8_outputs(8588) <= a xor b;
    layer8_outputs(8589) <= b;
    layer8_outputs(8590) <= a xor b;
    layer8_outputs(8591) <= not (a xor b);
    layer8_outputs(8592) <= b;
    layer8_outputs(8593) <= not (a and b);
    layer8_outputs(8594) <= a xor b;
    layer8_outputs(8595) <= a xor b;
    layer8_outputs(8596) <= not b or a;
    layer8_outputs(8597) <= not a;
    layer8_outputs(8598) <= not b;
    layer8_outputs(8599) <= not a or b;
    layer8_outputs(8600) <= b;
    layer8_outputs(8601) <= b and not a;
    layer8_outputs(8602) <= not a;
    layer8_outputs(8603) <= not a;
    layer8_outputs(8604) <= a xor b;
    layer8_outputs(8605) <= a xor b;
    layer8_outputs(8606) <= b;
    layer8_outputs(8607) <= a and b;
    layer8_outputs(8608) <= a xor b;
    layer8_outputs(8609) <= not b;
    layer8_outputs(8610) <= a or b;
    layer8_outputs(8611) <= a and not b;
    layer8_outputs(8612) <= a;
    layer8_outputs(8613) <= not (a xor b);
    layer8_outputs(8614) <= not (a or b);
    layer8_outputs(8615) <= b;
    layer8_outputs(8616) <= not (a xor b);
    layer8_outputs(8617) <= a;
    layer8_outputs(8618) <= a and not b;
    layer8_outputs(8619) <= not a;
    layer8_outputs(8620) <= not (a or b);
    layer8_outputs(8621) <= not b;
    layer8_outputs(8622) <= not (a or b);
    layer8_outputs(8623) <= a;
    layer8_outputs(8624) <= a xor b;
    layer8_outputs(8625) <= not b;
    layer8_outputs(8626) <= a;
    layer8_outputs(8627) <= a or b;
    layer8_outputs(8628) <= not a;
    layer8_outputs(8629) <= not b;
    layer8_outputs(8630) <= not a;
    layer8_outputs(8631) <= a;
    layer8_outputs(8632) <= not a or b;
    layer8_outputs(8633) <= 1'b0;
    layer8_outputs(8634) <= a;
    layer8_outputs(8635) <= a;
    layer8_outputs(8636) <= a;
    layer8_outputs(8637) <= not a;
    layer8_outputs(8638) <= not a;
    layer8_outputs(8639) <= not a;
    layer8_outputs(8640) <= a xor b;
    layer8_outputs(8641) <= not a;
    layer8_outputs(8642) <= a;
    layer8_outputs(8643) <= not b;
    layer8_outputs(8644) <= a and b;
    layer8_outputs(8645) <= not a or b;
    layer8_outputs(8646) <= not a or b;
    layer8_outputs(8647) <= a or b;
    layer8_outputs(8648) <= not b or a;
    layer8_outputs(8649) <= a;
    layer8_outputs(8650) <= a xor b;
    layer8_outputs(8651) <= a and b;
    layer8_outputs(8652) <= not a;
    layer8_outputs(8653) <= not a;
    layer8_outputs(8654) <= b;
    layer8_outputs(8655) <= not a or b;
    layer8_outputs(8656) <= not (a xor b);
    layer8_outputs(8657) <= a;
    layer8_outputs(8658) <= not (a and b);
    layer8_outputs(8659) <= b;
    layer8_outputs(8660) <= not a;
    layer8_outputs(8661) <= b;
    layer8_outputs(8662) <= not a;
    layer8_outputs(8663) <= not a;
    layer8_outputs(8664) <= not a;
    layer8_outputs(8665) <= b and not a;
    layer8_outputs(8666) <= not b;
    layer8_outputs(8667) <= not a;
    layer8_outputs(8668) <= not (a xor b);
    layer8_outputs(8669) <= b;
    layer8_outputs(8670) <= a and b;
    layer8_outputs(8671) <= not a or b;
    layer8_outputs(8672) <= a and b;
    layer8_outputs(8673) <= not a;
    layer8_outputs(8674) <= a;
    layer8_outputs(8675) <= not a or b;
    layer8_outputs(8676) <= b;
    layer8_outputs(8677) <= not b;
    layer8_outputs(8678) <= not (a or b);
    layer8_outputs(8679) <= not (a or b);
    layer8_outputs(8680) <= not a;
    layer8_outputs(8681) <= a and b;
    layer8_outputs(8682) <= a;
    layer8_outputs(8683) <= a and b;
    layer8_outputs(8684) <= not (a or b);
    layer8_outputs(8685) <= not b;
    layer8_outputs(8686) <= not a or b;
    layer8_outputs(8687) <= not (a xor b);
    layer8_outputs(8688) <= not a;
    layer8_outputs(8689) <= not (a xor b);
    layer8_outputs(8690) <= a;
    layer8_outputs(8691) <= not (a or b);
    layer8_outputs(8692) <= not b or a;
    layer8_outputs(8693) <= a;
    layer8_outputs(8694) <= b;
    layer8_outputs(8695) <= a xor b;
    layer8_outputs(8696) <= not a;
    layer8_outputs(8697) <= b;
    layer8_outputs(8698) <= not b or a;
    layer8_outputs(8699) <= b;
    layer8_outputs(8700) <= not (a xor b);
    layer8_outputs(8701) <= not a;
    layer8_outputs(8702) <= not b;
    layer8_outputs(8703) <= not a;
    layer8_outputs(8704) <= not (a or b);
    layer8_outputs(8705) <= not (a or b);
    layer8_outputs(8706) <= a or b;
    layer8_outputs(8707) <= not b;
    layer8_outputs(8708) <= a;
    layer8_outputs(8709) <= not (a xor b);
    layer8_outputs(8710) <= b and not a;
    layer8_outputs(8711) <= b and not a;
    layer8_outputs(8712) <= not (a or b);
    layer8_outputs(8713) <= not b;
    layer8_outputs(8714) <= a and b;
    layer8_outputs(8715) <= a;
    layer8_outputs(8716) <= a xor b;
    layer8_outputs(8717) <= b;
    layer8_outputs(8718) <= a or b;
    layer8_outputs(8719) <= b;
    layer8_outputs(8720) <= not (a xor b);
    layer8_outputs(8721) <= not a;
    layer8_outputs(8722) <= not (a or b);
    layer8_outputs(8723) <= not b;
    layer8_outputs(8724) <= a and not b;
    layer8_outputs(8725) <= not a;
    layer8_outputs(8726) <= b and not a;
    layer8_outputs(8727) <= b;
    layer8_outputs(8728) <= a and not b;
    layer8_outputs(8729) <= a;
    layer8_outputs(8730) <= not b;
    layer8_outputs(8731) <= not a or b;
    layer8_outputs(8732) <= b;
    layer8_outputs(8733) <= a xor b;
    layer8_outputs(8734) <= a or b;
    layer8_outputs(8735) <= a and not b;
    layer8_outputs(8736) <= not a;
    layer8_outputs(8737) <= not a;
    layer8_outputs(8738) <= b;
    layer8_outputs(8739) <= not (a and b);
    layer8_outputs(8740) <= a and not b;
    layer8_outputs(8741) <= not b;
    layer8_outputs(8742) <= not a;
    layer8_outputs(8743) <= b and not a;
    layer8_outputs(8744) <= not a;
    layer8_outputs(8745) <= not (a and b);
    layer8_outputs(8746) <= a and not b;
    layer8_outputs(8747) <= not a;
    layer8_outputs(8748) <= not a;
    layer8_outputs(8749) <= a xor b;
    layer8_outputs(8750) <= not (a xor b);
    layer8_outputs(8751) <= not (a and b);
    layer8_outputs(8752) <= a xor b;
    layer8_outputs(8753) <= a and b;
    layer8_outputs(8754) <= b;
    layer8_outputs(8755) <= not a;
    layer8_outputs(8756) <= a and not b;
    layer8_outputs(8757) <= not (a or b);
    layer8_outputs(8758) <= not a or b;
    layer8_outputs(8759) <= not b;
    layer8_outputs(8760) <= a;
    layer8_outputs(8761) <= a;
    layer8_outputs(8762) <= b;
    layer8_outputs(8763) <= not a or b;
    layer8_outputs(8764) <= not b;
    layer8_outputs(8765) <= a xor b;
    layer8_outputs(8766) <= not a;
    layer8_outputs(8767) <= a xor b;
    layer8_outputs(8768) <= not a;
    layer8_outputs(8769) <= a xor b;
    layer8_outputs(8770) <= 1'b1;
    layer8_outputs(8771) <= not a;
    layer8_outputs(8772) <= a and not b;
    layer8_outputs(8773) <= not b or a;
    layer8_outputs(8774) <= b;
    layer8_outputs(8775) <= not a or b;
    layer8_outputs(8776) <= b;
    layer8_outputs(8777) <= not a;
    layer8_outputs(8778) <= a xor b;
    layer8_outputs(8779) <= not b or a;
    layer8_outputs(8780) <= not (a and b);
    layer8_outputs(8781) <= not (a xor b);
    layer8_outputs(8782) <= not b or a;
    layer8_outputs(8783) <= b;
    layer8_outputs(8784) <= not b;
    layer8_outputs(8785) <= a;
    layer8_outputs(8786) <= a and b;
    layer8_outputs(8787) <= not b;
    layer8_outputs(8788) <= 1'b0;
    layer8_outputs(8789) <= not a;
    layer8_outputs(8790) <= a and not b;
    layer8_outputs(8791) <= b;
    layer8_outputs(8792) <= not a;
    layer8_outputs(8793) <= b;
    layer8_outputs(8794) <= not b;
    layer8_outputs(8795) <= not (a xor b);
    layer8_outputs(8796) <= a xor b;
    layer8_outputs(8797) <= b and not a;
    layer8_outputs(8798) <= a;
    layer8_outputs(8799) <= not a;
    layer8_outputs(8800) <= not (a and b);
    layer8_outputs(8801) <= a xor b;
    layer8_outputs(8802) <= a xor b;
    layer8_outputs(8803) <= not a;
    layer8_outputs(8804) <= a and not b;
    layer8_outputs(8805) <= not b;
    layer8_outputs(8806) <= not (a xor b);
    layer8_outputs(8807) <= a;
    layer8_outputs(8808) <= not (a and b);
    layer8_outputs(8809) <= a xor b;
    layer8_outputs(8810) <= b;
    layer8_outputs(8811) <= not b;
    layer8_outputs(8812) <= not b;
    layer8_outputs(8813) <= a;
    layer8_outputs(8814) <= not a;
    layer8_outputs(8815) <= a;
    layer8_outputs(8816) <= not a;
    layer8_outputs(8817) <= b and not a;
    layer8_outputs(8818) <= not b;
    layer8_outputs(8819) <= not b;
    layer8_outputs(8820) <= b;
    layer8_outputs(8821) <= a;
    layer8_outputs(8822) <= not b;
    layer8_outputs(8823) <= not b or a;
    layer8_outputs(8824) <= a xor b;
    layer8_outputs(8825) <= 1'b0;
    layer8_outputs(8826) <= b;
    layer8_outputs(8827) <= not b;
    layer8_outputs(8828) <= not (a and b);
    layer8_outputs(8829) <= a or b;
    layer8_outputs(8830) <= not a;
    layer8_outputs(8831) <= not a;
    layer8_outputs(8832) <= not (a xor b);
    layer8_outputs(8833) <= a;
    layer8_outputs(8834) <= a and not b;
    layer8_outputs(8835) <= a xor b;
    layer8_outputs(8836) <= not (a xor b);
    layer8_outputs(8837) <= a;
    layer8_outputs(8838) <= b and not a;
    layer8_outputs(8839) <= b;
    layer8_outputs(8840) <= not (a and b);
    layer8_outputs(8841) <= not (a xor b);
    layer8_outputs(8842) <= a and not b;
    layer8_outputs(8843) <= not (a or b);
    layer8_outputs(8844) <= not a;
    layer8_outputs(8845) <= a;
    layer8_outputs(8846) <= not (a xor b);
    layer8_outputs(8847) <= not b;
    layer8_outputs(8848) <= a;
    layer8_outputs(8849) <= not a;
    layer8_outputs(8850) <= a;
    layer8_outputs(8851) <= not a;
    layer8_outputs(8852) <= not a or b;
    layer8_outputs(8853) <= not b or a;
    layer8_outputs(8854) <= a xor b;
    layer8_outputs(8855) <= not b;
    layer8_outputs(8856) <= a;
    layer8_outputs(8857) <= a or b;
    layer8_outputs(8858) <= b;
    layer8_outputs(8859) <= a;
    layer8_outputs(8860) <= not (a xor b);
    layer8_outputs(8861) <= not (a xor b);
    layer8_outputs(8862) <= not (a or b);
    layer8_outputs(8863) <= not a;
    layer8_outputs(8864) <= not a;
    layer8_outputs(8865) <= not (a or b);
    layer8_outputs(8866) <= not (a and b);
    layer8_outputs(8867) <= b;
    layer8_outputs(8868) <= b and not a;
    layer8_outputs(8869) <= b;
    layer8_outputs(8870) <= a xor b;
    layer8_outputs(8871) <= a;
    layer8_outputs(8872) <= not b;
    layer8_outputs(8873) <= not b;
    layer8_outputs(8874) <= b;
    layer8_outputs(8875) <= not a;
    layer8_outputs(8876) <= not b or a;
    layer8_outputs(8877) <= a xor b;
    layer8_outputs(8878) <= not (a and b);
    layer8_outputs(8879) <= not (a xor b);
    layer8_outputs(8880) <= b and not a;
    layer8_outputs(8881) <= b and not a;
    layer8_outputs(8882) <= a xor b;
    layer8_outputs(8883) <= a and not b;
    layer8_outputs(8884) <= not a or b;
    layer8_outputs(8885) <= not b;
    layer8_outputs(8886) <= a or b;
    layer8_outputs(8887) <= a;
    layer8_outputs(8888) <= a or b;
    layer8_outputs(8889) <= not b or a;
    layer8_outputs(8890) <= not b;
    layer8_outputs(8891) <= not a or b;
    layer8_outputs(8892) <= not b;
    layer8_outputs(8893) <= a and not b;
    layer8_outputs(8894) <= b;
    layer8_outputs(8895) <= not (a xor b);
    layer8_outputs(8896) <= not a;
    layer8_outputs(8897) <= b;
    layer8_outputs(8898) <= not (a xor b);
    layer8_outputs(8899) <= not b;
    layer8_outputs(8900) <= a xor b;
    layer8_outputs(8901) <= not (a and b);
    layer8_outputs(8902) <= not (a xor b);
    layer8_outputs(8903) <= a xor b;
    layer8_outputs(8904) <= a or b;
    layer8_outputs(8905) <= a and b;
    layer8_outputs(8906) <= a;
    layer8_outputs(8907) <= b;
    layer8_outputs(8908) <= a xor b;
    layer8_outputs(8909) <= a and b;
    layer8_outputs(8910) <= a and b;
    layer8_outputs(8911) <= not a;
    layer8_outputs(8912) <= b;
    layer8_outputs(8913) <= not a;
    layer8_outputs(8914) <= b;
    layer8_outputs(8915) <= not (a xor b);
    layer8_outputs(8916) <= not (a xor b);
    layer8_outputs(8917) <= b;
    layer8_outputs(8918) <= not a;
    layer8_outputs(8919) <= not a;
    layer8_outputs(8920) <= not (a xor b);
    layer8_outputs(8921) <= a or b;
    layer8_outputs(8922) <= a and not b;
    layer8_outputs(8923) <= a xor b;
    layer8_outputs(8924) <= not a;
    layer8_outputs(8925) <= not b or a;
    layer8_outputs(8926) <= b;
    layer8_outputs(8927) <= not (a or b);
    layer8_outputs(8928) <= a and b;
    layer8_outputs(8929) <= a xor b;
    layer8_outputs(8930) <= a;
    layer8_outputs(8931) <= not a;
    layer8_outputs(8932) <= not (a xor b);
    layer8_outputs(8933) <= b;
    layer8_outputs(8934) <= not (a and b);
    layer8_outputs(8935) <= not a or b;
    layer8_outputs(8936) <= a;
    layer8_outputs(8937) <= a xor b;
    layer8_outputs(8938) <= not b or a;
    layer8_outputs(8939) <= not a;
    layer8_outputs(8940) <= not (a and b);
    layer8_outputs(8941) <= not a;
    layer8_outputs(8942) <= a and not b;
    layer8_outputs(8943) <= not a;
    layer8_outputs(8944) <= not a;
    layer8_outputs(8945) <= not (a and b);
    layer8_outputs(8946) <= a;
    layer8_outputs(8947) <= not a;
    layer8_outputs(8948) <= b;
    layer8_outputs(8949) <= b;
    layer8_outputs(8950) <= a;
    layer8_outputs(8951) <= a;
    layer8_outputs(8952) <= not (a xor b);
    layer8_outputs(8953) <= not b;
    layer8_outputs(8954) <= a;
    layer8_outputs(8955) <= b;
    layer8_outputs(8956) <= a;
    layer8_outputs(8957) <= a or b;
    layer8_outputs(8958) <= not (a xor b);
    layer8_outputs(8959) <= a and not b;
    layer8_outputs(8960) <= not (a xor b);
    layer8_outputs(8961) <= not (a xor b);
    layer8_outputs(8962) <= not a or b;
    layer8_outputs(8963) <= a;
    layer8_outputs(8964) <= not b;
    layer8_outputs(8965) <= not a;
    layer8_outputs(8966) <= not a;
    layer8_outputs(8967) <= b and not a;
    layer8_outputs(8968) <= not a;
    layer8_outputs(8969) <= a or b;
    layer8_outputs(8970) <= not b;
    layer8_outputs(8971) <= not a;
    layer8_outputs(8972) <= not a or b;
    layer8_outputs(8973) <= b;
    layer8_outputs(8974) <= a xor b;
    layer8_outputs(8975) <= not a;
    layer8_outputs(8976) <= a and not b;
    layer8_outputs(8977) <= b;
    layer8_outputs(8978) <= not a;
    layer8_outputs(8979) <= b;
    layer8_outputs(8980) <= b;
    layer8_outputs(8981) <= a xor b;
    layer8_outputs(8982) <= not a or b;
    layer8_outputs(8983) <= a;
    layer8_outputs(8984) <= not a;
    layer8_outputs(8985) <= b;
    layer8_outputs(8986) <= not b or a;
    layer8_outputs(8987) <= not (a xor b);
    layer8_outputs(8988) <= not a or b;
    layer8_outputs(8989) <= a;
    layer8_outputs(8990) <= not a;
    layer8_outputs(8991) <= b;
    layer8_outputs(8992) <= b and not a;
    layer8_outputs(8993) <= a;
    layer8_outputs(8994) <= a and not b;
    layer8_outputs(8995) <= a;
    layer8_outputs(8996) <= b;
    layer8_outputs(8997) <= not a;
    layer8_outputs(8998) <= not a;
    layer8_outputs(8999) <= not (a xor b);
    layer8_outputs(9000) <= 1'b0;
    layer8_outputs(9001) <= not b or a;
    layer8_outputs(9002) <= not (a xor b);
    layer8_outputs(9003) <= not a;
    layer8_outputs(9004) <= not (a xor b);
    layer8_outputs(9005) <= not a or b;
    layer8_outputs(9006) <= not (a or b);
    layer8_outputs(9007) <= b;
    layer8_outputs(9008) <= a xor b;
    layer8_outputs(9009) <= a xor b;
    layer8_outputs(9010) <= b and not a;
    layer8_outputs(9011) <= not (a xor b);
    layer8_outputs(9012) <= not (a or b);
    layer8_outputs(9013) <= 1'b0;
    layer8_outputs(9014) <= not a;
    layer8_outputs(9015) <= not a or b;
    layer8_outputs(9016) <= b and not a;
    layer8_outputs(9017) <= not b;
    layer8_outputs(9018) <= a;
    layer8_outputs(9019) <= not a;
    layer8_outputs(9020) <= not (a xor b);
    layer8_outputs(9021) <= a or b;
    layer8_outputs(9022) <= b;
    layer8_outputs(9023) <= not a;
    layer8_outputs(9024) <= not b or a;
    layer8_outputs(9025) <= not b or a;
    layer8_outputs(9026) <= a and not b;
    layer8_outputs(9027) <= not b or a;
    layer8_outputs(9028) <= a xor b;
    layer8_outputs(9029) <= b;
    layer8_outputs(9030) <= not (a xor b);
    layer8_outputs(9031) <= a and b;
    layer8_outputs(9032) <= a xor b;
    layer8_outputs(9033) <= not b;
    layer8_outputs(9034) <= not a;
    layer8_outputs(9035) <= a xor b;
    layer8_outputs(9036) <= not b;
    layer8_outputs(9037) <= not (a xor b);
    layer8_outputs(9038) <= a;
    layer8_outputs(9039) <= not b;
    layer8_outputs(9040) <= a;
    layer8_outputs(9041) <= not (a xor b);
    layer8_outputs(9042) <= not b or a;
    layer8_outputs(9043) <= a;
    layer8_outputs(9044) <= a or b;
    layer8_outputs(9045) <= b;
    layer8_outputs(9046) <= a;
    layer8_outputs(9047) <= a and b;
    layer8_outputs(9048) <= 1'b0;
    layer8_outputs(9049) <= b and not a;
    layer8_outputs(9050) <= a xor b;
    layer8_outputs(9051) <= not a;
    layer8_outputs(9052) <= not b or a;
    layer8_outputs(9053) <= not (a and b);
    layer8_outputs(9054) <= b;
    layer8_outputs(9055) <= not a;
    layer8_outputs(9056) <= not a;
    layer8_outputs(9057) <= b;
    layer8_outputs(9058) <= b;
    layer8_outputs(9059) <= a and b;
    layer8_outputs(9060) <= a and not b;
    layer8_outputs(9061) <= b;
    layer8_outputs(9062) <= not a;
    layer8_outputs(9063) <= b;
    layer8_outputs(9064) <= a;
    layer8_outputs(9065) <= a;
    layer8_outputs(9066) <= a xor b;
    layer8_outputs(9067) <= not b or a;
    layer8_outputs(9068) <= not (a xor b);
    layer8_outputs(9069) <= not (a xor b);
    layer8_outputs(9070) <= not a or b;
    layer8_outputs(9071) <= not (a xor b);
    layer8_outputs(9072) <= not (a or b);
    layer8_outputs(9073) <= not b;
    layer8_outputs(9074) <= not (a xor b);
    layer8_outputs(9075) <= a or b;
    layer8_outputs(9076) <= not (a and b);
    layer8_outputs(9077) <= not a;
    layer8_outputs(9078) <= b and not a;
    layer8_outputs(9079) <= not b or a;
    layer8_outputs(9080) <= a;
    layer8_outputs(9081) <= not (a or b);
    layer8_outputs(9082) <= b;
    layer8_outputs(9083) <= not a;
    layer8_outputs(9084) <= not b or a;
    layer8_outputs(9085) <= a and not b;
    layer8_outputs(9086) <= not (a and b);
    layer8_outputs(9087) <= a and b;
    layer8_outputs(9088) <= b and not a;
    layer8_outputs(9089) <= not b or a;
    layer8_outputs(9090) <= b;
    layer8_outputs(9091) <= a xor b;
    layer8_outputs(9092) <= not (a or b);
    layer8_outputs(9093) <= not a;
    layer8_outputs(9094) <= a;
    layer8_outputs(9095) <= a xor b;
    layer8_outputs(9096) <= not b;
    layer8_outputs(9097) <= not b;
    layer8_outputs(9098) <= b and not a;
    layer8_outputs(9099) <= not (a xor b);
    layer8_outputs(9100) <= a or b;
    layer8_outputs(9101) <= not b;
    layer8_outputs(9102) <= a xor b;
    layer8_outputs(9103) <= a or b;
    layer8_outputs(9104) <= not a;
    layer8_outputs(9105) <= b;
    layer8_outputs(9106) <= b;
    layer8_outputs(9107) <= a;
    layer8_outputs(9108) <= a or b;
    layer8_outputs(9109) <= a or b;
    layer8_outputs(9110) <= not a;
    layer8_outputs(9111) <= b and not a;
    layer8_outputs(9112) <= a xor b;
    layer8_outputs(9113) <= not a;
    layer8_outputs(9114) <= a or b;
    layer8_outputs(9115) <= not (a xor b);
    layer8_outputs(9116) <= a or b;
    layer8_outputs(9117) <= b;
    layer8_outputs(9118) <= a xor b;
    layer8_outputs(9119) <= b and not a;
    layer8_outputs(9120) <= a;
    layer8_outputs(9121) <= a xor b;
    layer8_outputs(9122) <= not a;
    layer8_outputs(9123) <= b;
    layer8_outputs(9124) <= not b;
    layer8_outputs(9125) <= not b;
    layer8_outputs(9126) <= not b;
    layer8_outputs(9127) <= a xor b;
    layer8_outputs(9128) <= not (a xor b);
    layer8_outputs(9129) <= a and not b;
    layer8_outputs(9130) <= b and not a;
    layer8_outputs(9131) <= a;
    layer8_outputs(9132) <= b;
    layer8_outputs(9133) <= not (a or b);
    layer8_outputs(9134) <= a;
    layer8_outputs(9135) <= not a;
    layer8_outputs(9136) <= a or b;
    layer8_outputs(9137) <= not a;
    layer8_outputs(9138) <= a;
    layer8_outputs(9139) <= a xor b;
    layer8_outputs(9140) <= a and not b;
    layer8_outputs(9141) <= not (a xor b);
    layer8_outputs(9142) <= not (a xor b);
    layer8_outputs(9143) <= not a;
    layer8_outputs(9144) <= b;
    layer8_outputs(9145) <= b;
    layer8_outputs(9146) <= a;
    layer8_outputs(9147) <= b;
    layer8_outputs(9148) <= 1'b1;
    layer8_outputs(9149) <= a xor b;
    layer8_outputs(9150) <= not a or b;
    layer8_outputs(9151) <= a xor b;
    layer8_outputs(9152) <= not a or b;
    layer8_outputs(9153) <= b;
    layer8_outputs(9154) <= a xor b;
    layer8_outputs(9155) <= not (a xor b);
    layer8_outputs(9156) <= b;
    layer8_outputs(9157) <= b;
    layer8_outputs(9158) <= a xor b;
    layer8_outputs(9159) <= b;
    layer8_outputs(9160) <= a;
    layer8_outputs(9161) <= not (a xor b);
    layer8_outputs(9162) <= not (a and b);
    layer8_outputs(9163) <= b;
    layer8_outputs(9164) <= a and not b;
    layer8_outputs(9165) <= b and not a;
    layer8_outputs(9166) <= not a;
    layer8_outputs(9167) <= a xor b;
    layer8_outputs(9168) <= not a;
    layer8_outputs(9169) <= a or b;
    layer8_outputs(9170) <= b and not a;
    layer8_outputs(9171) <= b;
    layer8_outputs(9172) <= not a or b;
    layer8_outputs(9173) <= not a or b;
    layer8_outputs(9174) <= a or b;
    layer8_outputs(9175) <= not (a xor b);
    layer8_outputs(9176) <= not b or a;
    layer8_outputs(9177) <= a;
    layer8_outputs(9178) <= not b or a;
    layer8_outputs(9179) <= not a;
    layer8_outputs(9180) <= not a;
    layer8_outputs(9181) <= a or b;
    layer8_outputs(9182) <= a and b;
    layer8_outputs(9183) <= not b;
    layer8_outputs(9184) <= not b;
    layer8_outputs(9185) <= not b;
    layer8_outputs(9186) <= b;
    layer8_outputs(9187) <= not a;
    layer8_outputs(9188) <= b;
    layer8_outputs(9189) <= not (a xor b);
    layer8_outputs(9190) <= a;
    layer8_outputs(9191) <= not (a xor b);
    layer8_outputs(9192) <= not b;
    layer8_outputs(9193) <= a;
    layer8_outputs(9194) <= b;
    layer8_outputs(9195) <= b;
    layer8_outputs(9196) <= not b;
    layer8_outputs(9197) <= not b or a;
    layer8_outputs(9198) <= not b;
    layer8_outputs(9199) <= not a;
    layer8_outputs(9200) <= not (a xor b);
    layer8_outputs(9201) <= b;
    layer8_outputs(9202) <= a;
    layer8_outputs(9203) <= not a;
    layer8_outputs(9204) <= a;
    layer8_outputs(9205) <= not (a or b);
    layer8_outputs(9206) <= not b;
    layer8_outputs(9207) <= a and b;
    layer8_outputs(9208) <= not a;
    layer8_outputs(9209) <= a xor b;
    layer8_outputs(9210) <= not (a and b);
    layer8_outputs(9211) <= a xor b;
    layer8_outputs(9212) <= b;
    layer8_outputs(9213) <= not (a xor b);
    layer8_outputs(9214) <= not (a xor b);
    layer8_outputs(9215) <= not a;
    layer8_outputs(9216) <= a;
    layer8_outputs(9217) <= not (a and b);
    layer8_outputs(9218) <= not a;
    layer8_outputs(9219) <= not a;
    layer8_outputs(9220) <= b;
    layer8_outputs(9221) <= not a;
    layer8_outputs(9222) <= a xor b;
    layer8_outputs(9223) <= not a;
    layer8_outputs(9224) <= a and not b;
    layer8_outputs(9225) <= not (a or b);
    layer8_outputs(9226) <= b;
    layer8_outputs(9227) <= a xor b;
    layer8_outputs(9228) <= not (a xor b);
    layer8_outputs(9229) <= not a;
    layer8_outputs(9230) <= b;
    layer8_outputs(9231) <= not (a and b);
    layer8_outputs(9232) <= b and not a;
    layer8_outputs(9233) <= not a;
    layer8_outputs(9234) <= not a or b;
    layer8_outputs(9235) <= not b or a;
    layer8_outputs(9236) <= a or b;
    layer8_outputs(9237) <= not b;
    layer8_outputs(9238) <= a and not b;
    layer8_outputs(9239) <= not a;
    layer8_outputs(9240) <= a and not b;
    layer8_outputs(9241) <= not (a xor b);
    layer8_outputs(9242) <= not (a and b);
    layer8_outputs(9243) <= b;
    layer8_outputs(9244) <= not b;
    layer8_outputs(9245) <= not a;
    layer8_outputs(9246) <= b;
    layer8_outputs(9247) <= a or b;
    layer8_outputs(9248) <= a or b;
    layer8_outputs(9249) <= a;
    layer8_outputs(9250) <= a xor b;
    layer8_outputs(9251) <= not (a xor b);
    layer8_outputs(9252) <= a and b;
    layer8_outputs(9253) <= not (a xor b);
    layer8_outputs(9254) <= not b;
    layer8_outputs(9255) <= not a;
    layer8_outputs(9256) <= a;
    layer8_outputs(9257) <= b;
    layer8_outputs(9258) <= a;
    layer8_outputs(9259) <= a or b;
    layer8_outputs(9260) <= b;
    layer8_outputs(9261) <= b;
    layer8_outputs(9262) <= b and not a;
    layer8_outputs(9263) <= b;
    layer8_outputs(9264) <= not b;
    layer8_outputs(9265) <= b and not a;
    layer8_outputs(9266) <= a or b;
    layer8_outputs(9267) <= b and not a;
    layer8_outputs(9268) <= a and b;
    layer8_outputs(9269) <= not b;
    layer8_outputs(9270) <= a xor b;
    layer8_outputs(9271) <= a;
    layer8_outputs(9272) <= not a;
    layer8_outputs(9273) <= not b;
    layer8_outputs(9274) <= not (a xor b);
    layer8_outputs(9275) <= not (a and b);
    layer8_outputs(9276) <= a and b;
    layer8_outputs(9277) <= not (a xor b);
    layer8_outputs(9278) <= b;
    layer8_outputs(9279) <= a or b;
    layer8_outputs(9280) <= not b;
    layer8_outputs(9281) <= not (a xor b);
    layer8_outputs(9282) <= a;
    layer8_outputs(9283) <= a xor b;
    layer8_outputs(9284) <= a and b;
    layer8_outputs(9285) <= a;
    layer8_outputs(9286) <= not b or a;
    layer8_outputs(9287) <= not a;
    layer8_outputs(9288) <= not b or a;
    layer8_outputs(9289) <= not a;
    layer8_outputs(9290) <= a xor b;
    layer8_outputs(9291) <= not (a xor b);
    layer8_outputs(9292) <= a and not b;
    layer8_outputs(9293) <= b and not a;
    layer8_outputs(9294) <= a;
    layer8_outputs(9295) <= a;
    layer8_outputs(9296) <= not a;
    layer8_outputs(9297) <= not a;
    layer8_outputs(9298) <= not b or a;
    layer8_outputs(9299) <= a or b;
    layer8_outputs(9300) <= b;
    layer8_outputs(9301) <= a xor b;
    layer8_outputs(9302) <= a or b;
    layer8_outputs(9303) <= not b;
    layer8_outputs(9304) <= b;
    layer8_outputs(9305) <= a xor b;
    layer8_outputs(9306) <= not (a xor b);
    layer8_outputs(9307) <= a;
    layer8_outputs(9308) <= b and not a;
    layer8_outputs(9309) <= a;
    layer8_outputs(9310) <= not (a xor b);
    layer8_outputs(9311) <= not b or a;
    layer8_outputs(9312) <= not a or b;
    layer8_outputs(9313) <= not b;
    layer8_outputs(9314) <= a;
    layer8_outputs(9315) <= not a;
    layer8_outputs(9316) <= a;
    layer8_outputs(9317) <= not a;
    layer8_outputs(9318) <= not a;
    layer8_outputs(9319) <= a xor b;
    layer8_outputs(9320) <= a xor b;
    layer8_outputs(9321) <= not b;
    layer8_outputs(9322) <= a and not b;
    layer8_outputs(9323) <= not (a and b);
    layer8_outputs(9324) <= not (a xor b);
    layer8_outputs(9325) <= not a;
    layer8_outputs(9326) <= b;
    layer8_outputs(9327) <= a and not b;
    layer8_outputs(9328) <= a or b;
    layer8_outputs(9329) <= a xor b;
    layer8_outputs(9330) <= a xor b;
    layer8_outputs(9331) <= not a;
    layer8_outputs(9332) <= a;
    layer8_outputs(9333) <= not b or a;
    layer8_outputs(9334) <= a xor b;
    layer8_outputs(9335) <= not b;
    layer8_outputs(9336) <= not a;
    layer8_outputs(9337) <= not b;
    layer8_outputs(9338) <= a;
    layer8_outputs(9339) <= not b;
    layer8_outputs(9340) <= not (a or b);
    layer8_outputs(9341) <= not a or b;
    layer8_outputs(9342) <= a;
    layer8_outputs(9343) <= b;
    layer8_outputs(9344) <= not a;
    layer8_outputs(9345) <= not a;
    layer8_outputs(9346) <= not (a and b);
    layer8_outputs(9347) <= not a;
    layer8_outputs(9348) <= not (a xor b);
    layer8_outputs(9349) <= not (a xor b);
    layer8_outputs(9350) <= a or b;
    layer8_outputs(9351) <= not a;
    layer8_outputs(9352) <= a or b;
    layer8_outputs(9353) <= b;
    layer8_outputs(9354) <= 1'b0;
    layer8_outputs(9355) <= not (a xor b);
    layer8_outputs(9356) <= not b;
    layer8_outputs(9357) <= not (a or b);
    layer8_outputs(9358) <= a and not b;
    layer8_outputs(9359) <= not (a xor b);
    layer8_outputs(9360) <= a;
    layer8_outputs(9361) <= not (a xor b);
    layer8_outputs(9362) <= b and not a;
    layer8_outputs(9363) <= b;
    layer8_outputs(9364) <= not b;
    layer8_outputs(9365) <= not b;
    layer8_outputs(9366) <= not (a and b);
    layer8_outputs(9367) <= not (a xor b);
    layer8_outputs(9368) <= 1'b1;
    layer8_outputs(9369) <= not (a xor b);
    layer8_outputs(9370) <= not (a xor b);
    layer8_outputs(9371) <= a xor b;
    layer8_outputs(9372) <= not b or a;
    layer8_outputs(9373) <= not a;
    layer8_outputs(9374) <= a and not b;
    layer8_outputs(9375) <= a xor b;
    layer8_outputs(9376) <= not (a and b);
    layer8_outputs(9377) <= not a;
    layer8_outputs(9378) <= b and not a;
    layer8_outputs(9379) <= not (a xor b);
    layer8_outputs(9380) <= a or b;
    layer8_outputs(9381) <= b and not a;
    layer8_outputs(9382) <= not (a xor b);
    layer8_outputs(9383) <= not b;
    layer8_outputs(9384) <= not b or a;
    layer8_outputs(9385) <= not b;
    layer8_outputs(9386) <= not a;
    layer8_outputs(9387) <= not (a and b);
    layer8_outputs(9388) <= b;
    layer8_outputs(9389) <= b;
    layer8_outputs(9390) <= a;
    layer8_outputs(9391) <= a xor b;
    layer8_outputs(9392) <= a xor b;
    layer8_outputs(9393) <= a xor b;
    layer8_outputs(9394) <= not b;
    layer8_outputs(9395) <= a xor b;
    layer8_outputs(9396) <= b;
    layer8_outputs(9397) <= not (a xor b);
    layer8_outputs(9398) <= not (a xor b);
    layer8_outputs(9399) <= a xor b;
    layer8_outputs(9400) <= not a;
    layer8_outputs(9401) <= not b;
    layer8_outputs(9402) <= not b or a;
    layer8_outputs(9403) <= b;
    layer8_outputs(9404) <= not b;
    layer8_outputs(9405) <= not b or a;
    layer8_outputs(9406) <= not (a and b);
    layer8_outputs(9407) <= not (a and b);
    layer8_outputs(9408) <= not b;
    layer8_outputs(9409) <= not a;
    layer8_outputs(9410) <= 1'b0;
    layer8_outputs(9411) <= b;
    layer8_outputs(9412) <= b;
    layer8_outputs(9413) <= a and not b;
    layer8_outputs(9414) <= not (a and b);
    layer8_outputs(9415) <= not b;
    layer8_outputs(9416) <= a or b;
    layer8_outputs(9417) <= a and b;
    layer8_outputs(9418) <= a xor b;
    layer8_outputs(9419) <= not a;
    layer8_outputs(9420) <= not (a and b);
    layer8_outputs(9421) <= not (a or b);
    layer8_outputs(9422) <= not a;
    layer8_outputs(9423) <= not a;
    layer8_outputs(9424) <= not a;
    layer8_outputs(9425) <= not a or b;
    layer8_outputs(9426) <= a or b;
    layer8_outputs(9427) <= not b;
    layer8_outputs(9428) <= not b or a;
    layer8_outputs(9429) <= not a;
    layer8_outputs(9430) <= not (a xor b);
    layer8_outputs(9431) <= not (a or b);
    layer8_outputs(9432) <= b;
    layer8_outputs(9433) <= a or b;
    layer8_outputs(9434) <= b and not a;
    layer8_outputs(9435) <= b;
    layer8_outputs(9436) <= not b;
    layer8_outputs(9437) <= a;
    layer8_outputs(9438) <= not (a xor b);
    layer8_outputs(9439) <= not a;
    layer8_outputs(9440) <= a;
    layer8_outputs(9441) <= not (a and b);
    layer8_outputs(9442) <= not (a or b);
    layer8_outputs(9443) <= a xor b;
    layer8_outputs(9444) <= not a or b;
    layer8_outputs(9445) <= a xor b;
    layer8_outputs(9446) <= b;
    layer8_outputs(9447) <= 1'b1;
    layer8_outputs(9448) <= a and b;
    layer8_outputs(9449) <= a and b;
    layer8_outputs(9450) <= not (a xor b);
    layer8_outputs(9451) <= not a;
    layer8_outputs(9452) <= b;
    layer8_outputs(9453) <= not (a xor b);
    layer8_outputs(9454) <= not (a or b);
    layer8_outputs(9455) <= b and not a;
    layer8_outputs(9456) <= not a;
    layer8_outputs(9457) <= b and not a;
    layer8_outputs(9458) <= not b;
    layer8_outputs(9459) <= not a;
    layer8_outputs(9460) <= not (a xor b);
    layer8_outputs(9461) <= a xor b;
    layer8_outputs(9462) <= a and not b;
    layer8_outputs(9463) <= a;
    layer8_outputs(9464) <= a xor b;
    layer8_outputs(9465) <= a;
    layer8_outputs(9466) <= a or b;
    layer8_outputs(9467) <= a xor b;
    layer8_outputs(9468) <= not (a or b);
    layer8_outputs(9469) <= not b;
    layer8_outputs(9470) <= a and not b;
    layer8_outputs(9471) <= not (a xor b);
    layer8_outputs(9472) <= not a;
    layer8_outputs(9473) <= not a;
    layer8_outputs(9474) <= not a;
    layer8_outputs(9475) <= a and b;
    layer8_outputs(9476) <= not a;
    layer8_outputs(9477) <= a;
    layer8_outputs(9478) <= a;
    layer8_outputs(9479) <= not a or b;
    layer8_outputs(9480) <= not a;
    layer8_outputs(9481) <= not b or a;
    layer8_outputs(9482) <= not b;
    layer8_outputs(9483) <= not (a xor b);
    layer8_outputs(9484) <= not (a or b);
    layer8_outputs(9485) <= a and not b;
    layer8_outputs(9486) <= a xor b;
    layer8_outputs(9487) <= a xor b;
    layer8_outputs(9488) <= not b or a;
    layer8_outputs(9489) <= b;
    layer8_outputs(9490) <= not b;
    layer8_outputs(9491) <= a and b;
    layer8_outputs(9492) <= not (a xor b);
    layer8_outputs(9493) <= b;
    layer8_outputs(9494) <= a xor b;
    layer8_outputs(9495) <= not (a xor b);
    layer8_outputs(9496) <= not a;
    layer8_outputs(9497) <= b;
    layer8_outputs(9498) <= not b;
    layer8_outputs(9499) <= not a or b;
    layer8_outputs(9500) <= not (a xor b);
    layer8_outputs(9501) <= not (a xor b);
    layer8_outputs(9502) <= not (a xor b);
    layer8_outputs(9503) <= not a;
    layer8_outputs(9504) <= not b;
    layer8_outputs(9505) <= not (a xor b);
    layer8_outputs(9506) <= not b;
    layer8_outputs(9507) <= a xor b;
    layer8_outputs(9508) <= b;
    layer8_outputs(9509) <= a;
    layer8_outputs(9510) <= not b or a;
    layer8_outputs(9511) <= a xor b;
    layer8_outputs(9512) <= not a;
    layer8_outputs(9513) <= a xor b;
    layer8_outputs(9514) <= a and b;
    layer8_outputs(9515) <= b;
    layer8_outputs(9516) <= a and not b;
    layer8_outputs(9517) <= not b;
    layer8_outputs(9518) <= not (a xor b);
    layer8_outputs(9519) <= not (a xor b);
    layer8_outputs(9520) <= not a;
    layer8_outputs(9521) <= not b;
    layer8_outputs(9522) <= a xor b;
    layer8_outputs(9523) <= not b;
    layer8_outputs(9524) <= not a or b;
    layer8_outputs(9525) <= a;
    layer8_outputs(9526) <= not a;
    layer8_outputs(9527) <= a and b;
    layer8_outputs(9528) <= not a;
    layer8_outputs(9529) <= not b or a;
    layer8_outputs(9530) <= b;
    layer8_outputs(9531) <= a and not b;
    layer8_outputs(9532) <= a;
    layer8_outputs(9533) <= not b or a;
    layer8_outputs(9534) <= not a;
    layer8_outputs(9535) <= a and b;
    layer8_outputs(9536) <= not (a or b);
    layer8_outputs(9537) <= not b;
    layer8_outputs(9538) <= b;
    layer8_outputs(9539) <= b and not a;
    layer8_outputs(9540) <= not b;
    layer8_outputs(9541) <= not a;
    layer8_outputs(9542) <= not (a and b);
    layer8_outputs(9543) <= b;
    layer8_outputs(9544) <= not (a xor b);
    layer8_outputs(9545) <= not a;
    layer8_outputs(9546) <= a;
    layer8_outputs(9547) <= b;
    layer8_outputs(9548) <= a and not b;
    layer8_outputs(9549) <= not a;
    layer8_outputs(9550) <= b;
    layer8_outputs(9551) <= not a;
    layer8_outputs(9552) <= not (a xor b);
    layer8_outputs(9553) <= not b;
    layer8_outputs(9554) <= not a or b;
    layer8_outputs(9555) <= a xor b;
    layer8_outputs(9556) <= not b or a;
    layer8_outputs(9557) <= a xor b;
    layer8_outputs(9558) <= not (a and b);
    layer8_outputs(9559) <= not (a xor b);
    layer8_outputs(9560) <= a and b;
    layer8_outputs(9561) <= not a or b;
    layer8_outputs(9562) <= a and b;
    layer8_outputs(9563) <= a xor b;
    layer8_outputs(9564) <= b;
    layer8_outputs(9565) <= a and b;
    layer8_outputs(9566) <= a and not b;
    layer8_outputs(9567) <= a and not b;
    layer8_outputs(9568) <= not b;
    layer8_outputs(9569) <= not (a xor b);
    layer8_outputs(9570) <= not (a and b);
    layer8_outputs(9571) <= a;
    layer8_outputs(9572) <= a xor b;
    layer8_outputs(9573) <= not (a or b);
    layer8_outputs(9574) <= a xor b;
    layer8_outputs(9575) <= a;
    layer8_outputs(9576) <= a and not b;
    layer8_outputs(9577) <= not (a xor b);
    layer8_outputs(9578) <= a and b;
    layer8_outputs(9579) <= a and b;
    layer8_outputs(9580) <= a and b;
    layer8_outputs(9581) <= not (a xor b);
    layer8_outputs(9582) <= a;
    layer8_outputs(9583) <= a and b;
    layer8_outputs(9584) <= a and not b;
    layer8_outputs(9585) <= a xor b;
    layer8_outputs(9586) <= a;
    layer8_outputs(9587) <= not (a xor b);
    layer8_outputs(9588) <= not a;
    layer8_outputs(9589) <= not (a and b);
    layer8_outputs(9590) <= not b or a;
    layer8_outputs(9591) <= a;
    layer8_outputs(9592) <= a and not b;
    layer8_outputs(9593) <= not b or a;
    layer8_outputs(9594) <= not b;
    layer8_outputs(9595) <= not b;
    layer8_outputs(9596) <= not b;
    layer8_outputs(9597) <= not (a xor b);
    layer8_outputs(9598) <= not a;
    layer8_outputs(9599) <= b;
    layer8_outputs(9600) <= not b;
    layer8_outputs(9601) <= b;
    layer8_outputs(9602) <= not a or b;
    layer8_outputs(9603) <= a xor b;
    layer8_outputs(9604) <= not a;
    layer8_outputs(9605) <= a xor b;
    layer8_outputs(9606) <= b;
    layer8_outputs(9607) <= b and not a;
    layer8_outputs(9608) <= a and b;
    layer8_outputs(9609) <= not b;
    layer8_outputs(9610) <= not a;
    layer8_outputs(9611) <= b and not a;
    layer8_outputs(9612) <= b and not a;
    layer8_outputs(9613) <= not b;
    layer8_outputs(9614) <= a xor b;
    layer8_outputs(9615) <= not (a xor b);
    layer8_outputs(9616) <= not (a xor b);
    layer8_outputs(9617) <= not (a xor b);
    layer8_outputs(9618) <= a xor b;
    layer8_outputs(9619) <= not (a or b);
    layer8_outputs(9620) <= not b or a;
    layer8_outputs(9621) <= a or b;
    layer8_outputs(9622) <= not (a xor b);
    layer8_outputs(9623) <= b;
    layer8_outputs(9624) <= a xor b;
    layer8_outputs(9625) <= not b;
    layer8_outputs(9626) <= not b or a;
    layer8_outputs(9627) <= not (a xor b);
    layer8_outputs(9628) <= a;
    layer8_outputs(9629) <= not b or a;
    layer8_outputs(9630) <= not (a xor b);
    layer8_outputs(9631) <= a;
    layer8_outputs(9632) <= not b;
    layer8_outputs(9633) <= b and not a;
    layer8_outputs(9634) <= b;
    layer8_outputs(9635) <= a xor b;
    layer8_outputs(9636) <= not a;
    layer8_outputs(9637) <= not (a xor b);
    layer8_outputs(9638) <= b and not a;
    layer8_outputs(9639) <= not a or b;
    layer8_outputs(9640) <= a;
    layer8_outputs(9641) <= b;
    layer8_outputs(9642) <= a xor b;
    layer8_outputs(9643) <= a;
    layer8_outputs(9644) <= a;
    layer8_outputs(9645) <= b and not a;
    layer8_outputs(9646) <= not a or b;
    layer8_outputs(9647) <= a or b;
    layer8_outputs(9648) <= not a;
    layer8_outputs(9649) <= not a or b;
    layer8_outputs(9650) <= a xor b;
    layer8_outputs(9651) <= not a or b;
    layer8_outputs(9652) <= a xor b;
    layer8_outputs(9653) <= not (a and b);
    layer8_outputs(9654) <= b;
    layer8_outputs(9655) <= a and not b;
    layer8_outputs(9656) <= not (a or b);
    layer8_outputs(9657) <= a;
    layer8_outputs(9658) <= b and not a;
    layer8_outputs(9659) <= b;
    layer8_outputs(9660) <= not (a or b);
    layer8_outputs(9661) <= b;
    layer8_outputs(9662) <= not (a or b);
    layer8_outputs(9663) <= not (a xor b);
    layer8_outputs(9664) <= not a;
    layer8_outputs(9665) <= not a or b;
    layer8_outputs(9666) <= not (a and b);
    layer8_outputs(9667) <= not (a xor b);
    layer8_outputs(9668) <= not b or a;
    layer8_outputs(9669) <= not b;
    layer8_outputs(9670) <= a;
    layer8_outputs(9671) <= not (a xor b);
    layer8_outputs(9672) <= b;
    layer8_outputs(9673) <= not a or b;
    layer8_outputs(9674) <= not (a or b);
    layer8_outputs(9675) <= a;
    layer8_outputs(9676) <= not b;
    layer8_outputs(9677) <= a or b;
    layer8_outputs(9678) <= b;
    layer8_outputs(9679) <= not (a or b);
    layer8_outputs(9680) <= a and not b;
    layer8_outputs(9681) <= b;
    layer8_outputs(9682) <= not b or a;
    layer8_outputs(9683) <= not b or a;
    layer8_outputs(9684) <= a xor b;
    layer8_outputs(9685) <= not (a xor b);
    layer8_outputs(9686) <= not b;
    layer8_outputs(9687) <= not (a xor b);
    layer8_outputs(9688) <= a xor b;
    layer8_outputs(9689) <= not b;
    layer8_outputs(9690) <= a;
    layer8_outputs(9691) <= a;
    layer8_outputs(9692) <= a and not b;
    layer8_outputs(9693) <= b and not a;
    layer8_outputs(9694) <= b;
    layer8_outputs(9695) <= a;
    layer8_outputs(9696) <= a and not b;
    layer8_outputs(9697) <= not a;
    layer8_outputs(9698) <= a xor b;
    layer8_outputs(9699) <= a xor b;
    layer8_outputs(9700) <= b;
    layer8_outputs(9701) <= a xor b;
    layer8_outputs(9702) <= b;
    layer8_outputs(9703) <= b and not a;
    layer8_outputs(9704) <= not b or a;
    layer8_outputs(9705) <= not a or b;
    layer8_outputs(9706) <= not b or a;
    layer8_outputs(9707) <= not (a xor b);
    layer8_outputs(9708) <= a or b;
    layer8_outputs(9709) <= not a;
    layer8_outputs(9710) <= b and not a;
    layer8_outputs(9711) <= a or b;
    layer8_outputs(9712) <= a or b;
    layer8_outputs(9713) <= a xor b;
    layer8_outputs(9714) <= a xor b;
    layer8_outputs(9715) <= a xor b;
    layer8_outputs(9716) <= not (a and b);
    layer8_outputs(9717) <= b;
    layer8_outputs(9718) <= a and not b;
    layer8_outputs(9719) <= a xor b;
    layer8_outputs(9720) <= not (a xor b);
    layer8_outputs(9721) <= not (a xor b);
    layer8_outputs(9722) <= not (a xor b);
    layer8_outputs(9723) <= b and not a;
    layer8_outputs(9724) <= not a;
    layer8_outputs(9725) <= a;
    layer8_outputs(9726) <= a;
    layer8_outputs(9727) <= b and not a;
    layer8_outputs(9728) <= a or b;
    layer8_outputs(9729) <= a;
    layer8_outputs(9730) <= not a;
    layer8_outputs(9731) <= a and not b;
    layer8_outputs(9732) <= not a;
    layer8_outputs(9733) <= a and b;
    layer8_outputs(9734) <= a and b;
    layer8_outputs(9735) <= a xor b;
    layer8_outputs(9736) <= b;
    layer8_outputs(9737) <= not b;
    layer8_outputs(9738) <= not (a xor b);
    layer8_outputs(9739) <= b;
    layer8_outputs(9740) <= not b;
    layer8_outputs(9741) <= not a;
    layer8_outputs(9742) <= not a or b;
    layer8_outputs(9743) <= not a or b;
    layer8_outputs(9744) <= b;
    layer8_outputs(9745) <= a or b;
    layer8_outputs(9746) <= b;
    layer8_outputs(9747) <= not (a or b);
    layer8_outputs(9748) <= a xor b;
    layer8_outputs(9749) <= not a;
    layer8_outputs(9750) <= a;
    layer8_outputs(9751) <= b and not a;
    layer8_outputs(9752) <= a or b;
    layer8_outputs(9753) <= b;
    layer8_outputs(9754) <= not (a and b);
    layer8_outputs(9755) <= b;
    layer8_outputs(9756) <= b;
    layer8_outputs(9757) <= not (a and b);
    layer8_outputs(9758) <= not a;
    layer8_outputs(9759) <= not a;
    layer8_outputs(9760) <= not (a xor b);
    layer8_outputs(9761) <= not b;
    layer8_outputs(9762) <= a and not b;
    layer8_outputs(9763) <= a xor b;
    layer8_outputs(9764) <= not (a or b);
    layer8_outputs(9765) <= not b;
    layer8_outputs(9766) <= not b;
    layer8_outputs(9767) <= not (a and b);
    layer8_outputs(9768) <= a;
    layer8_outputs(9769) <= not (a xor b);
    layer8_outputs(9770) <= not a or b;
    layer8_outputs(9771) <= not (a or b);
    layer8_outputs(9772) <= a xor b;
    layer8_outputs(9773) <= not (a and b);
    layer8_outputs(9774) <= not b or a;
    layer8_outputs(9775) <= a xor b;
    layer8_outputs(9776) <= a and b;
    layer8_outputs(9777) <= b;
    layer8_outputs(9778) <= a xor b;
    layer8_outputs(9779) <= not b;
    layer8_outputs(9780) <= b;
    layer8_outputs(9781) <= a xor b;
    layer8_outputs(9782) <= not (a and b);
    layer8_outputs(9783) <= b;
    layer8_outputs(9784) <= not (a xor b);
    layer8_outputs(9785) <= not b;
    layer8_outputs(9786) <= not a;
    layer8_outputs(9787) <= a xor b;
    layer8_outputs(9788) <= a xor b;
    layer8_outputs(9789) <= a and b;
    layer8_outputs(9790) <= not a;
    layer8_outputs(9791) <= not a or b;
    layer8_outputs(9792) <= not (a xor b);
    layer8_outputs(9793) <= a or b;
    layer8_outputs(9794) <= a;
    layer8_outputs(9795) <= not b;
    layer8_outputs(9796) <= b;
    layer8_outputs(9797) <= not b;
    layer8_outputs(9798) <= b and not a;
    layer8_outputs(9799) <= not (a xor b);
    layer8_outputs(9800) <= not a or b;
    layer8_outputs(9801) <= b;
    layer8_outputs(9802) <= not a or b;
    layer8_outputs(9803) <= not (a xor b);
    layer8_outputs(9804) <= a;
    layer8_outputs(9805) <= a;
    layer8_outputs(9806) <= not (a xor b);
    layer8_outputs(9807) <= a;
    layer8_outputs(9808) <= not (a xor b);
    layer8_outputs(9809) <= a;
    layer8_outputs(9810) <= not b;
    layer8_outputs(9811) <= not (a xor b);
    layer8_outputs(9812) <= a xor b;
    layer8_outputs(9813) <= b;
    layer8_outputs(9814) <= a;
    layer8_outputs(9815) <= b;
    layer8_outputs(9816) <= not (a or b);
    layer8_outputs(9817) <= b;
    layer8_outputs(9818) <= a or b;
    layer8_outputs(9819) <= not a;
    layer8_outputs(9820) <= not a or b;
    layer8_outputs(9821) <= b;
    layer8_outputs(9822) <= not a or b;
    layer8_outputs(9823) <= a xor b;
    layer8_outputs(9824) <= 1'b1;
    layer8_outputs(9825) <= a;
    layer8_outputs(9826) <= not (a xor b);
    layer8_outputs(9827) <= not (a or b);
    layer8_outputs(9828) <= b;
    layer8_outputs(9829) <= not (a and b);
    layer8_outputs(9830) <= a xor b;
    layer8_outputs(9831) <= a and b;
    layer8_outputs(9832) <= not (a xor b);
    layer8_outputs(9833) <= not (a xor b);
    layer8_outputs(9834) <= not b or a;
    layer8_outputs(9835) <= a and b;
    layer8_outputs(9836) <= not a or b;
    layer8_outputs(9837) <= a;
    layer8_outputs(9838) <= not b;
    layer8_outputs(9839) <= b and not a;
    layer8_outputs(9840) <= a xor b;
    layer8_outputs(9841) <= b;
    layer8_outputs(9842) <= not a or b;
    layer8_outputs(9843) <= not (a xor b);
    layer8_outputs(9844) <= a and not b;
    layer8_outputs(9845) <= b and not a;
    layer8_outputs(9846) <= a xor b;
    layer8_outputs(9847) <= not (a xor b);
    layer8_outputs(9848) <= a and b;
    layer8_outputs(9849) <= b;
    layer8_outputs(9850) <= not b;
    layer8_outputs(9851) <= a xor b;
    layer8_outputs(9852) <= a xor b;
    layer8_outputs(9853) <= not (a xor b);
    layer8_outputs(9854) <= a;
    layer8_outputs(9855) <= not b or a;
    layer8_outputs(9856) <= a;
    layer8_outputs(9857) <= a and not b;
    layer8_outputs(9858) <= a or b;
    layer8_outputs(9859) <= a xor b;
    layer8_outputs(9860) <= not a;
    layer8_outputs(9861) <= b;
    layer8_outputs(9862) <= a and b;
    layer8_outputs(9863) <= b;
    layer8_outputs(9864) <= a xor b;
    layer8_outputs(9865) <= not b;
    layer8_outputs(9866) <= b;
    layer8_outputs(9867) <= not a or b;
    layer8_outputs(9868) <= b and not a;
    layer8_outputs(9869) <= not a;
    layer8_outputs(9870) <= b and not a;
    layer8_outputs(9871) <= not b;
    layer8_outputs(9872) <= not b;
    layer8_outputs(9873) <= b;
    layer8_outputs(9874) <= a xor b;
    layer8_outputs(9875) <= not b;
    layer8_outputs(9876) <= a and b;
    layer8_outputs(9877) <= not (a xor b);
    layer8_outputs(9878) <= not a;
    layer8_outputs(9879) <= a and b;
    layer8_outputs(9880) <= not a;
    layer8_outputs(9881) <= b;
    layer8_outputs(9882) <= not b or a;
    layer8_outputs(9883) <= b;
    layer8_outputs(9884) <= not b;
    layer8_outputs(9885) <= a;
    layer8_outputs(9886) <= a or b;
    layer8_outputs(9887) <= not a;
    layer8_outputs(9888) <= b;
    layer8_outputs(9889) <= b and not a;
    layer8_outputs(9890) <= not (a xor b);
    layer8_outputs(9891) <= not (a and b);
    layer8_outputs(9892) <= a xor b;
    layer8_outputs(9893) <= not a or b;
    layer8_outputs(9894) <= not a;
    layer8_outputs(9895) <= not b;
    layer8_outputs(9896) <= not b;
    layer8_outputs(9897) <= not b or a;
    layer8_outputs(9898) <= a and not b;
    layer8_outputs(9899) <= a or b;
    layer8_outputs(9900) <= not b or a;
    layer8_outputs(9901) <= a xor b;
    layer8_outputs(9902) <= b and not a;
    layer8_outputs(9903) <= not b;
    layer8_outputs(9904) <= not b or a;
    layer8_outputs(9905) <= b and not a;
    layer8_outputs(9906) <= a xor b;
    layer8_outputs(9907) <= b;
    layer8_outputs(9908) <= not (a xor b);
    layer8_outputs(9909) <= not a;
    layer8_outputs(9910) <= b;
    layer8_outputs(9911) <= not (a xor b);
    layer8_outputs(9912) <= not b;
    layer8_outputs(9913) <= not (a xor b);
    layer8_outputs(9914) <= not b or a;
    layer8_outputs(9915) <= a and not b;
    layer8_outputs(9916) <= b;
    layer8_outputs(9917) <= b and not a;
    layer8_outputs(9918) <= not a or b;
    layer8_outputs(9919) <= not (a xor b);
    layer8_outputs(9920) <= not (a xor b);
    layer8_outputs(9921) <= not b;
    layer8_outputs(9922) <= b and not a;
    layer8_outputs(9923) <= b and not a;
    layer8_outputs(9924) <= not b;
    layer8_outputs(9925) <= b and not a;
    layer8_outputs(9926) <= not a;
    layer8_outputs(9927) <= a and b;
    layer8_outputs(9928) <= a and b;
    layer8_outputs(9929) <= a;
    layer8_outputs(9930) <= not (a xor b);
    layer8_outputs(9931) <= not (a xor b);
    layer8_outputs(9932) <= a;
    layer8_outputs(9933) <= a;
    layer8_outputs(9934) <= b;
    layer8_outputs(9935) <= b;
    layer8_outputs(9936) <= not (a xor b);
    layer8_outputs(9937) <= a;
    layer8_outputs(9938) <= not (a xor b);
    layer8_outputs(9939) <= a;
    layer8_outputs(9940) <= b;
    layer8_outputs(9941) <= a or b;
    layer8_outputs(9942) <= b and not a;
    layer8_outputs(9943) <= not b;
    layer8_outputs(9944) <= b;
    layer8_outputs(9945) <= not b;
    layer8_outputs(9946) <= not (a or b);
    layer8_outputs(9947) <= a or b;
    layer8_outputs(9948) <= a xor b;
    layer8_outputs(9949) <= not (a xor b);
    layer8_outputs(9950) <= not (a xor b);
    layer8_outputs(9951) <= b;
    layer8_outputs(9952) <= a xor b;
    layer8_outputs(9953) <= a or b;
    layer8_outputs(9954) <= a and not b;
    layer8_outputs(9955) <= not a;
    layer8_outputs(9956) <= a;
    layer8_outputs(9957) <= not a;
    layer8_outputs(9958) <= a xor b;
    layer8_outputs(9959) <= not b;
    layer8_outputs(9960) <= not b;
    layer8_outputs(9961) <= not a;
    layer8_outputs(9962) <= not b;
    layer8_outputs(9963) <= not (a xor b);
    layer8_outputs(9964) <= a xor b;
    layer8_outputs(9965) <= a or b;
    layer8_outputs(9966) <= not a or b;
    layer8_outputs(9967) <= not b;
    layer8_outputs(9968) <= b;
    layer8_outputs(9969) <= not (a and b);
    layer8_outputs(9970) <= not (a xor b);
    layer8_outputs(9971) <= a and not b;
    layer8_outputs(9972) <= b;
    layer8_outputs(9973) <= a and not b;
    layer8_outputs(9974) <= b and not a;
    layer8_outputs(9975) <= not b or a;
    layer8_outputs(9976) <= not a;
    layer8_outputs(9977) <= a or b;
    layer8_outputs(9978) <= a or b;
    layer8_outputs(9979) <= not a or b;
    layer8_outputs(9980) <= a xor b;
    layer8_outputs(9981) <= a and b;
    layer8_outputs(9982) <= not a;
    layer8_outputs(9983) <= not a;
    layer8_outputs(9984) <= not (a xor b);
    layer8_outputs(9985) <= b;
    layer8_outputs(9986) <= a or b;
    layer8_outputs(9987) <= a;
    layer8_outputs(9988) <= not a or b;
    layer8_outputs(9989) <= a;
    layer8_outputs(9990) <= not a;
    layer8_outputs(9991) <= not (a xor b);
    layer8_outputs(9992) <= a;
    layer8_outputs(9993) <= not (a or b);
    layer8_outputs(9994) <= a;
    layer8_outputs(9995) <= a xor b;
    layer8_outputs(9996) <= a xor b;
    layer8_outputs(9997) <= not (a xor b);
    layer8_outputs(9998) <= not (a xor b);
    layer8_outputs(9999) <= not a;
    layer8_outputs(10000) <= a;
    layer8_outputs(10001) <= a;
    layer8_outputs(10002) <= not a;
    layer8_outputs(10003) <= a or b;
    layer8_outputs(10004) <= b;
    layer8_outputs(10005) <= a xor b;
    layer8_outputs(10006) <= not b;
    layer8_outputs(10007) <= a xor b;
    layer8_outputs(10008) <= a xor b;
    layer8_outputs(10009) <= a and b;
    layer8_outputs(10010) <= a xor b;
    layer8_outputs(10011) <= a xor b;
    layer8_outputs(10012) <= a xor b;
    layer8_outputs(10013) <= a or b;
    layer8_outputs(10014) <= not a;
    layer8_outputs(10015) <= not a or b;
    layer8_outputs(10016) <= not (a xor b);
    layer8_outputs(10017) <= not b;
    layer8_outputs(10018) <= a xor b;
    layer8_outputs(10019) <= a and not b;
    layer8_outputs(10020) <= a and b;
    layer8_outputs(10021) <= not (a xor b);
    layer8_outputs(10022) <= not a;
    layer8_outputs(10023) <= not a;
    layer8_outputs(10024) <= not (a and b);
    layer8_outputs(10025) <= not b;
    layer8_outputs(10026) <= a;
    layer8_outputs(10027) <= a or b;
    layer8_outputs(10028) <= a;
    layer8_outputs(10029) <= b;
    layer8_outputs(10030) <= b;
    layer8_outputs(10031) <= a and b;
    layer8_outputs(10032) <= b and not a;
    layer8_outputs(10033) <= not a;
    layer8_outputs(10034) <= a and b;
    layer8_outputs(10035) <= a;
    layer8_outputs(10036) <= not (a or b);
    layer8_outputs(10037) <= a xor b;
    layer8_outputs(10038) <= not b or a;
    layer8_outputs(10039) <= not b;
    layer8_outputs(10040) <= not (a or b);
    layer8_outputs(10041) <= not b or a;
    layer8_outputs(10042) <= a;
    layer8_outputs(10043) <= a and b;
    layer8_outputs(10044) <= a and not b;
    layer8_outputs(10045) <= b;
    layer8_outputs(10046) <= not b;
    layer8_outputs(10047) <= not a;
    layer8_outputs(10048) <= not b;
    layer8_outputs(10049) <= b;
    layer8_outputs(10050) <= not (a xor b);
    layer8_outputs(10051) <= a;
    layer8_outputs(10052) <= not a;
    layer8_outputs(10053) <= a;
    layer8_outputs(10054) <= not (a xor b);
    layer8_outputs(10055) <= not b or a;
    layer8_outputs(10056) <= not b;
    layer8_outputs(10057) <= not a;
    layer8_outputs(10058) <= not a or b;
    layer8_outputs(10059) <= b and not a;
    layer8_outputs(10060) <= a xor b;
    layer8_outputs(10061) <= a;
    layer8_outputs(10062) <= b and not a;
    layer8_outputs(10063) <= a xor b;
    layer8_outputs(10064) <= a and b;
    layer8_outputs(10065) <= not a;
    layer8_outputs(10066) <= not b;
    layer8_outputs(10067) <= not b or a;
    layer8_outputs(10068) <= not a;
    layer8_outputs(10069) <= b;
    layer8_outputs(10070) <= 1'b1;
    layer8_outputs(10071) <= not (a and b);
    layer8_outputs(10072) <= a and not b;
    layer8_outputs(10073) <= b;
    layer8_outputs(10074) <= not b;
    layer8_outputs(10075) <= not b or a;
    layer8_outputs(10076) <= not (a and b);
    layer8_outputs(10077) <= not a;
    layer8_outputs(10078) <= a xor b;
    layer8_outputs(10079) <= not (a or b);
    layer8_outputs(10080) <= a xor b;
    layer8_outputs(10081) <= 1'b1;
    layer8_outputs(10082) <= not (a xor b);
    layer8_outputs(10083) <= a xor b;
    layer8_outputs(10084) <= b;
    layer8_outputs(10085) <= not b;
    layer8_outputs(10086) <= not a or b;
    layer8_outputs(10087) <= b and not a;
    layer8_outputs(10088) <= a;
    layer8_outputs(10089) <= not b or a;
    layer8_outputs(10090) <= not a;
    layer8_outputs(10091) <= not a;
    layer8_outputs(10092) <= a xor b;
    layer8_outputs(10093) <= not (a xor b);
    layer8_outputs(10094) <= not a;
    layer8_outputs(10095) <= a xor b;
    layer8_outputs(10096) <= not (a xor b);
    layer8_outputs(10097) <= a or b;
    layer8_outputs(10098) <= b;
    layer8_outputs(10099) <= b;
    layer8_outputs(10100) <= not (a xor b);
    layer8_outputs(10101) <= not b or a;
    layer8_outputs(10102) <= a xor b;
    layer8_outputs(10103) <= not (a or b);
    layer8_outputs(10104) <= a xor b;
    layer8_outputs(10105) <= b and not a;
    layer8_outputs(10106) <= not b or a;
    layer8_outputs(10107) <= b;
    layer8_outputs(10108) <= not (a xor b);
    layer8_outputs(10109) <= a;
    layer8_outputs(10110) <= not b;
    layer8_outputs(10111) <= a xor b;
    layer8_outputs(10112) <= not (a xor b);
    layer8_outputs(10113) <= not a;
    layer8_outputs(10114) <= a xor b;
    layer8_outputs(10115) <= b and not a;
    layer8_outputs(10116) <= not (a xor b);
    layer8_outputs(10117) <= a;
    layer8_outputs(10118) <= a or b;
    layer8_outputs(10119) <= b;
    layer8_outputs(10120) <= not a;
    layer8_outputs(10121) <= not (a or b);
    layer8_outputs(10122) <= not b;
    layer8_outputs(10123) <= not b or a;
    layer8_outputs(10124) <= 1'b1;
    layer8_outputs(10125) <= not b;
    layer8_outputs(10126) <= not b or a;
    layer8_outputs(10127) <= b;
    layer8_outputs(10128) <= not a;
    layer8_outputs(10129) <= a and b;
    layer8_outputs(10130) <= not (a and b);
    layer8_outputs(10131) <= not a;
    layer8_outputs(10132) <= not a;
    layer8_outputs(10133) <= not (a xor b);
    layer8_outputs(10134) <= not a;
    layer8_outputs(10135) <= not a or b;
    layer8_outputs(10136) <= not b;
    layer8_outputs(10137) <= a xor b;
    layer8_outputs(10138) <= a;
    layer8_outputs(10139) <= b;
    layer8_outputs(10140) <= not (a xor b);
    layer8_outputs(10141) <= not (a and b);
    layer8_outputs(10142) <= a;
    layer8_outputs(10143) <= a and not b;
    layer8_outputs(10144) <= a;
    layer8_outputs(10145) <= not a or b;
    layer8_outputs(10146) <= b;
    layer8_outputs(10147) <= a xor b;
    layer8_outputs(10148) <= not (a or b);
    layer8_outputs(10149) <= a;
    layer8_outputs(10150) <= a xor b;
    layer8_outputs(10151) <= not b;
    layer8_outputs(10152) <= a xor b;
    layer8_outputs(10153) <= not b or a;
    layer8_outputs(10154) <= a;
    layer8_outputs(10155) <= a;
    layer8_outputs(10156) <= b and not a;
    layer8_outputs(10157) <= a or b;
    layer8_outputs(10158) <= b;
    layer8_outputs(10159) <= not b;
    layer8_outputs(10160) <= b;
    layer8_outputs(10161) <= not a;
    layer8_outputs(10162) <= a or b;
    layer8_outputs(10163) <= a;
    layer8_outputs(10164) <= not b;
    layer8_outputs(10165) <= b;
    layer8_outputs(10166) <= a or b;
    layer8_outputs(10167) <= b;
    layer8_outputs(10168) <= b;
    layer8_outputs(10169) <= a;
    layer8_outputs(10170) <= b;
    layer8_outputs(10171) <= a;
    layer8_outputs(10172) <= a;
    layer8_outputs(10173) <= not a;
    layer8_outputs(10174) <= not (a and b);
    layer8_outputs(10175) <= not a;
    layer8_outputs(10176) <= not b or a;
    layer8_outputs(10177) <= not (a and b);
    layer8_outputs(10178) <= b;
    layer8_outputs(10179) <= not b;
    layer8_outputs(10180) <= a or b;
    layer8_outputs(10181) <= not a;
    layer8_outputs(10182) <= a xor b;
    layer8_outputs(10183) <= not b;
    layer8_outputs(10184) <= b;
    layer8_outputs(10185) <= not a;
    layer8_outputs(10186) <= not (a and b);
    layer8_outputs(10187) <= not a;
    layer8_outputs(10188) <= not a;
    layer8_outputs(10189) <= a xor b;
    layer8_outputs(10190) <= b and not a;
    layer8_outputs(10191) <= not b;
    layer8_outputs(10192) <= a and not b;
    layer8_outputs(10193) <= not a or b;
    layer8_outputs(10194) <= a xor b;
    layer8_outputs(10195) <= a xor b;
    layer8_outputs(10196) <= not b or a;
    layer8_outputs(10197) <= not b;
    layer8_outputs(10198) <= not (a or b);
    layer8_outputs(10199) <= b;
    layer8_outputs(10200) <= a xor b;
    layer8_outputs(10201) <= not a or b;
    layer8_outputs(10202) <= not a;
    layer8_outputs(10203) <= not (a and b);
    layer8_outputs(10204) <= not a or b;
    layer8_outputs(10205) <= not a;
    layer8_outputs(10206) <= not b;
    layer8_outputs(10207) <= not (a and b);
    layer8_outputs(10208) <= 1'b1;
    layer8_outputs(10209) <= not (a and b);
    layer8_outputs(10210) <= not (a xor b);
    layer8_outputs(10211) <= a;
    layer8_outputs(10212) <= b and not a;
    layer8_outputs(10213) <= b;
    layer8_outputs(10214) <= not a;
    layer8_outputs(10215) <= not b or a;
    layer8_outputs(10216) <= a and not b;
    layer8_outputs(10217) <= a and b;
    layer8_outputs(10218) <= b;
    layer8_outputs(10219) <= not b;
    layer8_outputs(10220) <= not (a xor b);
    layer8_outputs(10221) <= not (a or b);
    layer8_outputs(10222) <= not (a and b);
    layer8_outputs(10223) <= a;
    layer8_outputs(10224) <= not a or b;
    layer8_outputs(10225) <= not a;
    layer8_outputs(10226) <= b;
    layer8_outputs(10227) <= a and not b;
    layer8_outputs(10228) <= b;
    layer8_outputs(10229) <= not a;
    layer8_outputs(10230) <= not b or a;
    layer8_outputs(10231) <= a and not b;
    layer8_outputs(10232) <= not b;
    layer8_outputs(10233) <= not a;
    layer8_outputs(10234) <= b;
    layer8_outputs(10235) <= not b;
    layer8_outputs(10236) <= a and b;
    layer8_outputs(10237) <= b;
    layer8_outputs(10238) <= not b;
    layer8_outputs(10239) <= not b;
    outputs(0) <= b;
    outputs(1) <= not a;
    outputs(2) <= a;
    outputs(3) <= a xor b;
    outputs(4) <= not a or b;
    outputs(5) <= a xor b;
    outputs(6) <= not (a xor b);
    outputs(7) <= b;
    outputs(8) <= b;
    outputs(9) <= not (a xor b);
    outputs(10) <= a;
    outputs(11) <= not a;
    outputs(12) <= a and b;
    outputs(13) <= not b;
    outputs(14) <= not a;
    outputs(15) <= a xor b;
    outputs(16) <= not (a xor b);
    outputs(17) <= a xor b;
    outputs(18) <= not a;
    outputs(19) <= not a;
    outputs(20) <= a xor b;
    outputs(21) <= not b;
    outputs(22) <= b;
    outputs(23) <= not a;
    outputs(24) <= b;
    outputs(25) <= not (a xor b);
    outputs(26) <= not a;
    outputs(27) <= not b;
    outputs(28) <= a and not b;
    outputs(29) <= b and not a;
    outputs(30) <= not (a or b);
    outputs(31) <= b;
    outputs(32) <= b;
    outputs(33) <= not a;
    outputs(34) <= not a;
    outputs(35) <= b and not a;
    outputs(36) <= not a;
    outputs(37) <= not (a xor b);
    outputs(38) <= a and b;
    outputs(39) <= a;
    outputs(40) <= not a;
    outputs(41) <= not b;
    outputs(42) <= not a;
    outputs(43) <= a xor b;
    outputs(44) <= a and b;
    outputs(45) <= a;
    outputs(46) <= a xor b;
    outputs(47) <= not a;
    outputs(48) <= b;
    outputs(49) <= a;
    outputs(50) <= not b;
    outputs(51) <= not b;
    outputs(52) <= not a;
    outputs(53) <= b;
    outputs(54) <= not (a and b);
    outputs(55) <= a xor b;
    outputs(56) <= b and not a;
    outputs(57) <= a and not b;
    outputs(58) <= not a;
    outputs(59) <= a;
    outputs(60) <= not b;
    outputs(61) <= not b;
    outputs(62) <= b;
    outputs(63) <= a xor b;
    outputs(64) <= a;
    outputs(65) <= not (a xor b);
    outputs(66) <= a and not b;
    outputs(67) <= a and b;
    outputs(68) <= a xor b;
    outputs(69) <= not (a xor b);
    outputs(70) <= not a;
    outputs(71) <= not a;
    outputs(72) <= not b;
    outputs(73) <= a xor b;
    outputs(74) <= a;
    outputs(75) <= a and not b;
    outputs(76) <= not a;
    outputs(77) <= not b;
    outputs(78) <= b;
    outputs(79) <= a and not b;
    outputs(80) <= a xor b;
    outputs(81) <= not b;
    outputs(82) <= not b;
    outputs(83) <= a xor b;
    outputs(84) <= a;
    outputs(85) <= not b;
    outputs(86) <= a;
    outputs(87) <= b and not a;
    outputs(88) <= not b;
    outputs(89) <= not (a or b);
    outputs(90) <= a xor b;
    outputs(91) <= not b;
    outputs(92) <= not a;
    outputs(93) <= not (a xor b);
    outputs(94) <= b;
    outputs(95) <= not b or a;
    outputs(96) <= not b;
    outputs(97) <= not b or a;
    outputs(98) <= not a;
    outputs(99) <= a xor b;
    outputs(100) <= b;
    outputs(101) <= not (a xor b);
    outputs(102) <= a;
    outputs(103) <= not b;
    outputs(104) <= b and not a;
    outputs(105) <= not (a xor b);
    outputs(106) <= not (a or b);
    outputs(107) <= not (a xor b);
    outputs(108) <= a;
    outputs(109) <= not a;
    outputs(110) <= not a;
    outputs(111) <= a;
    outputs(112) <= not a;
    outputs(113) <= not b;
    outputs(114) <= b and not a;
    outputs(115) <= a xor b;
    outputs(116) <= not a;
    outputs(117) <= a;
    outputs(118) <= not (a xor b);
    outputs(119) <= not (a xor b);
    outputs(120) <= not b;
    outputs(121) <= not (a xor b);
    outputs(122) <= a;
    outputs(123) <= not (a or b);
    outputs(124) <= a xor b;
    outputs(125) <= a xor b;
    outputs(126) <= a xor b;
    outputs(127) <= not a;
    outputs(128) <= not b;
    outputs(129) <= not b;
    outputs(130) <= not (a xor b);
    outputs(131) <= not (a xor b);
    outputs(132) <= not b or a;
    outputs(133) <= b;
    outputs(134) <= not a;
    outputs(135) <= a xor b;
    outputs(136) <= not b;
    outputs(137) <= not a;
    outputs(138) <= not (a and b);
    outputs(139) <= not (a xor b);
    outputs(140) <= not (a xor b);
    outputs(141) <= a xor b;
    outputs(142) <= not (a xor b);
    outputs(143) <= not b or a;
    outputs(144) <= a xor b;
    outputs(145) <= a xor b;
    outputs(146) <= not b or a;
    outputs(147) <= a and not b;
    outputs(148) <= b;
    outputs(149) <= b;
    outputs(150) <= a xor b;
    outputs(151) <= b;
    outputs(152) <= a;
    outputs(153) <= a and b;
    outputs(154) <= not (a or b);
    outputs(155) <= not b;
    outputs(156) <= a;
    outputs(157) <= a;
    outputs(158) <= not a;
    outputs(159) <= b;
    outputs(160) <= not (a xor b);
    outputs(161) <= a xor b;
    outputs(162) <= not b or a;
    outputs(163) <= a xor b;
    outputs(164) <= not (a xor b);
    outputs(165) <= not (a xor b);
    outputs(166) <= a xor b;
    outputs(167) <= a xor b;
    outputs(168) <= a xor b;
    outputs(169) <= b;
    outputs(170) <= not a;
    outputs(171) <= b;
    outputs(172) <= b and not a;
    outputs(173) <= a and b;
    outputs(174) <= not b;
    outputs(175) <= not a;
    outputs(176) <= b;
    outputs(177) <= a xor b;
    outputs(178) <= a xor b;
    outputs(179) <= a;
    outputs(180) <= a xor b;
    outputs(181) <= b;
    outputs(182) <= b;
    outputs(183) <= a xor b;
    outputs(184) <= not a or b;
    outputs(185) <= a xor b;
    outputs(186) <= a;
    outputs(187) <= a;
    outputs(188) <= a and b;
    outputs(189) <= a xor b;
    outputs(190) <= b;
    outputs(191) <= a and b;
    outputs(192) <= a and b;
    outputs(193) <= a;
    outputs(194) <= not (a xor b);
    outputs(195) <= a and b;
    outputs(196) <= not b;
    outputs(197) <= a and not b;
    outputs(198) <= not a;
    outputs(199) <= not a;
    outputs(200) <= a xor b;
    outputs(201) <= a and not b;
    outputs(202) <= a;
    outputs(203) <= not (a xor b);
    outputs(204) <= not (a xor b);
    outputs(205) <= not b;
    outputs(206) <= a xor b;
    outputs(207) <= b and not a;
    outputs(208) <= not a;
    outputs(209) <= not a;
    outputs(210) <= not a;
    outputs(211) <= b;
    outputs(212) <= b;
    outputs(213) <= b and not a;
    outputs(214) <= not (a xor b);
    outputs(215) <= a xor b;
    outputs(216) <= a xor b;
    outputs(217) <= a and not b;
    outputs(218) <= a;
    outputs(219) <= a;
    outputs(220) <= a and b;
    outputs(221) <= not (a xor b);
    outputs(222) <= not (a xor b);
    outputs(223) <= not b;
    outputs(224) <= a xor b;
    outputs(225) <= a xor b;
    outputs(226) <= a;
    outputs(227) <= a and b;
    outputs(228) <= a or b;
    outputs(229) <= not a;
    outputs(230) <= not (a xor b);
    outputs(231) <= not b;
    outputs(232) <= not (a xor b);
    outputs(233) <= not (a xor b);
    outputs(234) <= not b or a;
    outputs(235) <= not (a xor b);
    outputs(236) <= not b;
    outputs(237) <= not b;
    outputs(238) <= b and not a;
    outputs(239) <= a or b;
    outputs(240) <= not (a xor b);
    outputs(241) <= not b or a;
    outputs(242) <= not b;
    outputs(243) <= b;
    outputs(244) <= not b or a;
    outputs(245) <= not b or a;
    outputs(246) <= not b;
    outputs(247) <= a xor b;
    outputs(248) <= a xor b;
    outputs(249) <= a or b;
    outputs(250) <= a;
    outputs(251) <= not a;
    outputs(252) <= not (a xor b);
    outputs(253) <= a xor b;
    outputs(254) <= not b;
    outputs(255) <= a xor b;
    outputs(256) <= not a;
    outputs(257) <= a;
    outputs(258) <= b;
    outputs(259) <= not (a and b);
    outputs(260) <= a;
    outputs(261) <= not a;
    outputs(262) <= a and b;
    outputs(263) <= not b;
    outputs(264) <= not (a xor b);
    outputs(265) <= not b;
    outputs(266) <= a and b;
    outputs(267) <= a;
    outputs(268) <= not a or b;
    outputs(269) <= b;
    outputs(270) <= a xor b;
    outputs(271) <= not (a or b);
    outputs(272) <= not a;
    outputs(273) <= not (a xor b);
    outputs(274) <= a or b;
    outputs(275) <= b;
    outputs(276) <= a;
    outputs(277) <= b;
    outputs(278) <= b;
    outputs(279) <= not (a xor b);
    outputs(280) <= not (a xor b);
    outputs(281) <= not (a or b);
    outputs(282) <= not b or a;
    outputs(283) <= not a;
    outputs(284) <= a xor b;
    outputs(285) <= a;
    outputs(286) <= not b or a;
    outputs(287) <= a and b;
    outputs(288) <= not a;
    outputs(289) <= not a;
    outputs(290) <= not (a xor b);
    outputs(291) <= a and not b;
    outputs(292) <= a and not b;
    outputs(293) <= not (a xor b);
    outputs(294) <= not (a and b);
    outputs(295) <= not b;
    outputs(296) <= b and not a;
    outputs(297) <= not a or b;
    outputs(298) <= not (a xor b);
    outputs(299) <= a and b;
    outputs(300) <= b;
    outputs(301) <= not b;
    outputs(302) <= not a;
    outputs(303) <= a;
    outputs(304) <= not a or b;
    outputs(305) <= not b;
    outputs(306) <= a xor b;
    outputs(307) <= b;
    outputs(308) <= not b;
    outputs(309) <= a;
    outputs(310) <= not (a and b);
    outputs(311) <= a xor b;
    outputs(312) <= not b;
    outputs(313) <= not (a xor b);
    outputs(314) <= a xor b;
    outputs(315) <= b;
    outputs(316) <= not (a or b);
    outputs(317) <= not (a xor b);
    outputs(318) <= a xor b;
    outputs(319) <= b;
    outputs(320) <= not b;
    outputs(321) <= a xor b;
    outputs(322) <= a xor b;
    outputs(323) <= a xor b;
    outputs(324) <= b;
    outputs(325) <= a xor b;
    outputs(326) <= a xor b;
    outputs(327) <= not b;
    outputs(328) <= not b;
    outputs(329) <= not (a xor b);
    outputs(330) <= not a;
    outputs(331) <= not (a or b);
    outputs(332) <= not a;
    outputs(333) <= a xor b;
    outputs(334) <= a;
    outputs(335) <= a xor b;
    outputs(336) <= not (a xor b);
    outputs(337) <= a;
    outputs(338) <= a;
    outputs(339) <= not (a xor b);
    outputs(340) <= a xor b;
    outputs(341) <= b;
    outputs(342) <= b;
    outputs(343) <= b;
    outputs(344) <= not a;
    outputs(345) <= b;
    outputs(346) <= not b;
    outputs(347) <= not (a xor b);
    outputs(348) <= a xor b;
    outputs(349) <= not b;
    outputs(350) <= not a;
    outputs(351) <= not a;
    outputs(352) <= a xor b;
    outputs(353) <= not a or b;
    outputs(354) <= a xor b;
    outputs(355) <= a xor b;
    outputs(356) <= not a;
    outputs(357) <= not b;
    outputs(358) <= not a;
    outputs(359) <= not b;
    outputs(360) <= not (a xor b);
    outputs(361) <= not b;
    outputs(362) <= not a;
    outputs(363) <= not b;
    outputs(364) <= not (a xor b);
    outputs(365) <= not b;
    outputs(366) <= a;
    outputs(367) <= a;
    outputs(368) <= b and not a;
    outputs(369) <= a or b;
    outputs(370) <= not b;
    outputs(371) <= not (a xor b);
    outputs(372) <= not a;
    outputs(373) <= not a;
    outputs(374) <= a xor b;
    outputs(375) <= a and b;
    outputs(376) <= not b;
    outputs(377) <= b;
    outputs(378) <= not a;
    outputs(379) <= not (a or b);
    outputs(380) <= not a or b;
    outputs(381) <= a and b;
    outputs(382) <= not a;
    outputs(383) <= not (a xor b);
    outputs(384) <= not (a xor b);
    outputs(385) <= b;
    outputs(386) <= a xor b;
    outputs(387) <= not a or b;
    outputs(388) <= a xor b;
    outputs(389) <= b and not a;
    outputs(390) <= a;
    outputs(391) <= a xor b;
    outputs(392) <= not b;
    outputs(393) <= not a;
    outputs(394) <= not (a or b);
    outputs(395) <= b;
    outputs(396) <= a xor b;
    outputs(397) <= not b;
    outputs(398) <= a;
    outputs(399) <= a xor b;
    outputs(400) <= b;
    outputs(401) <= not b;
    outputs(402) <= a;
    outputs(403) <= a and b;
    outputs(404) <= a xor b;
    outputs(405) <= b;
    outputs(406) <= a xor b;
    outputs(407) <= a xor b;
    outputs(408) <= b;
    outputs(409) <= not a;
    outputs(410) <= not (a or b);
    outputs(411) <= not (a or b);
    outputs(412) <= b and not a;
    outputs(413) <= not a;
    outputs(414) <= b;
    outputs(415) <= not (a xor b);
    outputs(416) <= a xor b;
    outputs(417) <= not a;
    outputs(418) <= not b;
    outputs(419) <= b;
    outputs(420) <= a xor b;
    outputs(421) <= not (a and b);
    outputs(422) <= a xor b;
    outputs(423) <= a and not b;
    outputs(424) <= not a;
    outputs(425) <= not (a xor b);
    outputs(426) <= not b;
    outputs(427) <= a xor b;
    outputs(428) <= b;
    outputs(429) <= not b;
    outputs(430) <= a xor b;
    outputs(431) <= not b or a;
    outputs(432) <= not a;
    outputs(433) <= not (a xor b);
    outputs(434) <= b and not a;
    outputs(435) <= not a;
    outputs(436) <= not (a xor b);
    outputs(437) <= not b;
    outputs(438) <= b;
    outputs(439) <= a xor b;
    outputs(440) <= b;
    outputs(441) <= b;
    outputs(442) <= a;
    outputs(443) <= not b;
    outputs(444) <= not b;
    outputs(445) <= a;
    outputs(446) <= b;
    outputs(447) <= not b;
    outputs(448) <= not b or a;
    outputs(449) <= not b;
    outputs(450) <= a xor b;
    outputs(451) <= not a;
    outputs(452) <= not a;
    outputs(453) <= a xor b;
    outputs(454) <= a;
    outputs(455) <= b and not a;
    outputs(456) <= b;
    outputs(457) <= a or b;
    outputs(458) <= not (a or b);
    outputs(459) <= b;
    outputs(460) <= a xor b;
    outputs(461) <= a and b;
    outputs(462) <= a and b;
    outputs(463) <= not a;
    outputs(464) <= not (a xor b);
    outputs(465) <= a and not b;
    outputs(466) <= a;
    outputs(467) <= not (a and b);
    outputs(468) <= not a;
    outputs(469) <= a;
    outputs(470) <= a xor b;
    outputs(471) <= not (a xor b);
    outputs(472) <= a;
    outputs(473) <= b and not a;
    outputs(474) <= a xor b;
    outputs(475) <= a xor b;
    outputs(476) <= not b or a;
    outputs(477) <= not b;
    outputs(478) <= b;
    outputs(479) <= b;
    outputs(480) <= not (a xor b);
    outputs(481) <= not b;
    outputs(482) <= not a;
    outputs(483) <= not b;
    outputs(484) <= b;
    outputs(485) <= not a or b;
    outputs(486) <= not (a xor b);
    outputs(487) <= not b;
    outputs(488) <= a;
    outputs(489) <= a and not b;
    outputs(490) <= not (a xor b);
    outputs(491) <= a and not b;
    outputs(492) <= not a;
    outputs(493) <= a and not b;
    outputs(494) <= not a;
    outputs(495) <= a xor b;
    outputs(496) <= not b;
    outputs(497) <= not b or a;
    outputs(498) <= a and b;
    outputs(499) <= not (a xor b);
    outputs(500) <= not (a xor b);
    outputs(501) <= a xor b;
    outputs(502) <= a or b;
    outputs(503) <= not b;
    outputs(504) <= not (a xor b);
    outputs(505) <= a;
    outputs(506) <= a;
    outputs(507) <= a;
    outputs(508) <= b and not a;
    outputs(509) <= not b;
    outputs(510) <= b and not a;
    outputs(511) <= not (a or b);
    outputs(512) <= not b;
    outputs(513) <= a xor b;
    outputs(514) <= not a;
    outputs(515) <= a;
    outputs(516) <= a or b;
    outputs(517) <= a xor b;
    outputs(518) <= a;
    outputs(519) <= a;
    outputs(520) <= not (a xor b);
    outputs(521) <= not (a xor b);
    outputs(522) <= a;
    outputs(523) <= not (a xor b);
    outputs(524) <= not a;
    outputs(525) <= a;
    outputs(526) <= not a;
    outputs(527) <= a;
    outputs(528) <= not a;
    outputs(529) <= a and not b;
    outputs(530) <= not b;
    outputs(531) <= not b;
    outputs(532) <= a xor b;
    outputs(533) <= a;
    outputs(534) <= a and not b;
    outputs(535) <= not (a xor b);
    outputs(536) <= not a;
    outputs(537) <= a xor b;
    outputs(538) <= not a or b;
    outputs(539) <= a xor b;
    outputs(540) <= not a or b;
    outputs(541) <= not (a or b);
    outputs(542) <= not (a xor b);
    outputs(543) <= not b;
    outputs(544) <= not (a xor b);
    outputs(545) <= not b;
    outputs(546) <= a xor b;
    outputs(547) <= a xor b;
    outputs(548) <= a;
    outputs(549) <= not (a xor b);
    outputs(550) <= a;
    outputs(551) <= b;
    outputs(552) <= a xor b;
    outputs(553) <= a;
    outputs(554) <= not (a xor b);
    outputs(555) <= not (a xor b);
    outputs(556) <= not (a or b);
    outputs(557) <= a;
    outputs(558) <= b;
    outputs(559) <= not b;
    outputs(560) <= a xor b;
    outputs(561) <= not b or a;
    outputs(562) <= not (a xor b);
    outputs(563) <= not a;
    outputs(564) <= not (a and b);
    outputs(565) <= a xor b;
    outputs(566) <= b;
    outputs(567) <= a;
    outputs(568) <= not (a xor b);
    outputs(569) <= a xor b;
    outputs(570) <= b;
    outputs(571) <= b;
    outputs(572) <= a xor b;
    outputs(573) <= a xor b;
    outputs(574) <= not b or a;
    outputs(575) <= not a;
    outputs(576) <= a;
    outputs(577) <= not b;
    outputs(578) <= a or b;
    outputs(579) <= not a;
    outputs(580) <= a;
    outputs(581) <= not b;
    outputs(582) <= b;
    outputs(583) <= a and b;
    outputs(584) <= not (a xor b);
    outputs(585) <= not (a xor b);
    outputs(586) <= not a or b;
    outputs(587) <= not a;
    outputs(588) <= a;
    outputs(589) <= not b;
    outputs(590) <= not a;
    outputs(591) <= not (a xor b);
    outputs(592) <= b;
    outputs(593) <= not b;
    outputs(594) <= not (a xor b);
    outputs(595) <= a or b;
    outputs(596) <= not (a xor b);
    outputs(597) <= b;
    outputs(598) <= not (a xor b);
    outputs(599) <= not a;
    outputs(600) <= a;
    outputs(601) <= a;
    outputs(602) <= b;
    outputs(603) <= not (a xor b);
    outputs(604) <= not (a or b);
    outputs(605) <= not a;
    outputs(606) <= a;
    outputs(607) <= a xor b;
    outputs(608) <= not a;
    outputs(609) <= not b;
    outputs(610) <= not a;
    outputs(611) <= b;
    outputs(612) <= not (a xor b);
    outputs(613) <= a xor b;
    outputs(614) <= not (a xor b);
    outputs(615) <= a and not b;
    outputs(616) <= not b;
    outputs(617) <= a xor b;
    outputs(618) <= not (a xor b);
    outputs(619) <= not b;
    outputs(620) <= a;
    outputs(621) <= not (a xor b);
    outputs(622) <= not b;
    outputs(623) <= a and b;
    outputs(624) <= a;
    outputs(625) <= not (a or b);
    outputs(626) <= not (a xor b);
    outputs(627) <= not b;
    outputs(628) <= b;
    outputs(629) <= not a;
    outputs(630) <= b;
    outputs(631) <= b and not a;
    outputs(632) <= not (a xor b);
    outputs(633) <= a;
    outputs(634) <= not a or b;
    outputs(635) <= a xor b;
    outputs(636) <= b and not a;
    outputs(637) <= not a;
    outputs(638) <= a xor b;
    outputs(639) <= not (a xor b);
    outputs(640) <= b;
    outputs(641) <= not a;
    outputs(642) <= not a or b;
    outputs(643) <= not a;
    outputs(644) <= a;
    outputs(645) <= a xor b;
    outputs(646) <= not a;
    outputs(647) <= b and not a;
    outputs(648) <= a;
    outputs(649) <= not (a xor b);
    outputs(650) <= b;
    outputs(651) <= a;
    outputs(652) <= b;
    outputs(653) <= not b;
    outputs(654) <= not (a xor b);
    outputs(655) <= not a;
    outputs(656) <= a;
    outputs(657) <= not (a xor b);
    outputs(658) <= a;
    outputs(659) <= not a;
    outputs(660) <= a;
    outputs(661) <= not b;
    outputs(662) <= not a;
    outputs(663) <= b;
    outputs(664) <= not a;
    outputs(665) <= b;
    outputs(666) <= a and not b;
    outputs(667) <= not (a xor b);
    outputs(668) <= a;
    outputs(669) <= not a;
    outputs(670) <= b;
    outputs(671) <= a;
    outputs(672) <= a;
    outputs(673) <= a xor b;
    outputs(674) <= a xor b;
    outputs(675) <= not b;
    outputs(676) <= not b;
    outputs(677) <= a;
    outputs(678) <= not a;
    outputs(679) <= not b;
    outputs(680) <= not a;
    outputs(681) <= not b;
    outputs(682) <= b;
    outputs(683) <= b;
    outputs(684) <= not a;
    outputs(685) <= not (a xor b);
    outputs(686) <= not (a xor b);
    outputs(687) <= a xor b;
    outputs(688) <= a;
    outputs(689) <= not (a or b);
    outputs(690) <= a xor b;
    outputs(691) <= b;
    outputs(692) <= not a;
    outputs(693) <= not (a xor b);
    outputs(694) <= not (a xor b);
    outputs(695) <= not b;
    outputs(696) <= b and not a;
    outputs(697) <= a;
    outputs(698) <= a xor b;
    outputs(699) <= not b;
    outputs(700) <= not (a xor b);
    outputs(701) <= not (a xor b);
    outputs(702) <= a and not b;
    outputs(703) <= a xor b;
    outputs(704) <= not (a xor b);
    outputs(705) <= not (a xor b);
    outputs(706) <= b;
    outputs(707) <= a;
    outputs(708) <= a;
    outputs(709) <= not (a xor b);
    outputs(710) <= a xor b;
    outputs(711) <= not a;
    outputs(712) <= a;
    outputs(713) <= not (a xor b);
    outputs(714) <= not (a xor b);
    outputs(715) <= not (a xor b);
    outputs(716) <= not a;
    outputs(717) <= not a;
    outputs(718) <= b;
    outputs(719) <= not a;
    outputs(720) <= not (a xor b);
    outputs(721) <= not (a xor b);
    outputs(722) <= not a;
    outputs(723) <= not (a xor b);
    outputs(724) <= not (a xor b);
    outputs(725) <= a xor b;
    outputs(726) <= b;
    outputs(727) <= b;
    outputs(728) <= a or b;
    outputs(729) <= b and not a;
    outputs(730) <= a;
    outputs(731) <= not b;
    outputs(732) <= b and not a;
    outputs(733) <= not b;
    outputs(734) <= not a or b;
    outputs(735) <= a xor b;
    outputs(736) <= a or b;
    outputs(737) <= b;
    outputs(738) <= not b or a;
    outputs(739) <= not a;
    outputs(740) <= not a;
    outputs(741) <= a xor b;
    outputs(742) <= a xor b;
    outputs(743) <= not (a or b);
    outputs(744) <= a xor b;
    outputs(745) <= a xor b;
    outputs(746) <= not b;
    outputs(747) <= a;
    outputs(748) <= a xor b;
    outputs(749) <= not (a xor b);
    outputs(750) <= not a;
    outputs(751) <= not a;
    outputs(752) <= a xor b;
    outputs(753) <= b;
    outputs(754) <= a or b;
    outputs(755) <= a and not b;
    outputs(756) <= a;
    outputs(757) <= not (a xor b);
    outputs(758) <= a xor b;
    outputs(759) <= a and b;
    outputs(760) <= not a;
    outputs(761) <= not (a xor b);
    outputs(762) <= not a or b;
    outputs(763) <= not (a or b);
    outputs(764) <= not (a and b);
    outputs(765) <= not a or b;
    outputs(766) <= b;
    outputs(767) <= not a;
    outputs(768) <= a;
    outputs(769) <= not a;
    outputs(770) <= a xor b;
    outputs(771) <= b;
    outputs(772) <= b;
    outputs(773) <= not (a xor b);
    outputs(774) <= a;
    outputs(775) <= not (a or b);
    outputs(776) <= not a;
    outputs(777) <= not b or a;
    outputs(778) <= a;
    outputs(779) <= b;
    outputs(780) <= b;
    outputs(781) <= not b;
    outputs(782) <= a;
    outputs(783) <= not (a or b);
    outputs(784) <= b;
    outputs(785) <= b and not a;
    outputs(786) <= a;
    outputs(787) <= a xor b;
    outputs(788) <= a;
    outputs(789) <= a xor b;
    outputs(790) <= not (a and b);
    outputs(791) <= a;
    outputs(792) <= not (a or b);
    outputs(793) <= a;
    outputs(794) <= not b;
    outputs(795) <= a;
    outputs(796) <= not (a xor b);
    outputs(797) <= a and b;
    outputs(798) <= not (a xor b);
    outputs(799) <= not (a xor b);
    outputs(800) <= a or b;
    outputs(801) <= a;
    outputs(802) <= not (a xor b);
    outputs(803) <= not b;
    outputs(804) <= a;
    outputs(805) <= not (a xor b);
    outputs(806) <= b;
    outputs(807) <= not a;
    outputs(808) <= not (a xor b);
    outputs(809) <= a;
    outputs(810) <= not a;
    outputs(811) <= a and not b;
    outputs(812) <= b and not a;
    outputs(813) <= b;
    outputs(814) <= b;
    outputs(815) <= not (a xor b);
    outputs(816) <= a;
    outputs(817) <= a;
    outputs(818) <= a xor b;
    outputs(819) <= b;
    outputs(820) <= not b;
    outputs(821) <= not (a xor b);
    outputs(822) <= a and b;
    outputs(823) <= a;
    outputs(824) <= a;
    outputs(825) <= b and not a;
    outputs(826) <= a xor b;
    outputs(827) <= a;
    outputs(828) <= a xor b;
    outputs(829) <= a;
    outputs(830) <= a xor b;
    outputs(831) <= not b;
    outputs(832) <= a or b;
    outputs(833) <= not b;
    outputs(834) <= not (a and b);
    outputs(835) <= a;
    outputs(836) <= a xor b;
    outputs(837) <= a xor b;
    outputs(838) <= not (a and b);
    outputs(839) <= a and b;
    outputs(840) <= not (a xor b);
    outputs(841) <= not b;
    outputs(842) <= not b;
    outputs(843) <= not (a xor b);
    outputs(844) <= a;
    outputs(845) <= not b;
    outputs(846) <= not b;
    outputs(847) <= not b;
    outputs(848) <= not b;
    outputs(849) <= not b;
    outputs(850) <= not a;
    outputs(851) <= a and b;
    outputs(852) <= not b or a;
    outputs(853) <= not (a xor b);
    outputs(854) <= not b;
    outputs(855) <= a;
    outputs(856) <= b and not a;
    outputs(857) <= b;
    outputs(858) <= not b;
    outputs(859) <= not (a xor b);
    outputs(860) <= b and not a;
    outputs(861) <= a xor b;
    outputs(862) <= not (a xor b);
    outputs(863) <= a;
    outputs(864) <= not a;
    outputs(865) <= a;
    outputs(866) <= a;
    outputs(867) <= a and not b;
    outputs(868) <= not a;
    outputs(869) <= b;
    outputs(870) <= a;
    outputs(871) <= not a;
    outputs(872) <= not a;
    outputs(873) <= not b;
    outputs(874) <= a or b;
    outputs(875) <= not b;
    outputs(876) <= a and b;
    outputs(877) <= not (a xor b);
    outputs(878) <= a and b;
    outputs(879) <= a xor b;
    outputs(880) <= b;
    outputs(881) <= a xor b;
    outputs(882) <= a and not b;
    outputs(883) <= a;
    outputs(884) <= not b;
    outputs(885) <= not b or a;
    outputs(886) <= a;
    outputs(887) <= b and not a;
    outputs(888) <= not (a xor b);
    outputs(889) <= a xor b;
    outputs(890) <= not (a and b);
    outputs(891) <= a xor b;
    outputs(892) <= b;
    outputs(893) <= b;
    outputs(894) <= not a or b;
    outputs(895) <= b;
    outputs(896) <= a;
    outputs(897) <= not (a or b);
    outputs(898) <= b;
    outputs(899) <= a and not b;
    outputs(900) <= a xor b;
    outputs(901) <= not b;
    outputs(902) <= not b or a;
    outputs(903) <= not (a xor b);
    outputs(904) <= not a;
    outputs(905) <= not a or b;
    outputs(906) <= a xor b;
    outputs(907) <= a;
    outputs(908) <= a;
    outputs(909) <= b;
    outputs(910) <= b and not a;
    outputs(911) <= not (a xor b);
    outputs(912) <= not (a xor b);
    outputs(913) <= b;
    outputs(914) <= b;
    outputs(915) <= b;
    outputs(916) <= not b;
    outputs(917) <= a xor b;
    outputs(918) <= 1'b0;
    outputs(919) <= a;
    outputs(920) <= not a;
    outputs(921) <= not b;
    outputs(922) <= not (a or b);
    outputs(923) <= a xor b;
    outputs(924) <= a xor b;
    outputs(925) <= not a or b;
    outputs(926) <= a xor b;
    outputs(927) <= a xor b;
    outputs(928) <= a xor b;
    outputs(929) <= a xor b;
    outputs(930) <= a xor b;
    outputs(931) <= not (a xor b);
    outputs(932) <= a;
    outputs(933) <= a;
    outputs(934) <= not b;
    outputs(935) <= b;
    outputs(936) <= not b;
    outputs(937) <= a xor b;
    outputs(938) <= a or b;
    outputs(939) <= b and not a;
    outputs(940) <= a and b;
    outputs(941) <= a;
    outputs(942) <= b and not a;
    outputs(943) <= not (a xor b);
    outputs(944) <= b;
    outputs(945) <= not (a xor b);
    outputs(946) <= a xor b;
    outputs(947) <= a xor b;
    outputs(948) <= not a;
    outputs(949) <= a xor b;
    outputs(950) <= not a;
    outputs(951) <= not (a xor b);
    outputs(952) <= not b;
    outputs(953) <= not a;
    outputs(954) <= b;
    outputs(955) <= b;
    outputs(956) <= not a or b;
    outputs(957) <= b;
    outputs(958) <= a xor b;
    outputs(959) <= b;
    outputs(960) <= not (a xor b);
    outputs(961) <= a;
    outputs(962) <= not (a xor b);
    outputs(963) <= a;
    outputs(964) <= b;
    outputs(965) <= not (a xor b);
    outputs(966) <= a xor b;
    outputs(967) <= a and not b;
    outputs(968) <= not (a xor b);
    outputs(969) <= a xor b;
    outputs(970) <= not a;
    outputs(971) <= not a;
    outputs(972) <= not (a xor b);
    outputs(973) <= not (a or b);
    outputs(974) <= not b;
    outputs(975) <= not a;
    outputs(976) <= not b;
    outputs(977) <= not b or a;
    outputs(978) <= not b;
    outputs(979) <= a;
    outputs(980) <= not b;
    outputs(981) <= a;
    outputs(982) <= not b;
    outputs(983) <= b and not a;
    outputs(984) <= not a;
    outputs(985) <= not a;
    outputs(986) <= not b;
    outputs(987) <= a;
    outputs(988) <= b;
    outputs(989) <= a and not b;
    outputs(990) <= a;
    outputs(991) <= not (a xor b);
    outputs(992) <= b;
    outputs(993) <= not (a xor b);
    outputs(994) <= a and not b;
    outputs(995) <= not a;
    outputs(996) <= a;
    outputs(997) <= not (a and b);
    outputs(998) <= a and b;
    outputs(999) <= not (a xor b);
    outputs(1000) <= not a;
    outputs(1001) <= not (a xor b);
    outputs(1002) <= not (a and b);
    outputs(1003) <= a or b;
    outputs(1004) <= b;
    outputs(1005) <= not a;
    outputs(1006) <= not b;
    outputs(1007) <= not (a xor b);
    outputs(1008) <= b;
    outputs(1009) <= b;
    outputs(1010) <= a and not b;
    outputs(1011) <= a xor b;
    outputs(1012) <= a xor b;
    outputs(1013) <= a;
    outputs(1014) <= a and b;
    outputs(1015) <= a xor b;
    outputs(1016) <= not (a xor b);
    outputs(1017) <= not (a xor b);
    outputs(1018) <= a xor b;
    outputs(1019) <= a;
    outputs(1020) <= not a;
    outputs(1021) <= not (a xor b);
    outputs(1022) <= a;
    outputs(1023) <= not b;
    outputs(1024) <= not (a and b);
    outputs(1025) <= not b;
    outputs(1026) <= not a;
    outputs(1027) <= not b;
    outputs(1028) <= not b;
    outputs(1029) <= a;
    outputs(1030) <= b;
    outputs(1031) <= a xor b;
    outputs(1032) <= a and not b;
    outputs(1033) <= a and b;
    outputs(1034) <= not (a or b);
    outputs(1035) <= not (a or b);
    outputs(1036) <= not (a xor b);
    outputs(1037) <= b;
    outputs(1038) <= a xor b;
    outputs(1039) <= not (a xor b);
    outputs(1040) <= not b;
    outputs(1041) <= a and b;
    outputs(1042) <= not (a xor b);
    outputs(1043) <= a and b;
    outputs(1044) <= a;
    outputs(1045) <= a and b;
    outputs(1046) <= a;
    outputs(1047) <= b and not a;
    outputs(1048) <= 1'b0;
    outputs(1049) <= not (a or b);
    outputs(1050) <= a and b;
    outputs(1051) <= a;
    outputs(1052) <= a xor b;
    outputs(1053) <= a xor b;
    outputs(1054) <= not (a xor b);
    outputs(1055) <= b;
    outputs(1056) <= a xor b;
    outputs(1057) <= a;
    outputs(1058) <= a xor b;
    outputs(1059) <= b;
    outputs(1060) <= a xor b;
    outputs(1061) <= not (a xor b);
    outputs(1062) <= a xor b;
    outputs(1063) <= a xor b;
    outputs(1064) <= not b;
    outputs(1065) <= not b or a;
    outputs(1066) <= not (a or b);
    outputs(1067) <= not b;
    outputs(1068) <= a;
    outputs(1069) <= b;
    outputs(1070) <= b;
    outputs(1071) <= b;
    outputs(1072) <= b and not a;
    outputs(1073) <= not b;
    outputs(1074) <= not a or b;
    outputs(1075) <= a and b;
    outputs(1076) <= not (a xor b);
    outputs(1077) <= not b;
    outputs(1078) <= not b;
    outputs(1079) <= b;
    outputs(1080) <= b and not a;
    outputs(1081) <= a xor b;
    outputs(1082) <= not b;
    outputs(1083) <= not (a xor b);
    outputs(1084) <= b and not a;
    outputs(1085) <= b and not a;
    outputs(1086) <= not a;
    outputs(1087) <= not (a xor b);
    outputs(1088) <= not a;
    outputs(1089) <= a and not b;
    outputs(1090) <= not (a xor b);
    outputs(1091) <= not (a xor b);
    outputs(1092) <= not a;
    outputs(1093) <= not b;
    outputs(1094) <= not a or b;
    outputs(1095) <= b;
    outputs(1096) <= a and not b;
    outputs(1097) <= a and b;
    outputs(1098) <= b and not a;
    outputs(1099) <= a;
    outputs(1100) <= not (a xor b);
    outputs(1101) <= not (a and b);
    outputs(1102) <= a xor b;
    outputs(1103) <= a xor b;
    outputs(1104) <= a xor b;
    outputs(1105) <= not (a and b);
    outputs(1106) <= a and not b;
    outputs(1107) <= b;
    outputs(1108) <= not (a and b);
    outputs(1109) <= a and b;
    outputs(1110) <= not (a or b);
    outputs(1111) <= b;
    outputs(1112) <= not (a xor b);
    outputs(1113) <= a xor b;
    outputs(1114) <= not b;
    outputs(1115) <= a xor b;
    outputs(1116) <= a;
    outputs(1117) <= a;
    outputs(1118) <= b and not a;
    outputs(1119) <= not (a or b);
    outputs(1120) <= b and not a;
    outputs(1121) <= b and not a;
    outputs(1122) <= not (a xor b);
    outputs(1123) <= a;
    outputs(1124) <= not (a xor b);
    outputs(1125) <= not (a or b);
    outputs(1126) <= a and b;
    outputs(1127) <= b;
    outputs(1128) <= b and not a;
    outputs(1129) <= not (a or b);
    outputs(1130) <= b;
    outputs(1131) <= a xor b;
    outputs(1132) <= a and not b;
    outputs(1133) <= not (a or b);
    outputs(1134) <= a and not b;
    outputs(1135) <= a xor b;
    outputs(1136) <= b;
    outputs(1137) <= b;
    outputs(1138) <= not b;
    outputs(1139) <= a;
    outputs(1140) <= not b or a;
    outputs(1141) <= a;
    outputs(1142) <= not (a or b);
    outputs(1143) <= a and b;
    outputs(1144) <= a xor b;
    outputs(1145) <= a;
    outputs(1146) <= not (a xor b);
    outputs(1147) <= a or b;
    outputs(1148) <= not b;
    outputs(1149) <= a xor b;
    outputs(1150) <= not (a xor b);
    outputs(1151) <= a;
    outputs(1152) <= not (a xor b);
    outputs(1153) <= not b;
    outputs(1154) <= b and not a;
    outputs(1155) <= not a;
    outputs(1156) <= not a or b;
    outputs(1157) <= a and not b;
    outputs(1158) <= a and b;
    outputs(1159) <= not a or b;
    outputs(1160) <= a and b;
    outputs(1161) <= a and not b;
    outputs(1162) <= a xor b;
    outputs(1163) <= a;
    outputs(1164) <= a and not b;
    outputs(1165) <= a xor b;
    outputs(1166) <= not (a and b);
    outputs(1167) <= a xor b;
    outputs(1168) <= b;
    outputs(1169) <= a;
    outputs(1170) <= a and b;
    outputs(1171) <= not a;
    outputs(1172) <= b;
    outputs(1173) <= not a;
    outputs(1174) <= a xor b;
    outputs(1175) <= a xor b;
    outputs(1176) <= not a;
    outputs(1177) <= not (a or b);
    outputs(1178) <= a xor b;
    outputs(1179) <= a and not b;
    outputs(1180) <= not b;
    outputs(1181) <= a and not b;
    outputs(1182) <= b;
    outputs(1183) <= not (a xor b);
    outputs(1184) <= not (a xor b);
    outputs(1185) <= b and not a;
    outputs(1186) <= not a;
    outputs(1187) <= a;
    outputs(1188) <= b;
    outputs(1189) <= not b;
    outputs(1190) <= not a or b;
    outputs(1191) <= not a;
    outputs(1192) <= not b;
    outputs(1193) <= a xor b;
    outputs(1194) <= not (a xor b);
    outputs(1195) <= not b;
    outputs(1196) <= not b;
    outputs(1197) <= not a;
    outputs(1198) <= a;
    outputs(1199) <= not (a or b);
    outputs(1200) <= not a;
    outputs(1201) <= a;
    outputs(1202) <= b and not a;
    outputs(1203) <= not b;
    outputs(1204) <= a and b;
    outputs(1205) <= a xor b;
    outputs(1206) <= b;
    outputs(1207) <= a xor b;
    outputs(1208) <= b and not a;
    outputs(1209) <= a xor b;
    outputs(1210) <= b;
    outputs(1211) <= not (a xor b);
    outputs(1212) <= not (a xor b);
    outputs(1213) <= a and not b;
    outputs(1214) <= not a;
    outputs(1215) <= a and not b;
    outputs(1216) <= b;
    outputs(1217) <= not (a xor b);
    outputs(1218) <= a;
    outputs(1219) <= a and not b;
    outputs(1220) <= a;
    outputs(1221) <= not (a xor b);
    outputs(1222) <= b and not a;
    outputs(1223) <= not (a xor b);
    outputs(1224) <= not (a or b);
    outputs(1225) <= a xor b;
    outputs(1226) <= a;
    outputs(1227) <= 1'b0;
    outputs(1228) <= not b;
    outputs(1229) <= not a;
    outputs(1230) <= not b;
    outputs(1231) <= a xor b;
    outputs(1232) <= a xor b;
    outputs(1233) <= not (a xor b);
    outputs(1234) <= b;
    outputs(1235) <= not (a or b);
    outputs(1236) <= a xor b;
    outputs(1237) <= a and b;
    outputs(1238) <= a xor b;
    outputs(1239) <= not a;
    outputs(1240) <= b and not a;
    outputs(1241) <= b;
    outputs(1242) <= a and not b;
    outputs(1243) <= b and not a;
    outputs(1244) <= a xor b;
    outputs(1245) <= 1'b0;
    outputs(1246) <= not b;
    outputs(1247) <= not b;
    outputs(1248) <= not b;
    outputs(1249) <= a and b;
    outputs(1250) <= a xor b;
    outputs(1251) <= 1'b0;
    outputs(1252) <= not b;
    outputs(1253) <= a xor b;
    outputs(1254) <= b and not a;
    outputs(1255) <= a;
    outputs(1256) <= a and b;
    outputs(1257) <= not (a and b);
    outputs(1258) <= b and not a;
    outputs(1259) <= b;
    outputs(1260) <= a xor b;
    outputs(1261) <= not b;
    outputs(1262) <= a xor b;
    outputs(1263) <= a;
    outputs(1264) <= b;
    outputs(1265) <= a and b;
    outputs(1266) <= a xor b;
    outputs(1267) <= not (a xor b);
    outputs(1268) <= a and b;
    outputs(1269) <= not a;
    outputs(1270) <= not a;
    outputs(1271) <= not (a xor b);
    outputs(1272) <= not (a xor b);
    outputs(1273) <= not b;
    outputs(1274) <= not (a or b);
    outputs(1275) <= not b;
    outputs(1276) <= not b;
    outputs(1277) <= not (a xor b);
    outputs(1278) <= not (a xor b);
    outputs(1279) <= a xor b;
    outputs(1280) <= not (a xor b);
    outputs(1281) <= a;
    outputs(1282) <= a;
    outputs(1283) <= b;
    outputs(1284) <= a xor b;
    outputs(1285) <= not a;
    outputs(1286) <= not (a xor b);
    outputs(1287) <= a;
    outputs(1288) <= not (a xor b);
    outputs(1289) <= b;
    outputs(1290) <= not (a or b);
    outputs(1291) <= not (a or b);
    outputs(1292) <= not (a or b);
    outputs(1293) <= b and not a;
    outputs(1294) <= b and not a;
    outputs(1295) <= not a;
    outputs(1296) <= a;
    outputs(1297) <= a xor b;
    outputs(1298) <= not (a xor b);
    outputs(1299) <= a;
    outputs(1300) <= not b;
    outputs(1301) <= not b;
    outputs(1302) <= b;
    outputs(1303) <= a xor b;
    outputs(1304) <= b;
    outputs(1305) <= not (a or b);
    outputs(1306) <= b and not a;
    outputs(1307) <= a;
    outputs(1308) <= a and b;
    outputs(1309) <= b;
    outputs(1310) <= not a;
    outputs(1311) <= not (a xor b);
    outputs(1312) <= a and not b;
    outputs(1313) <= not a;
    outputs(1314) <= b;
    outputs(1315) <= not b;
    outputs(1316) <= a and not b;
    outputs(1317) <= not a;
    outputs(1318) <= b and not a;
    outputs(1319) <= b;
    outputs(1320) <= a;
    outputs(1321) <= not a;
    outputs(1322) <= not (a xor b);
    outputs(1323) <= not a;
    outputs(1324) <= not (a and b);
    outputs(1325) <= not a;
    outputs(1326) <= not b;
    outputs(1327) <= b;
    outputs(1328) <= a;
    outputs(1329) <= a and b;
    outputs(1330) <= b;
    outputs(1331) <= not b;
    outputs(1332) <= not a;
    outputs(1333) <= a xor b;
    outputs(1334) <= a;
    outputs(1335) <= a xor b;
    outputs(1336) <= not (a xor b);
    outputs(1337) <= not (a or b);
    outputs(1338) <= not b;
    outputs(1339) <= a and b;
    outputs(1340) <= a xor b;
    outputs(1341) <= not (a xor b);
    outputs(1342) <= not (a xor b);
    outputs(1343) <= a;
    outputs(1344) <= b;
    outputs(1345) <= a xor b;
    outputs(1346) <= a and not b;
    outputs(1347) <= not (a and b);
    outputs(1348) <= b and not a;
    outputs(1349) <= not a or b;
    outputs(1350) <= a xor b;
    outputs(1351) <= not (a xor b);
    outputs(1352) <= not (a xor b);
    outputs(1353) <= not b;
    outputs(1354) <= not a;
    outputs(1355) <= b and not a;
    outputs(1356) <= not a;
    outputs(1357) <= not (a xor b);
    outputs(1358) <= not b;
    outputs(1359) <= a xor b;
    outputs(1360) <= b;
    outputs(1361) <= not (a or b);
    outputs(1362) <= not (a or b);
    outputs(1363) <= a xor b;
    outputs(1364) <= a xor b;
    outputs(1365) <= 1'b0;
    outputs(1366) <= not a;
    outputs(1367) <= a;
    outputs(1368) <= not (a xor b);
    outputs(1369) <= a xor b;
    outputs(1370) <= not b;
    outputs(1371) <= a and b;
    outputs(1372) <= a;
    outputs(1373) <= a;
    outputs(1374) <= not (a xor b);
    outputs(1375) <= not (a or b);
    outputs(1376) <= a and not b;
    outputs(1377) <= not (a xor b);
    outputs(1378) <= b;
    outputs(1379) <= a;
    outputs(1380) <= not b;
    outputs(1381) <= b and not a;
    outputs(1382) <= not a;
    outputs(1383) <= not b;
    outputs(1384) <= not (a xor b);
    outputs(1385) <= not a;
    outputs(1386) <= not b;
    outputs(1387) <= not (a or b);
    outputs(1388) <= not a;
    outputs(1389) <= not (a xor b);
    outputs(1390) <= a xor b;
    outputs(1391) <= b;
    outputs(1392) <= not (a xor b);
    outputs(1393) <= b;
    outputs(1394) <= not (a or b);
    outputs(1395) <= not (a xor b);
    outputs(1396) <= not b;
    outputs(1397) <= a;
    outputs(1398) <= a xor b;
    outputs(1399) <= b and not a;
    outputs(1400) <= not (a xor b);
    outputs(1401) <= b;
    outputs(1402) <= a and not b;
    outputs(1403) <= a;
    outputs(1404) <= not b;
    outputs(1405) <= a and b;
    outputs(1406) <= not (a xor b);
    outputs(1407) <= a xor b;
    outputs(1408) <= not (a or b);
    outputs(1409) <= a and b;
    outputs(1410) <= not b;
    outputs(1411) <= not (a xor b);
    outputs(1412) <= a and b;
    outputs(1413) <= a xor b;
    outputs(1414) <= not a or b;
    outputs(1415) <= a xor b;
    outputs(1416) <= not (a or b);
    outputs(1417) <= a xor b;
    outputs(1418) <= not a;
    outputs(1419) <= a or b;
    outputs(1420) <= not (a xor b);
    outputs(1421) <= not b;
    outputs(1422) <= a and not b;
    outputs(1423) <= a and b;
    outputs(1424) <= b and not a;
    outputs(1425) <= a xor b;
    outputs(1426) <= a and not b;
    outputs(1427) <= a xor b;
    outputs(1428) <= a;
    outputs(1429) <= not b;
    outputs(1430) <= not b;
    outputs(1431) <= not (a xor b);
    outputs(1432) <= a or b;
    outputs(1433) <= a xor b;
    outputs(1434) <= b and not a;
    outputs(1435) <= not (a or b);
    outputs(1436) <= not (a or b);
    outputs(1437) <= a and b;
    outputs(1438) <= a and not b;
    outputs(1439) <= not (a xor b);
    outputs(1440) <= not (a xor b);
    outputs(1441) <= b;
    outputs(1442) <= not a;
    outputs(1443) <= not a;
    outputs(1444) <= not b or a;
    outputs(1445) <= a xor b;
    outputs(1446) <= b;
    outputs(1447) <= b;
    outputs(1448) <= not a;
    outputs(1449) <= a xor b;
    outputs(1450) <= not (a or b);
    outputs(1451) <= a xor b;
    outputs(1452) <= not a;
    outputs(1453) <= b and not a;
    outputs(1454) <= a xor b;
    outputs(1455) <= not a or b;
    outputs(1456) <= a xor b;
    outputs(1457) <= not (a xor b);
    outputs(1458) <= a xor b;
    outputs(1459) <= a;
    outputs(1460) <= a xor b;
    outputs(1461) <= b and not a;
    outputs(1462) <= b;
    outputs(1463) <= b and not a;
    outputs(1464) <= b;
    outputs(1465) <= a xor b;
    outputs(1466) <= not b;
    outputs(1467) <= a;
    outputs(1468) <= not b;
    outputs(1469) <= not (a xor b);
    outputs(1470) <= not a;
    outputs(1471) <= not b or a;
    outputs(1472) <= a and not b;
    outputs(1473) <= b;
    outputs(1474) <= a xor b;
    outputs(1475) <= not b;
    outputs(1476) <= not (a xor b);
    outputs(1477) <= b;
    outputs(1478) <= not (a and b);
    outputs(1479) <= not b;
    outputs(1480) <= a and not b;
    outputs(1481) <= not b;
    outputs(1482) <= a and b;
    outputs(1483) <= not a;
    outputs(1484) <= not a;
    outputs(1485) <= not b;
    outputs(1486) <= not a;
    outputs(1487) <= a;
    outputs(1488) <= not b;
    outputs(1489) <= a xor b;
    outputs(1490) <= not (a xor b);
    outputs(1491) <= not a;
    outputs(1492) <= not b;
    outputs(1493) <= not b;
    outputs(1494) <= b and not a;
    outputs(1495) <= not b;
    outputs(1496) <= a and b;
    outputs(1497) <= not (a xor b);
    outputs(1498) <= not (a xor b);
    outputs(1499) <= a;
    outputs(1500) <= b;
    outputs(1501) <= a xor b;
    outputs(1502) <= not (a xor b);
    outputs(1503) <= a xor b;
    outputs(1504) <= a;
    outputs(1505) <= not a or b;
    outputs(1506) <= a xor b;
    outputs(1507) <= not a;
    outputs(1508) <= not a;
    outputs(1509) <= b and not a;
    outputs(1510) <= a xor b;
    outputs(1511) <= not a;
    outputs(1512) <= a;
    outputs(1513) <= a xor b;
    outputs(1514) <= not a;
    outputs(1515) <= not b;
    outputs(1516) <= b;
    outputs(1517) <= b;
    outputs(1518) <= b and not a;
    outputs(1519) <= a and not b;
    outputs(1520) <= a xor b;
    outputs(1521) <= a and not b;
    outputs(1522) <= b;
    outputs(1523) <= b;
    outputs(1524) <= not b;
    outputs(1525) <= not (a xor b);
    outputs(1526) <= not b;
    outputs(1527) <= not (a xor b);
    outputs(1528) <= b and not a;
    outputs(1529) <= a and not b;
    outputs(1530) <= not (a xor b);
    outputs(1531) <= not (a or b);
    outputs(1532) <= a;
    outputs(1533) <= not (a or b);
    outputs(1534) <= a xor b;
    outputs(1535) <= b and not a;
    outputs(1536) <= not b;
    outputs(1537) <= not (a or b);
    outputs(1538) <= a and not b;
    outputs(1539) <= a and not b;
    outputs(1540) <= a or b;
    outputs(1541) <= a and b;
    outputs(1542) <= not b or a;
    outputs(1543) <= a;
    outputs(1544) <= not (a xor b);
    outputs(1545) <= not b;
    outputs(1546) <= a and b;
    outputs(1547) <= not (a xor b);
    outputs(1548) <= not b;
    outputs(1549) <= not a;
    outputs(1550) <= a and not b;
    outputs(1551) <= not (a xor b);
    outputs(1552) <= a;
    outputs(1553) <= not (a xor b);
    outputs(1554) <= not (a xor b);
    outputs(1555) <= a and not b;
    outputs(1556) <= a and not b;
    outputs(1557) <= a xor b;
    outputs(1558) <= a;
    outputs(1559) <= b;
    outputs(1560) <= a;
    outputs(1561) <= b and not a;
    outputs(1562) <= a and b;
    outputs(1563) <= not a;
    outputs(1564) <= b and not a;
    outputs(1565) <= a;
    outputs(1566) <= a and not b;
    outputs(1567) <= a and not b;
    outputs(1568) <= not (a and b);
    outputs(1569) <= not (a or b);
    outputs(1570) <= not (a or b);
    outputs(1571) <= b;
    outputs(1572) <= a;
    outputs(1573) <= not (a xor b);
    outputs(1574) <= a xor b;
    outputs(1575) <= a;
    outputs(1576) <= not (a xor b);
    outputs(1577) <= not (a xor b);
    outputs(1578) <= not (a or b);
    outputs(1579) <= not b;
    outputs(1580) <= not (a xor b);
    outputs(1581) <= a and not b;
    outputs(1582) <= a and b;
    outputs(1583) <= not b;
    outputs(1584) <= a and not b;
    outputs(1585) <= not a;
    outputs(1586) <= a xor b;
    outputs(1587) <= not (a xor b);
    outputs(1588) <= a xor b;
    outputs(1589) <= a xor b;
    outputs(1590) <= not (a and b);
    outputs(1591) <= not a;
    outputs(1592) <= b and not a;
    outputs(1593) <= b and not a;
    outputs(1594) <= a and b;
    outputs(1595) <= not (a or b);
    outputs(1596) <= not (a or b);
    outputs(1597) <= b;
    outputs(1598) <= b and not a;
    outputs(1599) <= a;
    outputs(1600) <= not (a xor b);
    outputs(1601) <= not (a or b);
    outputs(1602) <= b and not a;
    outputs(1603) <= a and not b;
    outputs(1604) <= b;
    outputs(1605) <= a and b;
    outputs(1606) <= not (a xor b);
    outputs(1607) <= a and b;
    outputs(1608) <= b;
    outputs(1609) <= not a;
    outputs(1610) <= b and not a;
    outputs(1611) <= not (a or b);
    outputs(1612) <= a;
    outputs(1613) <= a and b;
    outputs(1614) <= b and not a;
    outputs(1615) <= a xor b;
    outputs(1616) <= not (a xor b);
    outputs(1617) <= 1'b0;
    outputs(1618) <= not a;
    outputs(1619) <= not b;
    outputs(1620) <= not a;
    outputs(1621) <= not (a xor b);
    outputs(1622) <= a and not b;
    outputs(1623) <= a and not b;
    outputs(1624) <= not b;
    outputs(1625) <= not b;
    outputs(1626) <= not (a xor b);
    outputs(1627) <= a and b;
    outputs(1628) <= a;
    outputs(1629) <= a xor b;
    outputs(1630) <= a and b;
    outputs(1631) <= a and b;
    outputs(1632) <= not (a or b);
    outputs(1633) <= a;
    outputs(1634) <= not (a xor b);
    outputs(1635) <= a and b;
    outputs(1636) <= b;
    outputs(1637) <= a xor b;
    outputs(1638) <= a xor b;
    outputs(1639) <= b and not a;
    outputs(1640) <= a and b;
    outputs(1641) <= a xor b;
    outputs(1642) <= b and not a;
    outputs(1643) <= a xor b;
    outputs(1644) <= not (a or b);
    outputs(1645) <= b;
    outputs(1646) <= b;
    outputs(1647) <= b;
    outputs(1648) <= a and b;
    outputs(1649) <= a and b;
    outputs(1650) <= a and b;
    outputs(1651) <= not (a xor b);
    outputs(1652) <= not (a xor b);
    outputs(1653) <= not b;
    outputs(1654) <= not a;
    outputs(1655) <= a xor b;
    outputs(1656) <= a xor b;
    outputs(1657) <= a and b;
    outputs(1658) <= a and not b;
    outputs(1659) <= b;
    outputs(1660) <= a;
    outputs(1661) <= not (a or b);
    outputs(1662) <= b and not a;
    outputs(1663) <= a xor b;
    outputs(1664) <= a and b;
    outputs(1665) <= not a;
    outputs(1666) <= not b;
    outputs(1667) <= not b;
    outputs(1668) <= a xor b;
    outputs(1669) <= a and b;
    outputs(1670) <= b;
    outputs(1671) <= a xor b;
    outputs(1672) <= not a;
    outputs(1673) <= not (a xor b);
    outputs(1674) <= a;
    outputs(1675) <= not b;
    outputs(1676) <= a;
    outputs(1677) <= b;
    outputs(1678) <= not (a xor b);
    outputs(1679) <= a;
    outputs(1680) <= a xor b;
    outputs(1681) <= b and not a;
    outputs(1682) <= not b;
    outputs(1683) <= b and not a;
    outputs(1684) <= not a;
    outputs(1685) <= not a;
    outputs(1686) <= not a or b;
    outputs(1687) <= not b;
    outputs(1688) <= a and b;
    outputs(1689) <= not (a xor b);
    outputs(1690) <= a xor b;
    outputs(1691) <= a xor b;
    outputs(1692) <= not a;
    outputs(1693) <= not (a xor b);
    outputs(1694) <= a xor b;
    outputs(1695) <= b and not a;
    outputs(1696) <= a;
    outputs(1697) <= a and not b;
    outputs(1698) <= not (a or b);
    outputs(1699) <= b and not a;
    outputs(1700) <= b and not a;
    outputs(1701) <= not (a xor b);
    outputs(1702) <= a and b;
    outputs(1703) <= a xor b;
    outputs(1704) <= a;
    outputs(1705) <= a and not b;
    outputs(1706) <= a xor b;
    outputs(1707) <= not (a xor b);
    outputs(1708) <= b;
    outputs(1709) <= b;
    outputs(1710) <= not (a and b);
    outputs(1711) <= a;
    outputs(1712) <= b and not a;
    outputs(1713) <= a and b;
    outputs(1714) <= not a;
    outputs(1715) <= not (a xor b);
    outputs(1716) <= b;
    outputs(1717) <= a xor b;
    outputs(1718) <= not b;
    outputs(1719) <= not (a xor b);
    outputs(1720) <= b;
    outputs(1721) <= not (a or b);
    outputs(1722) <= not a;
    outputs(1723) <= not a;
    outputs(1724) <= not (a and b);
    outputs(1725) <= not a;
    outputs(1726) <= a and b;
    outputs(1727) <= not (a or b);
    outputs(1728) <= not (a xor b);
    outputs(1729) <= a xor b;
    outputs(1730) <= b;
    outputs(1731) <= not (a or b);
    outputs(1732) <= a and not b;
    outputs(1733) <= b;
    outputs(1734) <= b;
    outputs(1735) <= not b;
    outputs(1736) <= not (a xor b);
    outputs(1737) <= a xor b;
    outputs(1738) <= not a;
    outputs(1739) <= b;
    outputs(1740) <= a;
    outputs(1741) <= not b;
    outputs(1742) <= not a or b;
    outputs(1743) <= not (a xor b);
    outputs(1744) <= not a;
    outputs(1745) <= not b;
    outputs(1746) <= not b;
    outputs(1747) <= not b;
    outputs(1748) <= not (a xor b);
    outputs(1749) <= not b;
    outputs(1750) <= not (a xor b);
    outputs(1751) <= a xor b;
    outputs(1752) <= a;
    outputs(1753) <= b;
    outputs(1754) <= a;
    outputs(1755) <= not (a or b);
    outputs(1756) <= not b;
    outputs(1757) <= a xor b;
    outputs(1758) <= a or b;
    outputs(1759) <= b;
    outputs(1760) <= a and not b;
    outputs(1761) <= not a;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= not (a xor b);
    outputs(1764) <= not a;
    outputs(1765) <= a and not b;
    outputs(1766) <= not b;
    outputs(1767) <= a xor b;
    outputs(1768) <= b;
    outputs(1769) <= b;
    outputs(1770) <= a;
    outputs(1771) <= a;
    outputs(1772) <= a xor b;
    outputs(1773) <= not (a or b);
    outputs(1774) <= a xor b;
    outputs(1775) <= b;
    outputs(1776) <= not b or a;
    outputs(1777) <= a;
    outputs(1778) <= a;
    outputs(1779) <= a;
    outputs(1780) <= a;
    outputs(1781) <= a xor b;
    outputs(1782) <= a and not b;
    outputs(1783) <= a and not b;
    outputs(1784) <= b and not a;
    outputs(1785) <= b;
    outputs(1786) <= not (a xor b);
    outputs(1787) <= a;
    outputs(1788) <= not b;
    outputs(1789) <= a and b;
    outputs(1790) <= a xor b;
    outputs(1791) <= not (a or b);
    outputs(1792) <= b and not a;
    outputs(1793) <= a;
    outputs(1794) <= not a;
    outputs(1795) <= a or b;
    outputs(1796) <= not b;
    outputs(1797) <= b;
    outputs(1798) <= not b;
    outputs(1799) <= a and not b;
    outputs(1800) <= a;
    outputs(1801) <= not a;
    outputs(1802) <= b;
    outputs(1803) <= a xor b;
    outputs(1804) <= not a;
    outputs(1805) <= not (a xor b);
    outputs(1806) <= not a;
    outputs(1807) <= b and not a;
    outputs(1808) <= b;
    outputs(1809) <= a xor b;
    outputs(1810) <= not (a xor b);
    outputs(1811) <= not (a or b);
    outputs(1812) <= not (a or b);
    outputs(1813) <= not (a xor b);
    outputs(1814) <= a or b;
    outputs(1815) <= b;
    outputs(1816) <= not (a xor b);
    outputs(1817) <= a;
    outputs(1818) <= b;
    outputs(1819) <= a and not b;
    outputs(1820) <= not (a or b);
    outputs(1821) <= not (a xor b);
    outputs(1822) <= not b;
    outputs(1823) <= b;
    outputs(1824) <= 1'b0;
    outputs(1825) <= not a;
    outputs(1826) <= a and b;
    outputs(1827) <= b and not a;
    outputs(1828) <= a and not b;
    outputs(1829) <= a;
    outputs(1830) <= not a;
    outputs(1831) <= a;
    outputs(1832) <= a xor b;
    outputs(1833) <= a xor b;
    outputs(1834) <= a and b;
    outputs(1835) <= b;
    outputs(1836) <= a and not b;
    outputs(1837) <= not (a xor b);
    outputs(1838) <= a xor b;
    outputs(1839) <= a xor b;
    outputs(1840) <= not b;
    outputs(1841) <= not b;
    outputs(1842) <= not (a xor b);
    outputs(1843) <= a and not b;
    outputs(1844) <= a;
    outputs(1845) <= not b;
    outputs(1846) <= a xor b;
    outputs(1847) <= not b;
    outputs(1848) <= a xor b;
    outputs(1849) <= b;
    outputs(1850) <= not (a or b);
    outputs(1851) <= a and not b;
    outputs(1852) <= a;
    outputs(1853) <= not b;
    outputs(1854) <= a and b;
    outputs(1855) <= not (a xor b);
    outputs(1856) <= b;
    outputs(1857) <= not (a xor b);
    outputs(1858) <= not (a xor b);
    outputs(1859) <= not (a or b);
    outputs(1860) <= a;
    outputs(1861) <= b and not a;
    outputs(1862) <= not (a xor b);
    outputs(1863) <= a;
    outputs(1864) <= a and b;
    outputs(1865) <= not a;
    outputs(1866) <= a xor b;
    outputs(1867) <= not a;
    outputs(1868) <= not a;
    outputs(1869) <= not (a xor b);
    outputs(1870) <= b and not a;
    outputs(1871) <= a;
    outputs(1872) <= b and not a;
    outputs(1873) <= not a;
    outputs(1874) <= not (a or b);
    outputs(1875) <= not (a xor b);
    outputs(1876) <= not b;
    outputs(1877) <= a and b;
    outputs(1878) <= a xor b;
    outputs(1879) <= a and b;
    outputs(1880) <= not (a xor b);
    outputs(1881) <= not (a xor b);
    outputs(1882) <= not a;
    outputs(1883) <= a and not b;
    outputs(1884) <= a and not b;
    outputs(1885) <= not (a or b);
    outputs(1886) <= a xor b;
    outputs(1887) <= a xor b;
    outputs(1888) <= not b;
    outputs(1889) <= not (a or b);
    outputs(1890) <= not a;
    outputs(1891) <= a or b;
    outputs(1892) <= a;
    outputs(1893) <= not a;
    outputs(1894) <= not (a xor b);
    outputs(1895) <= not (a xor b);
    outputs(1896) <= not (a xor b);
    outputs(1897) <= not (a xor b);
    outputs(1898) <= not (a xor b);
    outputs(1899) <= b and not a;
    outputs(1900) <= a and b;
    outputs(1901) <= not a;
    outputs(1902) <= a;
    outputs(1903) <= not (a or b);
    outputs(1904) <= not (a xor b);
    outputs(1905) <= not a;
    outputs(1906) <= a xor b;
    outputs(1907) <= b and not a;
    outputs(1908) <= a and b;
    outputs(1909) <= not (a or b);
    outputs(1910) <= not a;
    outputs(1911) <= a and not b;
    outputs(1912) <= not (a xor b);
    outputs(1913) <= a xor b;
    outputs(1914) <= not (a xor b);
    outputs(1915) <= a and not b;
    outputs(1916) <= a and b;
    outputs(1917) <= a and not b;
    outputs(1918) <= not b;
    outputs(1919) <= not (a xor b);
    outputs(1920) <= a xor b;
    outputs(1921) <= a and not b;
    outputs(1922) <= not (a xor b);
    outputs(1923) <= not a or b;
    outputs(1924) <= a and not b;
    outputs(1925) <= a;
    outputs(1926) <= not (a or b);
    outputs(1927) <= b;
    outputs(1928) <= a;
    outputs(1929) <= not b;
    outputs(1930) <= a and b;
    outputs(1931) <= b;
    outputs(1932) <= not (a xor b);
    outputs(1933) <= not b;
    outputs(1934) <= not a;
    outputs(1935) <= not b;
    outputs(1936) <= a;
    outputs(1937) <= not a;
    outputs(1938) <= not b or a;
    outputs(1939) <= a xor b;
    outputs(1940) <= not (a xor b);
    outputs(1941) <= not a;
    outputs(1942) <= a xor b;
    outputs(1943) <= not b or a;
    outputs(1944) <= not (a xor b);
    outputs(1945) <= a xor b;
    outputs(1946) <= a and b;
    outputs(1947) <= not a;
    outputs(1948) <= a and b;
    outputs(1949) <= a and not b;
    outputs(1950) <= a;
    outputs(1951) <= a or b;
    outputs(1952) <= b;
    outputs(1953) <= a;
    outputs(1954) <= a xor b;
    outputs(1955) <= a;
    outputs(1956) <= not (a xor b);
    outputs(1957) <= b and not a;
    outputs(1958) <= b;
    outputs(1959) <= b;
    outputs(1960) <= not (a or b);
    outputs(1961) <= a xor b;
    outputs(1962) <= not (a or b);
    outputs(1963) <= a and b;
    outputs(1964) <= b;
    outputs(1965) <= a xor b;
    outputs(1966) <= not (a or b);
    outputs(1967) <= not (a xor b);
    outputs(1968) <= not (a xor b);
    outputs(1969) <= b;
    outputs(1970) <= not (a xor b);
    outputs(1971) <= not b;
    outputs(1972) <= a and b;
    outputs(1973) <= not (a and b);
    outputs(1974) <= a xor b;
    outputs(1975) <= not (a and b);
    outputs(1976) <= not (a or b);
    outputs(1977) <= 1'b0;
    outputs(1978) <= not b;
    outputs(1979) <= not (a or b);
    outputs(1980) <= a xor b;
    outputs(1981) <= b and not a;
    outputs(1982) <= not a or b;
    outputs(1983) <= b;
    outputs(1984) <= not a;
    outputs(1985) <= not b;
    outputs(1986) <= a;
    outputs(1987) <= not (a or b);
    outputs(1988) <= a;
    outputs(1989) <= not (a or b);
    outputs(1990) <= a and not b;
    outputs(1991) <= a;
    outputs(1992) <= not (a xor b);
    outputs(1993) <= not b or a;
    outputs(1994) <= not (a or b);
    outputs(1995) <= not b or a;
    outputs(1996) <= a and not b;
    outputs(1997) <= a xor b;
    outputs(1998) <= a and b;
    outputs(1999) <= b;
    outputs(2000) <= a and b;
    outputs(2001) <= not a;
    outputs(2002) <= a and not b;
    outputs(2003) <= not (a xor b);
    outputs(2004) <= not (a or b);
    outputs(2005) <= a and b;
    outputs(2006) <= not b;
    outputs(2007) <= not b;
    outputs(2008) <= a xor b;
    outputs(2009) <= not b or a;
    outputs(2010) <= a xor b;
    outputs(2011) <= a;
    outputs(2012) <= not a;
    outputs(2013) <= a xor b;
    outputs(2014) <= not (a or b);
    outputs(2015) <= a;
    outputs(2016) <= b and not a;
    outputs(2017) <= not (a or b);
    outputs(2018) <= b and not a;
    outputs(2019) <= a and not b;
    outputs(2020) <= a and b;
    outputs(2021) <= a xor b;
    outputs(2022) <= not a;
    outputs(2023) <= not a;
    outputs(2024) <= not a;
    outputs(2025) <= a or b;
    outputs(2026) <= b;
    outputs(2027) <= a xor b;
    outputs(2028) <= not (a xor b);
    outputs(2029) <= a and b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= a and not b;
    outputs(2032) <= a and b;
    outputs(2033) <= a xor b;
    outputs(2034) <= not (a xor b);
    outputs(2035) <= not (a xor b);
    outputs(2036) <= not a;
    outputs(2037) <= b;
    outputs(2038) <= not b;
    outputs(2039) <= b and not a;
    outputs(2040) <= a;
    outputs(2041) <= a xor b;
    outputs(2042) <= b and not a;
    outputs(2043) <= not (a xor b);
    outputs(2044) <= b;
    outputs(2045) <= a xor b;
    outputs(2046) <= a xor b;
    outputs(2047) <= a and not b;
    outputs(2048) <= not b;
    outputs(2049) <= not b or a;
    outputs(2050) <= not (a xor b);
    outputs(2051) <= not (a and b);
    outputs(2052) <= b;
    outputs(2053) <= a;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= a xor b;
    outputs(2056) <= a xor b;
    outputs(2057) <= not b;
    outputs(2058) <= a;
    outputs(2059) <= not a;
    outputs(2060) <= not a or b;
    outputs(2061) <= not a;
    outputs(2062) <= not (a xor b);
    outputs(2063) <= not b or a;
    outputs(2064) <= a;
    outputs(2065) <= a xor b;
    outputs(2066) <= a or b;
    outputs(2067) <= not b;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= not b or a;
    outputs(2070) <= a;
    outputs(2071) <= a;
    outputs(2072) <= b;
    outputs(2073) <= a xor b;
    outputs(2074) <= a;
    outputs(2075) <= not (a xor b);
    outputs(2076) <= not (a xor b);
    outputs(2077) <= a and not b;
    outputs(2078) <= not (a xor b);
    outputs(2079) <= a;
    outputs(2080) <= not a or b;
    outputs(2081) <= a xor b;
    outputs(2082) <= a;
    outputs(2083) <= a or b;
    outputs(2084) <= not a;
    outputs(2085) <= a xor b;
    outputs(2086) <= not (a and b);
    outputs(2087) <= b;
    outputs(2088) <= not (a xor b);
    outputs(2089) <= not (a and b);
    outputs(2090) <= not a;
    outputs(2091) <= a and not b;
    outputs(2092) <= a;
    outputs(2093) <= not (a xor b);
    outputs(2094) <= not (a xor b);
    outputs(2095) <= a;
    outputs(2096) <= a xor b;
    outputs(2097) <= a and not b;
    outputs(2098) <= not (a xor b);
    outputs(2099) <= not (a xor b);
    outputs(2100) <= b;
    outputs(2101) <= not b;
    outputs(2102) <= not a or b;
    outputs(2103) <= a and b;
    outputs(2104) <= a or b;
    outputs(2105) <= not a;
    outputs(2106) <= not (a xor b);
    outputs(2107) <= a and not b;
    outputs(2108) <= a;
    outputs(2109) <= a or b;
    outputs(2110) <= a xor b;
    outputs(2111) <= b;
    outputs(2112) <= a xor b;
    outputs(2113) <= a and b;
    outputs(2114) <= not (a xor b);
    outputs(2115) <= not (a xor b);
    outputs(2116) <= a;
    outputs(2117) <= not (a and b);
    outputs(2118) <= b and not a;
    outputs(2119) <= not a;
    outputs(2120) <= b;
    outputs(2121) <= not b;
    outputs(2122) <= not a;
    outputs(2123) <= a xor b;
    outputs(2124) <= a xor b;
    outputs(2125) <= not b;
    outputs(2126) <= a xor b;
    outputs(2127) <= not (a and b);
    outputs(2128) <= a;
    outputs(2129) <= a xor b;
    outputs(2130) <= not a or b;
    outputs(2131) <= a or b;
    outputs(2132) <= b;
    outputs(2133) <= a;
    outputs(2134) <= b and not a;
    outputs(2135) <= a xor b;
    outputs(2136) <= not a;
    outputs(2137) <= not (a and b);
    outputs(2138) <= not (a xor b);
    outputs(2139) <= a xor b;
    outputs(2140) <= a xor b;
    outputs(2141) <= not (a xor b);
    outputs(2142) <= b;
    outputs(2143) <= not a;
    outputs(2144) <= not (a xor b);
    outputs(2145) <= b;
    outputs(2146) <= a;
    outputs(2147) <= a;
    outputs(2148) <= b;
    outputs(2149) <= not a;
    outputs(2150) <= not b or a;
    outputs(2151) <= not (a and b);
    outputs(2152) <= not b;
    outputs(2153) <= b;
    outputs(2154) <= not a;
    outputs(2155) <= not (a xor b);
    outputs(2156) <= not b;
    outputs(2157) <= not (a xor b);
    outputs(2158) <= a and b;
    outputs(2159) <= a xor b;
    outputs(2160) <= a and not b;
    outputs(2161) <= a;
    outputs(2162) <= not b or a;
    outputs(2163) <= not b or a;
    outputs(2164) <= a xor b;
    outputs(2165) <= a and not b;
    outputs(2166) <= not a;
    outputs(2167) <= not b;
    outputs(2168) <= not b or a;
    outputs(2169) <= not b;
    outputs(2170) <= b and not a;
    outputs(2171) <= b;
    outputs(2172) <= not (a xor b);
    outputs(2173) <= a;
    outputs(2174) <= not (a xor b);
    outputs(2175) <= not a;
    outputs(2176) <= a xor b;
    outputs(2177) <= not b;
    outputs(2178) <= a and b;
    outputs(2179) <= not (a or b);
    outputs(2180) <= a;
    outputs(2181) <= not b;
    outputs(2182) <= b;
    outputs(2183) <= a xor b;
    outputs(2184) <= a;
    outputs(2185) <= not (a xor b);
    outputs(2186) <= b;
    outputs(2187) <= a;
    outputs(2188) <= a xor b;
    outputs(2189) <= a;
    outputs(2190) <= b;
    outputs(2191) <= not a or b;
    outputs(2192) <= not b;
    outputs(2193) <= not (a and b);
    outputs(2194) <= not b or a;
    outputs(2195) <= not a;
    outputs(2196) <= not a or b;
    outputs(2197) <= not (a xor b);
    outputs(2198) <= not b;
    outputs(2199) <= not b or a;
    outputs(2200) <= a and b;
    outputs(2201) <= not (a xor b);
    outputs(2202) <= not (a xor b);
    outputs(2203) <= a xor b;
    outputs(2204) <= not a;
    outputs(2205) <= not (a xor b);
    outputs(2206) <= not (a xor b);
    outputs(2207) <= not (a or b);
    outputs(2208) <= not (a xor b);
    outputs(2209) <= not (a and b);
    outputs(2210) <= a;
    outputs(2211) <= not b;
    outputs(2212) <= not a;
    outputs(2213) <= not (a xor b);
    outputs(2214) <= not a;
    outputs(2215) <= not (a xor b);
    outputs(2216) <= not (a or b);
    outputs(2217) <= not a;
    outputs(2218) <= not (a xor b);
    outputs(2219) <= not a;
    outputs(2220) <= not (a xor b);
    outputs(2221) <= not a;
    outputs(2222) <= not (a xor b);
    outputs(2223) <= not b;
    outputs(2224) <= a and not b;
    outputs(2225) <= a;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= not (a xor b);
    outputs(2228) <= b and not a;
    outputs(2229) <= not (a xor b);
    outputs(2230) <= b and not a;
    outputs(2231) <= not a;
    outputs(2232) <= not a;
    outputs(2233) <= not b;
    outputs(2234) <= not b;
    outputs(2235) <= a or b;
    outputs(2236) <= a;
    outputs(2237) <= a xor b;
    outputs(2238) <= not (a xor b);
    outputs(2239) <= not (a and b);
    outputs(2240) <= a xor b;
    outputs(2241) <= not (a xor b);
    outputs(2242) <= b;
    outputs(2243) <= a and b;
    outputs(2244) <= not (a or b);
    outputs(2245) <= a xor b;
    outputs(2246) <= not (a xor b);
    outputs(2247) <= not (a xor b);
    outputs(2248) <= not (a or b);
    outputs(2249) <= b;
    outputs(2250) <= b;
    outputs(2251) <= a xor b;
    outputs(2252) <= a and b;
    outputs(2253) <= not a;
    outputs(2254) <= a;
    outputs(2255) <= not b;
    outputs(2256) <= b and not a;
    outputs(2257) <= b;
    outputs(2258) <= not a or b;
    outputs(2259) <= not b;
    outputs(2260) <= not b;
    outputs(2261) <= a or b;
    outputs(2262) <= not a;
    outputs(2263) <= a and not b;
    outputs(2264) <= not (a and b);
    outputs(2265) <= not b;
    outputs(2266) <= a and not b;
    outputs(2267) <= a xor b;
    outputs(2268) <= b;
    outputs(2269) <= not a;
    outputs(2270) <= not b or a;
    outputs(2271) <= not (a xor b);
    outputs(2272) <= a;
    outputs(2273) <= a xor b;
    outputs(2274) <= a xor b;
    outputs(2275) <= b;
    outputs(2276) <= not (a xor b);
    outputs(2277) <= a xor b;
    outputs(2278) <= not a or b;
    outputs(2279) <= b;
    outputs(2280) <= not (a xor b);
    outputs(2281) <= not b;
    outputs(2282) <= not a;
    outputs(2283) <= a;
    outputs(2284) <= not b;
    outputs(2285) <= not (a or b);
    outputs(2286) <= a or b;
    outputs(2287) <= a;
    outputs(2288) <= a;
    outputs(2289) <= not b;
    outputs(2290) <= not b;
    outputs(2291) <= b;
    outputs(2292) <= not b;
    outputs(2293) <= b;
    outputs(2294) <= not a;
    outputs(2295) <= a xor b;
    outputs(2296) <= not b or a;
    outputs(2297) <= a xor b;
    outputs(2298) <= a;
    outputs(2299) <= not (a xor b);
    outputs(2300) <= a xor b;
    outputs(2301) <= not b;
    outputs(2302) <= not (a or b);
    outputs(2303) <= not (a xor b);
    outputs(2304) <= a or b;
    outputs(2305) <= a xor b;
    outputs(2306) <= not (a xor b);
    outputs(2307) <= not (a or b);
    outputs(2308) <= not (a xor b);
    outputs(2309) <= not a;
    outputs(2310) <= not a;
    outputs(2311) <= a and not b;
    outputs(2312) <= a;
    outputs(2313) <= b;
    outputs(2314) <= b;
    outputs(2315) <= b;
    outputs(2316) <= a;
    outputs(2317) <= not (a xor b);
    outputs(2318) <= a xor b;
    outputs(2319) <= b;
    outputs(2320) <= a or b;
    outputs(2321) <= a xor b;
    outputs(2322) <= not b;
    outputs(2323) <= not (a xor b);
    outputs(2324) <= a and not b;
    outputs(2325) <= a and not b;
    outputs(2326) <= not a;
    outputs(2327) <= not b or a;
    outputs(2328) <= b;
    outputs(2329) <= a xor b;
    outputs(2330) <= not b;
    outputs(2331) <= not b or a;
    outputs(2332) <= b;
    outputs(2333) <= a xor b;
    outputs(2334) <= b;
    outputs(2335) <= not b or a;
    outputs(2336) <= a or b;
    outputs(2337) <= not (a and b);
    outputs(2338) <= not b;
    outputs(2339) <= a xor b;
    outputs(2340) <= not a;
    outputs(2341) <= a xor b;
    outputs(2342) <= not b;
    outputs(2343) <= not (a xor b);
    outputs(2344) <= a xor b;
    outputs(2345) <= a or b;
    outputs(2346) <= not a;
    outputs(2347) <= not a or b;
    outputs(2348) <= not (a or b);
    outputs(2349) <= not (a or b);
    outputs(2350) <= not (a xor b);
    outputs(2351) <= not b;
    outputs(2352) <= a xor b;
    outputs(2353) <= not b;
    outputs(2354) <= not (a or b);
    outputs(2355) <= a or b;
    outputs(2356) <= a and b;
    outputs(2357) <= not b;
    outputs(2358) <= a xor b;
    outputs(2359) <= not (a xor b);
    outputs(2360) <= a xor b;
    outputs(2361) <= b;
    outputs(2362) <= not a;
    outputs(2363) <= not (a xor b);
    outputs(2364) <= not a or b;
    outputs(2365) <= not (a and b);
    outputs(2366) <= not a or b;
    outputs(2367) <= not (a and b);
    outputs(2368) <= a;
    outputs(2369) <= not (a xor b);
    outputs(2370) <= not (a or b);
    outputs(2371) <= not (a xor b);
    outputs(2372) <= not b;
    outputs(2373) <= a xor b;
    outputs(2374) <= not b;
    outputs(2375) <= not b;
    outputs(2376) <= not (a xor b);
    outputs(2377) <= b;
    outputs(2378) <= a and not b;
    outputs(2379) <= a xor b;
    outputs(2380) <= a xor b;
    outputs(2381) <= a;
    outputs(2382) <= not (a xor b);
    outputs(2383) <= a and b;
    outputs(2384) <= not (a xor b);
    outputs(2385) <= not (a xor b);
    outputs(2386) <= not b;
    outputs(2387) <= a;
    outputs(2388) <= not (a and b);
    outputs(2389) <= a or b;
    outputs(2390) <= a;
    outputs(2391) <= not (a xor b);
    outputs(2392) <= not b;
    outputs(2393) <= a and not b;
    outputs(2394) <= b;
    outputs(2395) <= a xor b;
    outputs(2396) <= a xor b;
    outputs(2397) <= a xor b;
    outputs(2398) <= a xor b;
    outputs(2399) <= not (a xor b);
    outputs(2400) <= not a;
    outputs(2401) <= b;
    outputs(2402) <= not (a xor b);
    outputs(2403) <= a and not b;
    outputs(2404) <= not (a and b);
    outputs(2405) <= b;
    outputs(2406) <= b;
    outputs(2407) <= not b;
    outputs(2408) <= not (a and b);
    outputs(2409) <= not b;
    outputs(2410) <= not (a xor b);
    outputs(2411) <= not a or b;
    outputs(2412) <= a xor b;
    outputs(2413) <= a or b;
    outputs(2414) <= not b or a;
    outputs(2415) <= a xor b;
    outputs(2416) <= a;
    outputs(2417) <= a;
    outputs(2418) <= not a;
    outputs(2419) <= not (a xor b);
    outputs(2420) <= b;
    outputs(2421) <= not a;
    outputs(2422) <= b;
    outputs(2423) <= a xor b;
    outputs(2424) <= b;
    outputs(2425) <= a;
    outputs(2426) <= not a or b;
    outputs(2427) <= not (a and b);
    outputs(2428) <= not a;
    outputs(2429) <= not b or a;
    outputs(2430) <= not b;
    outputs(2431) <= not (a xor b);
    outputs(2432) <= a;
    outputs(2433) <= a xor b;
    outputs(2434) <= a xor b;
    outputs(2435) <= a;
    outputs(2436) <= a xor b;
    outputs(2437) <= b;
    outputs(2438) <= not (a xor b);
    outputs(2439) <= not (a xor b);
    outputs(2440) <= not (a xor b);
    outputs(2441) <= not b;
    outputs(2442) <= not (a xor b);
    outputs(2443) <= b;
    outputs(2444) <= not b or a;
    outputs(2445) <= not b;
    outputs(2446) <= a xor b;
    outputs(2447) <= b;
    outputs(2448) <= a xor b;
    outputs(2449) <= a xor b;
    outputs(2450) <= not b;
    outputs(2451) <= a xor b;
    outputs(2452) <= not a;
    outputs(2453) <= a;
    outputs(2454) <= a xor b;
    outputs(2455) <= not (a or b);
    outputs(2456) <= a and b;
    outputs(2457) <= a;
    outputs(2458) <= not a;
    outputs(2459) <= a xor b;
    outputs(2460) <= b;
    outputs(2461) <= not (a or b);
    outputs(2462) <= not a;
    outputs(2463) <= a;
    outputs(2464) <= a and b;
    outputs(2465) <= not (a xor b);
    outputs(2466) <= not a;
    outputs(2467) <= not a;
    outputs(2468) <= not b;
    outputs(2469) <= b;
    outputs(2470) <= not b;
    outputs(2471) <= a;
    outputs(2472) <= a or b;
    outputs(2473) <= b;
    outputs(2474) <= not a;
    outputs(2475) <= not a;
    outputs(2476) <= not (a xor b);
    outputs(2477) <= not b;
    outputs(2478) <= a or b;
    outputs(2479) <= a;
    outputs(2480) <= a;
    outputs(2481) <= not (a xor b);
    outputs(2482) <= not (a xor b);
    outputs(2483) <= b;
    outputs(2484) <= not b;
    outputs(2485) <= a xor b;
    outputs(2486) <= not (a and b);
    outputs(2487) <= not b;
    outputs(2488) <= a xor b;
    outputs(2489) <= not (a or b);
    outputs(2490) <= b;
    outputs(2491) <= not (a xor b);
    outputs(2492) <= not (a xor b);
    outputs(2493) <= a and not b;
    outputs(2494) <= not b or a;
    outputs(2495) <= not b;
    outputs(2496) <= b;
    outputs(2497) <= not (a or b);
    outputs(2498) <= not a;
    outputs(2499) <= b;
    outputs(2500) <= not (a xor b);
    outputs(2501) <= b;
    outputs(2502) <= not b;
    outputs(2503) <= a xor b;
    outputs(2504) <= b;
    outputs(2505) <= not (a and b);
    outputs(2506) <= not (a xor b);
    outputs(2507) <= a xor b;
    outputs(2508) <= b;
    outputs(2509) <= not (a or b);
    outputs(2510) <= b;
    outputs(2511) <= not b;
    outputs(2512) <= not (a or b);
    outputs(2513) <= b;
    outputs(2514) <= a;
    outputs(2515) <= a xor b;
    outputs(2516) <= b;
    outputs(2517) <= not b;
    outputs(2518) <= not b;
    outputs(2519) <= not (a xor b);
    outputs(2520) <= a;
    outputs(2521) <= a;
    outputs(2522) <= b;
    outputs(2523) <= not a;
    outputs(2524) <= a xor b;
    outputs(2525) <= a or b;
    outputs(2526) <= not a;
    outputs(2527) <= a and not b;
    outputs(2528) <= not b;
    outputs(2529) <= a xor b;
    outputs(2530) <= not b;
    outputs(2531) <= not (a and b);
    outputs(2532) <= not (a xor b);
    outputs(2533) <= b;
    outputs(2534) <= not (a xor b);
    outputs(2535) <= not b;
    outputs(2536) <= not b;
    outputs(2537) <= a xor b;
    outputs(2538) <= not (a xor b);
    outputs(2539) <= a xor b;
    outputs(2540) <= a and b;
    outputs(2541) <= a or b;
    outputs(2542) <= not (a xor b);
    outputs(2543) <= a;
    outputs(2544) <= a xor b;
    outputs(2545) <= b;
    outputs(2546) <= a xor b;
    outputs(2547) <= a and not b;
    outputs(2548) <= not (a xor b);
    outputs(2549) <= 1'b1;
    outputs(2550) <= b;
    outputs(2551) <= not a;
    outputs(2552) <= not (a xor b);
    outputs(2553) <= a xor b;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= a xor b;
    outputs(2556) <= not (a or b);
    outputs(2557) <= b and not a;
    outputs(2558) <= a and not b;
    outputs(2559) <= a xor b;
    outputs(2560) <= a and not b;
    outputs(2561) <= b;
    outputs(2562) <= b;
    outputs(2563) <= not (a xor b);
    outputs(2564) <= not b;
    outputs(2565) <= not a or b;
    outputs(2566) <= not b;
    outputs(2567) <= not b;
    outputs(2568) <= not a;
    outputs(2569) <= not b;
    outputs(2570) <= b;
    outputs(2571) <= b;
    outputs(2572) <= a and b;
    outputs(2573) <= a;
    outputs(2574) <= not a;
    outputs(2575) <= a xor b;
    outputs(2576) <= b;
    outputs(2577) <= not a;
    outputs(2578) <= not a;
    outputs(2579) <= a xor b;
    outputs(2580) <= not (a or b);
    outputs(2581) <= a xor b;
    outputs(2582) <= a xor b;
    outputs(2583) <= not a or b;
    outputs(2584) <= not (a xor b);
    outputs(2585) <= a xor b;
    outputs(2586) <= not a;
    outputs(2587) <= not (a or b);
    outputs(2588) <= not a;
    outputs(2589) <= not (a or b);
    outputs(2590) <= b;
    outputs(2591) <= not a;
    outputs(2592) <= not b;
    outputs(2593) <= a xor b;
    outputs(2594) <= not (a and b);
    outputs(2595) <= not (a or b);
    outputs(2596) <= b;
    outputs(2597) <= not b;
    outputs(2598) <= a xor b;
    outputs(2599) <= a xor b;
    outputs(2600) <= not a or b;
    outputs(2601) <= b;
    outputs(2602) <= not b;
    outputs(2603) <= a and not b;
    outputs(2604) <= a;
    outputs(2605) <= not a;
    outputs(2606) <= not (a xor b);
    outputs(2607) <= not a;
    outputs(2608) <= not a;
    outputs(2609) <= not a or b;
    outputs(2610) <= a xor b;
    outputs(2611) <= a;
    outputs(2612) <= not (a xor b);
    outputs(2613) <= not b;
    outputs(2614) <= b;
    outputs(2615) <= a;
    outputs(2616) <= a;
    outputs(2617) <= a;
    outputs(2618) <= not b;
    outputs(2619) <= not b;
    outputs(2620) <= a xor b;
    outputs(2621) <= not a or b;
    outputs(2622) <= a;
    outputs(2623) <= a;
    outputs(2624) <= not (a xor b);
    outputs(2625) <= a xor b;
    outputs(2626) <= a;
    outputs(2627) <= not a or b;
    outputs(2628) <= a;
    outputs(2629) <= not (a xor b);
    outputs(2630) <= not (a and b);
    outputs(2631) <= not a;
    outputs(2632) <= a and not b;
    outputs(2633) <= not a;
    outputs(2634) <= a or b;
    outputs(2635) <= b;
    outputs(2636) <= b and not a;
    outputs(2637) <= a and b;
    outputs(2638) <= a xor b;
    outputs(2639) <= a and b;
    outputs(2640) <= not (a and b);
    outputs(2641) <= not b;
    outputs(2642) <= a xor b;
    outputs(2643) <= b;
    outputs(2644) <= not a;
    outputs(2645) <= not (a xor b);
    outputs(2646) <= not b;
    outputs(2647) <= not a;
    outputs(2648) <= a xor b;
    outputs(2649) <= not a or b;
    outputs(2650) <= not (a and b);
    outputs(2651) <= not b or a;
    outputs(2652) <= not b;
    outputs(2653) <= b;
    outputs(2654) <= not (a and b);
    outputs(2655) <= not b;
    outputs(2656) <= a;
    outputs(2657) <= not (a xor b);
    outputs(2658) <= not a;
    outputs(2659) <= a and not b;
    outputs(2660) <= a;
    outputs(2661) <= a;
    outputs(2662) <= a and not b;
    outputs(2663) <= a or b;
    outputs(2664) <= a or b;
    outputs(2665) <= b;
    outputs(2666) <= a xor b;
    outputs(2667) <= a;
    outputs(2668) <= a xor b;
    outputs(2669) <= not b;
    outputs(2670) <= a;
    outputs(2671) <= not (a and b);
    outputs(2672) <= b;
    outputs(2673) <= b;
    outputs(2674) <= a and b;
    outputs(2675) <= not a;
    outputs(2676) <= not b;
    outputs(2677) <= a;
    outputs(2678) <= a xor b;
    outputs(2679) <= not (a xor b);
    outputs(2680) <= a xor b;
    outputs(2681) <= 1'b1;
    outputs(2682) <= not a;
    outputs(2683) <= not (a or b);
    outputs(2684) <= a;
    outputs(2685) <= a;
    outputs(2686) <= b;
    outputs(2687) <= a and b;
    outputs(2688) <= not b;
    outputs(2689) <= a xor b;
    outputs(2690) <= a xor b;
    outputs(2691) <= a xor b;
    outputs(2692) <= a;
    outputs(2693) <= not (a xor b);
    outputs(2694) <= b;
    outputs(2695) <= not a or b;
    outputs(2696) <= b and not a;
    outputs(2697) <= not a;
    outputs(2698) <= b and not a;
    outputs(2699) <= not b or a;
    outputs(2700) <= a xor b;
    outputs(2701) <= not (a and b);
    outputs(2702) <= not (a xor b);
    outputs(2703) <= not a;
    outputs(2704) <= a xor b;
    outputs(2705) <= not (a xor b);
    outputs(2706) <= not (a xor b);
    outputs(2707) <= not (a xor b);
    outputs(2708) <= a;
    outputs(2709) <= not a;
    outputs(2710) <= not b;
    outputs(2711) <= not b;
    outputs(2712) <= not (a or b);
    outputs(2713) <= not (a and b);
    outputs(2714) <= not b;
    outputs(2715) <= not (a xor b);
    outputs(2716) <= a xor b;
    outputs(2717) <= not a;
    outputs(2718) <= a xor b;
    outputs(2719) <= a xor b;
    outputs(2720) <= a;
    outputs(2721) <= not b or a;
    outputs(2722) <= a xor b;
    outputs(2723) <= not a;
    outputs(2724) <= not a or b;
    outputs(2725) <= not b;
    outputs(2726) <= b;
    outputs(2727) <= not (a xor b);
    outputs(2728) <= b;
    outputs(2729) <= a;
    outputs(2730) <= not (a or b);
    outputs(2731) <= not b;
    outputs(2732) <= not a;
    outputs(2733) <= not (a xor b);
    outputs(2734) <= a;
    outputs(2735) <= not b;
    outputs(2736) <= not (a xor b);
    outputs(2737) <= not a;
    outputs(2738) <= not (a or b);
    outputs(2739) <= a;
    outputs(2740) <= a xor b;
    outputs(2741) <= not b;
    outputs(2742) <= b;
    outputs(2743) <= b;
    outputs(2744) <= not (a xor b);
    outputs(2745) <= not b;
    outputs(2746) <= b and not a;
    outputs(2747) <= not (a and b);
    outputs(2748) <= not b;
    outputs(2749) <= b;
    outputs(2750) <= not b;
    outputs(2751) <= not a;
    outputs(2752) <= a xor b;
    outputs(2753) <= a xor b;
    outputs(2754) <= not a;
    outputs(2755) <= a;
    outputs(2756) <= not b;
    outputs(2757) <= not (a xor b);
    outputs(2758) <= b;
    outputs(2759) <= not (a or b);
    outputs(2760) <= a xor b;
    outputs(2761) <= a or b;
    outputs(2762) <= a and b;
    outputs(2763) <= not b or a;
    outputs(2764) <= not (a xor b);
    outputs(2765) <= b;
    outputs(2766) <= a xor b;
    outputs(2767) <= a and not b;
    outputs(2768) <= a;
    outputs(2769) <= a xor b;
    outputs(2770) <= a xor b;
    outputs(2771) <= b and not a;
    outputs(2772) <= a;
    outputs(2773) <= not a or b;
    outputs(2774) <= not (a and b);
    outputs(2775) <= not a;
    outputs(2776) <= b;
    outputs(2777) <= a xor b;
    outputs(2778) <= not b;
    outputs(2779) <= b;
    outputs(2780) <= a xor b;
    outputs(2781) <= not a;
    outputs(2782) <= a xor b;
    outputs(2783) <= not b;
    outputs(2784) <= not (a and b);
    outputs(2785) <= b;
    outputs(2786) <= not a;
    outputs(2787) <= a xor b;
    outputs(2788) <= not (a and b);
    outputs(2789) <= not b or a;
    outputs(2790) <= a and not b;
    outputs(2791) <= a xor b;
    outputs(2792) <= not (a xor b);
    outputs(2793) <= not a or b;
    outputs(2794) <= b;
    outputs(2795) <= not (a xor b);
    outputs(2796) <= not a;
    outputs(2797) <= not (a and b);
    outputs(2798) <= not b;
    outputs(2799) <= a and not b;
    outputs(2800) <= a xor b;
    outputs(2801) <= not a or b;
    outputs(2802) <= b;
    outputs(2803) <= a;
    outputs(2804) <= not b;
    outputs(2805) <= a xor b;
    outputs(2806) <= a or b;
    outputs(2807) <= not (a xor b);
    outputs(2808) <= b;
    outputs(2809) <= a xor b;
    outputs(2810) <= a;
    outputs(2811) <= b;
    outputs(2812) <= a;
    outputs(2813) <= not (a xor b);
    outputs(2814) <= b;
    outputs(2815) <= a;
    outputs(2816) <= not a;
    outputs(2817) <= a and not b;
    outputs(2818) <= b;
    outputs(2819) <= b;
    outputs(2820) <= a or b;
    outputs(2821) <= not (a xor b);
    outputs(2822) <= not (a xor b);
    outputs(2823) <= not a or b;
    outputs(2824) <= not b;
    outputs(2825) <= a or b;
    outputs(2826) <= a xor b;
    outputs(2827) <= a xor b;
    outputs(2828) <= a xor b;
    outputs(2829) <= not b;
    outputs(2830) <= not a;
    outputs(2831) <= b;
    outputs(2832) <= a xor b;
    outputs(2833) <= b;
    outputs(2834) <= a xor b;
    outputs(2835) <= not a;
    outputs(2836) <= not (a xor b);
    outputs(2837) <= a xor b;
    outputs(2838) <= b;
    outputs(2839) <= not b;
    outputs(2840) <= not a;
    outputs(2841) <= b;
    outputs(2842) <= a and not b;
    outputs(2843) <= not b;
    outputs(2844) <= a;
    outputs(2845) <= a;
    outputs(2846) <= not (a xor b);
    outputs(2847) <= a xor b;
    outputs(2848) <= a;
    outputs(2849) <= not a;
    outputs(2850) <= a;
    outputs(2851) <= a or b;
    outputs(2852) <= a;
    outputs(2853) <= a and b;
    outputs(2854) <= not (a xor b);
    outputs(2855) <= a xor b;
    outputs(2856) <= b and not a;
    outputs(2857) <= not a;
    outputs(2858) <= b;
    outputs(2859) <= not a or b;
    outputs(2860) <= a and not b;
    outputs(2861) <= not (a and b);
    outputs(2862) <= a or b;
    outputs(2863) <= a xor b;
    outputs(2864) <= a and not b;
    outputs(2865) <= not b;
    outputs(2866) <= a;
    outputs(2867) <= a xor b;
    outputs(2868) <= not (a and b);
    outputs(2869) <= a and not b;
    outputs(2870) <= not a;
    outputs(2871) <= b;
    outputs(2872) <= b;
    outputs(2873) <= a and b;
    outputs(2874) <= not (a and b);
    outputs(2875) <= b;
    outputs(2876) <= a and not b;
    outputs(2877) <= not a;
    outputs(2878) <= not (a xor b);
    outputs(2879) <= not (a xor b);
    outputs(2880) <= b;
    outputs(2881) <= not (a xor b);
    outputs(2882) <= not (a xor b);
    outputs(2883) <= a xor b;
    outputs(2884) <= a;
    outputs(2885) <= not b;
    outputs(2886) <= a and b;
    outputs(2887) <= a xor b;
    outputs(2888) <= b;
    outputs(2889) <= not a;
    outputs(2890) <= not b;
    outputs(2891) <= not a;
    outputs(2892) <= b;
    outputs(2893) <= not a;
    outputs(2894) <= not b;
    outputs(2895) <= not (a and b);
    outputs(2896) <= not (a xor b);
    outputs(2897) <= not (a xor b);
    outputs(2898) <= not a;
    outputs(2899) <= a and not b;
    outputs(2900) <= a;
    outputs(2901) <= a xor b;
    outputs(2902) <= not b or a;
    outputs(2903) <= not b;
    outputs(2904) <= a;
    outputs(2905) <= not (a and b);
    outputs(2906) <= not (a xor b);
    outputs(2907) <= not b;
    outputs(2908) <= not (a or b);
    outputs(2909) <= not (a xor b);
    outputs(2910) <= a xor b;
    outputs(2911) <= not b or a;
    outputs(2912) <= not a;
    outputs(2913) <= b;
    outputs(2914) <= not b;
    outputs(2915) <= not (a xor b);
    outputs(2916) <= a xor b;
    outputs(2917) <= not b or a;
    outputs(2918) <= not b;
    outputs(2919) <= not b;
    outputs(2920) <= a xor b;
    outputs(2921) <= not b;
    outputs(2922) <= not b or a;
    outputs(2923) <= a xor b;
    outputs(2924) <= a xor b;
    outputs(2925) <= not a;
    outputs(2926) <= not (a xor b);
    outputs(2927) <= not (a xor b);
    outputs(2928) <= a and b;
    outputs(2929) <= b and not a;
    outputs(2930) <= not b;
    outputs(2931) <= b;
    outputs(2932) <= a;
    outputs(2933) <= a xor b;
    outputs(2934) <= a or b;
    outputs(2935) <= not (a xor b);
    outputs(2936) <= not a or b;
    outputs(2937) <= b;
    outputs(2938) <= not (a xor b);
    outputs(2939) <= b;
    outputs(2940) <= a;
    outputs(2941) <= not (a and b);
    outputs(2942) <= not (a xor b);
    outputs(2943) <= not b or a;
    outputs(2944) <= b;
    outputs(2945) <= not (a xor b);
    outputs(2946) <= a xor b;
    outputs(2947) <= not (a xor b);
    outputs(2948) <= a or b;
    outputs(2949) <= not b;
    outputs(2950) <= not a or b;
    outputs(2951) <= b;
    outputs(2952) <= not b;
    outputs(2953) <= not a;
    outputs(2954) <= not (a and b);
    outputs(2955) <= a or b;
    outputs(2956) <= not b;
    outputs(2957) <= a or b;
    outputs(2958) <= a;
    outputs(2959) <= a xor b;
    outputs(2960) <= b;
    outputs(2961) <= b;
    outputs(2962) <= not b or a;
    outputs(2963) <= not a;
    outputs(2964) <= not (a xor b);
    outputs(2965) <= a and b;
    outputs(2966) <= b;
    outputs(2967) <= not b;
    outputs(2968) <= not a;
    outputs(2969) <= a xor b;
    outputs(2970) <= not (a xor b);
    outputs(2971) <= a;
    outputs(2972) <= a xor b;
    outputs(2973) <= not b or a;
    outputs(2974) <= not (a xor b);
    outputs(2975) <= a or b;
    outputs(2976) <= not a;
    outputs(2977) <= a;
    outputs(2978) <= a;
    outputs(2979) <= not (a xor b);
    outputs(2980) <= a xor b;
    outputs(2981) <= not a;
    outputs(2982) <= not b;
    outputs(2983) <= not b;
    outputs(2984) <= a or b;
    outputs(2985) <= a xor b;
    outputs(2986) <= not (a xor b);
    outputs(2987) <= a xor b;
    outputs(2988) <= not a;
    outputs(2989) <= a;
    outputs(2990) <= a or b;
    outputs(2991) <= a;
    outputs(2992) <= a;
    outputs(2993) <= not (a xor b);
    outputs(2994) <= not a;
    outputs(2995) <= not a;
    outputs(2996) <= not (a xor b);
    outputs(2997) <= a xor b;
    outputs(2998) <= b;
    outputs(2999) <= not a;
    outputs(3000) <= a;
    outputs(3001) <= not (a or b);
    outputs(3002) <= a;
    outputs(3003) <= not b;
    outputs(3004) <= a;
    outputs(3005) <= not b;
    outputs(3006) <= not a or b;
    outputs(3007) <= not a;
    outputs(3008) <= b;
    outputs(3009) <= not a;
    outputs(3010) <= a or b;
    outputs(3011) <= a xor b;
    outputs(3012) <= b;
    outputs(3013) <= not b;
    outputs(3014) <= b;
    outputs(3015) <= a or b;
    outputs(3016) <= a;
    outputs(3017) <= not b;
    outputs(3018) <= not b or a;
    outputs(3019) <= not b or a;
    outputs(3020) <= not (a and b);
    outputs(3021) <= not (a and b);
    outputs(3022) <= a and not b;
    outputs(3023) <= not b;
    outputs(3024) <= a or b;
    outputs(3025) <= a and b;
    outputs(3026) <= a xor b;
    outputs(3027) <= not b;
    outputs(3028) <= b;
    outputs(3029) <= b;
    outputs(3030) <= not a;
    outputs(3031) <= not b or a;
    outputs(3032) <= not (a and b);
    outputs(3033) <= not (a xor b);
    outputs(3034) <= a and b;
    outputs(3035) <= not (a xor b);
    outputs(3036) <= not b;
    outputs(3037) <= a and b;
    outputs(3038) <= not b;
    outputs(3039) <= not a or b;
    outputs(3040) <= not a;
    outputs(3041) <= not a;
    outputs(3042) <= b;
    outputs(3043) <= not (a xor b);
    outputs(3044) <= b;
    outputs(3045) <= a and b;
    outputs(3046) <= not b;
    outputs(3047) <= b;
    outputs(3048) <= a;
    outputs(3049) <= a;
    outputs(3050) <= not (a xor b);
    outputs(3051) <= not a;
    outputs(3052) <= not b;
    outputs(3053) <= not (a xor b);
    outputs(3054) <= a xor b;
    outputs(3055) <= not b;
    outputs(3056) <= b;
    outputs(3057) <= a;
    outputs(3058) <= not a or b;
    outputs(3059) <= b;
    outputs(3060) <= b and not a;
    outputs(3061) <= b;
    outputs(3062) <= a;
    outputs(3063) <= not a or b;
    outputs(3064) <= not b;
    outputs(3065) <= not a or b;
    outputs(3066) <= not b;
    outputs(3067) <= a or b;
    outputs(3068) <= b;
    outputs(3069) <= not a or b;
    outputs(3070) <= a or b;
    outputs(3071) <= b;
    outputs(3072) <= not b;
    outputs(3073) <= a xor b;
    outputs(3074) <= b;
    outputs(3075) <= b;
    outputs(3076) <= a xor b;
    outputs(3077) <= not b;
    outputs(3078) <= not b;
    outputs(3079) <= not b;
    outputs(3080) <= b;
    outputs(3081) <= not b;
    outputs(3082) <= a and b;
    outputs(3083) <= a xor b;
    outputs(3084) <= a;
    outputs(3085) <= a xor b;
    outputs(3086) <= a;
    outputs(3087) <= not (a or b);
    outputs(3088) <= not (a xor b);
    outputs(3089) <= b;
    outputs(3090) <= a xor b;
    outputs(3091) <= not b;
    outputs(3092) <= a or b;
    outputs(3093) <= not a;
    outputs(3094) <= not (a or b);
    outputs(3095) <= a;
    outputs(3096) <= b;
    outputs(3097) <= a or b;
    outputs(3098) <= a;
    outputs(3099) <= a xor b;
    outputs(3100) <= a;
    outputs(3101) <= a xor b;
    outputs(3102) <= b;
    outputs(3103) <= not b;
    outputs(3104) <= not (a or b);
    outputs(3105) <= a and not b;
    outputs(3106) <= not b or a;
    outputs(3107) <= not b or a;
    outputs(3108) <= not a;
    outputs(3109) <= not (a xor b);
    outputs(3110) <= not b;
    outputs(3111) <= a and not b;
    outputs(3112) <= a xor b;
    outputs(3113) <= a xor b;
    outputs(3114) <= not (a and b);
    outputs(3115) <= a and b;
    outputs(3116) <= a xor b;
    outputs(3117) <= not a;
    outputs(3118) <= b and not a;
    outputs(3119) <= not b;
    outputs(3120) <= not (a or b);
    outputs(3121) <= not (a xor b);
    outputs(3122) <= a;
    outputs(3123) <= a and b;
    outputs(3124) <= b and not a;
    outputs(3125) <= not b;
    outputs(3126) <= a;
    outputs(3127) <= a or b;
    outputs(3128) <= b;
    outputs(3129) <= a xor b;
    outputs(3130) <= b;
    outputs(3131) <= not (a xor b);
    outputs(3132) <= not a;
    outputs(3133) <= b;
    outputs(3134) <= not a;
    outputs(3135) <= a and not b;
    outputs(3136) <= not (a xor b);
    outputs(3137) <= a and not b;
    outputs(3138) <= not a or b;
    outputs(3139) <= not a;
    outputs(3140) <= b;
    outputs(3141) <= b;
    outputs(3142) <= not a;
    outputs(3143) <= not b;
    outputs(3144) <= not (a xor b);
    outputs(3145) <= not a or b;
    outputs(3146) <= b;
    outputs(3147) <= not b;
    outputs(3148) <= b;
    outputs(3149) <= a;
    outputs(3150) <= a xor b;
    outputs(3151) <= a;
    outputs(3152) <= not b;
    outputs(3153) <= b;
    outputs(3154) <= not b;
    outputs(3155) <= not (a xor b);
    outputs(3156) <= not (a xor b);
    outputs(3157) <= b;
    outputs(3158) <= a xor b;
    outputs(3159) <= a and not b;
    outputs(3160) <= not b or a;
    outputs(3161) <= a xor b;
    outputs(3162) <= a and not b;
    outputs(3163) <= a;
    outputs(3164) <= a xor b;
    outputs(3165) <= a xor b;
    outputs(3166) <= a and b;
    outputs(3167) <= not a;
    outputs(3168) <= not (a xor b);
    outputs(3169) <= not a;
    outputs(3170) <= b and not a;
    outputs(3171) <= b;
    outputs(3172) <= not b;
    outputs(3173) <= not a;
    outputs(3174) <= not a;
    outputs(3175) <= not (a xor b);
    outputs(3176) <= b;
    outputs(3177) <= a;
    outputs(3178) <= not b;
    outputs(3179) <= a xor b;
    outputs(3180) <= not (a and b);
    outputs(3181) <= not (a xor b);
    outputs(3182) <= a;
    outputs(3183) <= not b;
    outputs(3184) <= a;
    outputs(3185) <= b;
    outputs(3186) <= a;
    outputs(3187) <= not (a xor b);
    outputs(3188) <= not (a xor b);
    outputs(3189) <= a;
    outputs(3190) <= a and not b;
    outputs(3191) <= not (a xor b);
    outputs(3192) <= a and not b;
    outputs(3193) <= not (a xor b);
    outputs(3194) <= a xor b;
    outputs(3195) <= not a or b;
    outputs(3196) <= a xor b;
    outputs(3197) <= not (a xor b);
    outputs(3198) <= not a;
    outputs(3199) <= not (a xor b);
    outputs(3200) <= a;
    outputs(3201) <= a xor b;
    outputs(3202) <= b and not a;
    outputs(3203) <= b;
    outputs(3204) <= a and not b;
    outputs(3205) <= b;
    outputs(3206) <= a;
    outputs(3207) <= a;
    outputs(3208) <= a and b;
    outputs(3209) <= a xor b;
    outputs(3210) <= not (a xor b);
    outputs(3211) <= not (a xor b);
    outputs(3212) <= b;
    outputs(3213) <= not (a xor b);
    outputs(3214) <= a xor b;
    outputs(3215) <= a xor b;
    outputs(3216) <= not a;
    outputs(3217) <= not a;
    outputs(3218) <= b and not a;
    outputs(3219) <= a xor b;
    outputs(3220) <= a xor b;
    outputs(3221) <= a;
    outputs(3222) <= not (a or b);
    outputs(3223) <= not b;
    outputs(3224) <= not a;
    outputs(3225) <= not b;
    outputs(3226) <= b and not a;
    outputs(3227) <= not (a xor b);
    outputs(3228) <= not (a xor b);
    outputs(3229) <= not a;
    outputs(3230) <= not a;
    outputs(3231) <= not (a xor b);
    outputs(3232) <= a;
    outputs(3233) <= b;
    outputs(3234) <= a xor b;
    outputs(3235) <= a and not b;
    outputs(3236) <= b;
    outputs(3237) <= a;
    outputs(3238) <= not (a and b);
    outputs(3239) <= not a;
    outputs(3240) <= a;
    outputs(3241) <= not (a and b);
    outputs(3242) <= a xor b;
    outputs(3243) <= not b or a;
    outputs(3244) <= not b;
    outputs(3245) <= not (a and b);
    outputs(3246) <= b;
    outputs(3247) <= a or b;
    outputs(3248) <= not b;
    outputs(3249) <= a xor b;
    outputs(3250) <= a and b;
    outputs(3251) <= not b;
    outputs(3252) <= a xor b;
    outputs(3253) <= not (a xor b);
    outputs(3254) <= not (a xor b);
    outputs(3255) <= not b;
    outputs(3256) <= a;
    outputs(3257) <= not (a xor b);
    outputs(3258) <= not a;
    outputs(3259) <= not a;
    outputs(3260) <= not b or a;
    outputs(3261) <= not (a or b);
    outputs(3262) <= a xor b;
    outputs(3263) <= not (a xor b);
    outputs(3264) <= not a;
    outputs(3265) <= not (a or b);
    outputs(3266) <= not a;
    outputs(3267) <= not a;
    outputs(3268) <= b and not a;
    outputs(3269) <= b and not a;
    outputs(3270) <= not (a xor b);
    outputs(3271) <= a;
    outputs(3272) <= b;
    outputs(3273) <= not b or a;
    outputs(3274) <= a;
    outputs(3275) <= not (a xor b);
    outputs(3276) <= not b;
    outputs(3277) <= not (a or b);
    outputs(3278) <= a xor b;
    outputs(3279) <= a;
    outputs(3280) <= a xor b;
    outputs(3281) <= a;
    outputs(3282) <= not (a or b);
    outputs(3283) <= a xor b;
    outputs(3284) <= not a;
    outputs(3285) <= a xor b;
    outputs(3286) <= not b;
    outputs(3287) <= a xor b;
    outputs(3288) <= not a;
    outputs(3289) <= a xor b;
    outputs(3290) <= a;
    outputs(3291) <= b;
    outputs(3292) <= not (a or b);
    outputs(3293) <= a;
    outputs(3294) <= b and not a;
    outputs(3295) <= not b;
    outputs(3296) <= not (a xor b);
    outputs(3297) <= a and b;
    outputs(3298) <= not b;
    outputs(3299) <= not (a xor b);
    outputs(3300) <= a;
    outputs(3301) <= not a;
    outputs(3302) <= b;
    outputs(3303) <= a;
    outputs(3304) <= a;
    outputs(3305) <= a xor b;
    outputs(3306) <= not (a xor b);
    outputs(3307) <= a;
    outputs(3308) <= a;
    outputs(3309) <= b;
    outputs(3310) <= not a or b;
    outputs(3311) <= not (a xor b);
    outputs(3312) <= a and not b;
    outputs(3313) <= a or b;
    outputs(3314) <= a;
    outputs(3315) <= b and not a;
    outputs(3316) <= not (a xor b);
    outputs(3317) <= b;
    outputs(3318) <= a xor b;
    outputs(3319) <= a xor b;
    outputs(3320) <= not a;
    outputs(3321) <= not a or b;
    outputs(3322) <= a xor b;
    outputs(3323) <= a xor b;
    outputs(3324) <= b;
    outputs(3325) <= b and not a;
    outputs(3326) <= not (a or b);
    outputs(3327) <= not (a xor b);
    outputs(3328) <= not (a xor b);
    outputs(3329) <= b and not a;
    outputs(3330) <= a;
    outputs(3331) <= a xor b;
    outputs(3332) <= a xor b;
    outputs(3333) <= a xor b;
    outputs(3334) <= not a or b;
    outputs(3335) <= a xor b;
    outputs(3336) <= b;
    outputs(3337) <= not a;
    outputs(3338) <= not a;
    outputs(3339) <= b;
    outputs(3340) <= b;
    outputs(3341) <= a xor b;
    outputs(3342) <= a xor b;
    outputs(3343) <= not (a xor b);
    outputs(3344) <= a;
    outputs(3345) <= b;
    outputs(3346) <= a;
    outputs(3347) <= not a;
    outputs(3348) <= not (a xor b);
    outputs(3349) <= not (a xor b);
    outputs(3350) <= not b;
    outputs(3351) <= b;
    outputs(3352) <= a xor b;
    outputs(3353) <= not (a xor b);
    outputs(3354) <= b and not a;
    outputs(3355) <= not b;
    outputs(3356) <= not a;
    outputs(3357) <= a xor b;
    outputs(3358) <= not (a xor b);
    outputs(3359) <= a or b;
    outputs(3360) <= not (a xor b);
    outputs(3361) <= a xor b;
    outputs(3362) <= a xor b;
    outputs(3363) <= b;
    outputs(3364) <= a xor b;
    outputs(3365) <= not b;
    outputs(3366) <= not b;
    outputs(3367) <= not a;
    outputs(3368) <= not (a or b);
    outputs(3369) <= a xor b;
    outputs(3370) <= not b;
    outputs(3371) <= not b;
    outputs(3372) <= a xor b;
    outputs(3373) <= not (a xor b);
    outputs(3374) <= b;
    outputs(3375) <= not (a and b);
    outputs(3376) <= not (a xor b);
    outputs(3377) <= not (a or b);
    outputs(3378) <= not b;
    outputs(3379) <= a and b;
    outputs(3380) <= not a;
    outputs(3381) <= b;
    outputs(3382) <= not a;
    outputs(3383) <= not a;
    outputs(3384) <= not a;
    outputs(3385) <= a and not b;
    outputs(3386) <= not b;
    outputs(3387) <= b;
    outputs(3388) <= a;
    outputs(3389) <= a and not b;
    outputs(3390) <= a;
    outputs(3391) <= not b;
    outputs(3392) <= not a or b;
    outputs(3393) <= b;
    outputs(3394) <= a;
    outputs(3395) <= not b;
    outputs(3396) <= a xor b;
    outputs(3397) <= a or b;
    outputs(3398) <= not (a xor b);
    outputs(3399) <= a xor b;
    outputs(3400) <= not a;
    outputs(3401) <= a;
    outputs(3402) <= not a;
    outputs(3403) <= a;
    outputs(3404) <= a xor b;
    outputs(3405) <= a xor b;
    outputs(3406) <= a xor b;
    outputs(3407) <= a xor b;
    outputs(3408) <= b;
    outputs(3409) <= not (a xor b);
    outputs(3410) <= not b;
    outputs(3411) <= not a;
    outputs(3412) <= b;
    outputs(3413) <= not a;
    outputs(3414) <= not (a xor b);
    outputs(3415) <= not (a xor b);
    outputs(3416) <= not a;
    outputs(3417) <= not (a or b);
    outputs(3418) <= b;
    outputs(3419) <= a;
    outputs(3420) <= not (a and b);
    outputs(3421) <= not a;
    outputs(3422) <= not a;
    outputs(3423) <= a;
    outputs(3424) <= a and b;
    outputs(3425) <= a xor b;
    outputs(3426) <= not a;
    outputs(3427) <= a;
    outputs(3428) <= not a;
    outputs(3429) <= not (a xor b);
    outputs(3430) <= not (a xor b);
    outputs(3431) <= a or b;
    outputs(3432) <= not (a xor b);
    outputs(3433) <= not b;
    outputs(3434) <= a and not b;
    outputs(3435) <= not (a xor b);
    outputs(3436) <= b;
    outputs(3437) <= a xor b;
    outputs(3438) <= a;
    outputs(3439) <= not (a or b);
    outputs(3440) <= a xor b;
    outputs(3441) <= not (a xor b);
    outputs(3442) <= not b;
    outputs(3443) <= not b or a;
    outputs(3444) <= not (a and b);
    outputs(3445) <= a xor b;
    outputs(3446) <= b;
    outputs(3447) <= a and not b;
    outputs(3448) <= not a;
    outputs(3449) <= not (a xor b);
    outputs(3450) <= not b;
    outputs(3451) <= not (a or b);
    outputs(3452) <= not a;
    outputs(3453) <= not (a xor b);
    outputs(3454) <= not b;
    outputs(3455) <= b and not a;
    outputs(3456) <= a and not b;
    outputs(3457) <= a;
    outputs(3458) <= not (a and b);
    outputs(3459) <= b;
    outputs(3460) <= not (a xor b);
    outputs(3461) <= not (a xor b);
    outputs(3462) <= not (a xor b);
    outputs(3463) <= not (a or b);
    outputs(3464) <= a xor b;
    outputs(3465) <= not b;
    outputs(3466) <= a xor b;
    outputs(3467) <= not a;
    outputs(3468) <= not (a xor b);
    outputs(3469) <= a xor b;
    outputs(3470) <= not b or a;
    outputs(3471) <= not (a xor b);
    outputs(3472) <= a;
    outputs(3473) <= not a;
    outputs(3474) <= not b or a;
    outputs(3475) <= not a;
    outputs(3476) <= not a;
    outputs(3477) <= a xor b;
    outputs(3478) <= a;
    outputs(3479) <= not (a or b);
    outputs(3480) <= a xor b;
    outputs(3481) <= not b or a;
    outputs(3482) <= a and b;
    outputs(3483) <= not (a xor b);
    outputs(3484) <= a xor b;
    outputs(3485) <= not (a xor b);
    outputs(3486) <= not a;
    outputs(3487) <= not a or b;
    outputs(3488) <= b and not a;
    outputs(3489) <= not a;
    outputs(3490) <= not (a xor b);
    outputs(3491) <= b and not a;
    outputs(3492) <= not b;
    outputs(3493) <= a;
    outputs(3494) <= a xor b;
    outputs(3495) <= not (a xor b);
    outputs(3496) <= a or b;
    outputs(3497) <= not (a or b);
    outputs(3498) <= a xor b;
    outputs(3499) <= b;
    outputs(3500) <= a or b;
    outputs(3501) <= not (a xor b);
    outputs(3502) <= not b;
    outputs(3503) <= b;
    outputs(3504) <= not (a xor b);
    outputs(3505) <= not (a xor b);
    outputs(3506) <= a;
    outputs(3507) <= a and not b;
    outputs(3508) <= not (a xor b);
    outputs(3509) <= a;
    outputs(3510) <= not a;
    outputs(3511) <= not a;
    outputs(3512) <= b;
    outputs(3513) <= a and b;
    outputs(3514) <= not a;
    outputs(3515) <= not (a xor b);
    outputs(3516) <= b;
    outputs(3517) <= not b;
    outputs(3518) <= a xor b;
    outputs(3519) <= b;
    outputs(3520) <= a;
    outputs(3521) <= b;
    outputs(3522) <= a or b;
    outputs(3523) <= not a;
    outputs(3524) <= a xor b;
    outputs(3525) <= a xor b;
    outputs(3526) <= not a;
    outputs(3527) <= not (a or b);
    outputs(3528) <= not b;
    outputs(3529) <= a xor b;
    outputs(3530) <= a;
    outputs(3531) <= a xor b;
    outputs(3532) <= b;
    outputs(3533) <= a xor b;
    outputs(3534) <= b;
    outputs(3535) <= b;
    outputs(3536) <= a and not b;
    outputs(3537) <= a xor b;
    outputs(3538) <= b;
    outputs(3539) <= not b;
    outputs(3540) <= not (a xor b);
    outputs(3541) <= a;
    outputs(3542) <= not b or a;
    outputs(3543) <= a xor b;
    outputs(3544) <= not a;
    outputs(3545) <= not a or b;
    outputs(3546) <= not (a xor b);
    outputs(3547) <= not b;
    outputs(3548) <= a or b;
    outputs(3549) <= not a;
    outputs(3550) <= not a;
    outputs(3551) <= not (a xor b);
    outputs(3552) <= not b;
    outputs(3553) <= not b or a;
    outputs(3554) <= b;
    outputs(3555) <= a;
    outputs(3556) <= not b;
    outputs(3557) <= a xor b;
    outputs(3558) <= b and not a;
    outputs(3559) <= b;
    outputs(3560) <= not (a xor b);
    outputs(3561) <= not b;
    outputs(3562) <= not (a xor b);
    outputs(3563) <= not b;
    outputs(3564) <= not a;
    outputs(3565) <= not b or a;
    outputs(3566) <= a xor b;
    outputs(3567) <= b;
    outputs(3568) <= a;
    outputs(3569) <= b and not a;
    outputs(3570) <= not (a xor b);
    outputs(3571) <= a and b;
    outputs(3572) <= not (a or b);
    outputs(3573) <= not a or b;
    outputs(3574) <= a or b;
    outputs(3575) <= b;
    outputs(3576) <= a;
    outputs(3577) <= a;
    outputs(3578) <= not b or a;
    outputs(3579) <= b;
    outputs(3580) <= not (a xor b);
    outputs(3581) <= not (a xor b);
    outputs(3582) <= a;
    outputs(3583) <= not a;
    outputs(3584) <= not a;
    outputs(3585) <= not (a or b);
    outputs(3586) <= a;
    outputs(3587) <= a;
    outputs(3588) <= not a;
    outputs(3589) <= a and not b;
    outputs(3590) <= not (a or b);
    outputs(3591) <= not b or a;
    outputs(3592) <= not b;
    outputs(3593) <= a xor b;
    outputs(3594) <= a xor b;
    outputs(3595) <= a;
    outputs(3596) <= a xor b;
    outputs(3597) <= not a;
    outputs(3598) <= not b;
    outputs(3599) <= b;
    outputs(3600) <= not (a xor b);
    outputs(3601) <= b and not a;
    outputs(3602) <= not a;
    outputs(3603) <= b;
    outputs(3604) <= not a;
    outputs(3605) <= not a or b;
    outputs(3606) <= not (a or b);
    outputs(3607) <= not a;
    outputs(3608) <= b;
    outputs(3609) <= a;
    outputs(3610) <= not (a xor b);
    outputs(3611) <= not (a xor b);
    outputs(3612) <= a xor b;
    outputs(3613) <= a;
    outputs(3614) <= not (a or b);
    outputs(3615) <= not (a xor b);
    outputs(3616) <= not a;
    outputs(3617) <= not b or a;
    outputs(3618) <= a xor b;
    outputs(3619) <= not (a xor b);
    outputs(3620) <= a and b;
    outputs(3621) <= not b;
    outputs(3622) <= a xor b;
    outputs(3623) <= not b or a;
    outputs(3624) <= not (a xor b);
    outputs(3625) <= a xor b;
    outputs(3626) <= not b;
    outputs(3627) <= not (a and b);
    outputs(3628) <= b;
    outputs(3629) <= b and not a;
    outputs(3630) <= not (a xor b);
    outputs(3631) <= a xor b;
    outputs(3632) <= not (a xor b);
    outputs(3633) <= a or b;
    outputs(3634) <= not a;
    outputs(3635) <= not (a xor b);
    outputs(3636) <= not (a xor b);
    outputs(3637) <= not a;
    outputs(3638) <= b;
    outputs(3639) <= a;
    outputs(3640) <= not b or a;
    outputs(3641) <= a xor b;
    outputs(3642) <= not (a xor b);
    outputs(3643) <= not (a xor b);
    outputs(3644) <= not a;
    outputs(3645) <= not b;
    outputs(3646) <= not (a xor b);
    outputs(3647) <= a xor b;
    outputs(3648) <= b;
    outputs(3649) <= not a;
    outputs(3650) <= a and not b;
    outputs(3651) <= not b;
    outputs(3652) <= b;
    outputs(3653) <= a;
    outputs(3654) <= not (a or b);
    outputs(3655) <= a or b;
    outputs(3656) <= b;
    outputs(3657) <= a or b;
    outputs(3658) <= not b;
    outputs(3659) <= not b;
    outputs(3660) <= not b;
    outputs(3661) <= not (a xor b);
    outputs(3662) <= not b or a;
    outputs(3663) <= not b;
    outputs(3664) <= a;
    outputs(3665) <= not a;
    outputs(3666) <= not a or b;
    outputs(3667) <= b and not a;
    outputs(3668) <= not (a xor b);
    outputs(3669) <= a and b;
    outputs(3670) <= a xor b;
    outputs(3671) <= not (a or b);
    outputs(3672) <= a xor b;
    outputs(3673) <= a;
    outputs(3674) <= a;
    outputs(3675) <= not a;
    outputs(3676) <= not (a xor b);
    outputs(3677) <= not a or b;
    outputs(3678) <= not b;
    outputs(3679) <= b;
    outputs(3680) <= a xor b;
    outputs(3681) <= not b;
    outputs(3682) <= b;
    outputs(3683) <= a and b;
    outputs(3684) <= not b;
    outputs(3685) <= b;
    outputs(3686) <= a;
    outputs(3687) <= a xor b;
    outputs(3688) <= not (a or b);
    outputs(3689) <= not b;
    outputs(3690) <= not a;
    outputs(3691) <= a;
    outputs(3692) <= b;
    outputs(3693) <= a xor b;
    outputs(3694) <= not a;
    outputs(3695) <= not (a and b);
    outputs(3696) <= a;
    outputs(3697) <= not b;
    outputs(3698) <= b and not a;
    outputs(3699) <= a xor b;
    outputs(3700) <= a and b;
    outputs(3701) <= not (a and b);
    outputs(3702) <= a;
    outputs(3703) <= b;
    outputs(3704) <= a xor b;
    outputs(3705) <= not b;
    outputs(3706) <= not a;
    outputs(3707) <= a;
    outputs(3708) <= not (a and b);
    outputs(3709) <= not (a or b);
    outputs(3710) <= not (a or b);
    outputs(3711) <= not (a xor b);
    outputs(3712) <= not (a xor b);
    outputs(3713) <= a;
    outputs(3714) <= not b;
    outputs(3715) <= not b;
    outputs(3716) <= b;
    outputs(3717) <= a or b;
    outputs(3718) <= not (a xor b);
    outputs(3719) <= a;
    outputs(3720) <= a and not b;
    outputs(3721) <= a xor b;
    outputs(3722) <= a and b;
    outputs(3723) <= not a;
    outputs(3724) <= not (a xor b);
    outputs(3725) <= not (a xor b);
    outputs(3726) <= b;
    outputs(3727) <= not (a xor b);
    outputs(3728) <= b;
    outputs(3729) <= not (a xor b);
    outputs(3730) <= a or b;
    outputs(3731) <= not (a and b);
    outputs(3732) <= not b;
    outputs(3733) <= not a or b;
    outputs(3734) <= b;
    outputs(3735) <= not (a xor b);
    outputs(3736) <= not (a xor b);
    outputs(3737) <= not a or b;
    outputs(3738) <= b and not a;
    outputs(3739) <= a or b;
    outputs(3740) <= not a;
    outputs(3741) <= a xor b;
    outputs(3742) <= b;
    outputs(3743) <= a and b;
    outputs(3744) <= a;
    outputs(3745) <= b;
    outputs(3746) <= not a or b;
    outputs(3747) <= a and not b;
    outputs(3748) <= not b;
    outputs(3749) <= not (a xor b);
    outputs(3750) <= not a;
    outputs(3751) <= not b;
    outputs(3752) <= a xor b;
    outputs(3753) <= not a;
    outputs(3754) <= a;
    outputs(3755) <= not a;
    outputs(3756) <= a xor b;
    outputs(3757) <= a xor b;
    outputs(3758) <= b and not a;
    outputs(3759) <= b;
    outputs(3760) <= a xor b;
    outputs(3761) <= not (a xor b);
    outputs(3762) <= a xor b;
    outputs(3763) <= a and not b;
    outputs(3764) <= b;
    outputs(3765) <= not (a xor b);
    outputs(3766) <= a xor b;
    outputs(3767) <= not (a xor b);
    outputs(3768) <= not b;
    outputs(3769) <= not (a xor b);
    outputs(3770) <= a xor b;
    outputs(3771) <= not b;
    outputs(3772) <= not (a xor b);
    outputs(3773) <= not b;
    outputs(3774) <= b and not a;
    outputs(3775) <= a;
    outputs(3776) <= not (a or b);
    outputs(3777) <= a;
    outputs(3778) <= not (a xor b);
    outputs(3779) <= a;
    outputs(3780) <= not b;
    outputs(3781) <= not (a or b);
    outputs(3782) <= not b;
    outputs(3783) <= a xor b;
    outputs(3784) <= a or b;
    outputs(3785) <= not a;
    outputs(3786) <= not (a and b);
    outputs(3787) <= a;
    outputs(3788) <= not a or b;
    outputs(3789) <= b;
    outputs(3790) <= not (a xor b);
    outputs(3791) <= b;
    outputs(3792) <= a;
    outputs(3793) <= b;
    outputs(3794) <= b and not a;
    outputs(3795) <= a and b;
    outputs(3796) <= not a or b;
    outputs(3797) <= a xor b;
    outputs(3798) <= a xor b;
    outputs(3799) <= not (a xor b);
    outputs(3800) <= a xor b;
    outputs(3801) <= a and b;
    outputs(3802) <= b;
    outputs(3803) <= not (a xor b);
    outputs(3804) <= b;
    outputs(3805) <= not (a xor b);
    outputs(3806) <= not (a or b);
    outputs(3807) <= a xor b;
    outputs(3808) <= a and b;
    outputs(3809) <= not (a xor b);
    outputs(3810) <= b;
    outputs(3811) <= b;
    outputs(3812) <= a xor b;
    outputs(3813) <= a;
    outputs(3814) <= not b or a;
    outputs(3815) <= not b;
    outputs(3816) <= a xor b;
    outputs(3817) <= not (a and b);
    outputs(3818) <= a;
    outputs(3819) <= not a;
    outputs(3820) <= not (a xor b);
    outputs(3821) <= not (a xor b);
    outputs(3822) <= a xor b;
    outputs(3823) <= not (a xor b);
    outputs(3824) <= a xor b;
    outputs(3825) <= a;
    outputs(3826) <= b;
    outputs(3827) <= not (a xor b);
    outputs(3828) <= not b or a;
    outputs(3829) <= not a;
    outputs(3830) <= not b;
    outputs(3831) <= a;
    outputs(3832) <= a xor b;
    outputs(3833) <= not a;
    outputs(3834) <= b and not a;
    outputs(3835) <= not a or b;
    outputs(3836) <= not (a xor b);
    outputs(3837) <= a or b;
    outputs(3838) <= a xor b;
    outputs(3839) <= not (a xor b);
    outputs(3840) <= a xor b;
    outputs(3841) <= not a or b;
    outputs(3842) <= b;
    outputs(3843) <= b;
    outputs(3844) <= not (a or b);
    outputs(3845) <= not (a xor b);
    outputs(3846) <= not (a xor b);
    outputs(3847) <= b;
    outputs(3848) <= a;
    outputs(3849) <= b and not a;
    outputs(3850) <= b;
    outputs(3851) <= b;
    outputs(3852) <= not b or a;
    outputs(3853) <= a xor b;
    outputs(3854) <= not a;
    outputs(3855) <= not a;
    outputs(3856) <= not a;
    outputs(3857) <= not a;
    outputs(3858) <= not b;
    outputs(3859) <= a;
    outputs(3860) <= not (a xor b);
    outputs(3861) <= a;
    outputs(3862) <= not (a xor b);
    outputs(3863) <= b and not a;
    outputs(3864) <= not b;
    outputs(3865) <= not (a xor b);
    outputs(3866) <= not a or b;
    outputs(3867) <= not (a xor b);
    outputs(3868) <= a xor b;
    outputs(3869) <= not a;
    outputs(3870) <= a and not b;
    outputs(3871) <= not (a xor b);
    outputs(3872) <= b;
    outputs(3873) <= not b;
    outputs(3874) <= not (a xor b);
    outputs(3875) <= not (a xor b);
    outputs(3876) <= not a;
    outputs(3877) <= a and not b;
    outputs(3878) <= not (a and b);
    outputs(3879) <= b and not a;
    outputs(3880) <= a;
    outputs(3881) <= b;
    outputs(3882) <= not (a xor b);
    outputs(3883) <= not a;
    outputs(3884) <= not (a xor b);
    outputs(3885) <= a and b;
    outputs(3886) <= a xor b;
    outputs(3887) <= not (a xor b);
    outputs(3888) <= not (a xor b);
    outputs(3889) <= not (a or b);
    outputs(3890) <= a xor b;
    outputs(3891) <= not (a xor b);
    outputs(3892) <= a and b;
    outputs(3893) <= not b or a;
    outputs(3894) <= not (a xor b);
    outputs(3895) <= a and b;
    outputs(3896) <= a xor b;
    outputs(3897) <= not (a xor b);
    outputs(3898) <= a xor b;
    outputs(3899) <= a;
    outputs(3900) <= a;
    outputs(3901) <= a xor b;
    outputs(3902) <= not a or b;
    outputs(3903) <= a xor b;
    outputs(3904) <= b;
    outputs(3905) <= a and b;
    outputs(3906) <= b and not a;
    outputs(3907) <= b;
    outputs(3908) <= not a;
    outputs(3909) <= a xor b;
    outputs(3910) <= not a;
    outputs(3911) <= not (a xor b);
    outputs(3912) <= not b;
    outputs(3913) <= b;
    outputs(3914) <= b;
    outputs(3915) <= b;
    outputs(3916) <= a xor b;
    outputs(3917) <= b;
    outputs(3918) <= a and not b;
    outputs(3919) <= not (a xor b);
    outputs(3920) <= not a;
    outputs(3921) <= a and b;
    outputs(3922) <= a xor b;
    outputs(3923) <= a;
    outputs(3924) <= a xor b;
    outputs(3925) <= a xor b;
    outputs(3926) <= b;
    outputs(3927) <= b;
    outputs(3928) <= b;
    outputs(3929) <= not (a xor b);
    outputs(3930) <= not (a xor b);
    outputs(3931) <= a;
    outputs(3932) <= not a;
    outputs(3933) <= a;
    outputs(3934) <= a or b;
    outputs(3935) <= a;
    outputs(3936) <= not b;
    outputs(3937) <= a and not b;
    outputs(3938) <= a and not b;
    outputs(3939) <= a or b;
    outputs(3940) <= not (a xor b);
    outputs(3941) <= not (a and b);
    outputs(3942) <= b;
    outputs(3943) <= not (a xor b);
    outputs(3944) <= a and not b;
    outputs(3945) <= not b;
    outputs(3946) <= a xor b;
    outputs(3947) <= a or b;
    outputs(3948) <= not (a xor b);
    outputs(3949) <= not a;
    outputs(3950) <= not (a xor b);
    outputs(3951) <= a;
    outputs(3952) <= b and not a;
    outputs(3953) <= not b;
    outputs(3954) <= not a;
    outputs(3955) <= not b;
    outputs(3956) <= not a;
    outputs(3957) <= b;
    outputs(3958) <= not (a xor b);
    outputs(3959) <= a;
    outputs(3960) <= a or b;
    outputs(3961) <= not (a and b);
    outputs(3962) <= not (a or b);
    outputs(3963) <= not (a xor b);
    outputs(3964) <= not a;
    outputs(3965) <= not a;
    outputs(3966) <= not a or b;
    outputs(3967) <= b and not a;
    outputs(3968) <= not a;
    outputs(3969) <= not b or a;
    outputs(3970) <= not (a and b);
    outputs(3971) <= b and not a;
    outputs(3972) <= not (a or b);
    outputs(3973) <= a xor b;
    outputs(3974) <= a;
    outputs(3975) <= a and b;
    outputs(3976) <= not (a xor b);
    outputs(3977) <= b;
    outputs(3978) <= not a;
    outputs(3979) <= a and b;
    outputs(3980) <= a;
    outputs(3981) <= b;
    outputs(3982) <= not b;
    outputs(3983) <= a xor b;
    outputs(3984) <= a xor b;
    outputs(3985) <= not b;
    outputs(3986) <= b;
    outputs(3987) <= not (a or b);
    outputs(3988) <= not b;
    outputs(3989) <= a or b;
    outputs(3990) <= a and b;
    outputs(3991) <= not (a xor b);
    outputs(3992) <= not (a and b);
    outputs(3993) <= not (a xor b);
    outputs(3994) <= a;
    outputs(3995) <= not (a xor b);
    outputs(3996) <= not a;
    outputs(3997) <= a;
    outputs(3998) <= a xor b;
    outputs(3999) <= a;
    outputs(4000) <= not a;
    outputs(4001) <= not b;
    outputs(4002) <= not (a and b);
    outputs(4003) <= not b or a;
    outputs(4004) <= a xor b;
    outputs(4005) <= b;
    outputs(4006) <= b;
    outputs(4007) <= b and not a;
    outputs(4008) <= a;
    outputs(4009) <= not b;
    outputs(4010) <= a and not b;
    outputs(4011) <= a and not b;
    outputs(4012) <= not (a and b);
    outputs(4013) <= not a;
    outputs(4014) <= not b;
    outputs(4015) <= not b;
    outputs(4016) <= not (a xor b);
    outputs(4017) <= not a;
    outputs(4018) <= b and not a;
    outputs(4019) <= not b or a;
    outputs(4020) <= b;
    outputs(4021) <= b;
    outputs(4022) <= b;
    outputs(4023) <= a xor b;
    outputs(4024) <= a xor b;
    outputs(4025) <= b and not a;
    outputs(4026) <= not a;
    outputs(4027) <= a;
    outputs(4028) <= not a or b;
    outputs(4029) <= not (a xor b);
    outputs(4030) <= b;
    outputs(4031) <= not (a xor b);
    outputs(4032) <= a;
    outputs(4033) <= b;
    outputs(4034) <= not (a or b);
    outputs(4035) <= a and not b;
    outputs(4036) <= b;
    outputs(4037) <= a xor b;
    outputs(4038) <= a xor b;
    outputs(4039) <= not (a and b);
    outputs(4040) <= a xor b;
    outputs(4041) <= a xor b;
    outputs(4042) <= a xor b;
    outputs(4043) <= a xor b;
    outputs(4044) <= a xor b;
    outputs(4045) <= not b or a;
    outputs(4046) <= not a or b;
    outputs(4047) <= not b;
    outputs(4048) <= not (a xor b);
    outputs(4049) <= a xor b;
    outputs(4050) <= not a;
    outputs(4051) <= not (a and b);
    outputs(4052) <= a xor b;
    outputs(4053) <= not (a xor b);
    outputs(4054) <= a xor b;
    outputs(4055) <= a xor b;
    outputs(4056) <= not (a xor b);
    outputs(4057) <= not a;
    outputs(4058) <= not b;
    outputs(4059) <= not (a or b);
    outputs(4060) <= a;
    outputs(4061) <= a and not b;
    outputs(4062) <= b;
    outputs(4063) <= a and b;
    outputs(4064) <= b;
    outputs(4065) <= not b;
    outputs(4066) <= not b;
    outputs(4067) <= a;
    outputs(4068) <= b;
    outputs(4069) <= not a;
    outputs(4070) <= not b;
    outputs(4071) <= a or b;
    outputs(4072) <= b and not a;
    outputs(4073) <= not a;
    outputs(4074) <= a;
    outputs(4075) <= not (a xor b);
    outputs(4076) <= not (a xor b);
    outputs(4077) <= a;
    outputs(4078) <= not a;
    outputs(4079) <= a xor b;
    outputs(4080) <= not (a xor b);
    outputs(4081) <= a xor b;
    outputs(4082) <= not b;
    outputs(4083) <= b;
    outputs(4084) <= a xor b;
    outputs(4085) <= b;
    outputs(4086) <= not a or b;
    outputs(4087) <= not b or a;
    outputs(4088) <= a;
    outputs(4089) <= not a;
    outputs(4090) <= not a or b;
    outputs(4091) <= not a;
    outputs(4092) <= not b;
    outputs(4093) <= b;
    outputs(4094) <= b;
    outputs(4095) <= not a;
    outputs(4096) <= not (a xor b);
    outputs(4097) <= not b;
    outputs(4098) <= not (a xor b);
    outputs(4099) <= not b;
    outputs(4100) <= not a;
    outputs(4101) <= b;
    outputs(4102) <= a;
    outputs(4103) <= b and not a;
    outputs(4104) <= not a or b;
    outputs(4105) <= not (a and b);
    outputs(4106) <= a and not b;
    outputs(4107) <= a xor b;
    outputs(4108) <= not a;
    outputs(4109) <= a xor b;
    outputs(4110) <= not a;
    outputs(4111) <= a and b;
    outputs(4112) <= not a;
    outputs(4113) <= b;
    outputs(4114) <= a xor b;
    outputs(4115) <= not b;
    outputs(4116) <= a;
    outputs(4117) <= not a;
    outputs(4118) <= b;
    outputs(4119) <= b;
    outputs(4120) <= a and b;
    outputs(4121) <= b;
    outputs(4122) <= a xor b;
    outputs(4123) <= a;
    outputs(4124) <= not (a xor b);
    outputs(4125) <= a;
    outputs(4126) <= a;
    outputs(4127) <= a xor b;
    outputs(4128) <= not a;
    outputs(4129) <= not b;
    outputs(4130) <= not a;
    outputs(4131) <= a and not b;
    outputs(4132) <= a xor b;
    outputs(4133) <= a;
    outputs(4134) <= a xor b;
    outputs(4135) <= b;
    outputs(4136) <= not a;
    outputs(4137) <= a xor b;
    outputs(4138) <= a;
    outputs(4139) <= a xor b;
    outputs(4140) <= a;
    outputs(4141) <= a xor b;
    outputs(4142) <= a xor b;
    outputs(4143) <= not (a xor b);
    outputs(4144) <= b and not a;
    outputs(4145) <= not (a xor b);
    outputs(4146) <= not a;
    outputs(4147) <= a xor b;
    outputs(4148) <= not b or a;
    outputs(4149) <= not a;
    outputs(4150) <= a;
    outputs(4151) <= a;
    outputs(4152) <= b;
    outputs(4153) <= a;
    outputs(4154) <= a xor b;
    outputs(4155) <= not a;
    outputs(4156) <= a xor b;
    outputs(4157) <= not a;
    outputs(4158) <= a xor b;
    outputs(4159) <= a xor b;
    outputs(4160) <= not a;
    outputs(4161) <= not b;
    outputs(4162) <= b;
    outputs(4163) <= not a;
    outputs(4164) <= b;
    outputs(4165) <= a and not b;
    outputs(4166) <= not a;
    outputs(4167) <= not b;
    outputs(4168) <= b;
    outputs(4169) <= a xor b;
    outputs(4170) <= a and not b;
    outputs(4171) <= b;
    outputs(4172) <= not b;
    outputs(4173) <= not a;
    outputs(4174) <= not (a xor b);
    outputs(4175) <= not (a xor b);
    outputs(4176) <= a xor b;
    outputs(4177) <= not a;
    outputs(4178) <= a and b;
    outputs(4179) <= a xor b;
    outputs(4180) <= not b;
    outputs(4181) <= a xor b;
    outputs(4182) <= not (a xor b);
    outputs(4183) <= a or b;
    outputs(4184) <= not b;
    outputs(4185) <= not a;
    outputs(4186) <= a xor b;
    outputs(4187) <= a or b;
    outputs(4188) <= a;
    outputs(4189) <= not b;
    outputs(4190) <= not b;
    outputs(4191) <= b and not a;
    outputs(4192) <= not a;
    outputs(4193) <= a;
    outputs(4194) <= not a;
    outputs(4195) <= b;
    outputs(4196) <= a xor b;
    outputs(4197) <= not a;
    outputs(4198) <= not b;
    outputs(4199) <= not (a xor b);
    outputs(4200) <= not (a xor b);
    outputs(4201) <= not b;
    outputs(4202) <= not (a xor b);
    outputs(4203) <= not b;
    outputs(4204) <= not b;
    outputs(4205) <= not (a xor b);
    outputs(4206) <= not (a xor b);
    outputs(4207) <= a xor b;
    outputs(4208) <= not a;
    outputs(4209) <= not b;
    outputs(4210) <= a;
    outputs(4211) <= a xor b;
    outputs(4212) <= not b or a;
    outputs(4213) <= b;
    outputs(4214) <= not b;
    outputs(4215) <= not b or a;
    outputs(4216) <= not (a or b);
    outputs(4217) <= not b;
    outputs(4218) <= a;
    outputs(4219) <= b;
    outputs(4220) <= a xor b;
    outputs(4221) <= a xor b;
    outputs(4222) <= not b;
    outputs(4223) <= not a;
    outputs(4224) <= not (a xor b);
    outputs(4225) <= a xor b;
    outputs(4226) <= a xor b;
    outputs(4227) <= a or b;
    outputs(4228) <= a and not b;
    outputs(4229) <= a xor b;
    outputs(4230) <= a xor b;
    outputs(4231) <= not a;
    outputs(4232) <= a xor b;
    outputs(4233) <= a and not b;
    outputs(4234) <= not b;
    outputs(4235) <= not b;
    outputs(4236) <= not a;
    outputs(4237) <= not (a or b);
    outputs(4238) <= not a;
    outputs(4239) <= not b;
    outputs(4240) <= not b;
    outputs(4241) <= a xor b;
    outputs(4242) <= b;
    outputs(4243) <= not b;
    outputs(4244) <= not (a xor b);
    outputs(4245) <= not b;
    outputs(4246) <= a;
    outputs(4247) <= not (a xor b);
    outputs(4248) <= a xor b;
    outputs(4249) <= a xor b;
    outputs(4250) <= not (a xor b);
    outputs(4251) <= not b;
    outputs(4252) <= a xor b;
    outputs(4253) <= not (a xor b);
    outputs(4254) <= a xor b;
    outputs(4255) <= not b;
    outputs(4256) <= not b or a;
    outputs(4257) <= not (a xor b);
    outputs(4258) <= not a;
    outputs(4259) <= a and b;
    outputs(4260) <= a;
    outputs(4261) <= not (a and b);
    outputs(4262) <= not a;
    outputs(4263) <= not a or b;
    outputs(4264) <= a;
    outputs(4265) <= not a;
    outputs(4266) <= a xor b;
    outputs(4267) <= a or b;
    outputs(4268) <= not b;
    outputs(4269) <= not a;
    outputs(4270) <= a xor b;
    outputs(4271) <= not (a xor b);
    outputs(4272) <= b and not a;
    outputs(4273) <= b;
    outputs(4274) <= not a;
    outputs(4275) <= a and b;
    outputs(4276) <= a;
    outputs(4277) <= a xor b;
    outputs(4278) <= a or b;
    outputs(4279) <= a xor b;
    outputs(4280) <= b;
    outputs(4281) <= a xor b;
    outputs(4282) <= not b;
    outputs(4283) <= not a;
    outputs(4284) <= not (a and b);
    outputs(4285) <= not b;
    outputs(4286) <= not b or a;
    outputs(4287) <= b;
    outputs(4288) <= not (a xor b);
    outputs(4289) <= a or b;
    outputs(4290) <= not (a xor b);
    outputs(4291) <= not (a xor b);
    outputs(4292) <= not (a xor b);
    outputs(4293) <= not b;
    outputs(4294) <= a and not b;
    outputs(4295) <= b;
    outputs(4296) <= a and not b;
    outputs(4297) <= a xor b;
    outputs(4298) <= b;
    outputs(4299) <= not (a xor b);
    outputs(4300) <= a;
    outputs(4301) <= b and not a;
    outputs(4302) <= a and not b;
    outputs(4303) <= not a;
    outputs(4304) <= b and not a;
    outputs(4305) <= not a;
    outputs(4306) <= not a;
    outputs(4307) <= not a;
    outputs(4308) <= a and b;
    outputs(4309) <= a;
    outputs(4310) <= not (a and b);
    outputs(4311) <= not b or a;
    outputs(4312) <= b;
    outputs(4313) <= b;
    outputs(4314) <= not a;
    outputs(4315) <= not a or b;
    outputs(4316) <= not a or b;
    outputs(4317) <= not (a xor b);
    outputs(4318) <= not a;
    outputs(4319) <= not a or b;
    outputs(4320) <= a xor b;
    outputs(4321) <= not (a xor b);
    outputs(4322) <= not (a or b);
    outputs(4323) <= not b;
    outputs(4324) <= not (a or b);
    outputs(4325) <= a;
    outputs(4326) <= b;
    outputs(4327) <= not b;
    outputs(4328) <= not (a xor b);
    outputs(4329) <= not b or a;
    outputs(4330) <= not a or b;
    outputs(4331) <= b and not a;
    outputs(4332) <= a xor b;
    outputs(4333) <= a xor b;
    outputs(4334) <= not b;
    outputs(4335) <= not (a xor b);
    outputs(4336) <= not b;
    outputs(4337) <= not (a and b);
    outputs(4338) <= not b;
    outputs(4339) <= not (a xor b);
    outputs(4340) <= a xor b;
    outputs(4341) <= not b or a;
    outputs(4342) <= a and not b;
    outputs(4343) <= not a;
    outputs(4344) <= not (a or b);
    outputs(4345) <= not a or b;
    outputs(4346) <= not (a xor b);
    outputs(4347) <= a;
    outputs(4348) <= b;
    outputs(4349) <= b;
    outputs(4350) <= not a;
    outputs(4351) <= a xor b;
    outputs(4352) <= not a or b;
    outputs(4353) <= a;
    outputs(4354) <= a;
    outputs(4355) <= not (a xor b);
    outputs(4356) <= not (a xor b);
    outputs(4357) <= b;
    outputs(4358) <= b;
    outputs(4359) <= not (a xor b);
    outputs(4360) <= a;
    outputs(4361) <= a xor b;
    outputs(4362) <= not a;
    outputs(4363) <= a and b;
    outputs(4364) <= a or b;
    outputs(4365) <= a xor b;
    outputs(4366) <= b and not a;
    outputs(4367) <= a xor b;
    outputs(4368) <= a or b;
    outputs(4369) <= a xor b;
    outputs(4370) <= a xor b;
    outputs(4371) <= a and not b;
    outputs(4372) <= a xor b;
    outputs(4373) <= a and b;
    outputs(4374) <= not a;
    outputs(4375) <= a or b;
    outputs(4376) <= a xor b;
    outputs(4377) <= a;
    outputs(4378) <= a xor b;
    outputs(4379) <= a and b;
    outputs(4380) <= not (a xor b);
    outputs(4381) <= a;
    outputs(4382) <= b and not a;
    outputs(4383) <= a;
    outputs(4384) <= b;
    outputs(4385) <= not (a xor b);
    outputs(4386) <= not (a xor b);
    outputs(4387) <= b and not a;
    outputs(4388) <= b;
    outputs(4389) <= a and b;
    outputs(4390) <= a;
    outputs(4391) <= a and not b;
    outputs(4392) <= a xor b;
    outputs(4393) <= not b;
    outputs(4394) <= not a;
    outputs(4395) <= 1'b0;
    outputs(4396) <= b;
    outputs(4397) <= not b;
    outputs(4398) <= a;
    outputs(4399) <= not a;
    outputs(4400) <= a xor b;
    outputs(4401) <= not (a xor b);
    outputs(4402) <= not (a xor b);
    outputs(4403) <= not (a or b);
    outputs(4404) <= b;
    outputs(4405) <= not a;
    outputs(4406) <= b;
    outputs(4407) <= not (a xor b);
    outputs(4408) <= not (a or b);
    outputs(4409) <= b;
    outputs(4410) <= not (a or b);
    outputs(4411) <= a;
    outputs(4412) <= a xor b;
    outputs(4413) <= a;
    outputs(4414) <= not a;
    outputs(4415) <= a and not b;
    outputs(4416) <= not a;
    outputs(4417) <= a xor b;
    outputs(4418) <= a and b;
    outputs(4419) <= not b;
    outputs(4420) <= a xor b;
    outputs(4421) <= b;
    outputs(4422) <= not b;
    outputs(4423) <= a xor b;
    outputs(4424) <= not (a or b);
    outputs(4425) <= not (a xor b);
    outputs(4426) <= b;
    outputs(4427) <= b;
    outputs(4428) <= not a;
    outputs(4429) <= a xor b;
    outputs(4430) <= not a;
    outputs(4431) <= a and b;
    outputs(4432) <= b and not a;
    outputs(4433) <= not a;
    outputs(4434) <= a and not b;
    outputs(4435) <= not (a xor b);
    outputs(4436) <= a xor b;
    outputs(4437) <= not a;
    outputs(4438) <= a and not b;
    outputs(4439) <= not a or b;
    outputs(4440) <= b and not a;
    outputs(4441) <= not b;
    outputs(4442) <= a and not b;
    outputs(4443) <= a;
    outputs(4444) <= not a or b;
    outputs(4445) <= b;
    outputs(4446) <= b and not a;
    outputs(4447) <= not a;
    outputs(4448) <= not (a xor b);
    outputs(4449) <= not b;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= a and b;
    outputs(4452) <= not b;
    outputs(4453) <= a;
    outputs(4454) <= a or b;
    outputs(4455) <= not b;
    outputs(4456) <= b;
    outputs(4457) <= a xor b;
    outputs(4458) <= not a or b;
    outputs(4459) <= not b;
    outputs(4460) <= a;
    outputs(4461) <= not a;
    outputs(4462) <= not (a xor b);
    outputs(4463) <= a;
    outputs(4464) <= b;
    outputs(4465) <= not (a xor b);
    outputs(4466) <= a xor b;
    outputs(4467) <= b;
    outputs(4468) <= a xor b;
    outputs(4469) <= a;
    outputs(4470) <= a and not b;
    outputs(4471) <= a;
    outputs(4472) <= not a;
    outputs(4473) <= a and b;
    outputs(4474) <= a;
    outputs(4475) <= not a;
    outputs(4476) <= b;
    outputs(4477) <= b and not a;
    outputs(4478) <= not b;
    outputs(4479) <= not a;
    outputs(4480) <= not b;
    outputs(4481) <= not b;
    outputs(4482) <= a or b;
    outputs(4483) <= b;
    outputs(4484) <= a;
    outputs(4485) <= not a or b;
    outputs(4486) <= not b;
    outputs(4487) <= not a or b;
    outputs(4488) <= a and not b;
    outputs(4489) <= not a;
    outputs(4490) <= not (a xor b);
    outputs(4491) <= b;
    outputs(4492) <= not (a or b);
    outputs(4493) <= a xor b;
    outputs(4494) <= not (a xor b);
    outputs(4495) <= a and not b;
    outputs(4496) <= not (a or b);
    outputs(4497) <= not (a or b);
    outputs(4498) <= not a;
    outputs(4499) <= not (a or b);
    outputs(4500) <= not (a xor b);
    outputs(4501) <= not a;
    outputs(4502) <= not (a xor b);
    outputs(4503) <= not (a or b);
    outputs(4504) <= a and not b;
    outputs(4505) <= not (a xor b);
    outputs(4506) <= not a;
    outputs(4507) <= not (a and b);
    outputs(4508) <= b;
    outputs(4509) <= not a;
    outputs(4510) <= not (a xor b);
    outputs(4511) <= a xor b;
    outputs(4512) <= a and not b;
    outputs(4513) <= 1'b0;
    outputs(4514) <= b;
    outputs(4515) <= a xor b;
    outputs(4516) <= b;
    outputs(4517) <= not (a xor b);
    outputs(4518) <= a xor b;
    outputs(4519) <= a xor b;
    outputs(4520) <= not b;
    outputs(4521) <= not (a xor b);
    outputs(4522) <= not (a or b);
    outputs(4523) <= a;
    outputs(4524) <= not (a xor b);
    outputs(4525) <= a xor b;
    outputs(4526) <= a;
    outputs(4527) <= not a;
    outputs(4528) <= a;
    outputs(4529) <= a;
    outputs(4530) <= a xor b;
    outputs(4531) <= a and b;
    outputs(4532) <= not a;
    outputs(4533) <= not (a xor b);
    outputs(4534) <= a and b;
    outputs(4535) <= not (a or b);
    outputs(4536) <= a;
    outputs(4537) <= not (a xor b);
    outputs(4538) <= not (a or b);
    outputs(4539) <= a or b;
    outputs(4540) <= a or b;
    outputs(4541) <= a and not b;
    outputs(4542) <= a;
    outputs(4543) <= not (a xor b);
    outputs(4544) <= not (a and b);
    outputs(4545) <= not a;
    outputs(4546) <= not (a xor b);
    outputs(4547) <= not b;
    outputs(4548) <= not (a xor b);
    outputs(4549) <= a;
    outputs(4550) <= not (a or b);
    outputs(4551) <= b;
    outputs(4552) <= not (a xor b);
    outputs(4553) <= a xor b;
    outputs(4554) <= not a or b;
    outputs(4555) <= a;
    outputs(4556) <= b;
    outputs(4557) <= not b;
    outputs(4558) <= b;
    outputs(4559) <= not (a xor b);
    outputs(4560) <= not (a or b);
    outputs(4561) <= b;
    outputs(4562) <= b;
    outputs(4563) <= not a;
    outputs(4564) <= not (a xor b);
    outputs(4565) <= not a;
    outputs(4566) <= not (a xor b);
    outputs(4567) <= b;
    outputs(4568) <= a xor b;
    outputs(4569) <= a and not b;
    outputs(4570) <= not (a or b);
    outputs(4571) <= b;
    outputs(4572) <= not a or b;
    outputs(4573) <= b;
    outputs(4574) <= not a or b;
    outputs(4575) <= not (a xor b);
    outputs(4576) <= b;
    outputs(4577) <= a;
    outputs(4578) <= a xor b;
    outputs(4579) <= not (a xor b);
    outputs(4580) <= b;
    outputs(4581) <= not (a xor b);
    outputs(4582) <= not a;
    outputs(4583) <= not a;
    outputs(4584) <= a xor b;
    outputs(4585) <= b and not a;
    outputs(4586) <= b;
    outputs(4587) <= not a;
    outputs(4588) <= b;
    outputs(4589) <= not a;
    outputs(4590) <= not b;
    outputs(4591) <= a;
    outputs(4592) <= not a;
    outputs(4593) <= not (a or b);
    outputs(4594) <= a and b;
    outputs(4595) <= a;
    outputs(4596) <= a xor b;
    outputs(4597) <= not (a xor b);
    outputs(4598) <= not (a xor b);
    outputs(4599) <= not (a or b);
    outputs(4600) <= a and not b;
    outputs(4601) <= a;
    outputs(4602) <= b;
    outputs(4603) <= a;
    outputs(4604) <= a;
    outputs(4605) <= not a;
    outputs(4606) <= a or b;
    outputs(4607) <= not (a xor b);
    outputs(4608) <= not (a xor b);
    outputs(4609) <= b;
    outputs(4610) <= a;
    outputs(4611) <= not b;
    outputs(4612) <= a;
    outputs(4613) <= b;
    outputs(4614) <= a and b;
    outputs(4615) <= b;
    outputs(4616) <= not (a xor b);
    outputs(4617) <= not (a xor b);
    outputs(4618) <= a and not b;
    outputs(4619) <= not a;
    outputs(4620) <= not (a xor b);
    outputs(4621) <= not a;
    outputs(4622) <= not (a xor b);
    outputs(4623) <= a;
    outputs(4624) <= a xor b;
    outputs(4625) <= not a;
    outputs(4626) <= not b;
    outputs(4627) <= b;
    outputs(4628) <= not b;
    outputs(4629) <= b;
    outputs(4630) <= not a;
    outputs(4631) <= b;
    outputs(4632) <= b;
    outputs(4633) <= not a;
    outputs(4634) <= not (a or b);
    outputs(4635) <= a;
    outputs(4636) <= not (a xor b);
    outputs(4637) <= not a;
    outputs(4638) <= not (a xor b);
    outputs(4639) <= not (a or b);
    outputs(4640) <= not (a xor b);
    outputs(4641) <= b and not a;
    outputs(4642) <= not a;
    outputs(4643) <= not (a xor b);
    outputs(4644) <= a xor b;
    outputs(4645) <= b and not a;
    outputs(4646) <= a;
    outputs(4647) <= a xor b;
    outputs(4648) <= not b;
    outputs(4649) <= b;
    outputs(4650) <= not b;
    outputs(4651) <= not a;
    outputs(4652) <= a;
    outputs(4653) <= not (a xor b);
    outputs(4654) <= a xor b;
    outputs(4655) <= not (a xor b);
    outputs(4656) <= not b;
    outputs(4657) <= a;
    outputs(4658) <= not b;
    outputs(4659) <= not b;
    outputs(4660) <= not (a xor b);
    outputs(4661) <= not (a xor b);
    outputs(4662) <= a xor b;
    outputs(4663) <= a;
    outputs(4664) <= not b;
    outputs(4665) <= a and not b;
    outputs(4666) <= a and not b;
    outputs(4667) <= b;
    outputs(4668) <= a xor b;
    outputs(4669) <= not b;
    outputs(4670) <= a and not b;
    outputs(4671) <= a;
    outputs(4672) <= not (a xor b);
    outputs(4673) <= not b;
    outputs(4674) <= not b;
    outputs(4675) <= a and not b;
    outputs(4676) <= not (a or b);
    outputs(4677) <= not a;
    outputs(4678) <= a;
    outputs(4679) <= a xor b;
    outputs(4680) <= b;
    outputs(4681) <= not (a xor b);
    outputs(4682) <= b;
    outputs(4683) <= not (a xor b);
    outputs(4684) <= not b;
    outputs(4685) <= not (a xor b);
    outputs(4686) <= not (a xor b);
    outputs(4687) <= not (a xor b);
    outputs(4688) <= a xor b;
    outputs(4689) <= a or b;
    outputs(4690) <= a xor b;
    outputs(4691) <= not a;
    outputs(4692) <= b;
    outputs(4693) <= a xor b;
    outputs(4694) <= not a;
    outputs(4695) <= a;
    outputs(4696) <= a and b;
    outputs(4697) <= b and not a;
    outputs(4698) <= not a;
    outputs(4699) <= a;
    outputs(4700) <= b;
    outputs(4701) <= not a;
    outputs(4702) <= a;
    outputs(4703) <= b and not a;
    outputs(4704) <= a;
    outputs(4705) <= not b;
    outputs(4706) <= a xor b;
    outputs(4707) <= not (a or b);
    outputs(4708) <= not b;
    outputs(4709) <= not (a xor b);
    outputs(4710) <= not (a xor b);
    outputs(4711) <= a and b;
    outputs(4712) <= not b;
    outputs(4713) <= a xor b;
    outputs(4714) <= not (a xor b);
    outputs(4715) <= not a;
    outputs(4716) <= a xor b;
    outputs(4717) <= b and not a;
    outputs(4718) <= not (a or b);
    outputs(4719) <= a;
    outputs(4720) <= not (a or b);
    outputs(4721) <= not b;
    outputs(4722) <= not (a xor b);
    outputs(4723) <= a;
    outputs(4724) <= not (a xor b);
    outputs(4725) <= not b or a;
    outputs(4726) <= not (a xor b);
    outputs(4727) <= a;
    outputs(4728) <= a and not b;
    outputs(4729) <= a xor b;
    outputs(4730) <= not (a xor b);
    outputs(4731) <= a and not b;
    outputs(4732) <= not b;
    outputs(4733) <= not b or a;
    outputs(4734) <= a;
    outputs(4735) <= b;
    outputs(4736) <= not b or a;
    outputs(4737) <= not b;
    outputs(4738) <= a xor b;
    outputs(4739) <= a and not b;
    outputs(4740) <= b and not a;
    outputs(4741) <= not b or a;
    outputs(4742) <= b;
    outputs(4743) <= not a;
    outputs(4744) <= not b;
    outputs(4745) <= a;
    outputs(4746) <= a;
    outputs(4747) <= not b;
    outputs(4748) <= b;
    outputs(4749) <= a xor b;
    outputs(4750) <= b and not a;
    outputs(4751) <= b;
    outputs(4752) <= a;
    outputs(4753) <= b;
    outputs(4754) <= a xor b;
    outputs(4755) <= a xor b;
    outputs(4756) <= a;
    outputs(4757) <= not (a xor b);
    outputs(4758) <= a xor b;
    outputs(4759) <= not (a xor b);
    outputs(4760) <= not b;
    outputs(4761) <= not a;
    outputs(4762) <= not a;
    outputs(4763) <= not (a xor b);
    outputs(4764) <= not (a xor b);
    outputs(4765) <= not a;
    outputs(4766) <= a xor b;
    outputs(4767) <= b and not a;
    outputs(4768) <= a and b;
    outputs(4769) <= a;
    outputs(4770) <= b;
    outputs(4771) <= not (a xor b);
    outputs(4772) <= a and not b;
    outputs(4773) <= not (a and b);
    outputs(4774) <= not (a or b);
    outputs(4775) <= b;
    outputs(4776) <= a and b;
    outputs(4777) <= a xor b;
    outputs(4778) <= a xor b;
    outputs(4779) <= not a;
    outputs(4780) <= a xor b;
    outputs(4781) <= not (a or b);
    outputs(4782) <= not (a or b);
    outputs(4783) <= not (a xor b);
    outputs(4784) <= a xor b;
    outputs(4785) <= b and not a;
    outputs(4786) <= a;
    outputs(4787) <= not b or a;
    outputs(4788) <= b;
    outputs(4789) <= not (a xor b);
    outputs(4790) <= b;
    outputs(4791) <= not b;
    outputs(4792) <= a;
    outputs(4793) <= b and not a;
    outputs(4794) <= not (a xor b);
    outputs(4795) <= not b;
    outputs(4796) <= not a;
    outputs(4797) <= not (a xor b);
    outputs(4798) <= not a or b;
    outputs(4799) <= not (a or b);
    outputs(4800) <= a and b;
    outputs(4801) <= not a or b;
    outputs(4802) <= a;
    outputs(4803) <= b;
    outputs(4804) <= not a;
    outputs(4805) <= b;
    outputs(4806) <= not b;
    outputs(4807) <= not a;
    outputs(4808) <= not (a xor b);
    outputs(4809) <= a xor b;
    outputs(4810) <= a;
    outputs(4811) <= not a or b;
    outputs(4812) <= a and not b;
    outputs(4813) <= a;
    outputs(4814) <= not (a or b);
    outputs(4815) <= not a;
    outputs(4816) <= b;
    outputs(4817) <= not b;
    outputs(4818) <= not (a xor b);
    outputs(4819) <= a xor b;
    outputs(4820) <= a;
    outputs(4821) <= not (a xor b);
    outputs(4822) <= b;
    outputs(4823) <= not (a xor b);
    outputs(4824) <= b and not a;
    outputs(4825) <= b;
    outputs(4826) <= a;
    outputs(4827) <= a xor b;
    outputs(4828) <= not (a xor b);
    outputs(4829) <= b;
    outputs(4830) <= a and b;
    outputs(4831) <= not b;
    outputs(4832) <= a;
    outputs(4833) <= not a;
    outputs(4834) <= not (a or b);
    outputs(4835) <= not a;
    outputs(4836) <= not b;
    outputs(4837) <= not b;
    outputs(4838) <= not (a and b);
    outputs(4839) <= a and b;
    outputs(4840) <= a;
    outputs(4841) <= not b or a;
    outputs(4842) <= a xor b;
    outputs(4843) <= not a;
    outputs(4844) <= a;
    outputs(4845) <= not a;
    outputs(4846) <= not a;
    outputs(4847) <= not b;
    outputs(4848) <= not (a xor b);
    outputs(4849) <= not (a or b);
    outputs(4850) <= not (a xor b);
    outputs(4851) <= not b;
    outputs(4852) <= not a;
    outputs(4853) <= not (a or b);
    outputs(4854) <= not (a xor b);
    outputs(4855) <= not (a and b);
    outputs(4856) <= not (a and b);
    outputs(4857) <= a;
    outputs(4858) <= 1'b1;
    outputs(4859) <= a xor b;
    outputs(4860) <= b;
    outputs(4861) <= not (a or b);
    outputs(4862) <= b;
    outputs(4863) <= not b;
    outputs(4864) <= b;
    outputs(4865) <= not b;
    outputs(4866) <= a and b;
    outputs(4867) <= not (a and b);
    outputs(4868) <= not (a or b);
    outputs(4869) <= a xor b;
    outputs(4870) <= not a;
    outputs(4871) <= a;
    outputs(4872) <= a;
    outputs(4873) <= b and not a;
    outputs(4874) <= a and not b;
    outputs(4875) <= a and not b;
    outputs(4876) <= b;
    outputs(4877) <= not a;
    outputs(4878) <= a xor b;
    outputs(4879) <= b;
    outputs(4880) <= b;
    outputs(4881) <= not b;
    outputs(4882) <= not (a and b);
    outputs(4883) <= b and not a;
    outputs(4884) <= a xor b;
    outputs(4885) <= not (a xor b);
    outputs(4886) <= a xor b;
    outputs(4887) <= not (a xor b);
    outputs(4888) <= not (a and b);
    outputs(4889) <= not a or b;
    outputs(4890) <= not (a xor b);
    outputs(4891) <= not a;
    outputs(4892) <= a xor b;
    outputs(4893) <= not a;
    outputs(4894) <= a and b;
    outputs(4895) <= b;
    outputs(4896) <= b and not a;
    outputs(4897) <= a xor b;
    outputs(4898) <= a xor b;
    outputs(4899) <= b;
    outputs(4900) <= not a;
    outputs(4901) <= not a;
    outputs(4902) <= not (a xor b);
    outputs(4903) <= b;
    outputs(4904) <= a;
    outputs(4905) <= b and not a;
    outputs(4906) <= not (a xor b);
    outputs(4907) <= a;
    outputs(4908) <= a xor b;
    outputs(4909) <= not b or a;
    outputs(4910) <= a;
    outputs(4911) <= a and b;
    outputs(4912) <= b and not a;
    outputs(4913) <= a xor b;
    outputs(4914) <= not a;
    outputs(4915) <= not (a xor b);
    outputs(4916) <= not b;
    outputs(4917) <= not (a xor b);
    outputs(4918) <= a;
    outputs(4919) <= b;
    outputs(4920) <= not (a xor b);
    outputs(4921) <= a;
    outputs(4922) <= not a;
    outputs(4923) <= b;
    outputs(4924) <= a and not b;
    outputs(4925) <= a xor b;
    outputs(4926) <= a;
    outputs(4927) <= not (a xor b);
    outputs(4928) <= b and not a;
    outputs(4929) <= a xor b;
    outputs(4930) <= a and b;
    outputs(4931) <= a;
    outputs(4932) <= a and not b;
    outputs(4933) <= a and not b;
    outputs(4934) <= b and not a;
    outputs(4935) <= b;
    outputs(4936) <= not b;
    outputs(4937) <= b;
    outputs(4938) <= a and not b;
    outputs(4939) <= not b;
    outputs(4940) <= not a;
    outputs(4941) <= b;
    outputs(4942) <= a;
    outputs(4943) <= a and b;
    outputs(4944) <= a;
    outputs(4945) <= b;
    outputs(4946) <= a and not b;
    outputs(4947) <= a xor b;
    outputs(4948) <= not (a xor b);
    outputs(4949) <= not (a or b);
    outputs(4950) <= b;
    outputs(4951) <= b and not a;
    outputs(4952) <= b;
    outputs(4953) <= a;
    outputs(4954) <= a and b;
    outputs(4955) <= a;
    outputs(4956) <= a xor b;
    outputs(4957) <= a and not b;
    outputs(4958) <= a and not b;
    outputs(4959) <= a xor b;
    outputs(4960) <= not a;
    outputs(4961) <= not b;
    outputs(4962) <= b;
    outputs(4963) <= a and b;
    outputs(4964) <= a;
    outputs(4965) <= a and b;
    outputs(4966) <= a and b;
    outputs(4967) <= not (a xor b);
    outputs(4968) <= a and not b;
    outputs(4969) <= not a;
    outputs(4970) <= a and not b;
    outputs(4971) <= a;
    outputs(4972) <= not (a xor b);
    outputs(4973) <= not a;
    outputs(4974) <= b and not a;
    outputs(4975) <= not (a or b);
    outputs(4976) <= b;
    outputs(4977) <= not (a xor b);
    outputs(4978) <= b;
    outputs(4979) <= a;
    outputs(4980) <= a xor b;
    outputs(4981) <= b;
    outputs(4982) <= not (a xor b);
    outputs(4983) <= not b;
    outputs(4984) <= not (a or b);
    outputs(4985) <= not (a xor b);
    outputs(4986) <= a;
    outputs(4987) <= not (a and b);
    outputs(4988) <= not a;
    outputs(4989) <= not a;
    outputs(4990) <= b and not a;
    outputs(4991) <= not b;
    outputs(4992) <= b and not a;
    outputs(4993) <= a;
    outputs(4994) <= not a;
    outputs(4995) <= not (a xor b);
    outputs(4996) <= a xor b;
    outputs(4997) <= not b;
    outputs(4998) <= a xor b;
    outputs(4999) <= not (a xor b);
    outputs(5000) <= not b;
    outputs(5001) <= not (a xor b);
    outputs(5002) <= not b;
    outputs(5003) <= b;
    outputs(5004) <= b;
    outputs(5005) <= a xor b;
    outputs(5006) <= a xor b;
    outputs(5007) <= not b;
    outputs(5008) <= not b;
    outputs(5009) <= b and not a;
    outputs(5010) <= a xor b;
    outputs(5011) <= a and b;
    outputs(5012) <= b;
    outputs(5013) <= a xor b;
    outputs(5014) <= b;
    outputs(5015) <= not b;
    outputs(5016) <= a xor b;
    outputs(5017) <= a xor b;
    outputs(5018) <= not b or a;
    outputs(5019) <= a or b;
    outputs(5020) <= a;
    outputs(5021) <= not (a xor b);
    outputs(5022) <= b;
    outputs(5023) <= not b;
    outputs(5024) <= not b;
    outputs(5025) <= not b;
    outputs(5026) <= b;
    outputs(5027) <= a;
    outputs(5028) <= a and b;
    outputs(5029) <= a xor b;
    outputs(5030) <= a xor b;
    outputs(5031) <= a and b;
    outputs(5032) <= not b;
    outputs(5033) <= not (a xor b);
    outputs(5034) <= not (a xor b);
    outputs(5035) <= a;
    outputs(5036) <= not (a xor b);
    outputs(5037) <= a xor b;
    outputs(5038) <= a xor b;
    outputs(5039) <= a and not b;
    outputs(5040) <= a xor b;
    outputs(5041) <= b;
    outputs(5042) <= a;
    outputs(5043) <= not (a xor b);
    outputs(5044) <= b;
    outputs(5045) <= not a;
    outputs(5046) <= a xor b;
    outputs(5047) <= not (a or b);
    outputs(5048) <= not (a xor b);
    outputs(5049) <= a;
    outputs(5050) <= b;
    outputs(5051) <= a xor b;
    outputs(5052) <= a and b;
    outputs(5053) <= b and not a;
    outputs(5054) <= not (a or b);
    outputs(5055) <= a xor b;
    outputs(5056) <= not b;
    outputs(5057) <= not b;
    outputs(5058) <= not a;
    outputs(5059) <= not (a xor b);
    outputs(5060) <= a and b;
    outputs(5061) <= a;
    outputs(5062) <= not b;
    outputs(5063) <= a and b;
    outputs(5064) <= b and not a;
    outputs(5065) <= a;
    outputs(5066) <= a;
    outputs(5067) <= not b;
    outputs(5068) <= not (a or b);
    outputs(5069) <= a xor b;
    outputs(5070) <= b;
    outputs(5071) <= not (a xor b);
    outputs(5072) <= a and not b;
    outputs(5073) <= a xor b;
    outputs(5074) <= not (a xor b);
    outputs(5075) <= not (a xor b);
    outputs(5076) <= a and b;
    outputs(5077) <= a or b;
    outputs(5078) <= a or b;
    outputs(5079) <= a xor b;
    outputs(5080) <= not b;
    outputs(5081) <= not (a xor b);
    outputs(5082) <= b;
    outputs(5083) <= not b;
    outputs(5084) <= not b or a;
    outputs(5085) <= b;
    outputs(5086) <= a and not b;
    outputs(5087) <= b;
    outputs(5088) <= not a;
    outputs(5089) <= a;
    outputs(5090) <= a xor b;
    outputs(5091) <= b and not a;
    outputs(5092) <= not (a or b);
    outputs(5093) <= not b or a;
    outputs(5094) <= not (a xor b);
    outputs(5095) <= b;
    outputs(5096) <= a and not b;
    outputs(5097) <= b;
    outputs(5098) <= not b;
    outputs(5099) <= b and not a;
    outputs(5100) <= b;
    outputs(5101) <= a;
    outputs(5102) <= not (a xor b);
    outputs(5103) <= not a or b;
    outputs(5104) <= a and not b;
    outputs(5105) <= a xor b;
    outputs(5106) <= not (a xor b);
    outputs(5107) <= not b;
    outputs(5108) <= a and not b;
    outputs(5109) <= b and not a;
    outputs(5110) <= not a;
    outputs(5111) <= a xor b;
    outputs(5112) <= not a;
    outputs(5113) <= a xor b;
    outputs(5114) <= a;
    outputs(5115) <= b;
    outputs(5116) <= a xor b;
    outputs(5117) <= not a;
    outputs(5118) <= a and b;
    outputs(5119) <= not b;
    outputs(5120) <= a;
    outputs(5121) <= not a;
    outputs(5122) <= a xor b;
    outputs(5123) <= b and not a;
    outputs(5124) <= not a;
    outputs(5125) <= not (a xor b);
    outputs(5126) <= not b;
    outputs(5127) <= not b;
    outputs(5128) <= not a;
    outputs(5129) <= not (a xor b);
    outputs(5130) <= not (a xor b);
    outputs(5131) <= not (a xor b);
    outputs(5132) <= a;
    outputs(5133) <= a and not b;
    outputs(5134) <= not b;
    outputs(5135) <= a xor b;
    outputs(5136) <= not b or a;
    outputs(5137) <= not (a xor b);
    outputs(5138) <= a and b;
    outputs(5139) <= not b;
    outputs(5140) <= a;
    outputs(5141) <= not a;
    outputs(5142) <= not b;
    outputs(5143) <= a xor b;
    outputs(5144) <= not (a or b);
    outputs(5145) <= not a;
    outputs(5146) <= a xor b;
    outputs(5147) <= not a or b;
    outputs(5148) <= not (a xor b);
    outputs(5149) <= b;
    outputs(5150) <= b;
    outputs(5151) <= not a;
    outputs(5152) <= a xor b;
    outputs(5153) <= a;
    outputs(5154) <= not (a xor b);
    outputs(5155) <= a and b;
    outputs(5156) <= a and not b;
    outputs(5157) <= a and not b;
    outputs(5158) <= not (a xor b);
    outputs(5159) <= b;
    outputs(5160) <= a;
    outputs(5161) <= a xor b;
    outputs(5162) <= a xor b;
    outputs(5163) <= not b or a;
    outputs(5164) <= a xor b;
    outputs(5165) <= b and not a;
    outputs(5166) <= a xor b;
    outputs(5167) <= a;
    outputs(5168) <= not b;
    outputs(5169) <= not a;
    outputs(5170) <= not (a xor b);
    outputs(5171) <= a and b;
    outputs(5172) <= not (a and b);
    outputs(5173) <= a xor b;
    outputs(5174) <= a;
    outputs(5175) <= b;
    outputs(5176) <= a xor b;
    outputs(5177) <= b;
    outputs(5178) <= not b or a;
    outputs(5179) <= not (a and b);
    outputs(5180) <= not (a xor b);
    outputs(5181) <= not a;
    outputs(5182) <= b;
    outputs(5183) <= b;
    outputs(5184) <= not (a xor b);
    outputs(5185) <= not a;
    outputs(5186) <= not b;
    outputs(5187) <= not a;
    outputs(5188) <= a;
    outputs(5189) <= a xor b;
    outputs(5190) <= not b or a;
    outputs(5191) <= a xor b;
    outputs(5192) <= a and not b;
    outputs(5193) <= b;
    outputs(5194) <= b;
    outputs(5195) <= a xor b;
    outputs(5196) <= b and not a;
    outputs(5197) <= b;
    outputs(5198) <= b;
    outputs(5199) <= not a or b;
    outputs(5200) <= not (a xor b);
    outputs(5201) <= b and not a;
    outputs(5202) <= a xor b;
    outputs(5203) <= not a;
    outputs(5204) <= not b;
    outputs(5205) <= b and not a;
    outputs(5206) <= a;
    outputs(5207) <= a xor b;
    outputs(5208) <= a and not b;
    outputs(5209) <= not (a xor b);
    outputs(5210) <= not a;
    outputs(5211) <= not (a and b);
    outputs(5212) <= b;
    outputs(5213) <= b and not a;
    outputs(5214) <= not (a and b);
    outputs(5215) <= not a;
    outputs(5216) <= not b;
    outputs(5217) <= a xor b;
    outputs(5218) <= not a or b;
    outputs(5219) <= not (a xor b);
    outputs(5220) <= b;
    outputs(5221) <= a xor b;
    outputs(5222) <= not a;
    outputs(5223) <= not (a or b);
    outputs(5224) <= not b;
    outputs(5225) <= not b or a;
    outputs(5226) <= not a;
    outputs(5227) <= b;
    outputs(5228) <= not a;
    outputs(5229) <= not b;
    outputs(5230) <= not (a xor b);
    outputs(5231) <= a xor b;
    outputs(5232) <= not b or a;
    outputs(5233) <= not (a xor b);
    outputs(5234) <= not b;
    outputs(5235) <= not b;
    outputs(5236) <= not b or a;
    outputs(5237) <= b;
    outputs(5238) <= b;
    outputs(5239) <= a and not b;
    outputs(5240) <= not a;
    outputs(5241) <= not a or b;
    outputs(5242) <= b;
    outputs(5243) <= b;
    outputs(5244) <= not a;
    outputs(5245) <= a xor b;
    outputs(5246) <= a xor b;
    outputs(5247) <= a;
    outputs(5248) <= b;
    outputs(5249) <= b;
    outputs(5250) <= a xor b;
    outputs(5251) <= a;
    outputs(5252) <= not b;
    outputs(5253) <= a xor b;
    outputs(5254) <= b;
    outputs(5255) <= a xor b;
    outputs(5256) <= b;
    outputs(5257) <= not b or a;
    outputs(5258) <= not a;
    outputs(5259) <= not (a xor b);
    outputs(5260) <= not (a or b);
    outputs(5261) <= a;
    outputs(5262) <= b;
    outputs(5263) <= a xor b;
    outputs(5264) <= not (a xor b);
    outputs(5265) <= a xor b;
    outputs(5266) <= a or b;
    outputs(5267) <= b;
    outputs(5268) <= a xor b;
    outputs(5269) <= a xor b;
    outputs(5270) <= a and not b;
    outputs(5271) <= a and b;
    outputs(5272) <= a xor b;
    outputs(5273) <= b;
    outputs(5274) <= not b or a;
    outputs(5275) <= not b or a;
    outputs(5276) <= not a;
    outputs(5277) <= a xor b;
    outputs(5278) <= a xor b;
    outputs(5279) <= not a or b;
    outputs(5280) <= a;
    outputs(5281) <= not b;
    outputs(5282) <= a and not b;
    outputs(5283) <= not (a xor b);
    outputs(5284) <= a and not b;
    outputs(5285) <= b and not a;
    outputs(5286) <= not (a and b);
    outputs(5287) <= not (a xor b);
    outputs(5288) <= a xor b;
    outputs(5289) <= not a;
    outputs(5290) <= b and not a;
    outputs(5291) <= not b or a;
    outputs(5292) <= not a;
    outputs(5293) <= a xor b;
    outputs(5294) <= not b;
    outputs(5295) <= not (a xor b);
    outputs(5296) <= not a or b;
    outputs(5297) <= not a;
    outputs(5298) <= not (a xor b);
    outputs(5299) <= not (a xor b);
    outputs(5300) <= b;
    outputs(5301) <= a xor b;
    outputs(5302) <= not (a xor b);
    outputs(5303) <= a;
    outputs(5304) <= not b or a;
    outputs(5305) <= a xor b;
    outputs(5306) <= not (a or b);
    outputs(5307) <= a or b;
    outputs(5308) <= a xor b;
    outputs(5309) <= not a or b;
    outputs(5310) <= a xor b;
    outputs(5311) <= a xor b;
    outputs(5312) <= not b or a;
    outputs(5313) <= a xor b;
    outputs(5314) <= not (a xor b);
    outputs(5315) <= a xor b;
    outputs(5316) <= not b or a;
    outputs(5317) <= not a;
    outputs(5318) <= not (a xor b);
    outputs(5319) <= not a;
    outputs(5320) <= a and b;
    outputs(5321) <= b;
    outputs(5322) <= a;
    outputs(5323) <= a;
    outputs(5324) <= not a;
    outputs(5325) <= not (a xor b);
    outputs(5326) <= a xor b;
    outputs(5327) <= b;
    outputs(5328) <= a xor b;
    outputs(5329) <= a xor b;
    outputs(5330) <= b;
    outputs(5331) <= b;
    outputs(5332) <= not (a xor b);
    outputs(5333) <= not (a xor b);
    outputs(5334) <= a and not b;
    outputs(5335) <= not (a xor b);
    outputs(5336) <= a xor b;
    outputs(5337) <= not b;
    outputs(5338) <= not (a xor b);
    outputs(5339) <= a xor b;
    outputs(5340) <= a or b;
    outputs(5341) <= b;
    outputs(5342) <= a xor b;
    outputs(5343) <= not a or b;
    outputs(5344) <= not b;
    outputs(5345) <= b and not a;
    outputs(5346) <= not b or a;
    outputs(5347) <= not a;
    outputs(5348) <= a xor b;
    outputs(5349) <= not (a xor b);
    outputs(5350) <= a xor b;
    outputs(5351) <= a;
    outputs(5352) <= not (a xor b);
    outputs(5353) <= a;
    outputs(5354) <= not a;
    outputs(5355) <= not b;
    outputs(5356) <= b;
    outputs(5357) <= not a or b;
    outputs(5358) <= not a;
    outputs(5359) <= b;
    outputs(5360) <= a;
    outputs(5361) <= not b;
    outputs(5362) <= a;
    outputs(5363) <= not a;
    outputs(5364) <= a and not b;
    outputs(5365) <= b;
    outputs(5366) <= not a;
    outputs(5367) <= a;
    outputs(5368) <= not a or b;
    outputs(5369) <= not a;
    outputs(5370) <= b;
    outputs(5371) <= a;
    outputs(5372) <= b;
    outputs(5373) <= a;
    outputs(5374) <= a xor b;
    outputs(5375) <= b and not a;
    outputs(5376) <= a;
    outputs(5377) <= a xor b;
    outputs(5378) <= not a;
    outputs(5379) <= not (a xor b);
    outputs(5380) <= b;
    outputs(5381) <= b and not a;
    outputs(5382) <= not b;
    outputs(5383) <= b and not a;
    outputs(5384) <= a xor b;
    outputs(5385) <= not a;
    outputs(5386) <= b;
    outputs(5387) <= b;
    outputs(5388) <= not (a or b);
    outputs(5389) <= not b;
    outputs(5390) <= b and not a;
    outputs(5391) <= a;
    outputs(5392) <= not a;
    outputs(5393) <= not a;
    outputs(5394) <= a xor b;
    outputs(5395) <= not (a xor b);
    outputs(5396) <= a and not b;
    outputs(5397) <= a xor b;
    outputs(5398) <= not b;
    outputs(5399) <= b;
    outputs(5400) <= a xor b;
    outputs(5401) <= a xor b;
    outputs(5402) <= not a;
    outputs(5403) <= a xor b;
    outputs(5404) <= not b;
    outputs(5405) <= not b;
    outputs(5406) <= b;
    outputs(5407) <= a;
    outputs(5408) <= a;
    outputs(5409) <= not b;
    outputs(5410) <= a xor b;
    outputs(5411) <= a and b;
    outputs(5412) <= not (a xor b);
    outputs(5413) <= not (a xor b);
    outputs(5414) <= not a;
    outputs(5415) <= not (a xor b);
    outputs(5416) <= a and not b;
    outputs(5417) <= b;
    outputs(5418) <= not b;
    outputs(5419) <= b;
    outputs(5420) <= not (a xor b);
    outputs(5421) <= not a;
    outputs(5422) <= not a;
    outputs(5423) <= a xor b;
    outputs(5424) <= a and not b;
    outputs(5425) <= b;
    outputs(5426) <= not (a xor b);
    outputs(5427) <= a xor b;
    outputs(5428) <= not (a or b);
    outputs(5429) <= not b;
    outputs(5430) <= b;
    outputs(5431) <= not a or b;
    outputs(5432) <= a;
    outputs(5433) <= a and b;
    outputs(5434) <= a and b;
    outputs(5435) <= a;
    outputs(5436) <= not a or b;
    outputs(5437) <= b;
    outputs(5438) <= not (a xor b);
    outputs(5439) <= not b;
    outputs(5440) <= a xor b;
    outputs(5441) <= a;
    outputs(5442) <= not (a or b);
    outputs(5443) <= not (a or b);
    outputs(5444) <= a or b;
    outputs(5445) <= a;
    outputs(5446) <= a xor b;
    outputs(5447) <= not b or a;
    outputs(5448) <= not (a or b);
    outputs(5449) <= b;
    outputs(5450) <= a xor b;
    outputs(5451) <= not (a or b);
    outputs(5452) <= not a;
    outputs(5453) <= not b or a;
    outputs(5454) <= not (a and b);
    outputs(5455) <= not (a and b);
    outputs(5456) <= a or b;
    outputs(5457) <= not a;
    outputs(5458) <= a;
    outputs(5459) <= a xor b;
    outputs(5460) <= a xor b;
    outputs(5461) <= a xor b;
    outputs(5462) <= a xor b;
    outputs(5463) <= b;
    outputs(5464) <= not a;
    outputs(5465) <= b;
    outputs(5466) <= not (a xor b);
    outputs(5467) <= not (a and b);
    outputs(5468) <= a and b;
    outputs(5469) <= not b;
    outputs(5470) <= a xor b;
    outputs(5471) <= not (a xor b);
    outputs(5472) <= b;
    outputs(5473) <= not a or b;
    outputs(5474) <= a or b;
    outputs(5475) <= a;
    outputs(5476) <= not (a xor b);
    outputs(5477) <= not b;
    outputs(5478) <= b;
    outputs(5479) <= b;
    outputs(5480) <= a xor b;
    outputs(5481) <= not b;
    outputs(5482) <= not (a or b);
    outputs(5483) <= not a;
    outputs(5484) <= not (a xor b);
    outputs(5485) <= a xor b;
    outputs(5486) <= not b;
    outputs(5487) <= not (a or b);
    outputs(5488) <= not a;
    outputs(5489) <= not (a xor b);
    outputs(5490) <= a xor b;
    outputs(5491) <= b;
    outputs(5492) <= a;
    outputs(5493) <= a;
    outputs(5494) <= a;
    outputs(5495) <= not b;
    outputs(5496) <= a;
    outputs(5497) <= not b or a;
    outputs(5498) <= not (a and b);
    outputs(5499) <= b and not a;
    outputs(5500) <= not (a xor b);
    outputs(5501) <= not (a xor b);
    outputs(5502) <= a xor b;
    outputs(5503) <= b;
    outputs(5504) <= a xor b;
    outputs(5505) <= a xor b;
    outputs(5506) <= a xor b;
    outputs(5507) <= a xor b;
    outputs(5508) <= a xor b;
    outputs(5509) <= a xor b;
    outputs(5510) <= not a;
    outputs(5511) <= a and b;
    outputs(5512) <= a and not b;
    outputs(5513) <= a or b;
    outputs(5514) <= a;
    outputs(5515) <= a and not b;
    outputs(5516) <= not b;
    outputs(5517) <= a xor b;
    outputs(5518) <= a or b;
    outputs(5519) <= not (a xor b);
    outputs(5520) <= a xor b;
    outputs(5521) <= not (a xor b);
    outputs(5522) <= a or b;
    outputs(5523) <= b;
    outputs(5524) <= b;
    outputs(5525) <= a and not b;
    outputs(5526) <= not a;
    outputs(5527) <= b;
    outputs(5528) <= a or b;
    outputs(5529) <= not a or b;
    outputs(5530) <= not a;
    outputs(5531) <= a xor b;
    outputs(5532) <= b;
    outputs(5533) <= not b;
    outputs(5534) <= not (a xor b);
    outputs(5535) <= not b;
    outputs(5536) <= a xor b;
    outputs(5537) <= not b;
    outputs(5538) <= not (a xor b);
    outputs(5539) <= not (a xor b);
    outputs(5540) <= not (a xor b);
    outputs(5541) <= a or b;
    outputs(5542) <= not (a or b);
    outputs(5543) <= not b;
    outputs(5544) <= not b;
    outputs(5545) <= b;
    outputs(5546) <= a or b;
    outputs(5547) <= not a or b;
    outputs(5548) <= a xor b;
    outputs(5549) <= a xor b;
    outputs(5550) <= a and b;
    outputs(5551) <= not b or a;
    outputs(5552) <= a xor b;
    outputs(5553) <= a and not b;
    outputs(5554) <= a xor b;
    outputs(5555) <= not (a xor b);
    outputs(5556) <= b;
    outputs(5557) <= not (a xor b);
    outputs(5558) <= not a;
    outputs(5559) <= not a;
    outputs(5560) <= not (a xor b);
    outputs(5561) <= b;
    outputs(5562) <= not (a xor b);
    outputs(5563) <= not (a or b);
    outputs(5564) <= b;
    outputs(5565) <= not (a xor b);
    outputs(5566) <= not a;
    outputs(5567) <= a xor b;
    outputs(5568) <= a and not b;
    outputs(5569) <= not b or a;
    outputs(5570) <= not b;
    outputs(5571) <= b;
    outputs(5572) <= not b;
    outputs(5573) <= b;
    outputs(5574) <= not b;
    outputs(5575) <= not a;
    outputs(5576) <= not (a xor b);
    outputs(5577) <= not (a or b);
    outputs(5578) <= not a or b;
    outputs(5579) <= b;
    outputs(5580) <= not (a xor b);
    outputs(5581) <= a;
    outputs(5582) <= not (a xor b);
    outputs(5583) <= not b;
    outputs(5584) <= a xor b;
    outputs(5585) <= a xor b;
    outputs(5586) <= not a;
    outputs(5587) <= b and not a;
    outputs(5588) <= not (a or b);
    outputs(5589) <= not b;
    outputs(5590) <= not a;
    outputs(5591) <= not (a xor b);
    outputs(5592) <= not (a xor b);
    outputs(5593) <= not (a xor b);
    outputs(5594) <= not a or b;
    outputs(5595) <= not b;
    outputs(5596) <= not (a xor b);
    outputs(5597) <= b;
    outputs(5598) <= a and not b;
    outputs(5599) <= a xor b;
    outputs(5600) <= not b or a;
    outputs(5601) <= a or b;
    outputs(5602) <= not b;
    outputs(5603) <= not a;
    outputs(5604) <= b;
    outputs(5605) <= b;
    outputs(5606) <= not (a xor b);
    outputs(5607) <= a;
    outputs(5608) <= b;
    outputs(5609) <= not b;
    outputs(5610) <= not (a and b);
    outputs(5611) <= a xor b;
    outputs(5612) <= not (a xor b);
    outputs(5613) <= a xor b;
    outputs(5614) <= not a;
    outputs(5615) <= a xor b;
    outputs(5616) <= not a;
    outputs(5617) <= not b;
    outputs(5618) <= not b;
    outputs(5619) <= a and b;
    outputs(5620) <= a;
    outputs(5621) <= b;
    outputs(5622) <= not a;
    outputs(5623) <= b;
    outputs(5624) <= a;
    outputs(5625) <= a xor b;
    outputs(5626) <= not (a xor b);
    outputs(5627) <= b;
    outputs(5628) <= a xor b;
    outputs(5629) <= not b;
    outputs(5630) <= b;
    outputs(5631) <= not a;
    outputs(5632) <= a or b;
    outputs(5633) <= not (a xor b);
    outputs(5634) <= a;
    outputs(5635) <= a xor b;
    outputs(5636) <= a xor b;
    outputs(5637) <= a xor b;
    outputs(5638) <= a and b;
    outputs(5639) <= not b;
    outputs(5640) <= a xor b;
    outputs(5641) <= not b;
    outputs(5642) <= a xor b;
    outputs(5643) <= not b;
    outputs(5644) <= b;
    outputs(5645) <= not (a xor b);
    outputs(5646) <= not a;
    outputs(5647) <= a xor b;
    outputs(5648) <= a xor b;
    outputs(5649) <= not a;
    outputs(5650) <= not b;
    outputs(5651) <= not (a and b);
    outputs(5652) <= b and not a;
    outputs(5653) <= a xor b;
    outputs(5654) <= not a;
    outputs(5655) <= a and b;
    outputs(5656) <= b;
    outputs(5657) <= not a;
    outputs(5658) <= not a;
    outputs(5659) <= b;
    outputs(5660) <= not a;
    outputs(5661) <= not (a and b);
    outputs(5662) <= a xor b;
    outputs(5663) <= a xor b;
    outputs(5664) <= a xor b;
    outputs(5665) <= a and not b;
    outputs(5666) <= a or b;
    outputs(5667) <= not a;
    outputs(5668) <= not a or b;
    outputs(5669) <= a and b;
    outputs(5670) <= a or b;
    outputs(5671) <= not (a xor b);
    outputs(5672) <= a or b;
    outputs(5673) <= a;
    outputs(5674) <= b and not a;
    outputs(5675) <= b and not a;
    outputs(5676) <= not b;
    outputs(5677) <= not b or a;
    outputs(5678) <= not (a xor b);
    outputs(5679) <= not b;
    outputs(5680) <= b;
    outputs(5681) <= not (a xor b);
    outputs(5682) <= b;
    outputs(5683) <= a or b;
    outputs(5684) <= a xor b;
    outputs(5685) <= not (a and b);
    outputs(5686) <= not b;
    outputs(5687) <= a xor b;
    outputs(5688) <= a xor b;
    outputs(5689) <= b;
    outputs(5690) <= not (a xor b);
    outputs(5691) <= not a;
    outputs(5692) <= a;
    outputs(5693) <= not (a xor b);
    outputs(5694) <= not (a xor b);
    outputs(5695) <= a xor b;
    outputs(5696) <= not a;
    outputs(5697) <= not a or b;
    outputs(5698) <= a;
    outputs(5699) <= b;
    outputs(5700) <= not b or a;
    outputs(5701) <= not (a xor b);
    outputs(5702) <= a or b;
    outputs(5703) <= a and not b;
    outputs(5704) <= a;
    outputs(5705) <= not a;
    outputs(5706) <= not a;
    outputs(5707) <= a and b;
    outputs(5708) <= a xor b;
    outputs(5709) <= not (a xor b);
    outputs(5710) <= not a;
    outputs(5711) <= a and not b;
    outputs(5712) <= a and b;
    outputs(5713) <= not b;
    outputs(5714) <= a;
    outputs(5715) <= not a;
    outputs(5716) <= not (a xor b);
    outputs(5717) <= not a or b;
    outputs(5718) <= a xor b;
    outputs(5719) <= not (a xor b);
    outputs(5720) <= a xor b;
    outputs(5721) <= not (a xor b);
    outputs(5722) <= not (a xor b);
    outputs(5723) <= not (a xor b);
    outputs(5724) <= a or b;
    outputs(5725) <= not a or b;
    outputs(5726) <= b;
    outputs(5727) <= not (a and b);
    outputs(5728) <= b;
    outputs(5729) <= not a;
    outputs(5730) <= not b;
    outputs(5731) <= not a;
    outputs(5732) <= a and b;
    outputs(5733) <= not (a xor b);
    outputs(5734) <= a and b;
    outputs(5735) <= not b or a;
    outputs(5736) <= a and b;
    outputs(5737) <= b;
    outputs(5738) <= a xor b;
    outputs(5739) <= not b;
    outputs(5740) <= a and not b;
    outputs(5741) <= a;
    outputs(5742) <= not (a xor b);
    outputs(5743) <= not a;
    outputs(5744) <= not b;
    outputs(5745) <= a xor b;
    outputs(5746) <= b;
    outputs(5747) <= a;
    outputs(5748) <= a;
    outputs(5749) <= b;
    outputs(5750) <= not b;
    outputs(5751) <= not (a xor b);
    outputs(5752) <= a xor b;
    outputs(5753) <= not (a xor b);
    outputs(5754) <= a xor b;
    outputs(5755) <= not (a and b);
    outputs(5756) <= not b;
    outputs(5757) <= not (a xor b);
    outputs(5758) <= a and b;
    outputs(5759) <= not b;
    outputs(5760) <= a or b;
    outputs(5761) <= b;
    outputs(5762) <= not (a xor b);
    outputs(5763) <= not b or a;
    outputs(5764) <= b;
    outputs(5765) <= b and not a;
    outputs(5766) <= a;
    outputs(5767) <= not b;
    outputs(5768) <= a;
    outputs(5769) <= not a;
    outputs(5770) <= a;
    outputs(5771) <= not (a xor b);
    outputs(5772) <= a or b;
    outputs(5773) <= not (a xor b);
    outputs(5774) <= not a;
    outputs(5775) <= a xor b;
    outputs(5776) <= b;
    outputs(5777) <= not b;
    outputs(5778) <= not (a xor b);
    outputs(5779) <= a xor b;
    outputs(5780) <= not b;
    outputs(5781) <= not (a xor b);
    outputs(5782) <= a xor b;
    outputs(5783) <= b;
    outputs(5784) <= a;
    outputs(5785) <= b;
    outputs(5786) <= not a;
    outputs(5787) <= not b;
    outputs(5788) <= b;
    outputs(5789) <= a xor b;
    outputs(5790) <= a and not b;
    outputs(5791) <= not a or b;
    outputs(5792) <= not (a or b);
    outputs(5793) <= a xor b;
    outputs(5794) <= a xor b;
    outputs(5795) <= a or b;
    outputs(5796) <= not b;
    outputs(5797) <= b;
    outputs(5798) <= a or b;
    outputs(5799) <= not (a xor b);
    outputs(5800) <= not b;
    outputs(5801) <= not b or a;
    outputs(5802) <= not b;
    outputs(5803) <= not a or b;
    outputs(5804) <= not a or b;
    outputs(5805) <= not a;
    outputs(5806) <= not b;
    outputs(5807) <= not (a xor b);
    outputs(5808) <= a xor b;
    outputs(5809) <= b;
    outputs(5810) <= not b;
    outputs(5811) <= a or b;
    outputs(5812) <= a and b;
    outputs(5813) <= a;
    outputs(5814) <= not b;
    outputs(5815) <= b;
    outputs(5816) <= b;
    outputs(5817) <= a and b;
    outputs(5818) <= not a;
    outputs(5819) <= a;
    outputs(5820) <= not b;
    outputs(5821) <= a xor b;
    outputs(5822) <= not b;
    outputs(5823) <= not (a xor b);
    outputs(5824) <= b;
    outputs(5825) <= a xor b;
    outputs(5826) <= b and not a;
    outputs(5827) <= not (a xor b);
    outputs(5828) <= a;
    outputs(5829) <= not (a xor b);
    outputs(5830) <= a xor b;
    outputs(5831) <= a;
    outputs(5832) <= not (a xor b);
    outputs(5833) <= not b;
    outputs(5834) <= a xor b;
    outputs(5835) <= not b;
    outputs(5836) <= not b;
    outputs(5837) <= a;
    outputs(5838) <= a xor b;
    outputs(5839) <= a;
    outputs(5840) <= not a;
    outputs(5841) <= not a;
    outputs(5842) <= a and b;
    outputs(5843) <= not b;
    outputs(5844) <= a;
    outputs(5845) <= not (a xor b);
    outputs(5846) <= not b;
    outputs(5847) <= a xor b;
    outputs(5848) <= b and not a;
    outputs(5849) <= not a;
    outputs(5850) <= not (a xor b);
    outputs(5851) <= b;
    outputs(5852) <= a and not b;
    outputs(5853) <= not b;
    outputs(5854) <= a xor b;
    outputs(5855) <= a and not b;
    outputs(5856) <= not a;
    outputs(5857) <= a xor b;
    outputs(5858) <= not (a xor b);
    outputs(5859) <= not (a xor b);
    outputs(5860) <= a;
    outputs(5861) <= not (a xor b);
    outputs(5862) <= a xor b;
    outputs(5863) <= a xor b;
    outputs(5864) <= not b;
    outputs(5865) <= not a;
    outputs(5866) <= b;
    outputs(5867) <= not b;
    outputs(5868) <= not b;
    outputs(5869) <= a or b;
    outputs(5870) <= a and not b;
    outputs(5871) <= not (a xor b);
    outputs(5872) <= a xor b;
    outputs(5873) <= not b;
    outputs(5874) <= not a;
    outputs(5875) <= not a;
    outputs(5876) <= a xor b;
    outputs(5877) <= not a;
    outputs(5878) <= not (a xor b);
    outputs(5879) <= b and not a;
    outputs(5880) <= not b;
    outputs(5881) <= a and b;
    outputs(5882) <= not (a and b);
    outputs(5883) <= a;
    outputs(5884) <= not (a xor b);
    outputs(5885) <= not a;
    outputs(5886) <= a;
    outputs(5887) <= a xor b;
    outputs(5888) <= b;
    outputs(5889) <= a xor b;
    outputs(5890) <= not a;
    outputs(5891) <= not b;
    outputs(5892) <= not b;
    outputs(5893) <= a and b;
    outputs(5894) <= not (a xor b);
    outputs(5895) <= not (a xor b);
    outputs(5896) <= not (a xor b);
    outputs(5897) <= not (a and b);
    outputs(5898) <= not a;
    outputs(5899) <= a or b;
    outputs(5900) <= not (a or b);
    outputs(5901) <= not (a xor b);
    outputs(5902) <= b;
    outputs(5903) <= a and b;
    outputs(5904) <= a and b;
    outputs(5905) <= b;
    outputs(5906) <= not b or a;
    outputs(5907) <= not (a xor b);
    outputs(5908) <= not b or a;
    outputs(5909) <= b;
    outputs(5910) <= a or b;
    outputs(5911) <= a and not b;
    outputs(5912) <= a xor b;
    outputs(5913) <= b;
    outputs(5914) <= not a;
    outputs(5915) <= not (a xor b);
    outputs(5916) <= not a;
    outputs(5917) <= a or b;
    outputs(5918) <= a xor b;
    outputs(5919) <= not a or b;
    outputs(5920) <= not (a and b);
    outputs(5921) <= not a;
    outputs(5922) <= a xor b;
    outputs(5923) <= not (a xor b);
    outputs(5924) <= not b;
    outputs(5925) <= not (a xor b);
    outputs(5926) <= not b;
    outputs(5927) <= a xor b;
    outputs(5928) <= b;
    outputs(5929) <= not b;
    outputs(5930) <= not (a and b);
    outputs(5931) <= a xor b;
    outputs(5932) <= not b;
    outputs(5933) <= b;
    outputs(5934) <= a xor b;
    outputs(5935) <= a and b;
    outputs(5936) <= a and b;
    outputs(5937) <= not b;
    outputs(5938) <= not (a xor b);
    outputs(5939) <= a and not b;
    outputs(5940) <= not (a xor b);
    outputs(5941) <= not (a xor b);
    outputs(5942) <= not b;
    outputs(5943) <= not b;
    outputs(5944) <= a and not b;
    outputs(5945) <= a;
    outputs(5946) <= a xor b;
    outputs(5947) <= a;
    outputs(5948) <= not a;
    outputs(5949) <= a;
    outputs(5950) <= a;
    outputs(5951) <= a and not b;
    outputs(5952) <= not a;
    outputs(5953) <= a;
    outputs(5954) <= not a or b;
    outputs(5955) <= a xor b;
    outputs(5956) <= not (a xor b);
    outputs(5957) <= a xor b;
    outputs(5958) <= a xor b;
    outputs(5959) <= not a;
    outputs(5960) <= a xor b;
    outputs(5961) <= not b or a;
    outputs(5962) <= b;
    outputs(5963) <= not (a and b);
    outputs(5964) <= a and not b;
    outputs(5965) <= a and not b;
    outputs(5966) <= b and not a;
    outputs(5967) <= not (a xor b);
    outputs(5968) <= b and not a;
    outputs(5969) <= not (a and b);
    outputs(5970) <= not a or b;
    outputs(5971) <= b;
    outputs(5972) <= b;
    outputs(5973) <= b and not a;
    outputs(5974) <= a;
    outputs(5975) <= not (a xor b);
    outputs(5976) <= not (a xor b);
    outputs(5977) <= a xor b;
    outputs(5978) <= a;
    outputs(5979) <= b;
    outputs(5980) <= not a or b;
    outputs(5981) <= not b;
    outputs(5982) <= a and b;
    outputs(5983) <= not (a xor b);
    outputs(5984) <= a;
    outputs(5985) <= not b or a;
    outputs(5986) <= not (a xor b);
    outputs(5987) <= not a;
    outputs(5988) <= a and not b;
    outputs(5989) <= not b;
    outputs(5990) <= not (a xor b);
    outputs(5991) <= a;
    outputs(5992) <= b;
    outputs(5993) <= not a or b;
    outputs(5994) <= not b or a;
    outputs(5995) <= not a;
    outputs(5996) <= b;
    outputs(5997) <= a or b;
    outputs(5998) <= b;
    outputs(5999) <= a xor b;
    outputs(6000) <= not b or a;
    outputs(6001) <= not (a xor b);
    outputs(6002) <= not (a and b);
    outputs(6003) <= a;
    outputs(6004) <= a xor b;
    outputs(6005) <= not b or a;
    outputs(6006) <= a and not b;
    outputs(6007) <= not b;
    outputs(6008) <= a;
    outputs(6009) <= a xor b;
    outputs(6010) <= a;
    outputs(6011) <= b;
    outputs(6012) <= a xor b;
    outputs(6013) <= not a or b;
    outputs(6014) <= b;
    outputs(6015) <= not b;
    outputs(6016) <= a xor b;
    outputs(6017) <= a and not b;
    outputs(6018) <= not (a xor b);
    outputs(6019) <= not b;
    outputs(6020) <= not a;
    outputs(6021) <= a xor b;
    outputs(6022) <= not b;
    outputs(6023) <= b;
    outputs(6024) <= not a;
    outputs(6025) <= not b;
    outputs(6026) <= a xor b;
    outputs(6027) <= not (a xor b);
    outputs(6028) <= not a;
    outputs(6029) <= not (a xor b);
    outputs(6030) <= b;
    outputs(6031) <= not b;
    outputs(6032) <= not (a xor b);
    outputs(6033) <= b;
    outputs(6034) <= a xor b;
    outputs(6035) <= not (a and b);
    outputs(6036) <= a;
    outputs(6037) <= a;
    outputs(6038) <= a;
    outputs(6039) <= a;
    outputs(6040) <= not a;
    outputs(6041) <= b;
    outputs(6042) <= a xor b;
    outputs(6043) <= not b;
    outputs(6044) <= not a;
    outputs(6045) <= not (a xor b);
    outputs(6046) <= b;
    outputs(6047) <= not b;
    outputs(6048) <= a and b;
    outputs(6049) <= not (a xor b);
    outputs(6050) <= not (a xor b);
    outputs(6051) <= b;
    outputs(6052) <= not (a xor b);
    outputs(6053) <= not b;
    outputs(6054) <= not (a xor b);
    outputs(6055) <= not (a and b);
    outputs(6056) <= b and not a;
    outputs(6057) <= b;
    outputs(6058) <= not (a xor b);
    outputs(6059) <= b;
    outputs(6060) <= not (a xor b);
    outputs(6061) <= not b;
    outputs(6062) <= b;
    outputs(6063) <= b;
    outputs(6064) <= a xor b;
    outputs(6065) <= a xor b;
    outputs(6066) <= not (a or b);
    outputs(6067) <= a xor b;
    outputs(6068) <= a xor b;
    outputs(6069) <= not (a xor b);
    outputs(6070) <= not a;
    outputs(6071) <= b;
    outputs(6072) <= b;
    outputs(6073) <= b;
    outputs(6074) <= not (a or b);
    outputs(6075) <= not a;
    outputs(6076) <= a;
    outputs(6077) <= b;
    outputs(6078) <= a;
    outputs(6079) <= not (a and b);
    outputs(6080) <= not (a xor b);
    outputs(6081) <= a xor b;
    outputs(6082) <= not a;
    outputs(6083) <= a and not b;
    outputs(6084) <= a and not b;
    outputs(6085) <= a;
    outputs(6086) <= a;
    outputs(6087) <= not a;
    outputs(6088) <= b;
    outputs(6089) <= not (a xor b);
    outputs(6090) <= not (a and b);
    outputs(6091) <= not b;
    outputs(6092) <= b;
    outputs(6093) <= not a;
    outputs(6094) <= not (a xor b);
    outputs(6095) <= a xor b;
    outputs(6096) <= a or b;
    outputs(6097) <= b and not a;
    outputs(6098) <= not (a xor b);
    outputs(6099) <= not b or a;
    outputs(6100) <= b and not a;
    outputs(6101) <= a or b;
    outputs(6102) <= not a;
    outputs(6103) <= a;
    outputs(6104) <= not (a xor b);
    outputs(6105) <= not (a xor b);
    outputs(6106) <= a or b;
    outputs(6107) <= b;
    outputs(6108) <= b;
    outputs(6109) <= not (a or b);
    outputs(6110) <= b and not a;
    outputs(6111) <= not (a or b);
    outputs(6112) <= a xor b;
    outputs(6113) <= a;
    outputs(6114) <= a;
    outputs(6115) <= b;
    outputs(6116) <= not a;
    outputs(6117) <= a xor b;
    outputs(6118) <= not b or a;
    outputs(6119) <= not (a xor b);
    outputs(6120) <= a xor b;
    outputs(6121) <= a;
    outputs(6122) <= a;
    outputs(6123) <= not a;
    outputs(6124) <= a xor b;
    outputs(6125) <= not b;
    outputs(6126) <= not b or a;
    outputs(6127) <= not a;
    outputs(6128) <= b and not a;
    outputs(6129) <= not b;
    outputs(6130) <= a xor b;
    outputs(6131) <= a or b;
    outputs(6132) <= not (a xor b);
    outputs(6133) <= b;
    outputs(6134) <= not b;
    outputs(6135) <= b;
    outputs(6136) <= a xor b;
    outputs(6137) <= not (a xor b);
    outputs(6138) <= not a;
    outputs(6139) <= not (a xor b);
    outputs(6140) <= not a or b;
    outputs(6141) <= a;
    outputs(6142) <= a xor b;
    outputs(6143) <= a;
    outputs(6144) <= b and not a;
    outputs(6145) <= a and b;
    outputs(6146) <= a and not b;
    outputs(6147) <= a;
    outputs(6148) <= b;
    outputs(6149) <= not (a xor b);
    outputs(6150) <= a and b;
    outputs(6151) <= not a;
    outputs(6152) <= a and not b;
    outputs(6153) <= not b;
    outputs(6154) <= a xor b;
    outputs(6155) <= not b;
    outputs(6156) <= not b;
    outputs(6157) <= not (a xor b);
    outputs(6158) <= not (a xor b);
    outputs(6159) <= not a;
    outputs(6160) <= not b;
    outputs(6161) <= not b or a;
    outputs(6162) <= not (a xor b);
    outputs(6163) <= a;
    outputs(6164) <= a xor b;
    outputs(6165) <= not (a or b);
    outputs(6166) <= not (a xor b);
    outputs(6167) <= not b;
    outputs(6168) <= a;
    outputs(6169) <= not (a xor b);
    outputs(6170) <= a xor b;
    outputs(6171) <= not a;
    outputs(6172) <= a;
    outputs(6173) <= a;
    outputs(6174) <= not (a xor b);
    outputs(6175) <= a and b;
    outputs(6176) <= not a;
    outputs(6177) <= a and not b;
    outputs(6178) <= b;
    outputs(6179) <= b and not a;
    outputs(6180) <= not b;
    outputs(6181) <= b;
    outputs(6182) <= a xor b;
    outputs(6183) <= not (a or b);
    outputs(6184) <= b;
    outputs(6185) <= b;
    outputs(6186) <= not a;
    outputs(6187) <= not (a xor b);
    outputs(6188) <= a;
    outputs(6189) <= a and not b;
    outputs(6190) <= not (a xor b);
    outputs(6191) <= not (a xor b);
    outputs(6192) <= b;
    outputs(6193) <= a;
    outputs(6194) <= a and b;
    outputs(6195) <= b and not a;
    outputs(6196) <= not a;
    outputs(6197) <= not (a or b);
    outputs(6198) <= a xor b;
    outputs(6199) <= not b;
    outputs(6200) <= a;
    outputs(6201) <= b;
    outputs(6202) <= a and b;
    outputs(6203) <= a and not b;
    outputs(6204) <= a and b;
    outputs(6205) <= a and not b;
    outputs(6206) <= not (a and b);
    outputs(6207) <= not b;
    outputs(6208) <= a;
    outputs(6209) <= not b;
    outputs(6210) <= b;
    outputs(6211) <= not (a xor b);
    outputs(6212) <= a xor b;
    outputs(6213) <= a and not b;
    outputs(6214) <= a xor b;
    outputs(6215) <= a;
    outputs(6216) <= not b;
    outputs(6217) <= a;
    outputs(6218) <= a and not b;
    outputs(6219) <= b;
    outputs(6220) <= not (a xor b);
    outputs(6221) <= b;
    outputs(6222) <= not (a xor b);
    outputs(6223) <= b and not a;
    outputs(6224) <= a;
    outputs(6225) <= not b;
    outputs(6226) <= not a;
    outputs(6227) <= not b;
    outputs(6228) <= not (a xor b);
    outputs(6229) <= b;
    outputs(6230) <= a;
    outputs(6231) <= not (a xor b);
    outputs(6232) <= not b or a;
    outputs(6233) <= not b;
    outputs(6234) <= a xor b;
    outputs(6235) <= not b;
    outputs(6236) <= a xor b;
    outputs(6237) <= b and not a;
    outputs(6238) <= not b;
    outputs(6239) <= a;
    outputs(6240) <= a xor b;
    outputs(6241) <= b;
    outputs(6242) <= not a;
    outputs(6243) <= a;
    outputs(6244) <= b;
    outputs(6245) <= not (a xor b);
    outputs(6246) <= not a;
    outputs(6247) <= a or b;
    outputs(6248) <= not (a xor b);
    outputs(6249) <= not a;
    outputs(6250) <= a or b;
    outputs(6251) <= a;
    outputs(6252) <= b;
    outputs(6253) <= a;
    outputs(6254) <= not a;
    outputs(6255) <= b;
    outputs(6256) <= a;
    outputs(6257) <= not (a xor b);
    outputs(6258) <= b;
    outputs(6259) <= not (a and b);
    outputs(6260) <= not (a xor b);
    outputs(6261) <= a xor b;
    outputs(6262) <= not (a or b);
    outputs(6263) <= not a;
    outputs(6264) <= not b;
    outputs(6265) <= not b;
    outputs(6266) <= not (a xor b);
    outputs(6267) <= not b;
    outputs(6268) <= a xor b;
    outputs(6269) <= not a;
    outputs(6270) <= b;
    outputs(6271) <= a and b;
    outputs(6272) <= a xor b;
    outputs(6273) <= a xor b;
    outputs(6274) <= a;
    outputs(6275) <= not b;
    outputs(6276) <= a xor b;
    outputs(6277) <= a xor b;
    outputs(6278) <= not a;
    outputs(6279) <= a xor b;
    outputs(6280) <= not (a xor b);
    outputs(6281) <= a;
    outputs(6282) <= a;
    outputs(6283) <= not a;
    outputs(6284) <= not (a xor b);
    outputs(6285) <= not a;
    outputs(6286) <= not b;
    outputs(6287) <= not b;
    outputs(6288) <= b;
    outputs(6289) <= not a;
    outputs(6290) <= not a or b;
    outputs(6291) <= not b or a;
    outputs(6292) <= a xor b;
    outputs(6293) <= a and b;
    outputs(6294) <= a;
    outputs(6295) <= a;
    outputs(6296) <= b and not a;
    outputs(6297) <= a;
    outputs(6298) <= a xor b;
    outputs(6299) <= not a;
    outputs(6300) <= a xor b;
    outputs(6301) <= a xor b;
    outputs(6302) <= a or b;
    outputs(6303) <= not (a xor b);
    outputs(6304) <= a xor b;
    outputs(6305) <= a and b;
    outputs(6306) <= a;
    outputs(6307) <= not b;
    outputs(6308) <= a and not b;
    outputs(6309) <= a xor b;
    outputs(6310) <= a;
    outputs(6311) <= a xor b;
    outputs(6312) <= not b;
    outputs(6313) <= a xor b;
    outputs(6314) <= not (a xor b);
    outputs(6315) <= not (a xor b);
    outputs(6316) <= b;
    outputs(6317) <= b;
    outputs(6318) <= b;
    outputs(6319) <= a;
    outputs(6320) <= not b;
    outputs(6321) <= not a;
    outputs(6322) <= not (a and b);
    outputs(6323) <= not a;
    outputs(6324) <= not a;
    outputs(6325) <= not (a xor b);
    outputs(6326) <= b and not a;
    outputs(6327) <= not b;
    outputs(6328) <= not (a xor b);
    outputs(6329) <= not a;
    outputs(6330) <= a xor b;
    outputs(6331) <= not (a xor b);
    outputs(6332) <= a;
    outputs(6333) <= b;
    outputs(6334) <= b;
    outputs(6335) <= a xor b;
    outputs(6336) <= a xor b;
    outputs(6337) <= a xor b;
    outputs(6338) <= not a;
    outputs(6339) <= not a;
    outputs(6340) <= not (a and b);
    outputs(6341) <= a and not b;
    outputs(6342) <= not b;
    outputs(6343) <= a;
    outputs(6344) <= a xor b;
    outputs(6345) <= not (a xor b);
    outputs(6346) <= not (a xor b);
    outputs(6347) <= not (a or b);
    outputs(6348) <= not (a xor b);
    outputs(6349) <= b and not a;
    outputs(6350) <= not a or b;
    outputs(6351) <= not b;
    outputs(6352) <= not (a or b);
    outputs(6353) <= a xor b;
    outputs(6354) <= a and b;
    outputs(6355) <= not (a xor b);
    outputs(6356) <= not (a or b);
    outputs(6357) <= b;
    outputs(6358) <= not (a xor b);
    outputs(6359) <= not (a xor b);
    outputs(6360) <= not b;
    outputs(6361) <= not a;
    outputs(6362) <= b;
    outputs(6363) <= not (a xor b);
    outputs(6364) <= not (a xor b);
    outputs(6365) <= a;
    outputs(6366) <= not b;
    outputs(6367) <= a xor b;
    outputs(6368) <= a xor b;
    outputs(6369) <= a xor b;
    outputs(6370) <= b;
    outputs(6371) <= not (a or b);
    outputs(6372) <= b;
    outputs(6373) <= b;
    outputs(6374) <= not a;
    outputs(6375) <= a or b;
    outputs(6376) <= not (a xor b);
    outputs(6377) <= b;
    outputs(6378) <= b and not a;
    outputs(6379) <= not b;
    outputs(6380) <= a;
    outputs(6381) <= not (a xor b);
    outputs(6382) <= a or b;
    outputs(6383) <= not (a xor b);
    outputs(6384) <= not (a or b);
    outputs(6385) <= a and b;
    outputs(6386) <= not (a xor b);
    outputs(6387) <= not (a xor b);
    outputs(6388) <= not (a xor b);
    outputs(6389) <= not (a and b);
    outputs(6390) <= b;
    outputs(6391) <= not a;
    outputs(6392) <= b;
    outputs(6393) <= a and not b;
    outputs(6394) <= b and not a;
    outputs(6395) <= not a;
    outputs(6396) <= a;
    outputs(6397) <= not (a xor b);
    outputs(6398) <= not a;
    outputs(6399) <= b;
    outputs(6400) <= not (a or b);
    outputs(6401) <= not (a and b);
    outputs(6402) <= not a;
    outputs(6403) <= b;
    outputs(6404) <= not a;
    outputs(6405) <= not b;
    outputs(6406) <= a xor b;
    outputs(6407) <= a xor b;
    outputs(6408) <= not b or a;
    outputs(6409) <= not (a xor b);
    outputs(6410) <= a xor b;
    outputs(6411) <= a xor b;
    outputs(6412) <= not a or b;
    outputs(6413) <= a xor b;
    outputs(6414) <= b;
    outputs(6415) <= a xor b;
    outputs(6416) <= b;
    outputs(6417) <= not a;
    outputs(6418) <= not (a xor b);
    outputs(6419) <= b;
    outputs(6420) <= b;
    outputs(6421) <= a xor b;
    outputs(6422) <= not (a xor b);
    outputs(6423) <= a xor b;
    outputs(6424) <= a xor b;
    outputs(6425) <= not (a xor b);
    outputs(6426) <= b;
    outputs(6427) <= b and not a;
    outputs(6428) <= not (a xor b);
    outputs(6429) <= a xor b;
    outputs(6430) <= a or b;
    outputs(6431) <= not b;
    outputs(6432) <= not (a xor b);
    outputs(6433) <= a;
    outputs(6434) <= not a;
    outputs(6435) <= a or b;
    outputs(6436) <= not b;
    outputs(6437) <= not b;
    outputs(6438) <= not a;
    outputs(6439) <= not (a xor b);
    outputs(6440) <= b;
    outputs(6441) <= not b;
    outputs(6442) <= not b;
    outputs(6443) <= a;
    outputs(6444) <= not a;
    outputs(6445) <= a or b;
    outputs(6446) <= not (a xor b);
    outputs(6447) <= not b;
    outputs(6448) <= a and b;
    outputs(6449) <= not a;
    outputs(6450) <= a or b;
    outputs(6451) <= not a;
    outputs(6452) <= not (a xor b);
    outputs(6453) <= not (a or b);
    outputs(6454) <= not b;
    outputs(6455) <= not b;
    outputs(6456) <= a and b;
    outputs(6457) <= a;
    outputs(6458) <= b and not a;
    outputs(6459) <= b;
    outputs(6460) <= not a;
    outputs(6461) <= not (a xor b);
    outputs(6462) <= not b;
    outputs(6463) <= not a or b;
    outputs(6464) <= b;
    outputs(6465) <= a and b;
    outputs(6466) <= b and not a;
    outputs(6467) <= not a;
    outputs(6468) <= b;
    outputs(6469) <= b;
    outputs(6470) <= a;
    outputs(6471) <= not b;
    outputs(6472) <= not a or b;
    outputs(6473) <= not a;
    outputs(6474) <= a and b;
    outputs(6475) <= b;
    outputs(6476) <= not b;
    outputs(6477) <= a or b;
    outputs(6478) <= a or b;
    outputs(6479) <= b and not a;
    outputs(6480) <= not b;
    outputs(6481) <= not (a and b);
    outputs(6482) <= not (a xor b);
    outputs(6483) <= not b;
    outputs(6484) <= not a;
    outputs(6485) <= not (a xor b);
    outputs(6486) <= not b;
    outputs(6487) <= not (a or b);
    outputs(6488) <= b;
    outputs(6489) <= not a;
    outputs(6490) <= not (a xor b);
    outputs(6491) <= not (a and b);
    outputs(6492) <= not b;
    outputs(6493) <= not b;
    outputs(6494) <= b and not a;
    outputs(6495) <= a xor b;
    outputs(6496) <= not (a and b);
    outputs(6497) <= a;
    outputs(6498) <= not (a and b);
    outputs(6499) <= not a;
    outputs(6500) <= not a;
    outputs(6501) <= b;
    outputs(6502) <= not (a or b);
    outputs(6503) <= b;
    outputs(6504) <= not (a xor b);
    outputs(6505) <= not b;
    outputs(6506) <= not a or b;
    outputs(6507) <= not a;
    outputs(6508) <= a;
    outputs(6509) <= b and not a;
    outputs(6510) <= a xor b;
    outputs(6511) <= a;
    outputs(6512) <= not (a xor b);
    outputs(6513) <= b;
    outputs(6514) <= not a;
    outputs(6515) <= a xor b;
    outputs(6516) <= b and not a;
    outputs(6517) <= not (a and b);
    outputs(6518) <= a xor b;
    outputs(6519) <= a xor b;
    outputs(6520) <= not a;
    outputs(6521) <= b;
    outputs(6522) <= not a or b;
    outputs(6523) <= not b;
    outputs(6524) <= not (a xor b);
    outputs(6525) <= not b;
    outputs(6526) <= a xor b;
    outputs(6527) <= a xor b;
    outputs(6528) <= not b;
    outputs(6529) <= not b;
    outputs(6530) <= b;
    outputs(6531) <= b;
    outputs(6532) <= a and b;
    outputs(6533) <= b and not a;
    outputs(6534) <= b and not a;
    outputs(6535) <= b;
    outputs(6536) <= a and not b;
    outputs(6537) <= a xor b;
    outputs(6538) <= not a;
    outputs(6539) <= a;
    outputs(6540) <= not a or b;
    outputs(6541) <= not (a xor b);
    outputs(6542) <= a and b;
    outputs(6543) <= not a;
    outputs(6544) <= b;
    outputs(6545) <= not a;
    outputs(6546) <= a;
    outputs(6547) <= b;
    outputs(6548) <= not a or b;
    outputs(6549) <= a xor b;
    outputs(6550) <= not (a xor b);
    outputs(6551) <= not (a xor b);
    outputs(6552) <= b;
    outputs(6553) <= not b or a;
    outputs(6554) <= a;
    outputs(6555) <= b;
    outputs(6556) <= b;
    outputs(6557) <= not (a xor b);
    outputs(6558) <= a xor b;
    outputs(6559) <= not a or b;
    outputs(6560) <= a or b;
    outputs(6561) <= a;
    outputs(6562) <= not (a xor b);
    outputs(6563) <= a xor b;
    outputs(6564) <= not a;
    outputs(6565) <= b and not a;
    outputs(6566) <= not a;
    outputs(6567) <= a;
    outputs(6568) <= a and not b;
    outputs(6569) <= not (a or b);
    outputs(6570) <= not (a xor b);
    outputs(6571) <= b;
    outputs(6572) <= a and not b;
    outputs(6573) <= b;
    outputs(6574) <= b and not a;
    outputs(6575) <= not (a or b);
    outputs(6576) <= a xor b;
    outputs(6577) <= a xor b;
    outputs(6578) <= b;
    outputs(6579) <= a and not b;
    outputs(6580) <= not a;
    outputs(6581) <= a xor b;
    outputs(6582) <= a and b;
    outputs(6583) <= a xor b;
    outputs(6584) <= not a;
    outputs(6585) <= not (a xor b);
    outputs(6586) <= not b;
    outputs(6587) <= a;
    outputs(6588) <= a;
    outputs(6589) <= not (a xor b);
    outputs(6590) <= a and b;
    outputs(6591) <= b;
    outputs(6592) <= not b or a;
    outputs(6593) <= not a;
    outputs(6594) <= a;
    outputs(6595) <= not a;
    outputs(6596) <= b;
    outputs(6597) <= a xor b;
    outputs(6598) <= not b;
    outputs(6599) <= not b;
    outputs(6600) <= not b;
    outputs(6601) <= not (a or b);
    outputs(6602) <= not (a xor b);
    outputs(6603) <= not a;
    outputs(6604) <= not (a and b);
    outputs(6605) <= not (a and b);
    outputs(6606) <= a and not b;
    outputs(6607) <= a;
    outputs(6608) <= not b;
    outputs(6609) <= not b;
    outputs(6610) <= not b;
    outputs(6611) <= a xor b;
    outputs(6612) <= not b;
    outputs(6613) <= a;
    outputs(6614) <= not a;
    outputs(6615) <= a xor b;
    outputs(6616) <= not b;
    outputs(6617) <= not a;
    outputs(6618) <= a;
    outputs(6619) <= a and b;
    outputs(6620) <= b;
    outputs(6621) <= a xor b;
    outputs(6622) <= b;
    outputs(6623) <= not a;
    outputs(6624) <= a xor b;
    outputs(6625) <= not a;
    outputs(6626) <= a and b;
    outputs(6627) <= a;
    outputs(6628) <= not a;
    outputs(6629) <= a xor b;
    outputs(6630) <= not b;
    outputs(6631) <= not a;
    outputs(6632) <= not (a xor b);
    outputs(6633) <= not a or b;
    outputs(6634) <= not (a xor b);
    outputs(6635) <= a;
    outputs(6636) <= a or b;
    outputs(6637) <= a;
    outputs(6638) <= a xor b;
    outputs(6639) <= a;
    outputs(6640) <= b;
    outputs(6641) <= not (a and b);
    outputs(6642) <= not a or b;
    outputs(6643) <= not a;
    outputs(6644) <= a and b;
    outputs(6645) <= b;
    outputs(6646) <= not a or b;
    outputs(6647) <= a xor b;
    outputs(6648) <= b;
    outputs(6649) <= not a;
    outputs(6650) <= not (a xor b);
    outputs(6651) <= b;
    outputs(6652) <= a;
    outputs(6653) <= not a;
    outputs(6654) <= a;
    outputs(6655) <= b;
    outputs(6656) <= a and not b;
    outputs(6657) <= b;
    outputs(6658) <= not b;
    outputs(6659) <= a;
    outputs(6660) <= b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= a and not b;
    outputs(6663) <= not b or a;
    outputs(6664) <= not a;
    outputs(6665) <= b;
    outputs(6666) <= not (a xor b);
    outputs(6667) <= a xor b;
    outputs(6668) <= not a;
    outputs(6669) <= a and b;
    outputs(6670) <= not b;
    outputs(6671) <= a xor b;
    outputs(6672) <= not b;
    outputs(6673) <= not (a or b);
    outputs(6674) <= b;
    outputs(6675) <= not (a or b);
    outputs(6676) <= not b;
    outputs(6677) <= not a;
    outputs(6678) <= b and not a;
    outputs(6679) <= not (a xor b);
    outputs(6680) <= a xor b;
    outputs(6681) <= not b;
    outputs(6682) <= not (a xor b);
    outputs(6683) <= b;
    outputs(6684) <= a;
    outputs(6685) <= not b;
    outputs(6686) <= a xor b;
    outputs(6687) <= not (a xor b);
    outputs(6688) <= not b;
    outputs(6689) <= a xor b;
    outputs(6690) <= b;
    outputs(6691) <= a and b;
    outputs(6692) <= not a;
    outputs(6693) <= b;
    outputs(6694) <= a or b;
    outputs(6695) <= a and not b;
    outputs(6696) <= not b;
    outputs(6697) <= a and b;
    outputs(6698) <= not (a and b);
    outputs(6699) <= a;
    outputs(6700) <= not a;
    outputs(6701) <= not a or b;
    outputs(6702) <= not (a xor b);
    outputs(6703) <= not a;
    outputs(6704) <= not a;
    outputs(6705) <= a;
    outputs(6706) <= a xor b;
    outputs(6707) <= not (a xor b);
    outputs(6708) <= a;
    outputs(6709) <= not (a and b);
    outputs(6710) <= not b;
    outputs(6711) <= not (a xor b);
    outputs(6712) <= a and not b;
    outputs(6713) <= not b;
    outputs(6714) <= a or b;
    outputs(6715) <= not a;
    outputs(6716) <= a and b;
    outputs(6717) <= a xor b;
    outputs(6718) <= not (a xor b);
    outputs(6719) <= b;
    outputs(6720) <= a and b;
    outputs(6721) <= not a or b;
    outputs(6722) <= not b;
    outputs(6723) <= not (a and b);
    outputs(6724) <= not a;
    outputs(6725) <= a;
    outputs(6726) <= not b or a;
    outputs(6727) <= not b;
    outputs(6728) <= a;
    outputs(6729) <= a xor b;
    outputs(6730) <= b;
    outputs(6731) <= not (a or b);
    outputs(6732) <= a xor b;
    outputs(6733) <= a xor b;
    outputs(6734) <= not (a or b);
    outputs(6735) <= a xor b;
    outputs(6736) <= not (a xor b);
    outputs(6737) <= not a;
    outputs(6738) <= not (a or b);
    outputs(6739) <= not b or a;
    outputs(6740) <= not b;
    outputs(6741) <= a xor b;
    outputs(6742) <= not (a or b);
    outputs(6743) <= a;
    outputs(6744) <= b;
    outputs(6745) <= not a or b;
    outputs(6746) <= a and not b;
    outputs(6747) <= a xor b;
    outputs(6748) <= a;
    outputs(6749) <= not b;
    outputs(6750) <= b;
    outputs(6751) <= not (a xor b);
    outputs(6752) <= b;
    outputs(6753) <= not (a and b);
    outputs(6754) <= b;
    outputs(6755) <= a and b;
    outputs(6756) <= a and b;
    outputs(6757) <= a and not b;
    outputs(6758) <= a and b;
    outputs(6759) <= b;
    outputs(6760) <= not b;
    outputs(6761) <= a xor b;
    outputs(6762) <= a xor b;
    outputs(6763) <= a xor b;
    outputs(6764) <= a;
    outputs(6765) <= b;
    outputs(6766) <= a and b;
    outputs(6767) <= b;
    outputs(6768) <= b;
    outputs(6769) <= not b;
    outputs(6770) <= not a;
    outputs(6771) <= a xor b;
    outputs(6772) <= a or b;
    outputs(6773) <= not b or a;
    outputs(6774) <= not a;
    outputs(6775) <= b;
    outputs(6776) <= a;
    outputs(6777) <= b and not a;
    outputs(6778) <= a xor b;
    outputs(6779) <= a xor b;
    outputs(6780) <= b;
    outputs(6781) <= a and not b;
    outputs(6782) <= not (a xor b);
    outputs(6783) <= b;
    outputs(6784) <= a;
    outputs(6785) <= b;
    outputs(6786) <= a xor b;
    outputs(6787) <= a xor b;
    outputs(6788) <= a;
    outputs(6789) <= not (a and b);
    outputs(6790) <= a;
    outputs(6791) <= not b;
    outputs(6792) <= a xor b;
    outputs(6793) <= not b;
    outputs(6794) <= a and not b;
    outputs(6795) <= not b;
    outputs(6796) <= a;
    outputs(6797) <= not (a xor b);
    outputs(6798) <= not b;
    outputs(6799) <= b;
    outputs(6800) <= b;
    outputs(6801) <= not b;
    outputs(6802) <= not b;
    outputs(6803) <= b;
    outputs(6804) <= b;
    outputs(6805) <= not (a and b);
    outputs(6806) <= a xor b;
    outputs(6807) <= a and b;
    outputs(6808) <= a;
    outputs(6809) <= a and not b;
    outputs(6810) <= not (a or b);
    outputs(6811) <= a xor b;
    outputs(6812) <= a and b;
    outputs(6813) <= a;
    outputs(6814) <= not (a xor b);
    outputs(6815) <= a xor b;
    outputs(6816) <= not (a xor b);
    outputs(6817) <= not a;
    outputs(6818) <= b and not a;
    outputs(6819) <= a xor b;
    outputs(6820) <= not b;
    outputs(6821) <= not b;
    outputs(6822) <= b;
    outputs(6823) <= not b;
    outputs(6824) <= b;
    outputs(6825) <= not b;
    outputs(6826) <= a;
    outputs(6827) <= not a;
    outputs(6828) <= a and b;
    outputs(6829) <= b;
    outputs(6830) <= not (a xor b);
    outputs(6831) <= not b;
    outputs(6832) <= a;
    outputs(6833) <= not (a xor b);
    outputs(6834) <= not (a xor b);
    outputs(6835) <= a;
    outputs(6836) <= a xor b;
    outputs(6837) <= a;
    outputs(6838) <= not b;
    outputs(6839) <= not (a xor b);
    outputs(6840) <= b;
    outputs(6841) <= a and not b;
    outputs(6842) <= not a;
    outputs(6843) <= b;
    outputs(6844) <= a;
    outputs(6845) <= not b;
    outputs(6846) <= not b;
    outputs(6847) <= not (a xor b);
    outputs(6848) <= b;
    outputs(6849) <= not b or a;
    outputs(6850) <= 1'b0;
    outputs(6851) <= a xor b;
    outputs(6852) <= not a;
    outputs(6853) <= a;
    outputs(6854) <= b;
    outputs(6855) <= not (a xor b);
    outputs(6856) <= not b;
    outputs(6857) <= not b;
    outputs(6858) <= not (a xor b);
    outputs(6859) <= a;
    outputs(6860) <= not (a and b);
    outputs(6861) <= not (a xor b);
    outputs(6862) <= a xor b;
    outputs(6863) <= a;
    outputs(6864) <= b;
    outputs(6865) <= a and not b;
    outputs(6866) <= not a;
    outputs(6867) <= not b;
    outputs(6868) <= b;
    outputs(6869) <= not a;
    outputs(6870) <= a xor b;
    outputs(6871) <= not a;
    outputs(6872) <= a;
    outputs(6873) <= a and b;
    outputs(6874) <= a xor b;
    outputs(6875) <= a and b;
    outputs(6876) <= a;
    outputs(6877) <= not (a xor b);
    outputs(6878) <= not (a xor b);
    outputs(6879) <= a xor b;
    outputs(6880) <= b;
    outputs(6881) <= not a;
    outputs(6882) <= not a;
    outputs(6883) <= b;
    outputs(6884) <= not b;
    outputs(6885) <= b;
    outputs(6886) <= not b;
    outputs(6887) <= not a;
    outputs(6888) <= not (a xor b);
    outputs(6889) <= not a;
    outputs(6890) <= not a or b;
    outputs(6891) <= not a;
    outputs(6892) <= a xor b;
    outputs(6893) <= a xor b;
    outputs(6894) <= a and not b;
    outputs(6895) <= a xor b;
    outputs(6896) <= not b;
    outputs(6897) <= not b;
    outputs(6898) <= not a;
    outputs(6899) <= a;
    outputs(6900) <= a xor b;
    outputs(6901) <= not (a or b);
    outputs(6902) <= a xor b;
    outputs(6903) <= not a;
    outputs(6904) <= not a or b;
    outputs(6905) <= a and b;
    outputs(6906) <= not a;
    outputs(6907) <= a xor b;
    outputs(6908) <= b and not a;
    outputs(6909) <= b;
    outputs(6910) <= not (a xor b);
    outputs(6911) <= not a;
    outputs(6912) <= a xor b;
    outputs(6913) <= b;
    outputs(6914) <= not (a xor b);
    outputs(6915) <= not (a xor b);
    outputs(6916) <= not b;
    outputs(6917) <= not a;
    outputs(6918) <= not (a xor b);
    outputs(6919) <= a and b;
    outputs(6920) <= not b;
    outputs(6921) <= not (a xor b);
    outputs(6922) <= a;
    outputs(6923) <= a xor b;
    outputs(6924) <= a xor b;
    outputs(6925) <= b;
    outputs(6926) <= not a;
    outputs(6927) <= not (a xor b);
    outputs(6928) <= a;
    outputs(6929) <= not b or a;
    outputs(6930) <= a xor b;
    outputs(6931) <= b;
    outputs(6932) <= b;
    outputs(6933) <= not (a xor b);
    outputs(6934) <= not b;
    outputs(6935) <= a and not b;
    outputs(6936) <= not a;
    outputs(6937) <= not a;
    outputs(6938) <= a xor b;
    outputs(6939) <= a xor b;
    outputs(6940) <= not b;
    outputs(6941) <= a xor b;
    outputs(6942) <= b;
    outputs(6943) <= a;
    outputs(6944) <= a;
    outputs(6945) <= a xor b;
    outputs(6946) <= b;
    outputs(6947) <= a xor b;
    outputs(6948) <= a and not b;
    outputs(6949) <= not (a or b);
    outputs(6950) <= a xor b;
    outputs(6951) <= a;
    outputs(6952) <= a xor b;
    outputs(6953) <= a xor b;
    outputs(6954) <= not b;
    outputs(6955) <= a xor b;
    outputs(6956) <= not (a and b);
    outputs(6957) <= b;
    outputs(6958) <= not a;
    outputs(6959) <= b;
    outputs(6960) <= not b;
    outputs(6961) <= not b;
    outputs(6962) <= not b;
    outputs(6963) <= a xor b;
    outputs(6964) <= not (a or b);
    outputs(6965) <= not b;
    outputs(6966) <= a xor b;
    outputs(6967) <= b and not a;
    outputs(6968) <= a;
    outputs(6969) <= a or b;
    outputs(6970) <= a;
    outputs(6971) <= not a;
    outputs(6972) <= b and not a;
    outputs(6973) <= not (a xor b);
    outputs(6974) <= a xor b;
    outputs(6975) <= b;
    outputs(6976) <= a and not b;
    outputs(6977) <= not b;
    outputs(6978) <= a;
    outputs(6979) <= not (a xor b);
    outputs(6980) <= a or b;
    outputs(6981) <= not a or b;
    outputs(6982) <= a xor b;
    outputs(6983) <= a and b;
    outputs(6984) <= not b;
    outputs(6985) <= not b or a;
    outputs(6986) <= not b;
    outputs(6987) <= not a;
    outputs(6988) <= not (a xor b);
    outputs(6989) <= a and b;
    outputs(6990) <= not (a and b);
    outputs(6991) <= b;
    outputs(6992) <= a and b;
    outputs(6993) <= a xor b;
    outputs(6994) <= not b;
    outputs(6995) <= not (a xor b);
    outputs(6996) <= not (a xor b);
    outputs(6997) <= not (a and b);
    outputs(6998) <= a xor b;
    outputs(6999) <= a xor b;
    outputs(7000) <= not b;
    outputs(7001) <= a or b;
    outputs(7002) <= a xor b;
    outputs(7003) <= b;
    outputs(7004) <= a and not b;
    outputs(7005) <= not a;
    outputs(7006) <= a and not b;
    outputs(7007) <= a xor b;
    outputs(7008) <= not a;
    outputs(7009) <= not a;
    outputs(7010) <= b;
    outputs(7011) <= a xor b;
    outputs(7012) <= not a;
    outputs(7013) <= a;
    outputs(7014) <= b;
    outputs(7015) <= a xor b;
    outputs(7016) <= not b;
    outputs(7017) <= not (a xor b);
    outputs(7018) <= b;
    outputs(7019) <= a xor b;
    outputs(7020) <= not (a or b);
    outputs(7021) <= b;
    outputs(7022) <= a xor b;
    outputs(7023) <= not b;
    outputs(7024) <= b;
    outputs(7025) <= b;
    outputs(7026) <= b;
    outputs(7027) <= b and not a;
    outputs(7028) <= not b;
    outputs(7029) <= not (a xor b);
    outputs(7030) <= not b;
    outputs(7031) <= a and b;
    outputs(7032) <= not (a xor b);
    outputs(7033) <= a;
    outputs(7034) <= not a;
    outputs(7035) <= a and not b;
    outputs(7036) <= a;
    outputs(7037) <= a;
    outputs(7038) <= a or b;
    outputs(7039) <= not (a xor b);
    outputs(7040) <= b and not a;
    outputs(7041) <= not b;
    outputs(7042) <= a and b;
    outputs(7043) <= not a;
    outputs(7044) <= not a;
    outputs(7045) <= b;
    outputs(7046) <= a xor b;
    outputs(7047) <= not (a xor b);
    outputs(7048) <= a and not b;
    outputs(7049) <= a xor b;
    outputs(7050) <= not b;
    outputs(7051) <= not (a xor b);
    outputs(7052) <= b;
    outputs(7053) <= a xor b;
    outputs(7054) <= not a;
    outputs(7055) <= a xor b;
    outputs(7056) <= a and not b;
    outputs(7057) <= a xor b;
    outputs(7058) <= a xor b;
    outputs(7059) <= a and b;
    outputs(7060) <= b;
    outputs(7061) <= not (a and b);
    outputs(7062) <= a;
    outputs(7063) <= a and b;
    outputs(7064) <= not (a xor b);
    outputs(7065) <= not a;
    outputs(7066) <= not b;
    outputs(7067) <= not b;
    outputs(7068) <= a xor b;
    outputs(7069) <= not (a xor b);
    outputs(7070) <= not (a and b);
    outputs(7071) <= b;
    outputs(7072) <= a;
    outputs(7073) <= not b;
    outputs(7074) <= not (a or b);
    outputs(7075) <= a xor b;
    outputs(7076) <= b;
    outputs(7077) <= not b;
    outputs(7078) <= b and not a;
    outputs(7079) <= a xor b;
    outputs(7080) <= not (a or b);
    outputs(7081) <= b;
    outputs(7082) <= a;
    outputs(7083) <= a xor b;
    outputs(7084) <= not (a or b);
    outputs(7085) <= not (a xor b);
    outputs(7086) <= not a;
    outputs(7087) <= not a or b;
    outputs(7088) <= not a;
    outputs(7089) <= a;
    outputs(7090) <= not (a and b);
    outputs(7091) <= a and not b;
    outputs(7092) <= not (a xor b);
    outputs(7093) <= not (a xor b);
    outputs(7094) <= b and not a;
    outputs(7095) <= b;
    outputs(7096) <= not a;
    outputs(7097) <= not b or a;
    outputs(7098) <= a xor b;
    outputs(7099) <= a and not b;
    outputs(7100) <= b;
    outputs(7101) <= not (a xor b);
    outputs(7102) <= not b;
    outputs(7103) <= not a or b;
    outputs(7104) <= a;
    outputs(7105) <= b;
    outputs(7106) <= a and b;
    outputs(7107) <= not (a xor b);
    outputs(7108) <= a and b;
    outputs(7109) <= a;
    outputs(7110) <= a;
    outputs(7111) <= b;
    outputs(7112) <= a and not b;
    outputs(7113) <= not (a xor b);
    outputs(7114) <= not a or b;
    outputs(7115) <= not (a xor b);
    outputs(7116) <= a;
    outputs(7117) <= not (a xor b);
    outputs(7118) <= not (a xor b);
    outputs(7119) <= b;
    outputs(7120) <= not (a and b);
    outputs(7121) <= not b or a;
    outputs(7122) <= not b;
    outputs(7123) <= a and b;
    outputs(7124) <= b;
    outputs(7125) <= not (a xor b);
    outputs(7126) <= not (a xor b);
    outputs(7127) <= a;
    outputs(7128) <= not b;
    outputs(7129) <= a xor b;
    outputs(7130) <= not (a or b);
    outputs(7131) <= b;
    outputs(7132) <= a xor b;
    outputs(7133) <= not (a and b);
    outputs(7134) <= not b;
    outputs(7135) <= a xor b;
    outputs(7136) <= not b;
    outputs(7137) <= not b;
    outputs(7138) <= not b;
    outputs(7139) <= not a or b;
    outputs(7140) <= not a;
    outputs(7141) <= not (a xor b);
    outputs(7142) <= a xor b;
    outputs(7143) <= b;
    outputs(7144) <= not (a xor b);
    outputs(7145) <= a xor b;
    outputs(7146) <= b;
    outputs(7147) <= not b;
    outputs(7148) <= a;
    outputs(7149) <= a or b;
    outputs(7150) <= a xor b;
    outputs(7151) <= a and b;
    outputs(7152) <= a;
    outputs(7153) <= not a;
    outputs(7154) <= not a or b;
    outputs(7155) <= a xor b;
    outputs(7156) <= a;
    outputs(7157) <= not b or a;
    outputs(7158) <= not a;
    outputs(7159) <= not a;
    outputs(7160) <= a;
    outputs(7161) <= a and not b;
    outputs(7162) <= not a;
    outputs(7163) <= b;
    outputs(7164) <= not b;
    outputs(7165) <= b;
    outputs(7166) <= a;
    outputs(7167) <= b;
    outputs(7168) <= a xor b;
    outputs(7169) <= not b;
    outputs(7170) <= not b;
    outputs(7171) <= not b;
    outputs(7172) <= not (a and b);
    outputs(7173) <= not a;
    outputs(7174) <= b;
    outputs(7175) <= not a;
    outputs(7176) <= a xor b;
    outputs(7177) <= a or b;
    outputs(7178) <= b;
    outputs(7179) <= b and not a;
    outputs(7180) <= not b;
    outputs(7181) <= a;
    outputs(7182) <= a and b;
    outputs(7183) <= a and not b;
    outputs(7184) <= b;
    outputs(7185) <= a and not b;
    outputs(7186) <= a or b;
    outputs(7187) <= b;
    outputs(7188) <= a and b;
    outputs(7189) <= not b;
    outputs(7190) <= not (a xor b);
    outputs(7191) <= not a;
    outputs(7192) <= a and b;
    outputs(7193) <= not a;
    outputs(7194) <= b;
    outputs(7195) <= not a;
    outputs(7196) <= not b;
    outputs(7197) <= not (a xor b);
    outputs(7198) <= not (a xor b);
    outputs(7199) <= not (a xor b);
    outputs(7200) <= a;
    outputs(7201) <= not b;
    outputs(7202) <= a;
    outputs(7203) <= not b;
    outputs(7204) <= not a;
    outputs(7205) <= not b;
    outputs(7206) <= b and not a;
    outputs(7207) <= not (a xor b);
    outputs(7208) <= not a;
    outputs(7209) <= a xor b;
    outputs(7210) <= a and not b;
    outputs(7211) <= not (a and b);
    outputs(7212) <= a xor b;
    outputs(7213) <= a;
    outputs(7214) <= not b;
    outputs(7215) <= not b;
    outputs(7216) <= not (a xor b);
    outputs(7217) <= not (a or b);
    outputs(7218) <= not b;
    outputs(7219) <= a xor b;
    outputs(7220) <= not (a xor b);
    outputs(7221) <= not a;
    outputs(7222) <= not a;
    outputs(7223) <= b and not a;
    outputs(7224) <= a and not b;
    outputs(7225) <= b;
    outputs(7226) <= not (a xor b);
    outputs(7227) <= b;
    outputs(7228) <= a;
    outputs(7229) <= not a or b;
    outputs(7230) <= b and not a;
    outputs(7231) <= a xor b;
    outputs(7232) <= not (a or b);
    outputs(7233) <= a xor b;
    outputs(7234) <= b and not a;
    outputs(7235) <= a;
    outputs(7236) <= b;
    outputs(7237) <= not (a xor b);
    outputs(7238) <= a xor b;
    outputs(7239) <= not (a or b);
    outputs(7240) <= not (a or b);
    outputs(7241) <= not (a xor b);
    outputs(7242) <= a;
    outputs(7243) <= not a;
    outputs(7244) <= a or b;
    outputs(7245) <= a xor b;
    outputs(7246) <= not b;
    outputs(7247) <= not (a xor b);
    outputs(7248) <= b;
    outputs(7249) <= b and not a;
    outputs(7250) <= b;
    outputs(7251) <= not (a xor b);
    outputs(7252) <= not (a xor b);
    outputs(7253) <= not (a and b);
    outputs(7254) <= not b;
    outputs(7255) <= a;
    outputs(7256) <= not (a or b);
    outputs(7257) <= not b;
    outputs(7258) <= a and b;
    outputs(7259) <= a;
    outputs(7260) <= b;
    outputs(7261) <= not (a xor b);
    outputs(7262) <= a and b;
    outputs(7263) <= not a;
    outputs(7264) <= not (a or b);
    outputs(7265) <= a and b;
    outputs(7266) <= b;
    outputs(7267) <= b;
    outputs(7268) <= a and not b;
    outputs(7269) <= not b;
    outputs(7270) <= not a;
    outputs(7271) <= a;
    outputs(7272) <= not a or b;
    outputs(7273) <= not (a or b);
    outputs(7274) <= not a;
    outputs(7275) <= a and not b;
    outputs(7276) <= a xor b;
    outputs(7277) <= a and not b;
    outputs(7278) <= a;
    outputs(7279) <= not (a or b);
    outputs(7280) <= not a;
    outputs(7281) <= not (a xor b);
    outputs(7282) <= a;
    outputs(7283) <= not a;
    outputs(7284) <= not b;
    outputs(7285) <= a;
    outputs(7286) <= b and not a;
    outputs(7287) <= a xor b;
    outputs(7288) <= b;
    outputs(7289) <= b;
    outputs(7290) <= not b;
    outputs(7291) <= not (a xor b);
    outputs(7292) <= b;
    outputs(7293) <= not (a xor b);
    outputs(7294) <= a xor b;
    outputs(7295) <= not (a and b);
    outputs(7296) <= not (a or b);
    outputs(7297) <= a and b;
    outputs(7298) <= b and not a;
    outputs(7299) <= b;
    outputs(7300) <= a xor b;
    outputs(7301) <= not b or a;
    outputs(7302) <= a;
    outputs(7303) <= not (a xor b);
    outputs(7304) <= b and not a;
    outputs(7305) <= not (a xor b);
    outputs(7306) <= not (a xor b);
    outputs(7307) <= not a or b;
    outputs(7308) <= not a;
    outputs(7309) <= not a;
    outputs(7310) <= b;
    outputs(7311) <= not a;
    outputs(7312) <= not b;
    outputs(7313) <= a;
    outputs(7314) <= a xor b;
    outputs(7315) <= b;
    outputs(7316) <= not (a xor b);
    outputs(7317) <= not a;
    outputs(7318) <= not a;
    outputs(7319) <= not a;
    outputs(7320) <= not (a xor b);
    outputs(7321) <= a;
    outputs(7322) <= not (a xor b);
    outputs(7323) <= not b;
    outputs(7324) <= not (a xor b);
    outputs(7325) <= not (a xor b);
    outputs(7326) <= b;
    outputs(7327) <= not a or b;
    outputs(7328) <= a;
    outputs(7329) <= a xor b;
    outputs(7330) <= not a;
    outputs(7331) <= a;
    outputs(7332) <= b;
    outputs(7333) <= a;
    outputs(7334) <= not a or b;
    outputs(7335) <= a and not b;
    outputs(7336) <= not a;
    outputs(7337) <= b;
    outputs(7338) <= a;
    outputs(7339) <= not (a or b);
    outputs(7340) <= b;
    outputs(7341) <= not a;
    outputs(7342) <= a and b;
    outputs(7343) <= b;
    outputs(7344) <= not (a or b);
    outputs(7345) <= b;
    outputs(7346) <= a and b;
    outputs(7347) <= not a;
    outputs(7348) <= a xor b;
    outputs(7349) <= not (a or b);
    outputs(7350) <= not (a xor b);
    outputs(7351) <= b;
    outputs(7352) <= a xor b;
    outputs(7353) <= a xor b;
    outputs(7354) <= a;
    outputs(7355) <= not b;
    outputs(7356) <= b;
    outputs(7357) <= not a or b;
    outputs(7358) <= a xor b;
    outputs(7359) <= a xor b;
    outputs(7360) <= not b or a;
    outputs(7361) <= not (a or b);
    outputs(7362) <= not (a xor b);
    outputs(7363) <= a;
    outputs(7364) <= not b;
    outputs(7365) <= a;
    outputs(7366) <= not b;
    outputs(7367) <= a and b;
    outputs(7368) <= a;
    outputs(7369) <= not b;
    outputs(7370) <= not (a or b);
    outputs(7371) <= not b;
    outputs(7372) <= not (a xor b);
    outputs(7373) <= a xor b;
    outputs(7374) <= not (a or b);
    outputs(7375) <= not a;
    outputs(7376) <= b and not a;
    outputs(7377) <= a and not b;
    outputs(7378) <= a and not b;
    outputs(7379) <= not b;
    outputs(7380) <= a and not b;
    outputs(7381) <= a xor b;
    outputs(7382) <= not (a xor b);
    outputs(7383) <= a xor b;
    outputs(7384) <= not (a and b);
    outputs(7385) <= a and not b;
    outputs(7386) <= a;
    outputs(7387) <= a xor b;
    outputs(7388) <= a;
    outputs(7389) <= a and not b;
    outputs(7390) <= a;
    outputs(7391) <= not b;
    outputs(7392) <= not (a xor b);
    outputs(7393) <= not a;
    outputs(7394) <= b;
    outputs(7395) <= a;
    outputs(7396) <= a xor b;
    outputs(7397) <= a xor b;
    outputs(7398) <= a xor b;
    outputs(7399) <= not (a xor b);
    outputs(7400) <= a;
    outputs(7401) <= not a;
    outputs(7402) <= not (a xor b);
    outputs(7403) <= a xor b;
    outputs(7404) <= a xor b;
    outputs(7405) <= a xor b;
    outputs(7406) <= b;
    outputs(7407) <= a;
    outputs(7408) <= not b;
    outputs(7409) <= not a;
    outputs(7410) <= not a;
    outputs(7411) <= not b;
    outputs(7412) <= not (a xor b);
    outputs(7413) <= not b;
    outputs(7414) <= a and not b;
    outputs(7415) <= not (a or b);
    outputs(7416) <= not a;
    outputs(7417) <= not b;
    outputs(7418) <= a;
    outputs(7419) <= not b;
    outputs(7420) <= not a;
    outputs(7421) <= not (a and b);
    outputs(7422) <= a xor b;
    outputs(7423) <= not a;
    outputs(7424) <= not (a xor b);
    outputs(7425) <= not (a xor b);
    outputs(7426) <= b;
    outputs(7427) <= not (a xor b);
    outputs(7428) <= not b;
    outputs(7429) <= not b;
    outputs(7430) <= not (a or b);
    outputs(7431) <= b;
    outputs(7432) <= not (a xor b);
    outputs(7433) <= a xor b;
    outputs(7434) <= b and not a;
    outputs(7435) <= a or b;
    outputs(7436) <= not b;
    outputs(7437) <= not (a xor b);
    outputs(7438) <= b and not a;
    outputs(7439) <= b;
    outputs(7440) <= b;
    outputs(7441) <= b;
    outputs(7442) <= not b;
    outputs(7443) <= a or b;
    outputs(7444) <= not b;
    outputs(7445) <= not (a or b);
    outputs(7446) <= a or b;
    outputs(7447) <= b;
    outputs(7448) <= not (a xor b);
    outputs(7449) <= not (a or b);
    outputs(7450) <= a and not b;
    outputs(7451) <= b;
    outputs(7452) <= not (a xor b);
    outputs(7453) <= not (a or b);
    outputs(7454) <= a xor b;
    outputs(7455) <= b;
    outputs(7456) <= a and not b;
    outputs(7457) <= not a;
    outputs(7458) <= a and b;
    outputs(7459) <= b and not a;
    outputs(7460) <= not (a xor b);
    outputs(7461) <= not b or a;
    outputs(7462) <= not b;
    outputs(7463) <= not a;
    outputs(7464) <= a;
    outputs(7465) <= not (a xor b);
    outputs(7466) <= a;
    outputs(7467) <= not a;
    outputs(7468) <= not (a xor b);
    outputs(7469) <= not b;
    outputs(7470) <= a xor b;
    outputs(7471) <= not b;
    outputs(7472) <= not (a and b);
    outputs(7473) <= not b;
    outputs(7474) <= a;
    outputs(7475) <= a;
    outputs(7476) <= b;
    outputs(7477) <= a xor b;
    outputs(7478) <= a and b;
    outputs(7479) <= not (a xor b);
    outputs(7480) <= not b;
    outputs(7481) <= not (a or b);
    outputs(7482) <= a;
    outputs(7483) <= not a;
    outputs(7484) <= a and not b;
    outputs(7485) <= not (a or b);
    outputs(7486) <= a and not b;
    outputs(7487) <= a or b;
    outputs(7488) <= not (a xor b);
    outputs(7489) <= b and not a;
    outputs(7490) <= not (a and b);
    outputs(7491) <= not (a or b);
    outputs(7492) <= a xor b;
    outputs(7493) <= not a;
    outputs(7494) <= a;
    outputs(7495) <= not a;
    outputs(7496) <= a and b;
    outputs(7497) <= a;
    outputs(7498) <= b;
    outputs(7499) <= not (a xor b);
    outputs(7500) <= a xor b;
    outputs(7501) <= b;
    outputs(7502) <= not (a xor b);
    outputs(7503) <= not (a xor b);
    outputs(7504) <= b;
    outputs(7505) <= b and not a;
    outputs(7506) <= a xor b;
    outputs(7507) <= a and b;
    outputs(7508) <= b;
    outputs(7509) <= not b;
    outputs(7510) <= a xor b;
    outputs(7511) <= a xor b;
    outputs(7512) <= not (a xor b);
    outputs(7513) <= a xor b;
    outputs(7514) <= a or b;
    outputs(7515) <= b;
    outputs(7516) <= a;
    outputs(7517) <= a xor b;
    outputs(7518) <= a and b;
    outputs(7519) <= not a;
    outputs(7520) <= b and not a;
    outputs(7521) <= a and not b;
    outputs(7522) <= not b;
    outputs(7523) <= not a or b;
    outputs(7524) <= not (a xor b);
    outputs(7525) <= not a;
    outputs(7526) <= not a;
    outputs(7527) <= not (a or b);
    outputs(7528) <= a xor b;
    outputs(7529) <= not (a xor b);
    outputs(7530) <= a xor b;
    outputs(7531) <= not a;
    outputs(7532) <= not (a xor b);
    outputs(7533) <= not (a and b);
    outputs(7534) <= not (a xor b);
    outputs(7535) <= not b;
    outputs(7536) <= not b;
    outputs(7537) <= b;
    outputs(7538) <= a;
    outputs(7539) <= a xor b;
    outputs(7540) <= a xor b;
    outputs(7541) <= a;
    outputs(7542) <= a;
    outputs(7543) <= a xor b;
    outputs(7544) <= a xor b;
    outputs(7545) <= not (a or b);
    outputs(7546) <= a xor b;
    outputs(7547) <= a xor b;
    outputs(7548) <= b;
    outputs(7549) <= a xor b;
    outputs(7550) <= a and not b;
    outputs(7551) <= b and not a;
    outputs(7552) <= b;
    outputs(7553) <= a xor b;
    outputs(7554) <= not b;
    outputs(7555) <= not (a xor b);
    outputs(7556) <= not b;
    outputs(7557) <= a and not b;
    outputs(7558) <= a and not b;
    outputs(7559) <= a xor b;
    outputs(7560) <= a and b;
    outputs(7561) <= a;
    outputs(7562) <= not b or a;
    outputs(7563) <= a;
    outputs(7564) <= not (a or b);
    outputs(7565) <= b;
    outputs(7566) <= not b;
    outputs(7567) <= not a;
    outputs(7568) <= not a;
    outputs(7569) <= not a;
    outputs(7570) <= not b or a;
    outputs(7571) <= a xor b;
    outputs(7572) <= b and not a;
    outputs(7573) <= not (a xor b);
    outputs(7574) <= b and not a;
    outputs(7575) <= a;
    outputs(7576) <= a xor b;
    outputs(7577) <= not (a xor b);
    outputs(7578) <= a;
    outputs(7579) <= not (a xor b);
    outputs(7580) <= a xor b;
    outputs(7581) <= not a;
    outputs(7582) <= b and not a;
    outputs(7583) <= not b;
    outputs(7584) <= b and not a;
    outputs(7585) <= a xor b;
    outputs(7586) <= a xor b;
    outputs(7587) <= b and not a;
    outputs(7588) <= b;
    outputs(7589) <= b and not a;
    outputs(7590) <= not (a and b);
    outputs(7591) <= not a;
    outputs(7592) <= not (a xor b);
    outputs(7593) <= not (a xor b);
    outputs(7594) <= not a;
    outputs(7595) <= not a;
    outputs(7596) <= 1'b1;
    outputs(7597) <= a xor b;
    outputs(7598) <= a and b;
    outputs(7599) <= not (a xor b);
    outputs(7600) <= not a;
    outputs(7601) <= not b;
    outputs(7602) <= not b;
    outputs(7603) <= not a;
    outputs(7604) <= not (a xor b);
    outputs(7605) <= not a;
    outputs(7606) <= a;
    outputs(7607) <= not b;
    outputs(7608) <= not (a xor b);
    outputs(7609) <= a;
    outputs(7610) <= not b;
    outputs(7611) <= not b or a;
    outputs(7612) <= b and not a;
    outputs(7613) <= b;
    outputs(7614) <= not (a or b);
    outputs(7615) <= not (a xor b);
    outputs(7616) <= b;
    outputs(7617) <= not (a xor b);
    outputs(7618) <= not b;
    outputs(7619) <= a xor b;
    outputs(7620) <= a and not b;
    outputs(7621) <= not a;
    outputs(7622) <= a xor b;
    outputs(7623) <= not b;
    outputs(7624) <= not (a or b);
    outputs(7625) <= not (a xor b);
    outputs(7626) <= not a;
    outputs(7627) <= a xor b;
    outputs(7628) <= not a;
    outputs(7629) <= a;
    outputs(7630) <= a xor b;
    outputs(7631) <= not b or a;
    outputs(7632) <= not (a xor b);
    outputs(7633) <= a xor b;
    outputs(7634) <= not (a xor b);
    outputs(7635) <= not (a xor b);
    outputs(7636) <= a xor b;
    outputs(7637) <= a;
    outputs(7638) <= not a;
    outputs(7639) <= not b;
    outputs(7640) <= b and not a;
    outputs(7641) <= not a;
    outputs(7642) <= not (a or b);
    outputs(7643) <= a and b;
    outputs(7644) <= not (a or b);
    outputs(7645) <= not b;
    outputs(7646) <= not a;
    outputs(7647) <= not (a xor b);
    outputs(7648) <= a;
    outputs(7649) <= b and not a;
    outputs(7650) <= a xor b;
    outputs(7651) <= not (a or b);
    outputs(7652) <= a xor b;
    outputs(7653) <= not (a xor b);
    outputs(7654) <= a and not b;
    outputs(7655) <= b;
    outputs(7656) <= a xor b;
    outputs(7657) <= not (a xor b);
    outputs(7658) <= not b;
    outputs(7659) <= not (a xor b);
    outputs(7660) <= not (a xor b);
    outputs(7661) <= a xor b;
    outputs(7662) <= a;
    outputs(7663) <= not (a xor b);
    outputs(7664) <= not (a and b);
    outputs(7665) <= not (a xor b);
    outputs(7666) <= not a;
    outputs(7667) <= a xor b;
    outputs(7668) <= a;
    outputs(7669) <= a;
    outputs(7670) <= not (a xor b);
    outputs(7671) <= a xor b;
    outputs(7672) <= b;
    outputs(7673) <= a xor b;
    outputs(7674) <= b and not a;
    outputs(7675) <= b;
    outputs(7676) <= not b;
    outputs(7677) <= not b;
    outputs(7678) <= a xor b;
    outputs(7679) <= a xor b;
    outputs(7680) <= a xor b;
    outputs(7681) <= not a;
    outputs(7682) <= a and not b;
    outputs(7683) <= b;
    outputs(7684) <= b;
    outputs(7685) <= a and not b;
    outputs(7686) <= a and b;
    outputs(7687) <= a xor b;
    outputs(7688) <= a xor b;
    outputs(7689) <= not (a xor b);
    outputs(7690) <= a;
    outputs(7691) <= a xor b;
    outputs(7692) <= not (a xor b);
    outputs(7693) <= not (a xor b);
    outputs(7694) <= a;
    outputs(7695) <= not b;
    outputs(7696) <= b and not a;
    outputs(7697) <= not b;
    outputs(7698) <= a xor b;
    outputs(7699) <= not b or a;
    outputs(7700) <= not a;
    outputs(7701) <= a xor b;
    outputs(7702) <= not b;
    outputs(7703) <= not (a or b);
    outputs(7704) <= b;
    outputs(7705) <= not b;
    outputs(7706) <= not a;
    outputs(7707) <= a xor b;
    outputs(7708) <= a;
    outputs(7709) <= a xor b;
    outputs(7710) <= a and b;
    outputs(7711) <= not (a xor b);
    outputs(7712) <= b and not a;
    outputs(7713) <= b and not a;
    outputs(7714) <= a;
    outputs(7715) <= b;
    outputs(7716) <= b;
    outputs(7717) <= a and not b;
    outputs(7718) <= not (a xor b);
    outputs(7719) <= not (a xor b);
    outputs(7720) <= a and b;
    outputs(7721) <= a and b;
    outputs(7722) <= a;
    outputs(7723) <= a or b;
    outputs(7724) <= a xor b;
    outputs(7725) <= not (a xor b);
    outputs(7726) <= a and b;
    outputs(7727) <= b;
    outputs(7728) <= not (a xor b);
    outputs(7729) <= a xor b;
    outputs(7730) <= not b;
    outputs(7731) <= a and b;
    outputs(7732) <= a;
    outputs(7733) <= a xor b;
    outputs(7734) <= not b or a;
    outputs(7735) <= not b;
    outputs(7736) <= not (a or b);
    outputs(7737) <= not a;
    outputs(7738) <= not (a xor b);
    outputs(7739) <= not b;
    outputs(7740) <= a;
    outputs(7741) <= not b or a;
    outputs(7742) <= not a;
    outputs(7743) <= not b;
    outputs(7744) <= not (a or b);
    outputs(7745) <= not a;
    outputs(7746) <= not b;
    outputs(7747) <= not b;
    outputs(7748) <= a;
    outputs(7749) <= not a;
    outputs(7750) <= a xor b;
    outputs(7751) <= a and b;
    outputs(7752) <= a xor b;
    outputs(7753) <= a and not b;
    outputs(7754) <= not (a xor b);
    outputs(7755) <= not b or a;
    outputs(7756) <= not (a xor b);
    outputs(7757) <= not (a xor b);
    outputs(7758) <= b;
    outputs(7759) <= a xor b;
    outputs(7760) <= a;
    outputs(7761) <= a;
    outputs(7762) <= not b;
    outputs(7763) <= a and not b;
    outputs(7764) <= b and not a;
    outputs(7765) <= not a;
    outputs(7766) <= a and not b;
    outputs(7767) <= not (a or b);
    outputs(7768) <= not a;
    outputs(7769) <= b;
    outputs(7770) <= b;
    outputs(7771) <= a xor b;
    outputs(7772) <= a;
    outputs(7773) <= a xor b;
    outputs(7774) <= b;
    outputs(7775) <= b;
    outputs(7776) <= a xor b;
    outputs(7777) <= not b;
    outputs(7778) <= a xor b;
    outputs(7779) <= not (a xor b);
    outputs(7780) <= not b;
    outputs(7781) <= not (a xor b);
    outputs(7782) <= a xor b;
    outputs(7783) <= not b;
    outputs(7784) <= not (a xor b);
    outputs(7785) <= not b;
    outputs(7786) <= not b;
    outputs(7787) <= a and b;
    outputs(7788) <= not a;
    outputs(7789) <= not b;
    outputs(7790) <= not (a xor b);
    outputs(7791) <= b;
    outputs(7792) <= a xor b;
    outputs(7793) <= not (a xor b);
    outputs(7794) <= a xor b;
    outputs(7795) <= not b;
    outputs(7796) <= a and not b;
    outputs(7797) <= not a;
    outputs(7798) <= not (a xor b);
    outputs(7799) <= a;
    outputs(7800) <= a and not b;
    outputs(7801) <= not a or b;
    outputs(7802) <= a;
    outputs(7803) <= a;
    outputs(7804) <= b;
    outputs(7805) <= not b;
    outputs(7806) <= a xor b;
    outputs(7807) <= b;
    outputs(7808) <= not a;
    outputs(7809) <= a and b;
    outputs(7810) <= a xor b;
    outputs(7811) <= b;
    outputs(7812) <= b;
    outputs(7813) <= a and not b;
    outputs(7814) <= b;
    outputs(7815) <= b;
    outputs(7816) <= not (a xor b);
    outputs(7817) <= a xor b;
    outputs(7818) <= a and b;
    outputs(7819) <= b;
    outputs(7820) <= b;
    outputs(7821) <= not (a and b);
    outputs(7822) <= not a;
    outputs(7823) <= a;
    outputs(7824) <= not b;
    outputs(7825) <= b and not a;
    outputs(7826) <= not b;
    outputs(7827) <= a xor b;
    outputs(7828) <= a;
    outputs(7829) <= b;
    outputs(7830) <= a xor b;
    outputs(7831) <= b;
    outputs(7832) <= a and not b;
    outputs(7833) <= a xor b;
    outputs(7834) <= b;
    outputs(7835) <= a and b;
    outputs(7836) <= a;
    outputs(7837) <= a xor b;
    outputs(7838) <= not (a xor b);
    outputs(7839) <= a;
    outputs(7840) <= not a;
    outputs(7841) <= not (a and b);
    outputs(7842) <= a xor b;
    outputs(7843) <= a xor b;
    outputs(7844) <= not b;
    outputs(7845) <= b;
    outputs(7846) <= a;
    outputs(7847) <= not b;
    outputs(7848) <= b and not a;
    outputs(7849) <= not a;
    outputs(7850) <= b and not a;
    outputs(7851) <= a;
    outputs(7852) <= not (a xor b);
    outputs(7853) <= a xor b;
    outputs(7854) <= not a;
    outputs(7855) <= not a;
    outputs(7856) <= a xor b;
    outputs(7857) <= a and b;
    outputs(7858) <= a and b;
    outputs(7859) <= not (a xor b);
    outputs(7860) <= not (a or b);
    outputs(7861) <= not a or b;
    outputs(7862) <= not (a xor b);
    outputs(7863) <= not (a xor b);
    outputs(7864) <= a xor b;
    outputs(7865) <= a;
    outputs(7866) <= not (a xor b);
    outputs(7867) <= a xor b;
    outputs(7868) <= not (a xor b);
    outputs(7869) <= b and not a;
    outputs(7870) <= b and not a;
    outputs(7871) <= a;
    outputs(7872) <= b;
    outputs(7873) <= not b;
    outputs(7874) <= a;
    outputs(7875) <= a;
    outputs(7876) <= not (a xor b);
    outputs(7877) <= a xor b;
    outputs(7878) <= not (a xor b);
    outputs(7879) <= not a;
    outputs(7880) <= not a;
    outputs(7881) <= not (a and b);
    outputs(7882) <= a or b;
    outputs(7883) <= not (a xor b);
    outputs(7884) <= a;
    outputs(7885) <= not a or b;
    outputs(7886) <= a;
    outputs(7887) <= not a;
    outputs(7888) <= not b;
    outputs(7889) <= not (a xor b);
    outputs(7890) <= not a;
    outputs(7891) <= not (a xor b);
    outputs(7892) <= a and not b;
    outputs(7893) <= a;
    outputs(7894) <= b and not a;
    outputs(7895) <= a;
    outputs(7896) <= not a;
    outputs(7897) <= not b;
    outputs(7898) <= a and not b;
    outputs(7899) <= b and not a;
    outputs(7900) <= a;
    outputs(7901) <= not (a or b);
    outputs(7902) <= not a;
    outputs(7903) <= not b;
    outputs(7904) <= not a;
    outputs(7905) <= not (a xor b);
    outputs(7906) <= b and not a;
    outputs(7907) <= not a;
    outputs(7908) <= not (a xor b);
    outputs(7909) <= not a;
    outputs(7910) <= not b;
    outputs(7911) <= a xor b;
    outputs(7912) <= not a;
    outputs(7913) <= not b or a;
    outputs(7914) <= b;
    outputs(7915) <= not b;
    outputs(7916) <= not (a xor b);
    outputs(7917) <= not (a or b);
    outputs(7918) <= a;
    outputs(7919) <= a or b;
    outputs(7920) <= not (a xor b);
    outputs(7921) <= not (a or b);
    outputs(7922) <= b;
    outputs(7923) <= a xor b;
    outputs(7924) <= not b;
    outputs(7925) <= a;
    outputs(7926) <= b;
    outputs(7927) <= a xor b;
    outputs(7928) <= a xor b;
    outputs(7929) <= b;
    outputs(7930) <= b;
    outputs(7931) <= a xor b;
    outputs(7932) <= not b;
    outputs(7933) <= a and b;
    outputs(7934) <= not (a and b);
    outputs(7935) <= not b;
    outputs(7936) <= not a;
    outputs(7937) <= not a;
    outputs(7938) <= not a;
    outputs(7939) <= not b;
    outputs(7940) <= a and not b;
    outputs(7941) <= a xor b;
    outputs(7942) <= not a;
    outputs(7943) <= not (a or b);
    outputs(7944) <= b;
    outputs(7945) <= not (a xor b);
    outputs(7946) <= a and b;
    outputs(7947) <= a xor b;
    outputs(7948) <= not (a xor b);
    outputs(7949) <= b;
    outputs(7950) <= a xor b;
    outputs(7951) <= not (a and b);
    outputs(7952) <= not (a or b);
    outputs(7953) <= b and not a;
    outputs(7954) <= a and not b;
    outputs(7955) <= a;
    outputs(7956) <= a or b;
    outputs(7957) <= not (a xor b);
    outputs(7958) <= a and b;
    outputs(7959) <= not (a or b);
    outputs(7960) <= not (a or b);
    outputs(7961) <= not a;
    outputs(7962) <= a;
    outputs(7963) <= not b;
    outputs(7964) <= not (a or b);
    outputs(7965) <= not b;
    outputs(7966) <= a;
    outputs(7967) <= not b;
    outputs(7968) <= a and b;
    outputs(7969) <= not (a xor b);
    outputs(7970) <= b and not a;
    outputs(7971) <= not (a xor b);
    outputs(7972) <= a and b;
    outputs(7973) <= not a;
    outputs(7974) <= not (a xor b);
    outputs(7975) <= not (a or b);
    outputs(7976) <= a;
    outputs(7977) <= b and not a;
    outputs(7978) <= not b;
    outputs(7979) <= a;
    outputs(7980) <= a xor b;
    outputs(7981) <= a or b;
    outputs(7982) <= not a;
    outputs(7983) <= a xor b;
    outputs(7984) <= b and not a;
    outputs(7985) <= not a;
    outputs(7986) <= not b;
    outputs(7987) <= a;
    outputs(7988) <= a or b;
    outputs(7989) <= not (a xor b);
    outputs(7990) <= not b;
    outputs(7991) <= not b or a;
    outputs(7992) <= a;
    outputs(7993) <= not a;
    outputs(7994) <= not (a xor b);
    outputs(7995) <= a;
    outputs(7996) <= not a;
    outputs(7997) <= a and b;
    outputs(7998) <= not (a and b);
    outputs(7999) <= a;
    outputs(8000) <= not a;
    outputs(8001) <= not a;
    outputs(8002) <= a and b;
    outputs(8003) <= not b;
    outputs(8004) <= not a or b;
    outputs(8005) <= a or b;
    outputs(8006) <= a xor b;
    outputs(8007) <= not (a xor b);
    outputs(8008) <= not a;
    outputs(8009) <= not (a xor b);
    outputs(8010) <= not (a xor b);
    outputs(8011) <= not a or b;
    outputs(8012) <= a xor b;
    outputs(8013) <= a xor b;
    outputs(8014) <= b and not a;
    outputs(8015) <= a;
    outputs(8016) <= a and not b;
    outputs(8017) <= not a;
    outputs(8018) <= not (a and b);
    outputs(8019) <= a;
    outputs(8020) <= a xor b;
    outputs(8021) <= b and not a;
    outputs(8022) <= not (a and b);
    outputs(8023) <= a xor b;
    outputs(8024) <= b and not a;
    outputs(8025) <= not a;
    outputs(8026) <= not (a xor b);
    outputs(8027) <= not (a xor b);
    outputs(8028) <= b;
    outputs(8029) <= not b;
    outputs(8030) <= b;
    outputs(8031) <= not (a xor b);
    outputs(8032) <= not (a xor b);
    outputs(8033) <= a xor b;
    outputs(8034) <= a and not b;
    outputs(8035) <= not a;
    outputs(8036) <= not (a xor b);
    outputs(8037) <= not a;
    outputs(8038) <= not a;
    outputs(8039) <= a xor b;
    outputs(8040) <= a xor b;
    outputs(8041) <= not a;
    outputs(8042) <= not a;
    outputs(8043) <= not a;
    outputs(8044) <= not (a xor b);
    outputs(8045) <= not (a xor b);
    outputs(8046) <= a xor b;
    outputs(8047) <= b;
    outputs(8048) <= not (a xor b);
    outputs(8049) <= not (a xor b);
    outputs(8050) <= not (a xor b);
    outputs(8051) <= not b;
    outputs(8052) <= not (a xor b);
    outputs(8053) <= b;
    outputs(8054) <= a;
    outputs(8055) <= not (a and b);
    outputs(8056) <= a xor b;
    outputs(8057) <= not a;
    outputs(8058) <= not a;
    outputs(8059) <= a;
    outputs(8060) <= not b;
    outputs(8061) <= not a;
    outputs(8062) <= b and not a;
    outputs(8063) <= not (a xor b);
    outputs(8064) <= a;
    outputs(8065) <= not (a xor b);
    outputs(8066) <= a;
    outputs(8067) <= a;
    outputs(8068) <= not (a xor b);
    outputs(8069) <= not a;
    outputs(8070) <= not (a and b);
    outputs(8071) <= not a;
    outputs(8072) <= not (a xor b);
    outputs(8073) <= not a;
    outputs(8074) <= not b;
    outputs(8075) <= b;
    outputs(8076) <= a xor b;
    outputs(8077) <= not b;
    outputs(8078) <= not a;
    outputs(8079) <= a;
    outputs(8080) <= not (a xor b);
    outputs(8081) <= a xor b;
    outputs(8082) <= b;
    outputs(8083) <= b;
    outputs(8084) <= not b;
    outputs(8085) <= not b;
    outputs(8086) <= not b;
    outputs(8087) <= not a;
    outputs(8088) <= a xor b;
    outputs(8089) <= a and not b;
    outputs(8090) <= a;
    outputs(8091) <= a xor b;
    outputs(8092) <= b and not a;
    outputs(8093) <= b and not a;
    outputs(8094) <= a xor b;
    outputs(8095) <= a and not b;
    outputs(8096) <= not b;
    outputs(8097) <= not (a xor b);
    outputs(8098) <= b;
    outputs(8099) <= b and not a;
    outputs(8100) <= not (a xor b);
    outputs(8101) <= not b;
    outputs(8102) <= a and b;
    outputs(8103) <= not b or a;
    outputs(8104) <= not (a xor b);
    outputs(8105) <= not (a and b);
    outputs(8106) <= not b;
    outputs(8107) <= not a;
    outputs(8108) <= not a;
    outputs(8109) <= not (a xor b);
    outputs(8110) <= a;
    outputs(8111) <= not a;
    outputs(8112) <= not b;
    outputs(8113) <= b;
    outputs(8114) <= a;
    outputs(8115) <= not b;
    outputs(8116) <= a;
    outputs(8117) <= a;
    outputs(8118) <= not a;
    outputs(8119) <= b;
    outputs(8120) <= a;
    outputs(8121) <= b;
    outputs(8122) <= not (a xor b);
    outputs(8123) <= b and not a;
    outputs(8124) <= a or b;
    outputs(8125) <= a;
    outputs(8126) <= b;
    outputs(8127) <= a and not b;
    outputs(8128) <= not a;
    outputs(8129) <= b;
    outputs(8130) <= a and not b;
    outputs(8131) <= a and not b;
    outputs(8132) <= a and not b;
    outputs(8133) <= not b;
    outputs(8134) <= a;
    outputs(8135) <= not (a xor b);
    outputs(8136) <= not a;
    outputs(8137) <= not (a or b);
    outputs(8138) <= a;
    outputs(8139) <= b and not a;
    outputs(8140) <= not b;
    outputs(8141) <= not (a xor b);
    outputs(8142) <= b and not a;
    outputs(8143) <= a;
    outputs(8144) <= b;
    outputs(8145) <= a;
    outputs(8146) <= not a;
    outputs(8147) <= a and b;
    outputs(8148) <= b and not a;
    outputs(8149) <= not b;
    outputs(8150) <= not (a xor b);
    outputs(8151) <= b;
    outputs(8152) <= not b;
    outputs(8153) <= a xor b;
    outputs(8154) <= not (a and b);
    outputs(8155) <= b;
    outputs(8156) <= not a;
    outputs(8157) <= b;
    outputs(8158) <= b;
    outputs(8159) <= b and not a;
    outputs(8160) <= a;
    outputs(8161) <= not a;
    outputs(8162) <= a and b;
    outputs(8163) <= a;
    outputs(8164) <= not a;
    outputs(8165) <= not (a xor b);
    outputs(8166) <= b;
    outputs(8167) <= not b or a;
    outputs(8168) <= not (a or b);
    outputs(8169) <= not b;
    outputs(8170) <= a or b;
    outputs(8171) <= a and b;
    outputs(8172) <= not a;
    outputs(8173) <= a and not b;
    outputs(8174) <= b and not a;
    outputs(8175) <= not b;
    outputs(8176) <= b;
    outputs(8177) <= not a;
    outputs(8178) <= not (a xor b);
    outputs(8179) <= not (a xor b);
    outputs(8180) <= not a;
    outputs(8181) <= not a;
    outputs(8182) <= not a or b;
    outputs(8183) <= a xor b;
    outputs(8184) <= a or b;
    outputs(8185) <= not a;
    outputs(8186) <= b;
    outputs(8187) <= a xor b;
    outputs(8188) <= a or b;
    outputs(8189) <= not b;
    outputs(8190) <= a;
    outputs(8191) <= a xor b;
    outputs(8192) <= not a;
    outputs(8193) <= not (a xor b);
    outputs(8194) <= a xor b;
    outputs(8195) <= b;
    outputs(8196) <= b;
    outputs(8197) <= not (a xor b);
    outputs(8198) <= not a;
    outputs(8199) <= a;
    outputs(8200) <= not a;
    outputs(8201) <= a xor b;
    outputs(8202) <= not b or a;
    outputs(8203) <= a;
    outputs(8204) <= not b;
    outputs(8205) <= not b or a;
    outputs(8206) <= b;
    outputs(8207) <= b;
    outputs(8208) <= not b or a;
    outputs(8209) <= not (a or b);
    outputs(8210) <= not (a xor b);
    outputs(8211) <= a xor b;
    outputs(8212) <= not (a xor b);
    outputs(8213) <= not a or b;
    outputs(8214) <= a;
    outputs(8215) <= not (a xor b);
    outputs(8216) <= a;
    outputs(8217) <= b;
    outputs(8218) <= b;
    outputs(8219) <= not (a xor b);
    outputs(8220) <= not (a xor b);
    outputs(8221) <= not b;
    outputs(8222) <= not a;
    outputs(8223) <= a xor b;
    outputs(8224) <= not (a xor b);
    outputs(8225) <= a and b;
    outputs(8226) <= not (a xor b);
    outputs(8227) <= a xor b;
    outputs(8228) <= a xor b;
    outputs(8229) <= not a;
    outputs(8230) <= a xor b;
    outputs(8231) <= not (a and b);
    outputs(8232) <= b;
    outputs(8233) <= not b;
    outputs(8234) <= a xor b;
    outputs(8235) <= b;
    outputs(8236) <= a;
    outputs(8237) <= b;
    outputs(8238) <= not (a or b);
    outputs(8239) <= not (a or b);
    outputs(8240) <= not b;
    outputs(8241) <= a and not b;
    outputs(8242) <= not a or b;
    outputs(8243) <= not a;
    outputs(8244) <= b;
    outputs(8245) <= not b;
    outputs(8246) <= b;
    outputs(8247) <= not a;
    outputs(8248) <= a;
    outputs(8249) <= not b or a;
    outputs(8250) <= a and not b;
    outputs(8251) <= a;
    outputs(8252) <= not a;
    outputs(8253) <= not (a xor b);
    outputs(8254) <= a xor b;
    outputs(8255) <= b;
    outputs(8256) <= not a;
    outputs(8257) <= a xor b;
    outputs(8258) <= a or b;
    outputs(8259) <= not (a xor b);
    outputs(8260) <= not (a xor b);
    outputs(8261) <= not (a or b);
    outputs(8262) <= a and not b;
    outputs(8263) <= not b;
    outputs(8264) <= not b;
    outputs(8265) <= a xor b;
    outputs(8266) <= not (a xor b);
    outputs(8267) <= not (a xor b);
    outputs(8268) <= a xor b;
    outputs(8269) <= not a;
    outputs(8270) <= a;
    outputs(8271) <= not a;
    outputs(8272) <= not a;
    outputs(8273) <= not b or a;
    outputs(8274) <= a or b;
    outputs(8275) <= not (a xor b);
    outputs(8276) <= a xor b;
    outputs(8277) <= not (a xor b);
    outputs(8278) <= a and not b;
    outputs(8279) <= a;
    outputs(8280) <= not (a xor b);
    outputs(8281) <= a xor b;
    outputs(8282) <= not (a xor b);
    outputs(8283) <= not a;
    outputs(8284) <= a and not b;
    outputs(8285) <= not b;
    outputs(8286) <= b;
    outputs(8287) <= a xor b;
    outputs(8288) <= not a;
    outputs(8289) <= not a;
    outputs(8290) <= b;
    outputs(8291) <= a and not b;
    outputs(8292) <= a;
    outputs(8293) <= not a;
    outputs(8294) <= not a;
    outputs(8295) <= a;
    outputs(8296) <= not b;
    outputs(8297) <= a or b;
    outputs(8298) <= a and not b;
    outputs(8299) <= not (a xor b);
    outputs(8300) <= not (a xor b);
    outputs(8301) <= a;
    outputs(8302) <= b and not a;
    outputs(8303) <= not b;
    outputs(8304) <= not b;
    outputs(8305) <= a and b;
    outputs(8306) <= b;
    outputs(8307) <= not a;
    outputs(8308) <= not b;
    outputs(8309) <= not b;
    outputs(8310) <= b;
    outputs(8311) <= b;
    outputs(8312) <= not (a xor b);
    outputs(8313) <= not b;
    outputs(8314) <= a;
    outputs(8315) <= not b;
    outputs(8316) <= a xor b;
    outputs(8317) <= b;
    outputs(8318) <= not (a xor b);
    outputs(8319) <= not (a xor b);
    outputs(8320) <= a or b;
    outputs(8321) <= a and b;
    outputs(8322) <= not a;
    outputs(8323) <= not b or a;
    outputs(8324) <= b;
    outputs(8325) <= not (a xor b);
    outputs(8326) <= b;
    outputs(8327) <= b and not a;
    outputs(8328) <= not a;
    outputs(8329) <= a;
    outputs(8330) <= a xor b;
    outputs(8331) <= not (a xor b);
    outputs(8332) <= a or b;
    outputs(8333) <= not (a xor b);
    outputs(8334) <= not a or b;
    outputs(8335) <= not (a xor b);
    outputs(8336) <= not (a xor b);
    outputs(8337) <= not a or b;
    outputs(8338) <= a or b;
    outputs(8339) <= not a;
    outputs(8340) <= not b;
    outputs(8341) <= not (a xor b);
    outputs(8342) <= not a;
    outputs(8343) <= not (a xor b);
    outputs(8344) <= not (a xor b);
    outputs(8345) <= not a;
    outputs(8346) <= a or b;
    outputs(8347) <= b;
    outputs(8348) <= not (a or b);
    outputs(8349) <= b;
    outputs(8350) <= not b;
    outputs(8351) <= not a;
    outputs(8352) <= b;
    outputs(8353) <= not (a xor b);
    outputs(8354) <= not b;
    outputs(8355) <= not b;
    outputs(8356) <= not (a or b);
    outputs(8357) <= a and not b;
    outputs(8358) <= not a or b;
    outputs(8359) <= not b;
    outputs(8360) <= b;
    outputs(8361) <= not a;
    outputs(8362) <= a or b;
    outputs(8363) <= b;
    outputs(8364) <= a;
    outputs(8365) <= not (a xor b);
    outputs(8366) <= a and not b;
    outputs(8367) <= a xor b;
    outputs(8368) <= not a;
    outputs(8369) <= a xor b;
    outputs(8370) <= a or b;
    outputs(8371) <= a and b;
    outputs(8372) <= a xor b;
    outputs(8373) <= not a;
    outputs(8374) <= a xor b;
    outputs(8375) <= not b;
    outputs(8376) <= a xor b;
    outputs(8377) <= not (a xor b);
    outputs(8378) <= not a;
    outputs(8379) <= not (a xor b);
    outputs(8380) <= not (a xor b);
    outputs(8381) <= a or b;
    outputs(8382) <= b;
    outputs(8383) <= not (a xor b);
    outputs(8384) <= b and not a;
    outputs(8385) <= not a or b;
    outputs(8386) <= b;
    outputs(8387) <= a and b;
    outputs(8388) <= not b;
    outputs(8389) <= not b;
    outputs(8390) <= a xor b;
    outputs(8391) <= a xor b;
    outputs(8392) <= a and b;
    outputs(8393) <= a;
    outputs(8394) <= a xor b;
    outputs(8395) <= not a;
    outputs(8396) <= not (a xor b);
    outputs(8397) <= a xor b;
    outputs(8398) <= b;
    outputs(8399) <= not b;
    outputs(8400) <= a or b;
    outputs(8401) <= b;
    outputs(8402) <= a;
    outputs(8403) <= a xor b;
    outputs(8404) <= a;
    outputs(8405) <= a;
    outputs(8406) <= not b or a;
    outputs(8407) <= b;
    outputs(8408) <= a xor b;
    outputs(8409) <= not (a xor b);
    outputs(8410) <= not (a xor b);
    outputs(8411) <= not (a xor b);
    outputs(8412) <= b;
    outputs(8413) <= not b or a;
    outputs(8414) <= a xor b;
    outputs(8415) <= not b;
    outputs(8416) <= a xor b;
    outputs(8417) <= not b;
    outputs(8418) <= not b;
    outputs(8419) <= not (a xor b);
    outputs(8420) <= not a or b;
    outputs(8421) <= not a or b;
    outputs(8422) <= not b;
    outputs(8423) <= not b;
    outputs(8424) <= a xor b;
    outputs(8425) <= not b;
    outputs(8426) <= a xor b;
    outputs(8427) <= not a;
    outputs(8428) <= not (a xor b);
    outputs(8429) <= a xor b;
    outputs(8430) <= not a;
    outputs(8431) <= not b or a;
    outputs(8432) <= not a;
    outputs(8433) <= not b;
    outputs(8434) <= b;
    outputs(8435) <= a xor b;
    outputs(8436) <= not b;
    outputs(8437) <= not (a xor b);
    outputs(8438) <= b;
    outputs(8439) <= a xor b;
    outputs(8440) <= not (a xor b);
    outputs(8441) <= not (a xor b);
    outputs(8442) <= not a or b;
    outputs(8443) <= b;
    outputs(8444) <= not (a xor b);
    outputs(8445) <= not (a xor b);
    outputs(8446) <= not (a xor b);
    outputs(8447) <= not b;
    outputs(8448) <= a xor b;
    outputs(8449) <= a or b;
    outputs(8450) <= not (a xor b);
    outputs(8451) <= a and b;
    outputs(8452) <= not a or b;
    outputs(8453) <= not (a xor b);
    outputs(8454) <= a xor b;
    outputs(8455) <= a xor b;
    outputs(8456) <= not b;
    outputs(8457) <= a;
    outputs(8458) <= not a;
    outputs(8459) <= a or b;
    outputs(8460) <= a;
    outputs(8461) <= a and not b;
    outputs(8462) <= not a;
    outputs(8463) <= not (a or b);
    outputs(8464) <= not a;
    outputs(8465) <= a;
    outputs(8466) <= not a;
    outputs(8467) <= not b;
    outputs(8468) <= b;
    outputs(8469) <= a xor b;
    outputs(8470) <= not (a xor b);
    outputs(8471) <= not (a xor b);
    outputs(8472) <= not b or a;
    outputs(8473) <= not b;
    outputs(8474) <= a or b;
    outputs(8475) <= not a;
    outputs(8476) <= b and not a;
    outputs(8477) <= a;
    outputs(8478) <= not (a xor b);
    outputs(8479) <= not b;
    outputs(8480) <= not a;
    outputs(8481) <= a xor b;
    outputs(8482) <= not b;
    outputs(8483) <= not a;
    outputs(8484) <= not b;
    outputs(8485) <= not (a xor b);
    outputs(8486) <= a xor b;
    outputs(8487) <= a xor b;
    outputs(8488) <= a or b;
    outputs(8489) <= a or b;
    outputs(8490) <= not b or a;
    outputs(8491) <= a xor b;
    outputs(8492) <= a;
    outputs(8493) <= a xor b;
    outputs(8494) <= not a;
    outputs(8495) <= not (a xor b);
    outputs(8496) <= a xor b;
    outputs(8497) <= not b;
    outputs(8498) <= a;
    outputs(8499) <= a;
    outputs(8500) <= a and not b;
    outputs(8501) <= not (a xor b);
    outputs(8502) <= a xor b;
    outputs(8503) <= not (a xor b);
    outputs(8504) <= not b;
    outputs(8505) <= not (a and b);
    outputs(8506) <= a xor b;
    outputs(8507) <= a xor b;
    outputs(8508) <= a xor b;
    outputs(8509) <= not a;
    outputs(8510) <= not (a xor b);
    outputs(8511) <= not a;
    outputs(8512) <= not (a xor b);
    outputs(8513) <= not (a xor b);
    outputs(8514) <= a;
    outputs(8515) <= not b or a;
    outputs(8516) <= not (a xor b);
    outputs(8517) <= not b;
    outputs(8518) <= a xor b;
    outputs(8519) <= not b;
    outputs(8520) <= b;
    outputs(8521) <= a;
    outputs(8522) <= a xor b;
    outputs(8523) <= a;
    outputs(8524) <= not (a xor b);
    outputs(8525) <= not (a xor b);
    outputs(8526) <= b;
    outputs(8527) <= a;
    outputs(8528) <= a xor b;
    outputs(8529) <= a and b;
    outputs(8530) <= not b;
    outputs(8531) <= a xor b;
    outputs(8532) <= a;
    outputs(8533) <= not a or b;
    outputs(8534) <= not a;
    outputs(8535) <= not (a xor b);
    outputs(8536) <= a;
    outputs(8537) <= not b or a;
    outputs(8538) <= a xor b;
    outputs(8539) <= not (a xor b);
    outputs(8540) <= not b;
    outputs(8541) <= not (a xor b);
    outputs(8542) <= not a;
    outputs(8543) <= b;
    outputs(8544) <= a and b;
    outputs(8545) <= not b;
    outputs(8546) <= not b or a;
    outputs(8547) <= b;
    outputs(8548) <= not b;
    outputs(8549) <= not (a xor b);
    outputs(8550) <= b and not a;
    outputs(8551) <= b;
    outputs(8552) <= b;
    outputs(8553) <= b;
    outputs(8554) <= a or b;
    outputs(8555) <= not b or a;
    outputs(8556) <= not b;
    outputs(8557) <= not (a xor b);
    outputs(8558) <= not (a and b);
    outputs(8559) <= not (a or b);
    outputs(8560) <= a or b;
    outputs(8561) <= not b;
    outputs(8562) <= not a or b;
    outputs(8563) <= not b;
    outputs(8564) <= not b;
    outputs(8565) <= a;
    outputs(8566) <= a and b;
    outputs(8567) <= not b or a;
    outputs(8568) <= a;
    outputs(8569) <= not b;
    outputs(8570) <= a;
    outputs(8571) <= not a;
    outputs(8572) <= b and not a;
    outputs(8573) <= a and not b;
    outputs(8574) <= not b;
    outputs(8575) <= a xor b;
    outputs(8576) <= a xor b;
    outputs(8577) <= a xor b;
    outputs(8578) <= b;
    outputs(8579) <= not b;
    outputs(8580) <= not b;
    outputs(8581) <= not a or b;
    outputs(8582) <= not (a xor b);
    outputs(8583) <= b;
    outputs(8584) <= a xor b;
    outputs(8585) <= a;
    outputs(8586) <= not a;
    outputs(8587) <= not b;
    outputs(8588) <= not (a xor b);
    outputs(8589) <= not a or b;
    outputs(8590) <= not (a and b);
    outputs(8591) <= not b or a;
    outputs(8592) <= a and b;
    outputs(8593) <= a or b;
    outputs(8594) <= not (a xor b);
    outputs(8595) <= a and b;
    outputs(8596) <= b;
    outputs(8597) <= a xor b;
    outputs(8598) <= a xor b;
    outputs(8599) <= not (a and b);
    outputs(8600) <= not (a xor b);
    outputs(8601) <= b;
    outputs(8602) <= not (a xor b);
    outputs(8603) <= not a;
    outputs(8604) <= not a or b;
    outputs(8605) <= not (a xor b);
    outputs(8606) <= a xor b;
    outputs(8607) <= not (a xor b);
    outputs(8608) <= b;
    outputs(8609) <= not b;
    outputs(8610) <= a and b;
    outputs(8611) <= not a;
    outputs(8612) <= b and not a;
    outputs(8613) <= not (a xor b);
    outputs(8614) <= not a or b;
    outputs(8615) <= a or b;
    outputs(8616) <= b and not a;
    outputs(8617) <= a;
    outputs(8618) <= a;
    outputs(8619) <= a;
    outputs(8620) <= not (a xor b);
    outputs(8621) <= a xor b;
    outputs(8622) <= not b or a;
    outputs(8623) <= b;
    outputs(8624) <= a xor b;
    outputs(8625) <= not (a xor b);
    outputs(8626) <= not a or b;
    outputs(8627) <= not (a xor b);
    outputs(8628) <= not b;
    outputs(8629) <= not (a or b);
    outputs(8630) <= not (a or b);
    outputs(8631) <= not a;
    outputs(8632) <= a xor b;
    outputs(8633) <= a;
    outputs(8634) <= a xor b;
    outputs(8635) <= not a or b;
    outputs(8636) <= not (a and b);
    outputs(8637) <= not (a and b);
    outputs(8638) <= a;
    outputs(8639) <= b;
    outputs(8640) <= not b;
    outputs(8641) <= b;
    outputs(8642) <= a xor b;
    outputs(8643) <= not (a xor b);
    outputs(8644) <= not (a xor b);
    outputs(8645) <= not a or b;
    outputs(8646) <= b;
    outputs(8647) <= not (a xor b);
    outputs(8648) <= not a or b;
    outputs(8649) <= a xor b;
    outputs(8650) <= a or b;
    outputs(8651) <= a or b;
    outputs(8652) <= not a;
    outputs(8653) <= b;
    outputs(8654) <= a or b;
    outputs(8655) <= a xor b;
    outputs(8656) <= a;
    outputs(8657) <= not (a xor b);
    outputs(8658) <= a xor b;
    outputs(8659) <= not b;
    outputs(8660) <= not a;
    outputs(8661) <= not a;
    outputs(8662) <= not (a xor b);
    outputs(8663) <= a xor b;
    outputs(8664) <= not b;
    outputs(8665) <= not (a xor b);
    outputs(8666) <= a xor b;
    outputs(8667) <= not (a and b);
    outputs(8668) <= not (a xor b);
    outputs(8669) <= a xor b;
    outputs(8670) <= a xor b;
    outputs(8671) <= not (a xor b);
    outputs(8672) <= b;
    outputs(8673) <= b;
    outputs(8674) <= not (a xor b);
    outputs(8675) <= b;
    outputs(8676) <= b;
    outputs(8677) <= a xor b;
    outputs(8678) <= not a or b;
    outputs(8679) <= a;
    outputs(8680) <= a or b;
    outputs(8681) <= a or b;
    outputs(8682) <= a xor b;
    outputs(8683) <= not b;
    outputs(8684) <= not (a xor b);
    outputs(8685) <= not b or a;
    outputs(8686) <= not (a xor b);
    outputs(8687) <= not (a xor b);
    outputs(8688) <= b;
    outputs(8689) <= not (a xor b);
    outputs(8690) <= a;
    outputs(8691) <= a and b;
    outputs(8692) <= not (a and b);
    outputs(8693) <= a xor b;
    outputs(8694) <= not b or a;
    outputs(8695) <= a and not b;
    outputs(8696) <= a xor b;
    outputs(8697) <= b;
    outputs(8698) <= not (a xor b);
    outputs(8699) <= a and b;
    outputs(8700) <= b;
    outputs(8701) <= not b;
    outputs(8702) <= not (a xor b);
    outputs(8703) <= a or b;
    outputs(8704) <= a and not b;
    outputs(8705) <= not (a xor b);
    outputs(8706) <= a xor b;
    outputs(8707) <= b;
    outputs(8708) <= not b;
    outputs(8709) <= a;
    outputs(8710) <= a xor b;
    outputs(8711) <= not (a xor b);
    outputs(8712) <= not b or a;
    outputs(8713) <= not (a xor b);
    outputs(8714) <= not a;
    outputs(8715) <= a and not b;
    outputs(8716) <= a xor b;
    outputs(8717) <= not a;
    outputs(8718) <= not b or a;
    outputs(8719) <= not a;
    outputs(8720) <= not b;
    outputs(8721) <= b;
    outputs(8722) <= not b;
    outputs(8723) <= a and not b;
    outputs(8724) <= b;
    outputs(8725) <= not (a xor b);
    outputs(8726) <= b;
    outputs(8727) <= a xor b;
    outputs(8728) <= a;
    outputs(8729) <= b;
    outputs(8730) <= not a;
    outputs(8731) <= not a or b;
    outputs(8732) <= not a;
    outputs(8733) <= a;
    outputs(8734) <= not b or a;
    outputs(8735) <= not (a and b);
    outputs(8736) <= a xor b;
    outputs(8737) <= a xor b;
    outputs(8738) <= a xor b;
    outputs(8739) <= not b or a;
    outputs(8740) <= b;
    outputs(8741) <= a or b;
    outputs(8742) <= not (a xor b);
    outputs(8743) <= a;
    outputs(8744) <= not b;
    outputs(8745) <= a;
    outputs(8746) <= a and not b;
    outputs(8747) <= b and not a;
    outputs(8748) <= not (a xor b);
    outputs(8749) <= a and b;
    outputs(8750) <= not a or b;
    outputs(8751) <= a xor b;
    outputs(8752) <= a and not b;
    outputs(8753) <= a xor b;
    outputs(8754) <= a and not b;
    outputs(8755) <= not (a xor b);
    outputs(8756) <= b;
    outputs(8757) <= not (a xor b);
    outputs(8758) <= a or b;
    outputs(8759) <= a xor b;
    outputs(8760) <= a or b;
    outputs(8761) <= a;
    outputs(8762) <= a or b;
    outputs(8763) <= a;
    outputs(8764) <= a or b;
    outputs(8765) <= a and b;
    outputs(8766) <= not (a xor b);
    outputs(8767) <= a xor b;
    outputs(8768) <= b;
    outputs(8769) <= not (a xor b);
    outputs(8770) <= not (a xor b);
    outputs(8771) <= not (a xor b);
    outputs(8772) <= a or b;
    outputs(8773) <= not b or a;
    outputs(8774) <= not a;
    outputs(8775) <= a xor b;
    outputs(8776) <= a;
    outputs(8777) <= a xor b;
    outputs(8778) <= not b;
    outputs(8779) <= not a;
    outputs(8780) <= b and not a;
    outputs(8781) <= not (a xor b);
    outputs(8782) <= a xor b;
    outputs(8783) <= not b;
    outputs(8784) <= a and b;
    outputs(8785) <= a xor b;
    outputs(8786) <= a xor b;
    outputs(8787) <= a;
    outputs(8788) <= not b;
    outputs(8789) <= b;
    outputs(8790) <= a xor b;
    outputs(8791) <= not (a xor b);
    outputs(8792) <= a or b;
    outputs(8793) <= a xor b;
    outputs(8794) <= not (a or b);
    outputs(8795) <= a xor b;
    outputs(8796) <= not b;
    outputs(8797) <= a xor b;
    outputs(8798) <= a and not b;
    outputs(8799) <= a xor b;
    outputs(8800) <= not a;
    outputs(8801) <= a xor b;
    outputs(8802) <= not b or a;
    outputs(8803) <= b;
    outputs(8804) <= a;
    outputs(8805) <= not b;
    outputs(8806) <= a xor b;
    outputs(8807) <= a xor b;
    outputs(8808) <= not (a xor b);
    outputs(8809) <= a or b;
    outputs(8810) <= a xor b;
    outputs(8811) <= a xor b;
    outputs(8812) <= a;
    outputs(8813) <= a or b;
    outputs(8814) <= a;
    outputs(8815) <= b;
    outputs(8816) <= a and b;
    outputs(8817) <= b;
    outputs(8818) <= not b;
    outputs(8819) <= a xor b;
    outputs(8820) <= a xor b;
    outputs(8821) <= not a or b;
    outputs(8822) <= not (a xor b);
    outputs(8823) <= a;
    outputs(8824) <= not a;
    outputs(8825) <= a xor b;
    outputs(8826) <= not a;
    outputs(8827) <= a xor b;
    outputs(8828) <= a;
    outputs(8829) <= a;
    outputs(8830) <= not b;
    outputs(8831) <= a or b;
    outputs(8832) <= not b;
    outputs(8833) <= not a or b;
    outputs(8834) <= not b or a;
    outputs(8835) <= not b or a;
    outputs(8836) <= a xor b;
    outputs(8837) <= b and not a;
    outputs(8838) <= not (a and b);
    outputs(8839) <= a xor b;
    outputs(8840) <= a and b;
    outputs(8841) <= not (a and b);
    outputs(8842) <= a xor b;
    outputs(8843) <= b;
    outputs(8844) <= not (a xor b);
    outputs(8845) <= a and not b;
    outputs(8846) <= a xor b;
    outputs(8847) <= not (a xor b);
    outputs(8848) <= a xor b;
    outputs(8849) <= a;
    outputs(8850) <= a;
    outputs(8851) <= a;
    outputs(8852) <= a or b;
    outputs(8853) <= a xor b;
    outputs(8854) <= not b;
    outputs(8855) <= a or b;
    outputs(8856) <= a and b;
    outputs(8857) <= not b;
    outputs(8858) <= not (a or b);
    outputs(8859) <= not (a and b);
    outputs(8860) <= b;
    outputs(8861) <= a xor b;
    outputs(8862) <= b;
    outputs(8863) <= not a;
    outputs(8864) <= not (a xor b);
    outputs(8865) <= not a;
    outputs(8866) <= not b;
    outputs(8867) <= not (a xor b);
    outputs(8868) <= not a;
    outputs(8869) <= not b;
    outputs(8870) <= not (a and b);
    outputs(8871) <= a xor b;
    outputs(8872) <= b and not a;
    outputs(8873) <= b;
    outputs(8874) <= not a or b;
    outputs(8875) <= a and not b;
    outputs(8876) <= a and not b;
    outputs(8877) <= not a;
    outputs(8878) <= not b or a;
    outputs(8879) <= not a;
    outputs(8880) <= a;
    outputs(8881) <= a;
    outputs(8882) <= not a or b;
    outputs(8883) <= not (a xor b);
    outputs(8884) <= a and not b;
    outputs(8885) <= a xor b;
    outputs(8886) <= not (a xor b);
    outputs(8887) <= a xor b;
    outputs(8888) <= not b;
    outputs(8889) <= not b;
    outputs(8890) <= not b;
    outputs(8891) <= not (a xor b);
    outputs(8892) <= b;
    outputs(8893) <= not b or a;
    outputs(8894) <= not (a or b);
    outputs(8895) <= b and not a;
    outputs(8896) <= not a;
    outputs(8897) <= not b;
    outputs(8898) <= not (a or b);
    outputs(8899) <= not (a xor b);
    outputs(8900) <= b;
    outputs(8901) <= not b;
    outputs(8902) <= not (a and b);
    outputs(8903) <= a and b;
    outputs(8904) <= a xor b;
    outputs(8905) <= a xor b;
    outputs(8906) <= a;
    outputs(8907) <= not (a or b);
    outputs(8908) <= a xor b;
    outputs(8909) <= not (a and b);
    outputs(8910) <= not b or a;
    outputs(8911) <= a;
    outputs(8912) <= b;
    outputs(8913) <= a;
    outputs(8914) <= not a;
    outputs(8915) <= b;
    outputs(8916) <= not a;
    outputs(8917) <= a xor b;
    outputs(8918) <= not a or b;
    outputs(8919) <= a or b;
    outputs(8920) <= not a or b;
    outputs(8921) <= not b;
    outputs(8922) <= not b;
    outputs(8923) <= not (a xor b);
    outputs(8924) <= a or b;
    outputs(8925) <= b;
    outputs(8926) <= not b;
    outputs(8927) <= b;
    outputs(8928) <= not a;
    outputs(8929) <= a and not b;
    outputs(8930) <= b;
    outputs(8931) <= a or b;
    outputs(8932) <= not a;
    outputs(8933) <= b;
    outputs(8934) <= not (a and b);
    outputs(8935) <= not (a xor b);
    outputs(8936) <= not b;
    outputs(8937) <= not b;
    outputs(8938) <= a and b;
    outputs(8939) <= not (a xor b);
    outputs(8940) <= not a;
    outputs(8941) <= b;
    outputs(8942) <= b;
    outputs(8943) <= not (a xor b);
    outputs(8944) <= not b;
    outputs(8945) <= b and not a;
    outputs(8946) <= a xor b;
    outputs(8947) <= a;
    outputs(8948) <= b;
    outputs(8949) <= b;
    outputs(8950) <= not b or a;
    outputs(8951) <= not a;
    outputs(8952) <= not b or a;
    outputs(8953) <= b;
    outputs(8954) <= not (a xor b);
    outputs(8955) <= not (a and b);
    outputs(8956) <= b;
    outputs(8957) <= not (a and b);
    outputs(8958) <= not a;
    outputs(8959) <= not b;
    outputs(8960) <= not b or a;
    outputs(8961) <= a and not b;
    outputs(8962) <= a or b;
    outputs(8963) <= b;
    outputs(8964) <= not (a xor b);
    outputs(8965) <= a xor b;
    outputs(8966) <= a and not b;
    outputs(8967) <= a;
    outputs(8968) <= not (a or b);
    outputs(8969) <= a;
    outputs(8970) <= a;
    outputs(8971) <= not a or b;
    outputs(8972) <= a;
    outputs(8973) <= not b or a;
    outputs(8974) <= a;
    outputs(8975) <= not b;
    outputs(8976) <= not (a xor b);
    outputs(8977) <= a xor b;
    outputs(8978) <= b and not a;
    outputs(8979) <= not a or b;
    outputs(8980) <= not (a xor b);
    outputs(8981) <= not a or b;
    outputs(8982) <= a and not b;
    outputs(8983) <= not a;
    outputs(8984) <= not (a xor b);
    outputs(8985) <= b;
    outputs(8986) <= not a;
    outputs(8987) <= a xor b;
    outputs(8988) <= a xor b;
    outputs(8989) <= not a;
    outputs(8990) <= not a;
    outputs(8991) <= not a;
    outputs(8992) <= not (a xor b);
    outputs(8993) <= not (a xor b);
    outputs(8994) <= not a;
    outputs(8995) <= not a;
    outputs(8996) <= not a;
    outputs(8997) <= b;
    outputs(8998) <= not (a xor b);
    outputs(8999) <= b;
    outputs(9000) <= not (a or b);
    outputs(9001) <= a;
    outputs(9002) <= not (a xor b);
    outputs(9003) <= a or b;
    outputs(9004) <= not (a xor b);
    outputs(9005) <= b;
    outputs(9006) <= a xor b;
    outputs(9007) <= a xor b;
    outputs(9008) <= not (a xor b);
    outputs(9009) <= not b;
    outputs(9010) <= b;
    outputs(9011) <= not (a xor b);
    outputs(9012) <= a;
    outputs(9013) <= not b;
    outputs(9014) <= a xor b;
    outputs(9015) <= not a;
    outputs(9016) <= a xor b;
    outputs(9017) <= not (a xor b);
    outputs(9018) <= not a;
    outputs(9019) <= a and not b;
    outputs(9020) <= not a or b;
    outputs(9021) <= not a;
    outputs(9022) <= not (a xor b);
    outputs(9023) <= b;
    outputs(9024) <= a xor b;
    outputs(9025) <= not b or a;
    outputs(9026) <= b;
    outputs(9027) <= a;
    outputs(9028) <= not a;
    outputs(9029) <= not a or b;
    outputs(9030) <= b;
    outputs(9031) <= not b;
    outputs(9032) <= a;
    outputs(9033) <= a;
    outputs(9034) <= not b;
    outputs(9035) <= not (a xor b);
    outputs(9036) <= b and not a;
    outputs(9037) <= not a or b;
    outputs(9038) <= not (a and b);
    outputs(9039) <= not a or b;
    outputs(9040) <= not a or b;
    outputs(9041) <= a xor b;
    outputs(9042) <= not a;
    outputs(9043) <= not a or b;
    outputs(9044) <= b;
    outputs(9045) <= b;
    outputs(9046) <= not (a xor b);
    outputs(9047) <= a xor b;
    outputs(9048) <= not (a xor b);
    outputs(9049) <= b;
    outputs(9050) <= not (a xor b);
    outputs(9051) <= a xor b;
    outputs(9052) <= not (a and b);
    outputs(9053) <= a and b;
    outputs(9054) <= not b or a;
    outputs(9055) <= a and not b;
    outputs(9056) <= not b or a;
    outputs(9057) <= not b;
    outputs(9058) <= b;
    outputs(9059) <= a xor b;
    outputs(9060) <= a xor b;
    outputs(9061) <= b;
    outputs(9062) <= a;
    outputs(9063) <= not (a xor b);
    outputs(9064) <= not b or a;
    outputs(9065) <= a xor b;
    outputs(9066) <= not a;
    outputs(9067) <= not b;
    outputs(9068) <= not (a or b);
    outputs(9069) <= not a;
    outputs(9070) <= not (a xor b);
    outputs(9071) <= not (a or b);
    outputs(9072) <= a;
    outputs(9073) <= a;
    outputs(9074) <= a;
    outputs(9075) <= not a or b;
    outputs(9076) <= b;
    outputs(9077) <= not (a xor b);
    outputs(9078) <= a;
    outputs(9079) <= not (a or b);
    outputs(9080) <= a;
    outputs(9081) <= a xor b;
    outputs(9082) <= b;
    outputs(9083) <= not a;
    outputs(9084) <= a xor b;
    outputs(9085) <= not b or a;
    outputs(9086) <= b;
    outputs(9087) <= not b;
    outputs(9088) <= a and b;
    outputs(9089) <= not (a xor b);
    outputs(9090) <= not b;
    outputs(9091) <= a xor b;
    outputs(9092) <= not b;
    outputs(9093) <= a xor b;
    outputs(9094) <= a xor b;
    outputs(9095) <= a xor b;
    outputs(9096) <= not a;
    outputs(9097) <= not a or b;
    outputs(9098) <= not b or a;
    outputs(9099) <= a;
    outputs(9100) <= not b or a;
    outputs(9101) <= not (a xor b);
    outputs(9102) <= a xor b;
    outputs(9103) <= a xor b;
    outputs(9104) <= a xor b;
    outputs(9105) <= a and b;
    outputs(9106) <= a xor b;
    outputs(9107) <= not a;
    outputs(9108) <= not a;
    outputs(9109) <= not b;
    outputs(9110) <= not (a xor b);
    outputs(9111) <= not a or b;
    outputs(9112) <= not (a and b);
    outputs(9113) <= a and b;
    outputs(9114) <= a or b;
    outputs(9115) <= a xor b;
    outputs(9116) <= not b or a;
    outputs(9117) <= a;
    outputs(9118) <= not a;
    outputs(9119) <= not (a xor b);
    outputs(9120) <= not (a xor b);
    outputs(9121) <= not b;
    outputs(9122) <= a;
    outputs(9123) <= a xor b;
    outputs(9124) <= a xor b;
    outputs(9125) <= not (a xor b);
    outputs(9126) <= b;
    outputs(9127) <= not a;
    outputs(9128) <= not b or a;
    outputs(9129) <= not a or b;
    outputs(9130) <= not a;
    outputs(9131) <= a xor b;
    outputs(9132) <= not (a and b);
    outputs(9133) <= not (a xor b);
    outputs(9134) <= not (a xor b);
    outputs(9135) <= not b;
    outputs(9136) <= a xor b;
    outputs(9137) <= a;
    outputs(9138) <= a xor b;
    outputs(9139) <= not a;
    outputs(9140) <= not (a and b);
    outputs(9141) <= not (a xor b);
    outputs(9142) <= not a;
    outputs(9143) <= not (a xor b);
    outputs(9144) <= not (a and b);
    outputs(9145) <= not (a xor b);
    outputs(9146) <= not (a xor b);
    outputs(9147) <= b;
    outputs(9148) <= not (a xor b);
    outputs(9149) <= a;
    outputs(9150) <= not (a xor b);
    outputs(9151) <= a and not b;
    outputs(9152) <= a;
    outputs(9153) <= not (a xor b);
    outputs(9154) <= b;
    outputs(9155) <= not (a xor b);
    outputs(9156) <= a;
    outputs(9157) <= a xor b;
    outputs(9158) <= not b;
    outputs(9159) <= a xor b;
    outputs(9160) <= b;
    outputs(9161) <= a and not b;
    outputs(9162) <= a xor b;
    outputs(9163) <= not (a xor b);
    outputs(9164) <= a;
    outputs(9165) <= a;
    outputs(9166) <= not b;
    outputs(9167) <= a xor b;
    outputs(9168) <= not a;
    outputs(9169) <= a;
    outputs(9170) <= not (a xor b);
    outputs(9171) <= b;
    outputs(9172) <= b;
    outputs(9173) <= not (a xor b);
    outputs(9174) <= a;
    outputs(9175) <= a;
    outputs(9176) <= not (a xor b);
    outputs(9177) <= not (a xor b);
    outputs(9178) <= a;
    outputs(9179) <= not b;
    outputs(9180) <= b;
    outputs(9181) <= not (a xor b);
    outputs(9182) <= b;
    outputs(9183) <= not (a xor b);
    outputs(9184) <= not b;
    outputs(9185) <= not b;
    outputs(9186) <= b;
    outputs(9187) <= b;
    outputs(9188) <= not (a xor b);
    outputs(9189) <= a xor b;
    outputs(9190) <= a and not b;
    outputs(9191) <= not b;
    outputs(9192) <= not (a or b);
    outputs(9193) <= a;
    outputs(9194) <= not (a xor b);
    outputs(9195) <= not (a xor b);
    outputs(9196) <= b;
    outputs(9197) <= not (a xor b);
    outputs(9198) <= not a;
    outputs(9199) <= a and not b;
    outputs(9200) <= not b;
    outputs(9201) <= not (a xor b);
    outputs(9202) <= a;
    outputs(9203) <= b;
    outputs(9204) <= not (a xor b);
    outputs(9205) <= not (a xor b);
    outputs(9206) <= not b;
    outputs(9207) <= a;
    outputs(9208) <= a;
    outputs(9209) <= b;
    outputs(9210) <= b and not a;
    outputs(9211) <= not b;
    outputs(9212) <= a xor b;
    outputs(9213) <= not (a xor b);
    outputs(9214) <= b;
    outputs(9215) <= not a;
    outputs(9216) <= not (a xor b);
    outputs(9217) <= a;
    outputs(9218) <= not (a xor b);
    outputs(9219) <= b;
    outputs(9220) <= b and not a;
    outputs(9221) <= a;
    outputs(9222) <= not (a xor b);
    outputs(9223) <= not (a xor b);
    outputs(9224) <= not a;
    outputs(9225) <= a and b;
    outputs(9226) <= a;
    outputs(9227) <= not (a xor b);
    outputs(9228) <= not b;
    outputs(9229) <= not (a xor b);
    outputs(9230) <= not (a xor b);
    outputs(9231) <= not a;
    outputs(9232) <= a;
    outputs(9233) <= b;
    outputs(9234) <= a xor b;
    outputs(9235) <= a and not b;
    outputs(9236) <= b;
    outputs(9237) <= a xor b;
    outputs(9238) <= a and b;
    outputs(9239) <= a xor b;
    outputs(9240) <= a xor b;
    outputs(9241) <= not a;
    outputs(9242) <= a;
    outputs(9243) <= not a;
    outputs(9244) <= b;
    outputs(9245) <= not (a xor b);
    outputs(9246) <= b;
    outputs(9247) <= not (a xor b);
    outputs(9248) <= b;
    outputs(9249) <= a xor b;
    outputs(9250) <= not (a xor b);
    outputs(9251) <= a xor b;
    outputs(9252) <= not (a xor b);
    outputs(9253) <= not (a xor b);
    outputs(9254) <= a and b;
    outputs(9255) <= not b;
    outputs(9256) <= a xor b;
    outputs(9257) <= a;
    outputs(9258) <= a xor b;
    outputs(9259) <= not (a xor b);
    outputs(9260) <= b;
    outputs(9261) <= a;
    outputs(9262) <= not (a xor b);
    outputs(9263) <= a xor b;
    outputs(9264) <= not a;
    outputs(9265) <= not (a xor b);
    outputs(9266) <= a xor b;
    outputs(9267) <= not (a xor b);
    outputs(9268) <= not (a xor b);
    outputs(9269) <= not a;
    outputs(9270) <= not a;
    outputs(9271) <= not (a xor b);
    outputs(9272) <= b;
    outputs(9273) <= b and not a;
    outputs(9274) <= a and not b;
    outputs(9275) <= a;
    outputs(9276) <= not b;
    outputs(9277) <= a;
    outputs(9278) <= a and not b;
    outputs(9279) <= not (a xor b);
    outputs(9280) <= a and not b;
    outputs(9281) <= b and not a;
    outputs(9282) <= a and not b;
    outputs(9283) <= not a;
    outputs(9284) <= a;
    outputs(9285) <= not (a xor b);
    outputs(9286) <= not (a xor b);
    outputs(9287) <= not a;
    outputs(9288) <= not (a xor b);
    outputs(9289) <= a;
    outputs(9290) <= not a;
    outputs(9291) <= b;
    outputs(9292) <= not a;
    outputs(9293) <= a;
    outputs(9294) <= b;
    outputs(9295) <= a xor b;
    outputs(9296) <= a and not b;
    outputs(9297) <= a xor b;
    outputs(9298) <= not b;
    outputs(9299) <= not b;
    outputs(9300) <= a;
    outputs(9301) <= not b;
    outputs(9302) <= not (a xor b);
    outputs(9303) <= not b or a;
    outputs(9304) <= not (a xor b);
    outputs(9305) <= a;
    outputs(9306) <= a;
    outputs(9307) <= not b;
    outputs(9308) <= not b;
    outputs(9309) <= b and not a;
    outputs(9310) <= a xor b;
    outputs(9311) <= a and b;
    outputs(9312) <= b;
    outputs(9313) <= a;
    outputs(9314) <= a and b;
    outputs(9315) <= not (a xor b);
    outputs(9316) <= not b;
    outputs(9317) <= not (a and b);
    outputs(9318) <= not (a xor b);
    outputs(9319) <= 1'b0;
    outputs(9320) <= a xor b;
    outputs(9321) <= a xor b;
    outputs(9322) <= a xor b;
    outputs(9323) <= b and not a;
    outputs(9324) <= not b;
    outputs(9325) <= b;
    outputs(9326) <= not (a and b);
    outputs(9327) <= not (a xor b);
    outputs(9328) <= a;
    outputs(9329) <= a and b;
    outputs(9330) <= not b;
    outputs(9331) <= not b;
    outputs(9332) <= not (a xor b);
    outputs(9333) <= not (a xor b);
    outputs(9334) <= not (a xor b);
    outputs(9335) <= not a;
    outputs(9336) <= not (a xor b);
    outputs(9337) <= b;
    outputs(9338) <= a;
    outputs(9339) <= a xor b;
    outputs(9340) <= not (a xor b);
    outputs(9341) <= not a;
    outputs(9342) <= b;
    outputs(9343) <= b and not a;
    outputs(9344) <= b;
    outputs(9345) <= a xor b;
    outputs(9346) <= a xor b;
    outputs(9347) <= not (a and b);
    outputs(9348) <= not a;
    outputs(9349) <= not (a and b);
    outputs(9350) <= b;
    outputs(9351) <= a xor b;
    outputs(9352) <= a;
    outputs(9353) <= not a;
    outputs(9354) <= not (a xor b);
    outputs(9355) <= not (a or b);
    outputs(9356) <= not b;
    outputs(9357) <= not b;
    outputs(9358) <= a and not b;
    outputs(9359) <= not a;
    outputs(9360) <= b;
    outputs(9361) <= a;
    outputs(9362) <= b and not a;
    outputs(9363) <= not b;
    outputs(9364) <= not b;
    outputs(9365) <= a and b;
    outputs(9366) <= a xor b;
    outputs(9367) <= a and not b;
    outputs(9368) <= not (a xor b);
    outputs(9369) <= not b;
    outputs(9370) <= a xor b;
    outputs(9371) <= a;
    outputs(9372) <= b;
    outputs(9373) <= not a;
    outputs(9374) <= not a;
    outputs(9375) <= a xor b;
    outputs(9376) <= not b;
    outputs(9377) <= b and not a;
    outputs(9378) <= not a or b;
    outputs(9379) <= b;
    outputs(9380) <= not a;
    outputs(9381) <= a xor b;
    outputs(9382) <= not a;
    outputs(9383) <= not (a xor b);
    outputs(9384) <= b;
    outputs(9385) <= not b;
    outputs(9386) <= a xor b;
    outputs(9387) <= b;
    outputs(9388) <= not (a xor b);
    outputs(9389) <= b and not a;
    outputs(9390) <= not (a xor b);
    outputs(9391) <= not b;
    outputs(9392) <= not (a xor b);
    outputs(9393) <= not a;
    outputs(9394) <= a;
    outputs(9395) <= not b;
    outputs(9396) <= b and not a;
    outputs(9397) <= not a;
    outputs(9398) <= a xor b;
    outputs(9399) <= not (a and b);
    outputs(9400) <= not (a or b);
    outputs(9401) <= not a;
    outputs(9402) <= not a;
    outputs(9403) <= not (a or b);
    outputs(9404) <= not b;
    outputs(9405) <= not (a or b);
    outputs(9406) <= not (a xor b);
    outputs(9407) <= not (a xor b);
    outputs(9408) <= a and b;
    outputs(9409) <= not (a xor b);
    outputs(9410) <= not (a or b);
    outputs(9411) <= a;
    outputs(9412) <= not b or a;
    outputs(9413) <= b and not a;
    outputs(9414) <= a xor b;
    outputs(9415) <= not a;
    outputs(9416) <= not a;
    outputs(9417) <= b;
    outputs(9418) <= b;
    outputs(9419) <= not (a xor b);
    outputs(9420) <= a xor b;
    outputs(9421) <= b;
    outputs(9422) <= b and not a;
    outputs(9423) <= a xor b;
    outputs(9424) <= not (a xor b);
    outputs(9425) <= not a;
    outputs(9426) <= b;
    outputs(9427) <= a and b;
    outputs(9428) <= a;
    outputs(9429) <= a xor b;
    outputs(9430) <= not b;
    outputs(9431) <= not (a xor b);
    outputs(9432) <= b;
    outputs(9433) <= b;
    outputs(9434) <= a and b;
    outputs(9435) <= not (a xor b);
    outputs(9436) <= not a;
    outputs(9437) <= a and b;
    outputs(9438) <= a;
    outputs(9439) <= not (a xor b);
    outputs(9440) <= b and not a;
    outputs(9441) <= b;
    outputs(9442) <= b;
    outputs(9443) <= a xor b;
    outputs(9444) <= a xor b;
    outputs(9445) <= not (a or b);
    outputs(9446) <= a and b;
    outputs(9447) <= a and not b;
    outputs(9448) <= not (a or b);
    outputs(9449) <= not (a or b);
    outputs(9450) <= not (a xor b);
    outputs(9451) <= not b;
    outputs(9452) <= a xor b;
    outputs(9453) <= not (a xor b);
    outputs(9454) <= not a or b;
    outputs(9455) <= a;
    outputs(9456) <= a;
    outputs(9457) <= a xor b;
    outputs(9458) <= not b;
    outputs(9459) <= not a;
    outputs(9460) <= not (a xor b);
    outputs(9461) <= b and not a;
    outputs(9462) <= not a;
    outputs(9463) <= a and not b;
    outputs(9464) <= not b;
    outputs(9465) <= not a;
    outputs(9466) <= a;
    outputs(9467) <= a xor b;
    outputs(9468) <= a and b;
    outputs(9469) <= a;
    outputs(9470) <= not a;
    outputs(9471) <= not (a xor b);
    outputs(9472) <= not b;
    outputs(9473) <= not (a xor b);
    outputs(9474) <= a xor b;
    outputs(9475) <= a xor b;
    outputs(9476) <= not (a xor b);
    outputs(9477) <= b;
    outputs(9478) <= a xor b;
    outputs(9479) <= not a;
    outputs(9480) <= b and not a;
    outputs(9481) <= b and not a;
    outputs(9482) <= not (a xor b);
    outputs(9483) <= not (a xor b);
    outputs(9484) <= a and not b;
    outputs(9485) <= b and not a;
    outputs(9486) <= a xor b;
    outputs(9487) <= a xor b;
    outputs(9488) <= not a;
    outputs(9489) <= not a;
    outputs(9490) <= not b or a;
    outputs(9491) <= a;
    outputs(9492) <= a;
    outputs(9493) <= not a;
    outputs(9494) <= not a;
    outputs(9495) <= not (a and b);
    outputs(9496) <= not a or b;
    outputs(9497) <= not (a xor b);
    outputs(9498) <= not b;
    outputs(9499) <= not (a or b);
    outputs(9500) <= a and not b;
    outputs(9501) <= not (a xor b);
    outputs(9502) <= a;
    outputs(9503) <= a xor b;
    outputs(9504) <= b and not a;
    outputs(9505) <= not a;
    outputs(9506) <= 1'b1;
    outputs(9507) <= a;
    outputs(9508) <= not (a xor b);
    outputs(9509) <= not (a xor b);
    outputs(9510) <= not a;
    outputs(9511) <= a and b;
    outputs(9512) <= a;
    outputs(9513) <= not (a xor b);
    outputs(9514) <= not (a xor b);
    outputs(9515) <= a xor b;
    outputs(9516) <= a xor b;
    outputs(9517) <= a xor b;
    outputs(9518) <= a;
    outputs(9519) <= a;
    outputs(9520) <= a and not b;
    outputs(9521) <= a;
    outputs(9522) <= a and b;
    outputs(9523) <= not b;
    outputs(9524) <= b;
    outputs(9525) <= a xor b;
    outputs(9526) <= not (a or b);
    outputs(9527) <= a xor b;
    outputs(9528) <= not (a xor b);
    outputs(9529) <= a xor b;
    outputs(9530) <= a;
    outputs(9531) <= not (a or b);
    outputs(9532) <= a;
    outputs(9533) <= not (a xor b);
    outputs(9534) <= a;
    outputs(9535) <= a xor b;
    outputs(9536) <= not b;
    outputs(9537) <= a or b;
    outputs(9538) <= not (a and b);
    outputs(9539) <= a and not b;
    outputs(9540) <= a xor b;
    outputs(9541) <= not b;
    outputs(9542) <= a xor b;
    outputs(9543) <= a xor b;
    outputs(9544) <= a and not b;
    outputs(9545) <= not b or a;
    outputs(9546) <= b and not a;
    outputs(9547) <= not b;
    outputs(9548) <= not b;
    outputs(9549) <= a xor b;
    outputs(9550) <= b;
    outputs(9551) <= not (a xor b);
    outputs(9552) <= a;
    outputs(9553) <= not b;
    outputs(9554) <= not (a xor b);
    outputs(9555) <= not (a xor b);
    outputs(9556) <= a xor b;
    outputs(9557) <= a;
    outputs(9558) <= not (a xor b);
    outputs(9559) <= not (a xor b);
    outputs(9560) <= a xor b;
    outputs(9561) <= not (a xor b);
    outputs(9562) <= not b;
    outputs(9563) <= not b;
    outputs(9564) <= a xor b;
    outputs(9565) <= a xor b;
    outputs(9566) <= not a;
    outputs(9567) <= a xor b;
    outputs(9568) <= b;
    outputs(9569) <= a xor b;
    outputs(9570) <= not a;
    outputs(9571) <= a;
    outputs(9572) <= b;
    outputs(9573) <= not a;
    outputs(9574) <= a xor b;
    outputs(9575) <= a;
    outputs(9576) <= a;
    outputs(9577) <= b and not a;
    outputs(9578) <= a;
    outputs(9579) <= a or b;
    outputs(9580) <= not a;
    outputs(9581) <= not (a xor b);
    outputs(9582) <= not (a or b);
    outputs(9583) <= not b;
    outputs(9584) <= a;
    outputs(9585) <= b;
    outputs(9586) <= not a;
    outputs(9587) <= not (a xor b);
    outputs(9588) <= a;
    outputs(9589) <= a or b;
    outputs(9590) <= not (a xor b);
    outputs(9591) <= a xor b;
    outputs(9592) <= a xor b;
    outputs(9593) <= not b;
    outputs(9594) <= not a or b;
    outputs(9595) <= a and b;
    outputs(9596) <= not b;
    outputs(9597) <= a;
    outputs(9598) <= b;
    outputs(9599) <= not (a or b);
    outputs(9600) <= a;
    outputs(9601) <= b;
    outputs(9602) <= not a;
    outputs(9603) <= a;
    outputs(9604) <= not (a xor b);
    outputs(9605) <= not (a xor b);
    outputs(9606) <= a;
    outputs(9607) <= not a;
    outputs(9608) <= a xor b;
    outputs(9609) <= b;
    outputs(9610) <= not a;
    outputs(9611) <= a xor b;
    outputs(9612) <= not a;
    outputs(9613) <= b;
    outputs(9614) <= a and not b;
    outputs(9615) <= not a;
    outputs(9616) <= a xor b;
    outputs(9617) <= a xor b;
    outputs(9618) <= a xor b;
    outputs(9619) <= a and not b;
    outputs(9620) <= a xor b;
    outputs(9621) <= a xor b;
    outputs(9622) <= a and not b;
    outputs(9623) <= a and b;
    outputs(9624) <= not b;
    outputs(9625) <= not b;
    outputs(9626) <= not (a and b);
    outputs(9627) <= b;
    outputs(9628) <= a xor b;
    outputs(9629) <= not (a or b);
    outputs(9630) <= not a;
    outputs(9631) <= not (a xor b);
    outputs(9632) <= not (a xor b);
    outputs(9633) <= b;
    outputs(9634) <= a or b;
    outputs(9635) <= not (a xor b);
    outputs(9636) <= not (a and b);
    outputs(9637) <= b and not a;
    outputs(9638) <= not (a xor b);
    outputs(9639) <= not a;
    outputs(9640) <= b and not a;
    outputs(9641) <= not a;
    outputs(9642) <= not (a or b);
    outputs(9643) <= a xor b;
    outputs(9644) <= a xor b;
    outputs(9645) <= a;
    outputs(9646) <= a xor b;
    outputs(9647) <= b;
    outputs(9648) <= not (a xor b);
    outputs(9649) <= a xor b;
    outputs(9650) <= a and not b;
    outputs(9651) <= not b;
    outputs(9652) <= a and b;
    outputs(9653) <= a and b;
    outputs(9654) <= a;
    outputs(9655) <= a xor b;
    outputs(9656) <= not (a xor b);
    outputs(9657) <= a;
    outputs(9658) <= a;
    outputs(9659) <= a xor b;
    outputs(9660) <= a xor b;
    outputs(9661) <= not b;
    outputs(9662) <= not a;
    outputs(9663) <= not b;
    outputs(9664) <= a xor b;
    outputs(9665) <= a and b;
    outputs(9666) <= a;
    outputs(9667) <= b;
    outputs(9668) <= a;
    outputs(9669) <= not (a xor b);
    outputs(9670) <= b and not a;
    outputs(9671) <= a and not b;
    outputs(9672) <= a and b;
    outputs(9673) <= 1'b0;
    outputs(9674) <= a and not b;
    outputs(9675) <= not a;
    outputs(9676) <= b;
    outputs(9677) <= b and not a;
    outputs(9678) <= b;
    outputs(9679) <= b;
    outputs(9680) <= a;
    outputs(9681) <= a;
    outputs(9682) <= a and b;
    outputs(9683) <= a and b;
    outputs(9684) <= a xor b;
    outputs(9685) <= not a;
    outputs(9686) <= not (a xor b);
    outputs(9687) <= not b;
    outputs(9688) <= not b;
    outputs(9689) <= a xor b;
    outputs(9690) <= a xor b;
    outputs(9691) <= a;
    outputs(9692) <= b;
    outputs(9693) <= b;
    outputs(9694) <= a xor b;
    outputs(9695) <= a xor b;
    outputs(9696) <= a;
    outputs(9697) <= not (a xor b);
    outputs(9698) <= b;
    outputs(9699) <= not b;
    outputs(9700) <= not b;
    outputs(9701) <= b;
    outputs(9702) <= b;
    outputs(9703) <= not b;
    outputs(9704) <= a;
    outputs(9705) <= a xor b;
    outputs(9706) <= a xor b;
    outputs(9707) <= a;
    outputs(9708) <= a xor b;
    outputs(9709) <= a xor b;
    outputs(9710) <= not b;
    outputs(9711) <= not (a xor b);
    outputs(9712) <= b;
    outputs(9713) <= not (a xor b);
    outputs(9714) <= not a;
    outputs(9715) <= not (a and b);
    outputs(9716) <= not b;
    outputs(9717) <= a;
    outputs(9718) <= a;
    outputs(9719) <= b;
    outputs(9720) <= a xor b;
    outputs(9721) <= not b;
    outputs(9722) <= not (a xor b);
    outputs(9723) <= not a;
    outputs(9724) <= a xor b;
    outputs(9725) <= a and not b;
    outputs(9726) <= not (a xor b);
    outputs(9727) <= a xor b;
    outputs(9728) <= b;
    outputs(9729) <= a xor b;
    outputs(9730) <= a xor b;
    outputs(9731) <= b and not a;
    outputs(9732) <= a xor b;
    outputs(9733) <= b;
    outputs(9734) <= a xor b;
    outputs(9735) <= not a or b;
    outputs(9736) <= a;
    outputs(9737) <= not (a xor b);
    outputs(9738) <= not (a xor b);
    outputs(9739) <= not b;
    outputs(9740) <= b and not a;
    outputs(9741) <= not (a xor b);
    outputs(9742) <= not (a or b);
    outputs(9743) <= a and not b;
    outputs(9744) <= not b or a;
    outputs(9745) <= b;
    outputs(9746) <= a xor b;
    outputs(9747) <= b and not a;
    outputs(9748) <= not (a xor b);
    outputs(9749) <= a;
    outputs(9750) <= not a;
    outputs(9751) <= a;
    outputs(9752) <= not b;
    outputs(9753) <= b;
    outputs(9754) <= not (a xor b);
    outputs(9755) <= a xor b;
    outputs(9756) <= a xor b;
    outputs(9757) <= a and not b;
    outputs(9758) <= not (a xor b);
    outputs(9759) <= not (a xor b);
    outputs(9760) <= a;
    outputs(9761) <= a;
    outputs(9762) <= not (a or b);
    outputs(9763) <= not (a xor b);
    outputs(9764) <= a;
    outputs(9765) <= a xor b;
    outputs(9766) <= not a;
    outputs(9767) <= not a;
    outputs(9768) <= not a;
    outputs(9769) <= not b;
    outputs(9770) <= not a;
    outputs(9771) <= not (a and b);
    outputs(9772) <= b;
    outputs(9773) <= not a;
    outputs(9774) <= b and not a;
    outputs(9775) <= a and not b;
    outputs(9776) <= not b;
    outputs(9777) <= not (a xor b);
    outputs(9778) <= a;
    outputs(9779) <= a xor b;
    outputs(9780) <= b;
    outputs(9781) <= not b;
    outputs(9782) <= not a;
    outputs(9783) <= a xor b;
    outputs(9784) <= not b;
    outputs(9785) <= not b;
    outputs(9786) <= b;
    outputs(9787) <= not a;
    outputs(9788) <= a xor b;
    outputs(9789) <= not (a xor b);
    outputs(9790) <= a;
    outputs(9791) <= not (a or b);
    outputs(9792) <= a and not b;
    outputs(9793) <= not a;
    outputs(9794) <= a xor b;
    outputs(9795) <= not (a xor b);
    outputs(9796) <= a and b;
    outputs(9797) <= a xor b;
    outputs(9798) <= b;
    outputs(9799) <= b;
    outputs(9800) <= not (a and b);
    outputs(9801) <= not b;
    outputs(9802) <= a;
    outputs(9803) <= b;
    outputs(9804) <= not b;
    outputs(9805) <= a;
    outputs(9806) <= a;
    outputs(9807) <= a xor b;
    outputs(9808) <= a or b;
    outputs(9809) <= not (a xor b);
    outputs(9810) <= a xor b;
    outputs(9811) <= a and not b;
    outputs(9812) <= a and b;
    outputs(9813) <= not a;
    outputs(9814) <= not (a xor b);
    outputs(9815) <= b;
    outputs(9816) <= a xor b;
    outputs(9817) <= not b;
    outputs(9818) <= b;
    outputs(9819) <= b;
    outputs(9820) <= not b or a;
    outputs(9821) <= not (a xor b);
    outputs(9822) <= a and b;
    outputs(9823) <= not (a xor b);
    outputs(9824) <= b and not a;
    outputs(9825) <= not (a xor b);
    outputs(9826) <= a and not b;
    outputs(9827) <= b;
    outputs(9828) <= a;
    outputs(9829) <= not a;
    outputs(9830) <= a and not b;
    outputs(9831) <= a and not b;
    outputs(9832) <= b and not a;
    outputs(9833) <= b;
    outputs(9834) <= not a or b;
    outputs(9835) <= not a;
    outputs(9836) <= not (a and b);
    outputs(9837) <= b and not a;
    outputs(9838) <= not (a xor b);
    outputs(9839) <= b;
    outputs(9840) <= not b;
    outputs(9841) <= not (a xor b);
    outputs(9842) <= b;
    outputs(9843) <= a;
    outputs(9844) <= a xor b;
    outputs(9845) <= a;
    outputs(9846) <= not (a xor b);
    outputs(9847) <= a xor b;
    outputs(9848) <= not (a xor b);
    outputs(9849) <= a and not b;
    outputs(9850) <= not a or b;
    outputs(9851) <= a;
    outputs(9852) <= a xor b;
    outputs(9853) <= not (a xor b);
    outputs(9854) <= a;
    outputs(9855) <= b and not a;
    outputs(9856) <= b;
    outputs(9857) <= a xor b;
    outputs(9858) <= b;
    outputs(9859) <= b and not a;
    outputs(9860) <= a;
    outputs(9861) <= a xor b;
    outputs(9862) <= a and not b;
    outputs(9863) <= a xor b;
    outputs(9864) <= a;
    outputs(9865) <= not (a xor b);
    outputs(9866) <= b;
    outputs(9867) <= a xor b;
    outputs(9868) <= b;
    outputs(9869) <= b and not a;
    outputs(9870) <= not (a xor b);
    outputs(9871) <= not (a xor b);
    outputs(9872) <= not a or b;
    outputs(9873) <= a;
    outputs(9874) <= a xor b;
    outputs(9875) <= not b;
    outputs(9876) <= b;
    outputs(9877) <= a;
    outputs(9878) <= b;
    outputs(9879) <= not a;
    outputs(9880) <= b;
    outputs(9881) <= a xor b;
    outputs(9882) <= not b;
    outputs(9883) <= not b;
    outputs(9884) <= a;
    outputs(9885) <= not b or a;
    outputs(9886) <= a and b;
    outputs(9887) <= a;
    outputs(9888) <= a or b;
    outputs(9889) <= not b or a;
    outputs(9890) <= a xor b;
    outputs(9891) <= a and not b;
    outputs(9892) <= not (a xor b);
    outputs(9893) <= not b;
    outputs(9894) <= not a;
    outputs(9895) <= not b;
    outputs(9896) <= a and b;
    outputs(9897) <= not (a or b);
    outputs(9898) <= a xor b;
    outputs(9899) <= b;
    outputs(9900) <= a and not b;
    outputs(9901) <= not b;
    outputs(9902) <= not b;
    outputs(9903) <= a xor b;
    outputs(9904) <= a or b;
    outputs(9905) <= a xor b;
    outputs(9906) <= not a;
    outputs(9907) <= b and not a;
    outputs(9908) <= not (a or b);
    outputs(9909) <= not b or a;
    outputs(9910) <= b;
    outputs(9911) <= b;
    outputs(9912) <= not (a xor b);
    outputs(9913) <= not b;
    outputs(9914) <= a;
    outputs(9915) <= not (a xor b);
    outputs(9916) <= not b;
    outputs(9917) <= b;
    outputs(9918) <= not b;
    outputs(9919) <= a xor b;
    outputs(9920) <= a xor b;
    outputs(9921) <= a xor b;
    outputs(9922) <= not a;
    outputs(9923) <= not (a xor b);
    outputs(9924) <= not b;
    outputs(9925) <= not (a xor b);
    outputs(9926) <= not (a xor b);
    outputs(9927) <= not (a and b);
    outputs(9928) <= not b;
    outputs(9929) <= a and not b;
    outputs(9930) <= a xor b;
    outputs(9931) <= a xor b;
    outputs(9932) <= not (a or b);
    outputs(9933) <= not (a or b);
    outputs(9934) <= not b;
    outputs(9935) <= not (a xor b);
    outputs(9936) <= not (a xor b);
    outputs(9937) <= b and not a;
    outputs(9938) <= not (a xor b);
    outputs(9939) <= a xor b;
    outputs(9940) <= not a or b;
    outputs(9941) <= not (a xor b);
    outputs(9942) <= a xor b;
    outputs(9943) <= not a;
    outputs(9944) <= not (a or b);
    outputs(9945) <= a;
    outputs(9946) <= not (a or b);
    outputs(9947) <= not (a xor b);
    outputs(9948) <= a and not b;
    outputs(9949) <= b;
    outputs(9950) <= not (a xor b);
    outputs(9951) <= not (a or b);
    outputs(9952) <= not b;
    outputs(9953) <= a xor b;
    outputs(9954) <= a;
    outputs(9955) <= b and not a;
    outputs(9956) <= a xor b;
    outputs(9957) <= a and not b;
    outputs(9958) <= a xor b;
    outputs(9959) <= a xor b;
    outputs(9960) <= not (a xor b);
    outputs(9961) <= a;
    outputs(9962) <= not b;
    outputs(9963) <= a and b;
    outputs(9964) <= a xor b;
    outputs(9965) <= a;
    outputs(9966) <= not (a xor b);
    outputs(9967) <= a;
    outputs(9968) <= a xor b;
    outputs(9969) <= a and not b;
    outputs(9970) <= a;
    outputs(9971) <= not a;
    outputs(9972) <= b and not a;
    outputs(9973) <= not (a xor b);
    outputs(9974) <= b;
    outputs(9975) <= a;
    outputs(9976) <= b;
    outputs(9977) <= not (a and b);
    outputs(9978) <= a xor b;
    outputs(9979) <= not (a xor b);
    outputs(9980) <= not b;
    outputs(9981) <= a xor b;
    outputs(9982) <= a xor b;
    outputs(9983) <= a;
    outputs(9984) <= not a;
    outputs(9985) <= a and b;
    outputs(9986) <= b;
    outputs(9987) <= not a;
    outputs(9988) <= b;
    outputs(9989) <= a xor b;
    outputs(9990) <= a and not b;
    outputs(9991) <= a xor b;
    outputs(9992) <= b;
    outputs(9993) <= not b or a;
    outputs(9994) <= not (a or b);
    outputs(9995) <= a;
    outputs(9996) <= not b;
    outputs(9997) <= a and b;
    outputs(9998) <= a;
    outputs(9999) <= not b or a;
    outputs(10000) <= not a;
    outputs(10001) <= a xor b;
    outputs(10002) <= a xor b;
    outputs(10003) <= not b;
    outputs(10004) <= b;
    outputs(10005) <= not (a xor b);
    outputs(10006) <= not (a xor b);
    outputs(10007) <= not (a xor b);
    outputs(10008) <= b;
    outputs(10009) <= not a or b;
    outputs(10010) <= a;
    outputs(10011) <= not a;
    outputs(10012) <= not b or a;
    outputs(10013) <= b and not a;
    outputs(10014) <= a xor b;
    outputs(10015) <= not (a xor b);
    outputs(10016) <= not (a xor b);
    outputs(10017) <= b;
    outputs(10018) <= b;
    outputs(10019) <= a xor b;
    outputs(10020) <= not (a xor b);
    outputs(10021) <= not (a xor b);
    outputs(10022) <= a and not b;
    outputs(10023) <= a xor b;
    outputs(10024) <= a xor b;
    outputs(10025) <= a xor b;
    outputs(10026) <= not a or b;
    outputs(10027) <= b;
    outputs(10028) <= not b;
    outputs(10029) <= not b or a;
    outputs(10030) <= not (a or b);
    outputs(10031) <= a xor b;
    outputs(10032) <= a xor b;
    outputs(10033) <= not b or a;
    outputs(10034) <= a;
    outputs(10035) <= not a;
    outputs(10036) <= b;
    outputs(10037) <= a xor b;
    outputs(10038) <= a xor b;
    outputs(10039) <= not b;
    outputs(10040) <= not a or b;
    outputs(10041) <= not b;
    outputs(10042) <= b;
    outputs(10043) <= b;
    outputs(10044) <= not a;
    outputs(10045) <= not (a xor b);
    outputs(10046) <= not a;
    outputs(10047) <= not a;
    outputs(10048) <= not (a xor b);
    outputs(10049) <= not (a xor b);
    outputs(10050) <= not (a xor b);
    outputs(10051) <= a;
    outputs(10052) <= a xor b;
    outputs(10053) <= not (a xor b);
    outputs(10054) <= a and not b;
    outputs(10055) <= a;
    outputs(10056) <= a;
    outputs(10057) <= a;
    outputs(10058) <= not b;
    outputs(10059) <= b;
    outputs(10060) <= not (a xor b);
    outputs(10061) <= a;
    outputs(10062) <= a;
    outputs(10063) <= not a;
    outputs(10064) <= a;
    outputs(10065) <= not (a xor b);
    outputs(10066) <= b;
    outputs(10067) <= not (a or b);
    outputs(10068) <= not b;
    outputs(10069) <= b;
    outputs(10070) <= b;
    outputs(10071) <= b;
    outputs(10072) <= not (a and b);
    outputs(10073) <= not b;
    outputs(10074) <= a and not b;
    outputs(10075) <= not (a xor b);
    outputs(10076) <= not a;
    outputs(10077) <= a and not b;
    outputs(10078) <= not a or b;
    outputs(10079) <= b and not a;
    outputs(10080) <= a;
    outputs(10081) <= not a;
    outputs(10082) <= b;
    outputs(10083) <= not (a xor b);
    outputs(10084) <= not b;
    outputs(10085) <= not a;
    outputs(10086) <= not (a or b);
    outputs(10087) <= not (a xor b);
    outputs(10088) <= not b;
    outputs(10089) <= not (a xor b);
    outputs(10090) <= not a or b;
    outputs(10091) <= a and not b;
    outputs(10092) <= a xor b;
    outputs(10093) <= a xor b;
    outputs(10094) <= a xor b;
    outputs(10095) <= not (a xor b);
    outputs(10096) <= a xor b;
    outputs(10097) <= not (a or b);
    outputs(10098) <= a;
    outputs(10099) <= a;
    outputs(10100) <= a and b;
    outputs(10101) <= not b;
    outputs(10102) <= a xor b;
    outputs(10103) <= a xor b;
    outputs(10104) <= not b;
    outputs(10105) <= a xor b;
    outputs(10106) <= a;
    outputs(10107) <= not (a xor b);
    outputs(10108) <= b;
    outputs(10109) <= a or b;
    outputs(10110) <= not (a or b);
    outputs(10111) <= b and not a;
    outputs(10112) <= not (a and b);
    outputs(10113) <= a;
    outputs(10114) <= a xor b;
    outputs(10115) <= b and not a;
    outputs(10116) <= not b or a;
    outputs(10117) <= a or b;
    outputs(10118) <= a xor b;
    outputs(10119) <= not (a or b);
    outputs(10120) <= a or b;
    outputs(10121) <= not a;
    outputs(10122) <= b;
    outputs(10123) <= not b or a;
    outputs(10124) <= not b;
    outputs(10125) <= a xor b;
    outputs(10126) <= b;
    outputs(10127) <= a xor b;
    outputs(10128) <= not (a xor b);
    outputs(10129) <= a xor b;
    outputs(10130) <= a xor b;
    outputs(10131) <= a xor b;
    outputs(10132) <= not a;
    outputs(10133) <= not (a xor b);
    outputs(10134) <= a;
    outputs(10135) <= a and b;
    outputs(10136) <= b and not a;
    outputs(10137) <= not (a xor b);
    outputs(10138) <= not (a xor b);
    outputs(10139) <= b;
    outputs(10140) <= not b;
    outputs(10141) <= a xor b;
    outputs(10142) <= not a;
    outputs(10143) <= not a;
    outputs(10144) <= a and b;
    outputs(10145) <= not (a xor b);
    outputs(10146) <= not (a and b);
    outputs(10147) <= b;
    outputs(10148) <= a;
    outputs(10149) <= not a;
    outputs(10150) <= b and not a;
    outputs(10151) <= b;
    outputs(10152) <= not (a or b);
    outputs(10153) <= b;
    outputs(10154) <= a;
    outputs(10155) <= a xor b;
    outputs(10156) <= not a;
    outputs(10157) <= a xor b;
    outputs(10158) <= not (a xor b);
    outputs(10159) <= not (a xor b);
    outputs(10160) <= a xor b;
    outputs(10161) <= a and not b;
    outputs(10162) <= not b or a;
    outputs(10163) <= not b;
    outputs(10164) <= a and not b;
    outputs(10165) <= a;
    outputs(10166) <= not (a xor b);
    outputs(10167) <= a xor b;
    outputs(10168) <= not a or b;
    outputs(10169) <= a xor b;
    outputs(10170) <= b;
    outputs(10171) <= not (a xor b);
    outputs(10172) <= not a;
    outputs(10173) <= a xor b;
    outputs(10174) <= b;
    outputs(10175) <= not (a xor b);
    outputs(10176) <= not b;
    outputs(10177) <= a or b;
    outputs(10178) <= not (a xor b);
    outputs(10179) <= a or b;
    outputs(10180) <= a xor b;
    outputs(10181) <= a xor b;
    outputs(10182) <= not b;
    outputs(10183) <= a xor b;
    outputs(10184) <= not (a and b);
    outputs(10185) <= not a;
    outputs(10186) <= b;
    outputs(10187) <= b and not a;
    outputs(10188) <= b;
    outputs(10189) <= a and b;
    outputs(10190) <= not (a xor b);
    outputs(10191) <= a xor b;
    outputs(10192) <= a xor b;
    outputs(10193) <= not (a xor b);
    outputs(10194) <= not a;
    outputs(10195) <= not a;
    outputs(10196) <= a xor b;
    outputs(10197) <= not (a xor b);
    outputs(10198) <= not (a and b);
    outputs(10199) <= a;
    outputs(10200) <= a and b;
    outputs(10201) <= not (a xor b);
    outputs(10202) <= not b;
    outputs(10203) <= a;
    outputs(10204) <= not a;
    outputs(10205) <= a xor b;
    outputs(10206) <= a;
    outputs(10207) <= a xor b;
    outputs(10208) <= not b;
    outputs(10209) <= a;
    outputs(10210) <= not (a and b);
    outputs(10211) <= a xor b;
    outputs(10212) <= not a or b;
    outputs(10213) <= not a;
    outputs(10214) <= b;
    outputs(10215) <= a xor b;
    outputs(10216) <= a and not b;
    outputs(10217) <= not (a xor b);
    outputs(10218) <= a xor b;
    outputs(10219) <= a xor b;
    outputs(10220) <= a xor b;
    outputs(10221) <= b and not a;
    outputs(10222) <= not (a xor b);
    outputs(10223) <= not b;
    outputs(10224) <= not (a xor b);
    outputs(10225) <= a xor b;
    outputs(10226) <= a xor b;
    outputs(10227) <= b;
    outputs(10228) <= b and not a;
    outputs(10229) <= not a or b;
    outputs(10230) <= not a;
    outputs(10231) <= not b;
    outputs(10232) <= not b;
    outputs(10233) <= b;
    outputs(10234) <= not b or a;
    outputs(10235) <= not b;
    outputs(10236) <= not (a and b);
    outputs(10237) <= not (a xor b);
    outputs(10238) <= not (a xor b);
    outputs(10239) <= a and not b;
end Behavioral;
