module dummy_network(
    input wire [255:0] inputs,
    output wire [2559:0] outputs
);

    assign outputs = 2560'b0;
endmodule