library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);
    signal layer1_outputs : std_logic_vector(2559 downto 0);
    signal layer2_outputs : std_logic_vector(2559 downto 0);
    signal layer3_outputs : std_logic_vector(2559 downto 0);
    signal layer4_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= '1';
    layer0_outputs(1) <= (inputs(36)) and not (inputs(76));
    layer0_outputs(2) <= not(inputs(227));
    layer0_outputs(3) <= '1';
    layer0_outputs(4) <= '0';
    layer0_outputs(5) <= not(inputs(100));
    layer0_outputs(6) <= '1';
    layer0_outputs(7) <= not(inputs(127)) or (inputs(136));
    layer0_outputs(8) <= (inputs(63)) or (inputs(62));
    layer0_outputs(9) <= '0';
    layer0_outputs(10) <= not(inputs(112));
    layer0_outputs(11) <= inputs(75);
    layer0_outputs(12) <= inputs(81);
    layer0_outputs(13) <= inputs(82);
    layer0_outputs(14) <= '1';
    layer0_outputs(15) <= not(inputs(200)) or (inputs(102));
    layer0_outputs(16) <= '0';
    layer0_outputs(17) <= (inputs(91)) or (inputs(58));
    layer0_outputs(18) <= (inputs(45)) xor (inputs(92));
    layer0_outputs(19) <= inputs(147);
    layer0_outputs(20) <= not(inputs(57)) or (inputs(116));
    layer0_outputs(21) <= not(inputs(151)) or (inputs(240));
    layer0_outputs(22) <= not(inputs(186));
    layer0_outputs(23) <= (inputs(110)) or (inputs(8));
    layer0_outputs(24) <= not((inputs(133)) or (inputs(218)));
    layer0_outputs(25) <= '1';
    layer0_outputs(26) <= '1';
    layer0_outputs(27) <= (inputs(156)) and (inputs(187));
    layer0_outputs(28) <= not((inputs(83)) or (inputs(84)));
    layer0_outputs(29) <= not(inputs(248)) or (inputs(85));
    layer0_outputs(30) <= not(inputs(246));
    layer0_outputs(31) <= not(inputs(31)) or (inputs(63));
    layer0_outputs(32) <= not(inputs(151));
    layer0_outputs(33) <= not(inputs(184)) or (inputs(133));
    layer0_outputs(34) <= not((inputs(252)) xor (inputs(95)));
    layer0_outputs(35) <= not(inputs(231));
    layer0_outputs(36) <= not(inputs(179));
    layer0_outputs(37) <= not(inputs(76));
    layer0_outputs(38) <= not(inputs(109));
    layer0_outputs(39) <= not(inputs(144));
    layer0_outputs(40) <= inputs(213);
    layer0_outputs(41) <= (inputs(250)) and not (inputs(8));
    layer0_outputs(42) <= (inputs(121)) or (inputs(183));
    layer0_outputs(43) <= '0';
    layer0_outputs(44) <= '0';
    layer0_outputs(45) <= inputs(107);
    layer0_outputs(46) <= not(inputs(180));
    layer0_outputs(47) <= (inputs(56)) xor (inputs(56));
    layer0_outputs(48) <= inputs(242);
    layer0_outputs(49) <= (inputs(175)) and (inputs(138));
    layer0_outputs(50) <= (inputs(160)) and not (inputs(218));
    layer0_outputs(51) <= (inputs(160)) and (inputs(209));
    layer0_outputs(52) <= not((inputs(211)) or (inputs(63)));
    layer0_outputs(53) <= (inputs(157)) and (inputs(45));
    layer0_outputs(54) <= inputs(245);
    layer0_outputs(55) <= not((inputs(213)) xor (inputs(197)));
    layer0_outputs(56) <= (inputs(63)) or (inputs(129));
    layer0_outputs(57) <= inputs(228);
    layer0_outputs(58) <= not((inputs(24)) or (inputs(197)));
    layer0_outputs(59) <= not(inputs(167)) or (inputs(105));
    layer0_outputs(60) <= '1';
    layer0_outputs(61) <= not((inputs(65)) xor (inputs(20)));
    layer0_outputs(62) <= inputs(33);
    layer0_outputs(63) <= not(inputs(97)) or (inputs(118));
    layer0_outputs(64) <= inputs(83);
    layer0_outputs(65) <= not((inputs(139)) or (inputs(251)));
    layer0_outputs(66) <= not(inputs(42));
    layer0_outputs(67) <= inputs(114);
    layer0_outputs(68) <= not(inputs(173));
    layer0_outputs(69) <= inputs(205);
    layer0_outputs(70) <= not(inputs(99)) or (inputs(61));
    layer0_outputs(71) <= not(inputs(248)) or (inputs(32));
    layer0_outputs(72) <= not(inputs(1)) or (inputs(166));
    layer0_outputs(73) <= inputs(131);
    layer0_outputs(74) <= inputs(115);
    layer0_outputs(75) <= '0';
    layer0_outputs(76) <= (inputs(199)) or (inputs(197));
    layer0_outputs(77) <= not(inputs(79));
    layer0_outputs(78) <= inputs(61);
    layer0_outputs(79) <= not((inputs(79)) or (inputs(101)));
    layer0_outputs(80) <= (inputs(95)) and not (inputs(218));
    layer0_outputs(81) <= '0';
    layer0_outputs(82) <= not((inputs(138)) and (inputs(242)));
    layer0_outputs(83) <= inputs(226);
    layer0_outputs(84) <= '1';
    layer0_outputs(85) <= inputs(196);
    layer0_outputs(86) <= inputs(123);
    layer0_outputs(87) <= not(inputs(181));
    layer0_outputs(88) <= not(inputs(234));
    layer0_outputs(89) <= not(inputs(34)) or (inputs(15));
    layer0_outputs(90) <= not((inputs(144)) or (inputs(100)));
    layer0_outputs(91) <= not((inputs(98)) or (inputs(96)));
    layer0_outputs(92) <= (inputs(118)) and not (inputs(155));
    layer0_outputs(93) <= inputs(228);
    layer0_outputs(94) <= inputs(210);
    layer0_outputs(95) <= '1';
    layer0_outputs(96) <= not(inputs(173));
    layer0_outputs(97) <= not(inputs(136)) or (inputs(192));
    layer0_outputs(98) <= (inputs(111)) or (inputs(140));
    layer0_outputs(99) <= inputs(220);
    layer0_outputs(100) <= inputs(188);
    layer0_outputs(101) <= inputs(106);
    layer0_outputs(102) <= not((inputs(253)) or (inputs(106)));
    layer0_outputs(103) <= not(inputs(62)) or (inputs(66));
    layer0_outputs(104) <= not(inputs(89));
    layer0_outputs(105) <= '0';
    layer0_outputs(106) <= (inputs(212)) xor (inputs(178));
    layer0_outputs(107) <= (inputs(198)) and (inputs(34));
    layer0_outputs(108) <= not((inputs(84)) xor (inputs(81)));
    layer0_outputs(109) <= not((inputs(56)) xor (inputs(42)));
    layer0_outputs(110) <= inputs(134);
    layer0_outputs(111) <= '1';
    layer0_outputs(112) <= not(inputs(83)) or (inputs(247));
    layer0_outputs(113) <= not((inputs(39)) xor (inputs(148)));
    layer0_outputs(114) <= not(inputs(163));
    layer0_outputs(115) <= (inputs(140)) and not (inputs(240));
    layer0_outputs(116) <= '1';
    layer0_outputs(117) <= '1';
    layer0_outputs(118) <= not((inputs(59)) or (inputs(50)));
    layer0_outputs(119) <= not(inputs(22)) or (inputs(152));
    layer0_outputs(120) <= (inputs(46)) or (inputs(32));
    layer0_outputs(121) <= not((inputs(143)) and (inputs(243)));
    layer0_outputs(122) <= '0';
    layer0_outputs(123) <= not(inputs(190)) or (inputs(3));
    layer0_outputs(124) <= (inputs(53)) xor (inputs(115));
    layer0_outputs(125) <= not(inputs(248));
    layer0_outputs(126) <= (inputs(17)) and (inputs(58));
    layer0_outputs(127) <= inputs(13);
    layer0_outputs(128) <= (inputs(172)) and not (inputs(71));
    layer0_outputs(129) <= not(inputs(138));
    layer0_outputs(130) <= not((inputs(55)) and (inputs(21)));
    layer0_outputs(131) <= (inputs(117)) and not (inputs(158));
    layer0_outputs(132) <= (inputs(103)) or (inputs(162));
    layer0_outputs(133) <= (inputs(102)) and not (inputs(223));
    layer0_outputs(134) <= not(inputs(221)) or (inputs(236));
    layer0_outputs(135) <= inputs(193);
    layer0_outputs(136) <= '0';
    layer0_outputs(137) <= (inputs(60)) and not (inputs(96));
    layer0_outputs(138) <= (inputs(21)) or (inputs(249));
    layer0_outputs(139) <= not(inputs(64)) or (inputs(126));
    layer0_outputs(140) <= not((inputs(172)) and (inputs(19)));
    layer0_outputs(141) <= (inputs(143)) and (inputs(3));
    layer0_outputs(142) <= inputs(113);
    layer0_outputs(143) <= not((inputs(65)) or (inputs(99)));
    layer0_outputs(144) <= not(inputs(167));
    layer0_outputs(145) <= not(inputs(156));
    layer0_outputs(146) <= not((inputs(128)) or (inputs(211)));
    layer0_outputs(147) <= inputs(167);
    layer0_outputs(148) <= '1';
    layer0_outputs(149) <= not(inputs(100));
    layer0_outputs(150) <= (inputs(124)) or (inputs(114));
    layer0_outputs(151) <= (inputs(142)) and not (inputs(252));
    layer0_outputs(152) <= (inputs(202)) and not (inputs(30));
    layer0_outputs(153) <= inputs(129);
    layer0_outputs(154) <= not(inputs(210));
    layer0_outputs(155) <= not((inputs(235)) and (inputs(225)));
    layer0_outputs(156) <= (inputs(83)) or (inputs(214));
    layer0_outputs(157) <= (inputs(125)) or (inputs(132));
    layer0_outputs(158) <= (inputs(230)) and not (inputs(195));
    layer0_outputs(159) <= not(inputs(53)) or (inputs(248));
    layer0_outputs(160) <= (inputs(38)) or (inputs(143));
    layer0_outputs(161) <= '0';
    layer0_outputs(162) <= not(inputs(145));
    layer0_outputs(163) <= (inputs(207)) or (inputs(125));
    layer0_outputs(164) <= not(inputs(230)) or (inputs(190));
    layer0_outputs(165) <= not(inputs(179));
    layer0_outputs(166) <= not((inputs(84)) and (inputs(77)));
    layer0_outputs(167) <= inputs(2);
    layer0_outputs(168) <= (inputs(43)) or (inputs(129));
    layer0_outputs(169) <= not((inputs(146)) and (inputs(216)));
    layer0_outputs(170) <= '0';
    layer0_outputs(171) <= '0';
    layer0_outputs(172) <= not((inputs(240)) and (inputs(7)));
    layer0_outputs(173) <= not(inputs(158));
    layer0_outputs(174) <= not((inputs(91)) or (inputs(91)));
    layer0_outputs(175) <= not((inputs(103)) or (inputs(10)));
    layer0_outputs(176) <= not(inputs(29));
    layer0_outputs(177) <= '0';
    layer0_outputs(178) <= (inputs(176)) and (inputs(126));
    layer0_outputs(179) <= not((inputs(125)) or (inputs(39)));
    layer0_outputs(180) <= not(inputs(198));
    layer0_outputs(181) <= (inputs(186)) or (inputs(16));
    layer0_outputs(182) <= not((inputs(160)) and (inputs(69)));
    layer0_outputs(183) <= not((inputs(250)) and (inputs(165)));
    layer0_outputs(184) <= '1';
    layer0_outputs(185) <= not(inputs(129)) or (inputs(34));
    layer0_outputs(186) <= not(inputs(106));
    layer0_outputs(187) <= inputs(167);
    layer0_outputs(188) <= not((inputs(95)) and (inputs(83)));
    layer0_outputs(189) <= '1';
    layer0_outputs(190) <= not((inputs(102)) or (inputs(13)));
    layer0_outputs(191) <= not(inputs(225));
    layer0_outputs(192) <= not(inputs(101));
    layer0_outputs(193) <= (inputs(94)) or (inputs(21));
    layer0_outputs(194) <= (inputs(223)) or (inputs(24));
    layer0_outputs(195) <= (inputs(141)) and not (inputs(169));
    layer0_outputs(196) <= not(inputs(183)) or (inputs(244));
    layer0_outputs(197) <= not((inputs(191)) xor (inputs(56)));
    layer0_outputs(198) <= (inputs(209)) xor (inputs(191));
    layer0_outputs(199) <= inputs(75);
    layer0_outputs(200) <= inputs(154);
    layer0_outputs(201) <= not(inputs(179));
    layer0_outputs(202) <= (inputs(175)) and not (inputs(71));
    layer0_outputs(203) <= (inputs(184)) and not (inputs(133));
    layer0_outputs(204) <= (inputs(12)) or (inputs(212));
    layer0_outputs(205) <= (inputs(150)) and not (inputs(174));
    layer0_outputs(206) <= (inputs(242)) and (inputs(66));
    layer0_outputs(207) <= '1';
    layer0_outputs(208) <= (inputs(103)) and not (inputs(64));
    layer0_outputs(209) <= not((inputs(120)) or (inputs(14)));
    layer0_outputs(210) <= (inputs(66)) and not (inputs(206));
    layer0_outputs(211) <= (inputs(20)) and not (inputs(102));
    layer0_outputs(212) <= not(inputs(167));
    layer0_outputs(213) <= inputs(60);
    layer0_outputs(214) <= (inputs(52)) xor (inputs(176));
    layer0_outputs(215) <= not(inputs(31)) or (inputs(151));
    layer0_outputs(216) <= (inputs(221)) and not (inputs(253));
    layer0_outputs(217) <= '0';
    layer0_outputs(218) <= inputs(33);
    layer0_outputs(219) <= (inputs(246)) and not (inputs(20));
    layer0_outputs(220) <= (inputs(6)) xor (inputs(62));
    layer0_outputs(221) <= (inputs(205)) and not (inputs(78));
    layer0_outputs(222) <= not(inputs(165));
    layer0_outputs(223) <= inputs(201);
    layer0_outputs(224) <= inputs(93);
    layer0_outputs(225) <= not(inputs(233)) or (inputs(9));
    layer0_outputs(226) <= inputs(39);
    layer0_outputs(227) <= (inputs(206)) and (inputs(200));
    layer0_outputs(228) <= not(inputs(196));
    layer0_outputs(229) <= not((inputs(111)) and (inputs(141)));
    layer0_outputs(230) <= (inputs(196)) or (inputs(249));
    layer0_outputs(231) <= '1';
    layer0_outputs(232) <= not((inputs(140)) or (inputs(170)));
    layer0_outputs(233) <= '0';
    layer0_outputs(234) <= not((inputs(207)) and (inputs(208)));
    layer0_outputs(235) <= not(inputs(2));
    layer0_outputs(236) <= (inputs(115)) or (inputs(246));
    layer0_outputs(237) <= not(inputs(227)) or (inputs(136));
    layer0_outputs(238) <= not((inputs(9)) xor (inputs(1)));
    layer0_outputs(239) <= not(inputs(169)) or (inputs(5));
    layer0_outputs(240) <= '1';
    layer0_outputs(241) <= not(inputs(164));
    layer0_outputs(242) <= inputs(82);
    layer0_outputs(243) <= not((inputs(91)) or (inputs(45)));
    layer0_outputs(244) <= (inputs(90)) and not (inputs(144));
    layer0_outputs(245) <= (inputs(195)) and (inputs(19));
    layer0_outputs(246) <= not(inputs(87)) or (inputs(180));
    layer0_outputs(247) <= inputs(147);
    layer0_outputs(248) <= not(inputs(24));
    layer0_outputs(249) <= not(inputs(94));
    layer0_outputs(250) <= not(inputs(105));
    layer0_outputs(251) <= not((inputs(222)) or (inputs(23)));
    layer0_outputs(252) <= not(inputs(171));
    layer0_outputs(253) <= (inputs(113)) and not (inputs(43));
    layer0_outputs(254) <= not((inputs(100)) or (inputs(29)));
    layer0_outputs(255) <= '0';
    layer0_outputs(256) <= (inputs(40)) or (inputs(70));
    layer0_outputs(257) <= not(inputs(151));
    layer0_outputs(258) <= not((inputs(88)) and (inputs(158)));
    layer0_outputs(259) <= inputs(90);
    layer0_outputs(260) <= '0';
    layer0_outputs(261) <= inputs(134);
    layer0_outputs(262) <= not(inputs(158));
    layer0_outputs(263) <= (inputs(56)) and not (inputs(213));
    layer0_outputs(264) <= inputs(52);
    layer0_outputs(265) <= (inputs(170)) and not (inputs(118));
    layer0_outputs(266) <= inputs(138);
    layer0_outputs(267) <= not(inputs(26));
    layer0_outputs(268) <= inputs(247);
    layer0_outputs(269) <= (inputs(189)) and not (inputs(101));
    layer0_outputs(270) <= inputs(210);
    layer0_outputs(271) <= (inputs(233)) and (inputs(230));
    layer0_outputs(272) <= not(inputs(103));
    layer0_outputs(273) <= (inputs(234)) or (inputs(205));
    layer0_outputs(274) <= '1';
    layer0_outputs(275) <= not((inputs(5)) or (inputs(28)));
    layer0_outputs(276) <= (inputs(205)) and not (inputs(144));
    layer0_outputs(277) <= '1';
    layer0_outputs(278) <= not((inputs(167)) and (inputs(27)));
    layer0_outputs(279) <= not((inputs(8)) or (inputs(158)));
    layer0_outputs(280) <= not(inputs(194));
    layer0_outputs(281) <= not(inputs(105));
    layer0_outputs(282) <= not(inputs(35)) or (inputs(14));
    layer0_outputs(283) <= (inputs(203)) xor (inputs(236));
    layer0_outputs(284) <= not(inputs(172)) or (inputs(80));
    layer0_outputs(285) <= (inputs(202)) or (inputs(2));
    layer0_outputs(286) <= not((inputs(74)) and (inputs(252)));
    layer0_outputs(287) <= (inputs(138)) and not (inputs(56));
    layer0_outputs(288) <= inputs(104);
    layer0_outputs(289) <= not((inputs(33)) or (inputs(123)));
    layer0_outputs(290) <= '0';
    layer0_outputs(291) <= not(inputs(33));
    layer0_outputs(292) <= not(inputs(72));
    layer0_outputs(293) <= not(inputs(238));
    layer0_outputs(294) <= (inputs(235)) or (inputs(183));
    layer0_outputs(295) <= inputs(210);
    layer0_outputs(296) <= not(inputs(38)) or (inputs(126));
    layer0_outputs(297) <= inputs(64);
    layer0_outputs(298) <= inputs(100);
    layer0_outputs(299) <= not(inputs(204)) or (inputs(99));
    layer0_outputs(300) <= not(inputs(87));
    layer0_outputs(301) <= (inputs(18)) or (inputs(136));
    layer0_outputs(302) <= not(inputs(234)) or (inputs(120));
    layer0_outputs(303) <= inputs(122);
    layer0_outputs(304) <= '1';
    layer0_outputs(305) <= '1';
    layer0_outputs(306) <= (inputs(71)) or (inputs(196));
    layer0_outputs(307) <= not(inputs(6));
    layer0_outputs(308) <= not(inputs(57));
    layer0_outputs(309) <= (inputs(183)) and not (inputs(122));
    layer0_outputs(310) <= inputs(180);
    layer0_outputs(311) <= not(inputs(246));
    layer0_outputs(312) <= inputs(133);
    layer0_outputs(313) <= not(inputs(31));
    layer0_outputs(314) <= not(inputs(0)) or (inputs(44));
    layer0_outputs(315) <= not(inputs(156));
    layer0_outputs(316) <= inputs(213);
    layer0_outputs(317) <= inputs(129);
    layer0_outputs(318) <= (inputs(253)) or (inputs(81));
    layer0_outputs(319) <= (inputs(202)) or (inputs(138));
    layer0_outputs(320) <= inputs(87);
    layer0_outputs(321) <= not(inputs(79));
    layer0_outputs(322) <= (inputs(132)) and not (inputs(240));
    layer0_outputs(323) <= inputs(180);
    layer0_outputs(324) <= inputs(188);
    layer0_outputs(325) <= inputs(67);
    layer0_outputs(326) <= (inputs(98)) or (inputs(173));
    layer0_outputs(327) <= not((inputs(166)) or (inputs(179)));
    layer0_outputs(328) <= (inputs(114)) or (inputs(219));
    layer0_outputs(329) <= (inputs(16)) and not (inputs(105));
    layer0_outputs(330) <= not((inputs(157)) and (inputs(9)));
    layer0_outputs(331) <= inputs(161);
    layer0_outputs(332) <= not(inputs(95));
    layer0_outputs(333) <= inputs(55);
    layer0_outputs(334) <= not((inputs(85)) or (inputs(226)));
    layer0_outputs(335) <= '1';
    layer0_outputs(336) <= not((inputs(193)) or (inputs(133)));
    layer0_outputs(337) <= (inputs(26)) and not (inputs(176));
    layer0_outputs(338) <= '0';
    layer0_outputs(339) <= '1';
    layer0_outputs(340) <= not(inputs(9));
    layer0_outputs(341) <= '1';
    layer0_outputs(342) <= (inputs(49)) and (inputs(160));
    layer0_outputs(343) <= not((inputs(235)) or (inputs(90)));
    layer0_outputs(344) <= (inputs(98)) or (inputs(163));
    layer0_outputs(345) <= not(inputs(16));
    layer0_outputs(346) <= not(inputs(112));
    layer0_outputs(347) <= not(inputs(124)) or (inputs(99));
    layer0_outputs(348) <= not((inputs(203)) or (inputs(4)));
    layer0_outputs(349) <= inputs(17);
    layer0_outputs(350) <= not(inputs(137));
    layer0_outputs(351) <= (inputs(193)) or (inputs(60));
    layer0_outputs(352) <= inputs(53);
    layer0_outputs(353) <= not((inputs(198)) or (inputs(216)));
    layer0_outputs(354) <= (inputs(157)) and (inputs(68));
    layer0_outputs(355) <= '1';
    layer0_outputs(356) <= (inputs(7)) and (inputs(123));
    layer0_outputs(357) <= not(inputs(83));
    layer0_outputs(358) <= not((inputs(191)) or (inputs(209)));
    layer0_outputs(359) <= not(inputs(53));
    layer0_outputs(360) <= not(inputs(19));
    layer0_outputs(361) <= (inputs(88)) and not (inputs(64));
    layer0_outputs(362) <= (inputs(5)) or (inputs(171));
    layer0_outputs(363) <= not(inputs(50));
    layer0_outputs(364) <= '1';
    layer0_outputs(365) <= not(inputs(109));
    layer0_outputs(366) <= (inputs(14)) or (inputs(128));
    layer0_outputs(367) <= (inputs(38)) and (inputs(52));
    layer0_outputs(368) <= (inputs(230)) and (inputs(229));
    layer0_outputs(369) <= (inputs(112)) and not (inputs(152));
    layer0_outputs(370) <= not(inputs(231));
    layer0_outputs(371) <= not(inputs(0));
    layer0_outputs(372) <= not(inputs(37));
    layer0_outputs(373) <= inputs(54);
    layer0_outputs(374) <= not(inputs(150));
    layer0_outputs(375) <= not(inputs(210));
    layer0_outputs(376) <= not((inputs(120)) or (inputs(11)));
    layer0_outputs(377) <= not(inputs(134)) or (inputs(48));
    layer0_outputs(378) <= not(inputs(162));
    layer0_outputs(379) <= '0';
    layer0_outputs(380) <= not(inputs(21));
    layer0_outputs(381) <= inputs(197);
    layer0_outputs(382) <= '1';
    layer0_outputs(383) <= not(inputs(118));
    layer0_outputs(384) <= inputs(119);
    layer0_outputs(385) <= (inputs(16)) and not (inputs(29));
    layer0_outputs(386) <= inputs(19);
    layer0_outputs(387) <= (inputs(73)) and not (inputs(234));
    layer0_outputs(388) <= inputs(217);
    layer0_outputs(389) <= inputs(150);
    layer0_outputs(390) <= (inputs(58)) or (inputs(154));
    layer0_outputs(391) <= '0';
    layer0_outputs(392) <= not(inputs(167));
    layer0_outputs(393) <= (inputs(72)) and (inputs(89));
    layer0_outputs(394) <= inputs(148);
    layer0_outputs(395) <= (inputs(40)) or (inputs(243));
    layer0_outputs(396) <= (inputs(123)) and (inputs(42));
    layer0_outputs(397) <= inputs(104);
    layer0_outputs(398) <= not(inputs(162));
    layer0_outputs(399) <= not(inputs(36));
    layer0_outputs(400) <= inputs(163);
    layer0_outputs(401) <= not(inputs(146));
    layer0_outputs(402) <= not(inputs(165));
    layer0_outputs(403) <= inputs(37);
    layer0_outputs(404) <= (inputs(23)) and not (inputs(178));
    layer0_outputs(405) <= not((inputs(108)) or (inputs(161)));
    layer0_outputs(406) <= not(inputs(91));
    layer0_outputs(407) <= not(inputs(132));
    layer0_outputs(408) <= not(inputs(152));
    layer0_outputs(409) <= not((inputs(230)) or (inputs(46)));
    layer0_outputs(410) <= inputs(99);
    layer0_outputs(411) <= not(inputs(237));
    layer0_outputs(412) <= not(inputs(164));
    layer0_outputs(413) <= not((inputs(96)) or (inputs(68)));
    layer0_outputs(414) <= not(inputs(214)) or (inputs(165));
    layer0_outputs(415) <= inputs(188);
    layer0_outputs(416) <= '0';
    layer0_outputs(417) <= '0';
    layer0_outputs(418) <= inputs(106);
    layer0_outputs(419) <= not(inputs(226)) or (inputs(152));
    layer0_outputs(420) <= '0';
    layer0_outputs(421) <= (inputs(203)) or (inputs(210));
    layer0_outputs(422) <= inputs(75);
    layer0_outputs(423) <= '0';
    layer0_outputs(424) <= inputs(91);
    layer0_outputs(425) <= (inputs(16)) or (inputs(205));
    layer0_outputs(426) <= not(inputs(111));
    layer0_outputs(427) <= inputs(6);
    layer0_outputs(428) <= '0';
    layer0_outputs(429) <= '0';
    layer0_outputs(430) <= (inputs(146)) and not (inputs(13));
    layer0_outputs(431) <= '1';
    layer0_outputs(432) <= not(inputs(219));
    layer0_outputs(433) <= not((inputs(28)) and (inputs(182)));
    layer0_outputs(434) <= (inputs(31)) and (inputs(1));
    layer0_outputs(435) <= '0';
    layer0_outputs(436) <= inputs(180);
    layer0_outputs(437) <= (inputs(98)) and not (inputs(168));
    layer0_outputs(438) <= not((inputs(76)) and (inputs(41)));
    layer0_outputs(439) <= '0';
    layer0_outputs(440) <= inputs(47);
    layer0_outputs(441) <= inputs(0);
    layer0_outputs(442) <= inputs(231);
    layer0_outputs(443) <= not((inputs(125)) or (inputs(43)));
    layer0_outputs(444) <= (inputs(132)) and (inputs(226));
    layer0_outputs(445) <= inputs(192);
    layer0_outputs(446) <= '1';
    layer0_outputs(447) <= not((inputs(254)) and (inputs(199)));
    layer0_outputs(448) <= not((inputs(105)) or (inputs(68)));
    layer0_outputs(449) <= not(inputs(192));
    layer0_outputs(450) <= (inputs(5)) and not (inputs(96));
    layer0_outputs(451) <= not(inputs(78));
    layer0_outputs(452) <= (inputs(115)) and not (inputs(222));
    layer0_outputs(453) <= not(inputs(67));
    layer0_outputs(454) <= (inputs(67)) or (inputs(171));
    layer0_outputs(455) <= not((inputs(171)) or (inputs(162)));
    layer0_outputs(456) <= (inputs(125)) and not (inputs(147));
    layer0_outputs(457) <= '1';
    layer0_outputs(458) <= not(inputs(72)) or (inputs(83));
    layer0_outputs(459) <= not(inputs(106));
    layer0_outputs(460) <= '0';
    layer0_outputs(461) <= inputs(47);
    layer0_outputs(462) <= not(inputs(155));
    layer0_outputs(463) <= not((inputs(178)) or (inputs(143)));
    layer0_outputs(464) <= inputs(213);
    layer0_outputs(465) <= '1';
    layer0_outputs(466) <= not(inputs(247));
    layer0_outputs(467) <= (inputs(110)) and not (inputs(34));
    layer0_outputs(468) <= not(inputs(218));
    layer0_outputs(469) <= (inputs(255)) and not (inputs(34));
    layer0_outputs(470) <= (inputs(244)) xor (inputs(199));
    layer0_outputs(471) <= not((inputs(208)) or (inputs(104)));
    layer0_outputs(472) <= '1';
    layer0_outputs(473) <= inputs(180);
    layer0_outputs(474) <= (inputs(92)) and (inputs(108));
    layer0_outputs(475) <= not(inputs(110));
    layer0_outputs(476) <= not((inputs(221)) or (inputs(99)));
    layer0_outputs(477) <= inputs(25);
    layer0_outputs(478) <= not((inputs(189)) or (inputs(222)));
    layer0_outputs(479) <= not(inputs(175));
    layer0_outputs(480) <= (inputs(82)) or (inputs(81));
    layer0_outputs(481) <= '1';
    layer0_outputs(482) <= '0';
    layer0_outputs(483) <= inputs(91);
    layer0_outputs(484) <= inputs(207);
    layer0_outputs(485) <= '0';
    layer0_outputs(486) <= not(inputs(101));
    layer0_outputs(487) <= not(inputs(194));
    layer0_outputs(488) <= '0';
    layer0_outputs(489) <= not((inputs(186)) or (inputs(162)));
    layer0_outputs(490) <= '1';
    layer0_outputs(491) <= inputs(4);
    layer0_outputs(492) <= '0';
    layer0_outputs(493) <= (inputs(15)) and not (inputs(8));
    layer0_outputs(494) <= '1';
    layer0_outputs(495) <= not(inputs(144));
    layer0_outputs(496) <= not(inputs(61)) or (inputs(190));
    layer0_outputs(497) <= (inputs(18)) and not (inputs(164));
    layer0_outputs(498) <= not(inputs(56));
    layer0_outputs(499) <= not(inputs(103));
    layer0_outputs(500) <= not(inputs(123)) or (inputs(33));
    layer0_outputs(501) <= '0';
    layer0_outputs(502) <= not((inputs(47)) and (inputs(244)));
    layer0_outputs(503) <= not(inputs(89));
    layer0_outputs(504) <= inputs(134);
    layer0_outputs(505) <= (inputs(213)) and (inputs(148));
    layer0_outputs(506) <= not((inputs(172)) or (inputs(148)));
    layer0_outputs(507) <= not((inputs(88)) and (inputs(33)));
    layer0_outputs(508) <= (inputs(220)) and (inputs(3));
    layer0_outputs(509) <= (inputs(163)) and not (inputs(157));
    layer0_outputs(510) <= inputs(194);
    layer0_outputs(511) <= not(inputs(165));
    layer0_outputs(512) <= not(inputs(174));
    layer0_outputs(513) <= '1';
    layer0_outputs(514) <= inputs(118);
    layer0_outputs(515) <= not((inputs(193)) or (inputs(173)));
    layer0_outputs(516) <= (inputs(196)) or (inputs(88));
    layer0_outputs(517) <= not((inputs(113)) or (inputs(124)));
    layer0_outputs(518) <= not(inputs(160));
    layer0_outputs(519) <= not(inputs(156));
    layer0_outputs(520) <= inputs(56);
    layer0_outputs(521) <= (inputs(82)) and not (inputs(200));
    layer0_outputs(522) <= not((inputs(188)) or (inputs(201)));
    layer0_outputs(523) <= (inputs(129)) and (inputs(200));
    layer0_outputs(524) <= not(inputs(126)) or (inputs(254));
    layer0_outputs(525) <= not((inputs(232)) and (inputs(123)));
    layer0_outputs(526) <= not(inputs(106));
    layer0_outputs(527) <= inputs(205);
    layer0_outputs(528) <= inputs(236);
    layer0_outputs(529) <= inputs(193);
    layer0_outputs(530) <= not(inputs(138)) or (inputs(93));
    layer0_outputs(531) <= not(inputs(129));
    layer0_outputs(532) <= inputs(117);
    layer0_outputs(533) <= not(inputs(241)) or (inputs(63));
    layer0_outputs(534) <= (inputs(211)) and not (inputs(4));
    layer0_outputs(535) <= not(inputs(165));
    layer0_outputs(536) <= (inputs(117)) or (inputs(174));
    layer0_outputs(537) <= not(inputs(93));
    layer0_outputs(538) <= '0';
    layer0_outputs(539) <= not((inputs(130)) or (inputs(203)));
    layer0_outputs(540) <= '0';
    layer0_outputs(541) <= not(inputs(119));
    layer0_outputs(542) <= inputs(177);
    layer0_outputs(543) <= inputs(216);
    layer0_outputs(544) <= not(inputs(40));
    layer0_outputs(545) <= (inputs(99)) or (inputs(80));
    layer0_outputs(546) <= not(inputs(95)) or (inputs(255));
    layer0_outputs(547) <= not((inputs(193)) or (inputs(80)));
    layer0_outputs(548) <= inputs(121);
    layer0_outputs(549) <= not(inputs(181));
    layer0_outputs(550) <= not(inputs(194)) or (inputs(127));
    layer0_outputs(551) <= inputs(214);
    layer0_outputs(552) <= not((inputs(140)) and (inputs(161)));
    layer0_outputs(553) <= not((inputs(229)) or (inputs(185)));
    layer0_outputs(554) <= (inputs(209)) and not (inputs(194));
    layer0_outputs(555) <= (inputs(175)) or (inputs(56));
    layer0_outputs(556) <= (inputs(27)) xor (inputs(105));
    layer0_outputs(557) <= not((inputs(189)) or (inputs(201)));
    layer0_outputs(558) <= inputs(183);
    layer0_outputs(559) <= (inputs(242)) and not (inputs(144));
    layer0_outputs(560) <= inputs(136);
    layer0_outputs(561) <= '0';
    layer0_outputs(562) <= (inputs(212)) or (inputs(131));
    layer0_outputs(563) <= '1';
    layer0_outputs(564) <= (inputs(24)) and not (inputs(128));
    layer0_outputs(565) <= not(inputs(72));
    layer0_outputs(566) <= inputs(130);
    layer0_outputs(567) <= (inputs(154)) and not (inputs(108));
    layer0_outputs(568) <= not((inputs(23)) or (inputs(84)));
    layer0_outputs(569) <= (inputs(158)) or (inputs(0));
    layer0_outputs(570) <= (inputs(112)) or (inputs(232));
    layer0_outputs(571) <= not(inputs(199)) or (inputs(77));
    layer0_outputs(572) <= not((inputs(28)) xor (inputs(223)));
    layer0_outputs(573) <= (inputs(51)) or (inputs(84));
    layer0_outputs(574) <= (inputs(125)) or (inputs(32));
    layer0_outputs(575) <= (inputs(53)) and not (inputs(189));
    layer0_outputs(576) <= not((inputs(52)) or (inputs(60)));
    layer0_outputs(577) <= not((inputs(151)) or (inputs(227)));
    layer0_outputs(578) <= (inputs(44)) and not (inputs(254));
    layer0_outputs(579) <= not((inputs(23)) or (inputs(220)));
    layer0_outputs(580) <= inputs(98);
    layer0_outputs(581) <= (inputs(188)) and not (inputs(15));
    layer0_outputs(582) <= (inputs(171)) and not (inputs(15));
    layer0_outputs(583) <= not(inputs(119)) or (inputs(60));
    layer0_outputs(584) <= inputs(52);
    layer0_outputs(585) <= not((inputs(217)) and (inputs(43)));
    layer0_outputs(586) <= inputs(3);
    layer0_outputs(587) <= not((inputs(32)) or (inputs(164)));
    layer0_outputs(588) <= '0';
    layer0_outputs(589) <= (inputs(82)) or (inputs(97));
    layer0_outputs(590) <= not((inputs(141)) xor (inputs(94)));
    layer0_outputs(591) <= (inputs(255)) or (inputs(188));
    layer0_outputs(592) <= (inputs(242)) and (inputs(131));
    layer0_outputs(593) <= not(inputs(139));
    layer0_outputs(594) <= not(inputs(130));
    layer0_outputs(595) <= inputs(83);
    layer0_outputs(596) <= not(inputs(187)) or (inputs(182));
    layer0_outputs(597) <= inputs(147);
    layer0_outputs(598) <= (inputs(133)) and not (inputs(153));
    layer0_outputs(599) <= not((inputs(43)) or (inputs(208)));
    layer0_outputs(600) <= (inputs(16)) and not (inputs(94));
    layer0_outputs(601) <= (inputs(62)) xor (inputs(148));
    layer0_outputs(602) <= (inputs(136)) and not (inputs(247));
    layer0_outputs(603) <= not((inputs(137)) and (inputs(70)));
    layer0_outputs(604) <= not((inputs(22)) or (inputs(168)));
    layer0_outputs(605) <= not(inputs(149));
    layer0_outputs(606) <= inputs(93);
    layer0_outputs(607) <= '1';
    layer0_outputs(608) <= not((inputs(26)) or (inputs(255)));
    layer0_outputs(609) <= not(inputs(58)) or (inputs(54));
    layer0_outputs(610) <= inputs(228);
    layer0_outputs(611) <= (inputs(169)) or (inputs(135));
    layer0_outputs(612) <= (inputs(107)) and not (inputs(239));
    layer0_outputs(613) <= not(inputs(153));
    layer0_outputs(614) <= inputs(98);
    layer0_outputs(615) <= (inputs(206)) and (inputs(165));
    layer0_outputs(616) <= (inputs(49)) xor (inputs(122));
    layer0_outputs(617) <= (inputs(10)) and (inputs(11));
    layer0_outputs(618) <= (inputs(142)) and (inputs(253));
    layer0_outputs(619) <= (inputs(199)) and (inputs(240));
    layer0_outputs(620) <= inputs(72);
    layer0_outputs(621) <= (inputs(66)) and not (inputs(212));
    layer0_outputs(622) <= (inputs(98)) and not (inputs(168));
    layer0_outputs(623) <= not(inputs(132)) or (inputs(76));
    layer0_outputs(624) <= '1';
    layer0_outputs(625) <= (inputs(37)) and not (inputs(4));
    layer0_outputs(626) <= (inputs(80)) or (inputs(78));
    layer0_outputs(627) <= not(inputs(25));
    layer0_outputs(628) <= (inputs(127)) or (inputs(21));
    layer0_outputs(629) <= '0';
    layer0_outputs(630) <= inputs(132);
    layer0_outputs(631) <= not(inputs(23));
    layer0_outputs(632) <= inputs(104);
    layer0_outputs(633) <= (inputs(85)) and (inputs(246));
    layer0_outputs(634) <= not(inputs(61));
    layer0_outputs(635) <= '1';
    layer0_outputs(636) <= not(inputs(73)) or (inputs(79));
    layer0_outputs(637) <= (inputs(154)) and not (inputs(132));
    layer0_outputs(638) <= not(inputs(207));
    layer0_outputs(639) <= not(inputs(209)) or (inputs(136));
    layer0_outputs(640) <= inputs(74);
    layer0_outputs(641) <= (inputs(115)) and not (inputs(63));
    layer0_outputs(642) <= (inputs(64)) and not (inputs(162));
    layer0_outputs(643) <= not(inputs(138));
    layer0_outputs(644) <= not(inputs(243)) or (inputs(121));
    layer0_outputs(645) <= not((inputs(54)) and (inputs(229)));
    layer0_outputs(646) <= (inputs(160)) and not (inputs(155));
    layer0_outputs(647) <= (inputs(210)) or (inputs(197));
    layer0_outputs(648) <= not(inputs(140));
    layer0_outputs(649) <= not(inputs(116));
    layer0_outputs(650) <= (inputs(121)) and not (inputs(175));
    layer0_outputs(651) <= not((inputs(101)) or (inputs(130)));
    layer0_outputs(652) <= not((inputs(191)) xor (inputs(90)));
    layer0_outputs(653) <= (inputs(253)) or (inputs(56));
    layer0_outputs(654) <= inputs(29);
    layer0_outputs(655) <= '0';
    layer0_outputs(656) <= '0';
    layer0_outputs(657) <= not(inputs(133)) or (inputs(240));
    layer0_outputs(658) <= (inputs(190)) and not (inputs(82));
    layer0_outputs(659) <= (inputs(185)) and not (inputs(247));
    layer0_outputs(660) <= '0';
    layer0_outputs(661) <= not(inputs(145));
    layer0_outputs(662) <= '1';
    layer0_outputs(663) <= not((inputs(139)) or (inputs(208)));
    layer0_outputs(664) <= not((inputs(62)) or (inputs(36)));
    layer0_outputs(665) <= (inputs(142)) or (inputs(227));
    layer0_outputs(666) <= not(inputs(236));
    layer0_outputs(667) <= '1';
    layer0_outputs(668) <= not(inputs(104));
    layer0_outputs(669) <= not(inputs(226));
    layer0_outputs(670) <= not((inputs(40)) and (inputs(88)));
    layer0_outputs(671) <= not(inputs(70)) or (inputs(136));
    layer0_outputs(672) <= inputs(121);
    layer0_outputs(673) <= inputs(232);
    layer0_outputs(674) <= (inputs(165)) xor (inputs(88));
    layer0_outputs(675) <= inputs(52);
    layer0_outputs(676) <= not(inputs(219));
    layer0_outputs(677) <= not(inputs(206)) or (inputs(128));
    layer0_outputs(678) <= '1';
    layer0_outputs(679) <= (inputs(77)) and not (inputs(105));
    layer0_outputs(680) <= not((inputs(241)) or (inputs(136)));
    layer0_outputs(681) <= not((inputs(146)) or (inputs(181)));
    layer0_outputs(682) <= not((inputs(11)) or (inputs(169)));
    layer0_outputs(683) <= (inputs(251)) and not (inputs(204));
    layer0_outputs(684) <= (inputs(65)) or (inputs(63));
    layer0_outputs(685) <= inputs(96);
    layer0_outputs(686) <= not(inputs(75)) or (inputs(47));
    layer0_outputs(687) <= '0';
    layer0_outputs(688) <= (inputs(45)) and (inputs(201));
    layer0_outputs(689) <= (inputs(213)) or (inputs(0));
    layer0_outputs(690) <= not(inputs(176));
    layer0_outputs(691) <= not((inputs(220)) or (inputs(222)));
    layer0_outputs(692) <= inputs(197);
    layer0_outputs(693) <= '1';
    layer0_outputs(694) <= '0';
    layer0_outputs(695) <= inputs(114);
    layer0_outputs(696) <= not(inputs(207)) or (inputs(46));
    layer0_outputs(697) <= not((inputs(225)) xor (inputs(33)));
    layer0_outputs(698) <= not(inputs(90));
    layer0_outputs(699) <= (inputs(48)) or (inputs(235));
    layer0_outputs(700) <= (inputs(51)) or (inputs(206));
    layer0_outputs(701) <= inputs(162);
    layer0_outputs(702) <= not(inputs(67));
    layer0_outputs(703) <= (inputs(165)) and not (inputs(35));
    layer0_outputs(704) <= not(inputs(20));
    layer0_outputs(705) <= inputs(22);
    layer0_outputs(706) <= not((inputs(176)) or (inputs(197)));
    layer0_outputs(707) <= (inputs(103)) and (inputs(136));
    layer0_outputs(708) <= not(inputs(59));
    layer0_outputs(709) <= inputs(124);
    layer0_outputs(710) <= not((inputs(171)) and (inputs(110)));
    layer0_outputs(711) <= '1';
    layer0_outputs(712) <= '0';
    layer0_outputs(713) <= '0';
    layer0_outputs(714) <= (inputs(209)) and not (inputs(183));
    layer0_outputs(715) <= not(inputs(179)) or (inputs(112));
    layer0_outputs(716) <= (inputs(213)) and (inputs(199));
    layer0_outputs(717) <= not(inputs(108)) or (inputs(252));
    layer0_outputs(718) <= inputs(170);
    layer0_outputs(719) <= (inputs(87)) and not (inputs(241));
    layer0_outputs(720) <= '1';
    layer0_outputs(721) <= not(inputs(229));
    layer0_outputs(722) <= (inputs(196)) and not (inputs(114));
    layer0_outputs(723) <= not(inputs(181));
    layer0_outputs(724) <= inputs(230);
    layer0_outputs(725) <= inputs(113);
    layer0_outputs(726) <= (inputs(49)) and not (inputs(146));
    layer0_outputs(727) <= '1';
    layer0_outputs(728) <= not((inputs(47)) or (inputs(139)));
    layer0_outputs(729) <= (inputs(209)) and not (inputs(89));
    layer0_outputs(730) <= not((inputs(88)) or (inputs(135)));
    layer0_outputs(731) <= (inputs(135)) and not (inputs(117));
    layer0_outputs(732) <= not((inputs(27)) or (inputs(31)));
    layer0_outputs(733) <= '1';
    layer0_outputs(734) <= inputs(255);
    layer0_outputs(735) <= '0';
    layer0_outputs(736) <= (inputs(126)) or (inputs(211));
    layer0_outputs(737) <= not(inputs(78));
    layer0_outputs(738) <= inputs(208);
    layer0_outputs(739) <= (inputs(116)) and not (inputs(32));
    layer0_outputs(740) <= '0';
    layer0_outputs(741) <= (inputs(192)) or (inputs(214));
    layer0_outputs(742) <= (inputs(190)) and not (inputs(159));
    layer0_outputs(743) <= not(inputs(157)) or (inputs(79));
    layer0_outputs(744) <= not(inputs(121));
    layer0_outputs(745) <= (inputs(160)) or (inputs(169));
    layer0_outputs(746) <= (inputs(41)) and not (inputs(73));
    layer0_outputs(747) <= (inputs(29)) or (inputs(100));
    layer0_outputs(748) <= '0';
    layer0_outputs(749) <= inputs(245);
    layer0_outputs(750) <= (inputs(113)) or (inputs(101));
    layer0_outputs(751) <= inputs(93);
    layer0_outputs(752) <= inputs(103);
    layer0_outputs(753) <= '0';
    layer0_outputs(754) <= not(inputs(193));
    layer0_outputs(755) <= not(inputs(125)) or (inputs(150));
    layer0_outputs(756) <= not((inputs(61)) or (inputs(35)));
    layer0_outputs(757) <= '0';
    layer0_outputs(758) <= not(inputs(85)) or (inputs(197));
    layer0_outputs(759) <= not(inputs(187)) or (inputs(20));
    layer0_outputs(760) <= not(inputs(145));
    layer0_outputs(761) <= '1';
    layer0_outputs(762) <= (inputs(171)) or (inputs(37));
    layer0_outputs(763) <= not((inputs(5)) and (inputs(120)));
    layer0_outputs(764) <= inputs(206);
    layer0_outputs(765) <= not((inputs(13)) and (inputs(51)));
    layer0_outputs(766) <= inputs(194);
    layer0_outputs(767) <= (inputs(127)) or (inputs(110));
    layer0_outputs(768) <= (inputs(35)) and not (inputs(161));
    layer0_outputs(769) <= (inputs(238)) xor (inputs(135));
    layer0_outputs(770) <= not(inputs(161)) or (inputs(237));
    layer0_outputs(771) <= not((inputs(57)) xor (inputs(148)));
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= (inputs(70)) and not (inputs(1));
    layer0_outputs(774) <= inputs(10);
    layer0_outputs(775) <= inputs(33);
    layer0_outputs(776) <= not((inputs(113)) and (inputs(110)));
    layer0_outputs(777) <= inputs(20);
    layer0_outputs(778) <= inputs(37);
    layer0_outputs(779) <= (inputs(76)) or (inputs(123));
    layer0_outputs(780) <= inputs(234);
    layer0_outputs(781) <= not(inputs(163)) or (inputs(176));
    layer0_outputs(782) <= (inputs(198)) or (inputs(198));
    layer0_outputs(783) <= (inputs(157)) or (inputs(253));
    layer0_outputs(784) <= (inputs(195)) and not (inputs(113));
    layer0_outputs(785) <= (inputs(26)) and not (inputs(17));
    layer0_outputs(786) <= '0';
    layer0_outputs(787) <= not((inputs(203)) or (inputs(220)));
    layer0_outputs(788) <= not(inputs(219));
    layer0_outputs(789) <= inputs(139);
    layer0_outputs(790) <= inputs(179);
    layer0_outputs(791) <= inputs(217);
    layer0_outputs(792) <= not(inputs(129)) or (inputs(161));
    layer0_outputs(793) <= (inputs(151)) and not (inputs(73));
    layer0_outputs(794) <= not((inputs(171)) or (inputs(116)));
    layer0_outputs(795) <= inputs(89);
    layer0_outputs(796) <= (inputs(20)) and not (inputs(113));
    layer0_outputs(797) <= (inputs(122)) and not (inputs(90));
    layer0_outputs(798) <= not(inputs(217)) or (inputs(154));
    layer0_outputs(799) <= inputs(192);
    layer0_outputs(800) <= inputs(204);
    layer0_outputs(801) <= '1';
    layer0_outputs(802) <= '0';
    layer0_outputs(803) <= '0';
    layer0_outputs(804) <= not(inputs(232));
    layer0_outputs(805) <= (inputs(90)) or (inputs(141));
    layer0_outputs(806) <= not((inputs(228)) or (inputs(33)));
    layer0_outputs(807) <= inputs(94);
    layer0_outputs(808) <= (inputs(227)) and not (inputs(89));
    layer0_outputs(809) <= not((inputs(38)) and (inputs(117)));
    layer0_outputs(810) <= '1';
    layer0_outputs(811) <= not(inputs(4)) or (inputs(28));
    layer0_outputs(812) <= inputs(25);
    layer0_outputs(813) <= not((inputs(129)) xor (inputs(112)));
    layer0_outputs(814) <= not(inputs(180)) or (inputs(109));
    layer0_outputs(815) <= (inputs(47)) or (inputs(111));
    layer0_outputs(816) <= not((inputs(223)) xor (inputs(84)));
    layer0_outputs(817) <= (inputs(151)) and (inputs(10));
    layer0_outputs(818) <= inputs(154);
    layer0_outputs(819) <= (inputs(185)) and (inputs(231));
    layer0_outputs(820) <= not(inputs(182));
    layer0_outputs(821) <= (inputs(135)) and (inputs(186));
    layer0_outputs(822) <= '0';
    layer0_outputs(823) <= inputs(132);
    layer0_outputs(824) <= not((inputs(246)) or (inputs(162)));
    layer0_outputs(825) <= not(inputs(198)) or (inputs(197));
    layer0_outputs(826) <= not(inputs(202)) or (inputs(46));
    layer0_outputs(827) <= (inputs(153)) and not (inputs(55));
    layer0_outputs(828) <= inputs(169);
    layer0_outputs(829) <= (inputs(198)) and not (inputs(30));
    layer0_outputs(830) <= '0';
    layer0_outputs(831) <= not((inputs(152)) xor (inputs(181)));
    layer0_outputs(832) <= (inputs(53)) xor (inputs(237));
    layer0_outputs(833) <= inputs(182);
    layer0_outputs(834) <= (inputs(226)) and not (inputs(29));
    layer0_outputs(835) <= not((inputs(130)) or (inputs(149)));
    layer0_outputs(836) <= not(inputs(133));
    layer0_outputs(837) <= inputs(254);
    layer0_outputs(838) <= (inputs(107)) and not (inputs(167));
    layer0_outputs(839) <= '0';
    layer0_outputs(840) <= (inputs(89)) or (inputs(190));
    layer0_outputs(841) <= not(inputs(105));
    layer0_outputs(842) <= '0';
    layer0_outputs(843) <= (inputs(166)) or (inputs(255));
    layer0_outputs(844) <= (inputs(155)) or (inputs(145));
    layer0_outputs(845) <= (inputs(228)) and not (inputs(109));
    layer0_outputs(846) <= (inputs(17)) and not (inputs(206));
    layer0_outputs(847) <= (inputs(22)) and not (inputs(113));
    layer0_outputs(848) <= not((inputs(93)) or (inputs(205)));
    layer0_outputs(849) <= not((inputs(218)) and (inputs(253)));
    layer0_outputs(850) <= '1';
    layer0_outputs(851) <= not(inputs(71)) or (inputs(163));
    layer0_outputs(852) <= not(inputs(169));
    layer0_outputs(853) <= (inputs(3)) and not (inputs(19));
    layer0_outputs(854) <= (inputs(142)) and not (inputs(201));
    layer0_outputs(855) <= not(inputs(210));
    layer0_outputs(856) <= not(inputs(131)) or (inputs(32));
    layer0_outputs(857) <= inputs(155);
    layer0_outputs(858) <= not(inputs(245));
    layer0_outputs(859) <= (inputs(197)) and not (inputs(131));
    layer0_outputs(860) <= not(inputs(243));
    layer0_outputs(861) <= not((inputs(148)) or (inputs(68)));
    layer0_outputs(862) <= '0';
    layer0_outputs(863) <= (inputs(99)) or (inputs(113));
    layer0_outputs(864) <= not(inputs(91));
    layer0_outputs(865) <= inputs(45);
    layer0_outputs(866) <= (inputs(66)) and (inputs(139));
    layer0_outputs(867) <= not(inputs(168));
    layer0_outputs(868) <= (inputs(39)) and (inputs(134));
    layer0_outputs(869) <= '0';
    layer0_outputs(870) <= (inputs(186)) or (inputs(140));
    layer0_outputs(871) <= not((inputs(67)) or (inputs(129)));
    layer0_outputs(872) <= not(inputs(133)) or (inputs(238));
    layer0_outputs(873) <= '0';
    layer0_outputs(874) <= not(inputs(111)) or (inputs(1));
    layer0_outputs(875) <= not(inputs(107)) or (inputs(224));
    layer0_outputs(876) <= inputs(121);
    layer0_outputs(877) <= (inputs(247)) or (inputs(190));
    layer0_outputs(878) <= (inputs(65)) and (inputs(184));
    layer0_outputs(879) <= (inputs(104)) or (inputs(252));
    layer0_outputs(880) <= not(inputs(216));
    layer0_outputs(881) <= not(inputs(191));
    layer0_outputs(882) <= not(inputs(142));
    layer0_outputs(883) <= not(inputs(141));
    layer0_outputs(884) <= not((inputs(227)) or (inputs(241)));
    layer0_outputs(885) <= '1';
    layer0_outputs(886) <= inputs(151);
    layer0_outputs(887) <= not((inputs(62)) and (inputs(58)));
    layer0_outputs(888) <= (inputs(224)) and (inputs(94));
    layer0_outputs(889) <= not(inputs(197)) or (inputs(32));
    layer0_outputs(890) <= '1';
    layer0_outputs(891) <= not((inputs(29)) and (inputs(67)));
    layer0_outputs(892) <= (inputs(24)) and (inputs(228));
    layer0_outputs(893) <= not((inputs(188)) and (inputs(153)));
    layer0_outputs(894) <= not(inputs(76));
    layer0_outputs(895) <= inputs(21);
    layer0_outputs(896) <= not((inputs(176)) or (inputs(109)));
    layer0_outputs(897) <= inputs(253);
    layer0_outputs(898) <= (inputs(7)) xor (inputs(82));
    layer0_outputs(899) <= not((inputs(107)) and (inputs(17)));
    layer0_outputs(900) <= (inputs(19)) and not (inputs(177));
    layer0_outputs(901) <= not(inputs(150));
    layer0_outputs(902) <= (inputs(207)) or (inputs(209));
    layer0_outputs(903) <= inputs(219);
    layer0_outputs(904) <= (inputs(11)) or (inputs(203));
    layer0_outputs(905) <= (inputs(193)) and not (inputs(42));
    layer0_outputs(906) <= not((inputs(182)) or (inputs(254)));
    layer0_outputs(907) <= not(inputs(157)) or (inputs(7));
    layer0_outputs(908) <= '1';
    layer0_outputs(909) <= not(inputs(74));
    layer0_outputs(910) <= inputs(45);
    layer0_outputs(911) <= not(inputs(26));
    layer0_outputs(912) <= not((inputs(202)) or (inputs(1)));
    layer0_outputs(913) <= not(inputs(182)) or (inputs(20));
    layer0_outputs(914) <= not(inputs(13));
    layer0_outputs(915) <= inputs(23);
    layer0_outputs(916) <= inputs(75);
    layer0_outputs(917) <= not((inputs(101)) or (inputs(117)));
    layer0_outputs(918) <= '0';
    layer0_outputs(919) <= not((inputs(194)) or (inputs(33)));
    layer0_outputs(920) <= not(inputs(174));
    layer0_outputs(921) <= inputs(37);
    layer0_outputs(922) <= (inputs(24)) or (inputs(35));
    layer0_outputs(923) <= '0';
    layer0_outputs(924) <= not((inputs(78)) and (inputs(211)));
    layer0_outputs(925) <= not((inputs(87)) and (inputs(130)));
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= not((inputs(127)) or (inputs(59)));
    layer0_outputs(928) <= (inputs(195)) and not (inputs(51));
    layer0_outputs(929) <= inputs(154);
    layer0_outputs(930) <= not(inputs(206)) or (inputs(215));
    layer0_outputs(931) <= not((inputs(69)) or (inputs(64)));
    layer0_outputs(932) <= not((inputs(73)) or (inputs(111)));
    layer0_outputs(933) <= inputs(67);
    layer0_outputs(934) <= (inputs(37)) or (inputs(75));
    layer0_outputs(935) <= not(inputs(160));
    layer0_outputs(936) <= '1';
    layer0_outputs(937) <= (inputs(67)) and not (inputs(182));
    layer0_outputs(938) <= not((inputs(151)) and (inputs(142)));
    layer0_outputs(939) <= not((inputs(44)) or (inputs(49)));
    layer0_outputs(940) <= not(inputs(155)) or (inputs(32));
    layer0_outputs(941) <= inputs(76);
    layer0_outputs(942) <= inputs(160);
    layer0_outputs(943) <= '0';
    layer0_outputs(944) <= inputs(66);
    layer0_outputs(945) <= inputs(144);
    layer0_outputs(946) <= not(inputs(254));
    layer0_outputs(947) <= '1';
    layer0_outputs(948) <= '0';
    layer0_outputs(949) <= not(inputs(121));
    layer0_outputs(950) <= not((inputs(232)) or (inputs(161)));
    layer0_outputs(951) <= (inputs(17)) and (inputs(238));
    layer0_outputs(952) <= (inputs(235)) or (inputs(208));
    layer0_outputs(953) <= not(inputs(37));
    layer0_outputs(954) <= not(inputs(91)) or (inputs(129));
    layer0_outputs(955) <= not((inputs(19)) and (inputs(17)));
    layer0_outputs(956) <= '1';
    layer0_outputs(957) <= not(inputs(221)) or (inputs(160));
    layer0_outputs(958) <= '0';
    layer0_outputs(959) <= (inputs(149)) or (inputs(71));
    layer0_outputs(960) <= not((inputs(43)) or (inputs(132)));
    layer0_outputs(961) <= not((inputs(63)) xor (inputs(167)));
    layer0_outputs(962) <= (inputs(237)) or (inputs(123));
    layer0_outputs(963) <= '1';
    layer0_outputs(964) <= not(inputs(128));
    layer0_outputs(965) <= inputs(109);
    layer0_outputs(966) <= (inputs(162)) and not (inputs(49));
    layer0_outputs(967) <= (inputs(93)) xor (inputs(123));
    layer0_outputs(968) <= (inputs(116)) and not (inputs(127));
    layer0_outputs(969) <= inputs(43);
    layer0_outputs(970) <= not(inputs(156));
    layer0_outputs(971) <= (inputs(40)) and (inputs(182));
    layer0_outputs(972) <= not(inputs(131));
    layer0_outputs(973) <= not(inputs(154));
    layer0_outputs(974) <= (inputs(244)) and not (inputs(51));
    layer0_outputs(975) <= '0';
    layer0_outputs(976) <= '1';
    layer0_outputs(977) <= not(inputs(109));
    layer0_outputs(978) <= not((inputs(179)) and (inputs(48)));
    layer0_outputs(979) <= '0';
    layer0_outputs(980) <= not(inputs(179));
    layer0_outputs(981) <= '0';
    layer0_outputs(982) <= '0';
    layer0_outputs(983) <= not(inputs(214)) or (inputs(122));
    layer0_outputs(984) <= not(inputs(102)) or (inputs(238));
    layer0_outputs(985) <= inputs(65);
    layer0_outputs(986) <= not(inputs(173));
    layer0_outputs(987) <= not(inputs(187));
    layer0_outputs(988) <= (inputs(157)) or (inputs(3));
    layer0_outputs(989) <= (inputs(36)) and (inputs(16));
    layer0_outputs(990) <= not(inputs(68));
    layer0_outputs(991) <= not((inputs(110)) and (inputs(222)));
    layer0_outputs(992) <= inputs(166);
    layer0_outputs(993) <= inputs(240);
    layer0_outputs(994) <= not(inputs(90));
    layer0_outputs(995) <= inputs(121);
    layer0_outputs(996) <= '1';
    layer0_outputs(997) <= not((inputs(206)) xor (inputs(157)));
    layer0_outputs(998) <= not(inputs(69)) or (inputs(159));
    layer0_outputs(999) <= (inputs(48)) and (inputs(123));
    layer0_outputs(1000) <= '1';
    layer0_outputs(1001) <= (inputs(145)) and not (inputs(133));
    layer0_outputs(1002) <= (inputs(245)) and not (inputs(105));
    layer0_outputs(1003) <= '0';
    layer0_outputs(1004) <= '0';
    layer0_outputs(1005) <= (inputs(28)) or (inputs(16));
    layer0_outputs(1006) <= inputs(184);
    layer0_outputs(1007) <= '0';
    layer0_outputs(1008) <= not(inputs(115));
    layer0_outputs(1009) <= not(inputs(186));
    layer0_outputs(1010) <= not(inputs(209));
    layer0_outputs(1011) <= (inputs(34)) or (inputs(229));
    layer0_outputs(1012) <= inputs(168);
    layer0_outputs(1013) <= (inputs(9)) and not (inputs(241));
    layer0_outputs(1014) <= not(inputs(204)) or (inputs(178));
    layer0_outputs(1015) <= not(inputs(35));
    layer0_outputs(1016) <= inputs(215);
    layer0_outputs(1017) <= (inputs(163)) and not (inputs(37));
    layer0_outputs(1018) <= (inputs(109)) and not (inputs(11));
    layer0_outputs(1019) <= not(inputs(151)) or (inputs(226));
    layer0_outputs(1020) <= not((inputs(58)) or (inputs(245)));
    layer0_outputs(1021) <= '1';
    layer0_outputs(1022) <= inputs(128);
    layer0_outputs(1023) <= '1';
    layer0_outputs(1024) <= not(inputs(182));
    layer0_outputs(1025) <= not(inputs(199)) or (inputs(106));
    layer0_outputs(1026) <= not(inputs(152));
    layer0_outputs(1027) <= inputs(122);
    layer0_outputs(1028) <= (inputs(208)) or (inputs(48));
    layer0_outputs(1029) <= (inputs(125)) or (inputs(10));
    layer0_outputs(1030) <= '1';
    layer0_outputs(1031) <= not(inputs(103));
    layer0_outputs(1032) <= (inputs(230)) or (inputs(206));
    layer0_outputs(1033) <= (inputs(73)) and not (inputs(217));
    layer0_outputs(1034) <= '0';
    layer0_outputs(1035) <= not(inputs(82));
    layer0_outputs(1036) <= inputs(59);
    layer0_outputs(1037) <= not((inputs(199)) and (inputs(110)));
    layer0_outputs(1038) <= not((inputs(137)) or (inputs(148)));
    layer0_outputs(1039) <= inputs(228);
    layer0_outputs(1040) <= not(inputs(164));
    layer0_outputs(1041) <= inputs(18);
    layer0_outputs(1042) <= not((inputs(61)) or (inputs(207)));
    layer0_outputs(1043) <= not(inputs(215));
    layer0_outputs(1044) <= not((inputs(198)) or (inputs(85)));
    layer0_outputs(1045) <= (inputs(83)) and not (inputs(27));
    layer0_outputs(1046) <= not(inputs(208)) or (inputs(227));
    layer0_outputs(1047) <= not(inputs(155)) or (inputs(101));
    layer0_outputs(1048) <= not(inputs(59)) or (inputs(214));
    layer0_outputs(1049) <= '0';
    layer0_outputs(1050) <= not(inputs(87)) or (inputs(48));
    layer0_outputs(1051) <= not(inputs(122)) or (inputs(16));
    layer0_outputs(1052) <= (inputs(1)) and not (inputs(80));
    layer0_outputs(1053) <= inputs(74);
    layer0_outputs(1054) <= (inputs(143)) xor (inputs(125));
    layer0_outputs(1055) <= not((inputs(236)) or (inputs(60)));
    layer0_outputs(1056) <= (inputs(96)) xor (inputs(181));
    layer0_outputs(1057) <= not((inputs(2)) or (inputs(4)));
    layer0_outputs(1058) <= inputs(239);
    layer0_outputs(1059) <= inputs(213);
    layer0_outputs(1060) <= not((inputs(26)) and (inputs(66)));
    layer0_outputs(1061) <= not(inputs(44));
    layer0_outputs(1062) <= (inputs(117)) or (inputs(133));
    layer0_outputs(1063) <= not((inputs(164)) or (inputs(237)));
    layer0_outputs(1064) <= not(inputs(115));
    layer0_outputs(1065) <= not(inputs(132));
    layer0_outputs(1066) <= (inputs(156)) and not (inputs(96));
    layer0_outputs(1067) <= not(inputs(82)) or (inputs(239));
    layer0_outputs(1068) <= inputs(82);
    layer0_outputs(1069) <= (inputs(56)) and (inputs(216));
    layer0_outputs(1070) <= (inputs(142)) and not (inputs(95));
    layer0_outputs(1071) <= inputs(72);
    layer0_outputs(1072) <= inputs(200);
    layer0_outputs(1073) <= not(inputs(233));
    layer0_outputs(1074) <= '1';
    layer0_outputs(1075) <= inputs(104);
    layer0_outputs(1076) <= '1';
    layer0_outputs(1077) <= not(inputs(119));
    layer0_outputs(1078) <= not(inputs(114));
    layer0_outputs(1079) <= inputs(90);
    layer0_outputs(1080) <= '1';
    layer0_outputs(1081) <= inputs(90);
    layer0_outputs(1082) <= not((inputs(214)) or (inputs(78)));
    layer0_outputs(1083) <= not(inputs(241));
    layer0_outputs(1084) <= not((inputs(75)) or (inputs(115)));
    layer0_outputs(1085) <= '0';
    layer0_outputs(1086) <= (inputs(22)) and not (inputs(179));
    layer0_outputs(1087) <= '0';
    layer0_outputs(1088) <= inputs(121);
    layer0_outputs(1089) <= (inputs(125)) and not (inputs(221));
    layer0_outputs(1090) <= (inputs(234)) or (inputs(227));
    layer0_outputs(1091) <= not((inputs(70)) or (inputs(83)));
    layer0_outputs(1092) <= not(inputs(195));
    layer0_outputs(1093) <= (inputs(2)) or (inputs(164));
    layer0_outputs(1094) <= inputs(20);
    layer0_outputs(1095) <= inputs(249);
    layer0_outputs(1096) <= not(inputs(119));
    layer0_outputs(1097) <= not((inputs(168)) or (inputs(137)));
    layer0_outputs(1098) <= not(inputs(167));
    layer0_outputs(1099) <= not(inputs(37));
    layer0_outputs(1100) <= '1';
    layer0_outputs(1101) <= (inputs(182)) and (inputs(147));
    layer0_outputs(1102) <= inputs(132);
    layer0_outputs(1103) <= '0';
    layer0_outputs(1104) <= (inputs(195)) or (inputs(98));
    layer0_outputs(1105) <= not((inputs(252)) or (inputs(166)));
    layer0_outputs(1106) <= (inputs(51)) and (inputs(168));
    layer0_outputs(1107) <= inputs(168);
    layer0_outputs(1108) <= (inputs(159)) and not (inputs(191));
    layer0_outputs(1109) <= '0';
    layer0_outputs(1110) <= not(inputs(17));
    layer0_outputs(1111) <= not((inputs(115)) or (inputs(113)));
    layer0_outputs(1112) <= (inputs(153)) and not (inputs(235));
    layer0_outputs(1113) <= (inputs(103)) or (inputs(30));
    layer0_outputs(1114) <= inputs(142);
    layer0_outputs(1115) <= not(inputs(59));
    layer0_outputs(1116) <= not(inputs(46)) or (inputs(251));
    layer0_outputs(1117) <= (inputs(71)) xor (inputs(224));
    layer0_outputs(1118) <= not(inputs(24));
    layer0_outputs(1119) <= (inputs(165)) or (inputs(101));
    layer0_outputs(1120) <= inputs(246);
    layer0_outputs(1121) <= not(inputs(82)) or (inputs(170));
    layer0_outputs(1122) <= '1';
    layer0_outputs(1123) <= not((inputs(178)) xor (inputs(131)));
    layer0_outputs(1124) <= not((inputs(180)) or (inputs(162)));
    layer0_outputs(1125) <= not(inputs(205)) or (inputs(81));
    layer0_outputs(1126) <= (inputs(224)) and (inputs(170));
    layer0_outputs(1127) <= not(inputs(179)) or (inputs(39));
    layer0_outputs(1128) <= not(inputs(232)) or (inputs(168));
    layer0_outputs(1129) <= inputs(106);
    layer0_outputs(1130) <= (inputs(147)) and not (inputs(108));
    layer0_outputs(1131) <= not(inputs(253));
    layer0_outputs(1132) <= not(inputs(233)) or (inputs(61));
    layer0_outputs(1133) <= (inputs(171)) and (inputs(88));
    layer0_outputs(1134) <= not((inputs(117)) and (inputs(153)));
    layer0_outputs(1135) <= not(inputs(109));
    layer0_outputs(1136) <= not((inputs(71)) xor (inputs(148)));
    layer0_outputs(1137) <= inputs(29);
    layer0_outputs(1138) <= not(inputs(179));
    layer0_outputs(1139) <= not((inputs(112)) or (inputs(247)));
    layer0_outputs(1140) <= not(inputs(241));
    layer0_outputs(1141) <= '0';
    layer0_outputs(1142) <= inputs(43);
    layer0_outputs(1143) <= (inputs(243)) and (inputs(190));
    layer0_outputs(1144) <= not(inputs(79));
    layer0_outputs(1145) <= (inputs(72)) and (inputs(216));
    layer0_outputs(1146) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(1147) <= not(inputs(239)) or (inputs(175));
    layer0_outputs(1148) <= not((inputs(86)) or (inputs(191)));
    layer0_outputs(1149) <= (inputs(76)) and not (inputs(58));
    layer0_outputs(1150) <= (inputs(107)) xor (inputs(111));
    layer0_outputs(1151) <= (inputs(96)) or (inputs(42));
    layer0_outputs(1152) <= not(inputs(26)) or (inputs(88));
    layer0_outputs(1153) <= not(inputs(158)) or (inputs(185));
    layer0_outputs(1154) <= not((inputs(202)) and (inputs(199)));
    layer0_outputs(1155) <= (inputs(245)) or (inputs(192));
    layer0_outputs(1156) <= (inputs(165)) and (inputs(185));
    layer0_outputs(1157) <= '1';
    layer0_outputs(1158) <= '0';
    layer0_outputs(1159) <= '0';
    layer0_outputs(1160) <= inputs(150);
    layer0_outputs(1161) <= not(inputs(117));
    layer0_outputs(1162) <= not((inputs(210)) or (inputs(126)));
    layer0_outputs(1163) <= (inputs(204)) or (inputs(133));
    layer0_outputs(1164) <= not((inputs(108)) and (inputs(213)));
    layer0_outputs(1165) <= inputs(199);
    layer0_outputs(1166) <= '1';
    layer0_outputs(1167) <= inputs(73);
    layer0_outputs(1168) <= '0';
    layer0_outputs(1169) <= inputs(163);
    layer0_outputs(1170) <= (inputs(38)) xor (inputs(6));
    layer0_outputs(1171) <= not((inputs(30)) and (inputs(95)));
    layer0_outputs(1172) <= '0';
    layer0_outputs(1173) <= (inputs(191)) or (inputs(143));
    layer0_outputs(1174) <= '0';
    layer0_outputs(1175) <= not((inputs(112)) and (inputs(83)));
    layer0_outputs(1176) <= (inputs(232)) and (inputs(204));
    layer0_outputs(1177) <= inputs(61);
    layer0_outputs(1178) <= '1';
    layer0_outputs(1179) <= not(inputs(115));
    layer0_outputs(1180) <= inputs(201);
    layer0_outputs(1181) <= (inputs(188)) and not (inputs(46));
    layer0_outputs(1182) <= not(inputs(192));
    layer0_outputs(1183) <= '0';
    layer0_outputs(1184) <= not(inputs(89));
    layer0_outputs(1185) <= inputs(18);
    layer0_outputs(1186) <= not((inputs(19)) or (inputs(227)));
    layer0_outputs(1187) <= (inputs(206)) and not (inputs(214));
    layer0_outputs(1188) <= '1';
    layer0_outputs(1189) <= '0';
    layer0_outputs(1190) <= inputs(50);
    layer0_outputs(1191) <= not((inputs(198)) and (inputs(166)));
    layer0_outputs(1192) <= not((inputs(191)) xor (inputs(89)));
    layer0_outputs(1193) <= not(inputs(169));
    layer0_outputs(1194) <= (inputs(39)) and not (inputs(150));
    layer0_outputs(1195) <= '1';
    layer0_outputs(1196) <= not(inputs(215)) or (inputs(18));
    layer0_outputs(1197) <= not((inputs(123)) and (inputs(105)));
    layer0_outputs(1198) <= not(inputs(196));
    layer0_outputs(1199) <= (inputs(126)) and not (inputs(124));
    layer0_outputs(1200) <= (inputs(29)) and not (inputs(244));
    layer0_outputs(1201) <= not(inputs(193));
    layer0_outputs(1202) <= (inputs(92)) and (inputs(132));
    layer0_outputs(1203) <= inputs(108);
    layer0_outputs(1204) <= inputs(201);
    layer0_outputs(1205) <= inputs(3);
    layer0_outputs(1206) <= '1';
    layer0_outputs(1207) <= (inputs(231)) and (inputs(234));
    layer0_outputs(1208) <= (inputs(238)) or (inputs(20));
    layer0_outputs(1209) <= inputs(194);
    layer0_outputs(1210) <= (inputs(121)) and (inputs(152));
    layer0_outputs(1211) <= not(inputs(252));
    layer0_outputs(1212) <= not(inputs(48)) or (inputs(140));
    layer0_outputs(1213) <= (inputs(24)) and not (inputs(15));
    layer0_outputs(1214) <= '1';
    layer0_outputs(1215) <= (inputs(23)) and not (inputs(184));
    layer0_outputs(1216) <= not(inputs(68));
    layer0_outputs(1217) <= not(inputs(161)) or (inputs(166));
    layer0_outputs(1218) <= not(inputs(215));
    layer0_outputs(1219) <= (inputs(213)) and not (inputs(237));
    layer0_outputs(1220) <= not((inputs(86)) and (inputs(27)));
    layer0_outputs(1221) <= inputs(62);
    layer0_outputs(1222) <= not((inputs(98)) and (inputs(242)));
    layer0_outputs(1223) <= (inputs(130)) or (inputs(61));
    layer0_outputs(1224) <= '1';
    layer0_outputs(1225) <= inputs(188);
    layer0_outputs(1226) <= not(inputs(224));
    layer0_outputs(1227) <= '0';
    layer0_outputs(1228) <= '1';
    layer0_outputs(1229) <= (inputs(117)) or (inputs(96));
    layer0_outputs(1230) <= inputs(121);
    layer0_outputs(1231) <= not(inputs(128)) or (inputs(90));
    layer0_outputs(1232) <= not(inputs(62)) or (inputs(101));
    layer0_outputs(1233) <= not((inputs(113)) or (inputs(142)));
    layer0_outputs(1234) <= not(inputs(93)) or (inputs(203));
    layer0_outputs(1235) <= (inputs(172)) and (inputs(231));
    layer0_outputs(1236) <= inputs(97);
    layer0_outputs(1237) <= not(inputs(194));
    layer0_outputs(1238) <= not((inputs(162)) or (inputs(73)));
    layer0_outputs(1239) <= '1';
    layer0_outputs(1240) <= (inputs(223)) or (inputs(114));
    layer0_outputs(1241) <= inputs(130);
    layer0_outputs(1242) <= not((inputs(36)) or (inputs(39)));
    layer0_outputs(1243) <= not(inputs(232));
    layer0_outputs(1244) <= (inputs(13)) or (inputs(160));
    layer0_outputs(1245) <= (inputs(233)) or (inputs(139));
    layer0_outputs(1246) <= not(inputs(209)) or (inputs(33));
    layer0_outputs(1247) <= (inputs(170)) or (inputs(255));
    layer0_outputs(1248) <= inputs(171);
    layer0_outputs(1249) <= not((inputs(232)) and (inputs(1)));
    layer0_outputs(1250) <= (inputs(224)) or (inputs(204));
    layer0_outputs(1251) <= inputs(177);
    layer0_outputs(1252) <= not((inputs(175)) xor (inputs(53)));
    layer0_outputs(1253) <= (inputs(75)) and not (inputs(178));
    layer0_outputs(1254) <= not(inputs(170)) or (inputs(208));
    layer0_outputs(1255) <= (inputs(122)) or (inputs(160));
    layer0_outputs(1256) <= '0';
    layer0_outputs(1257) <= not(inputs(128));
    layer0_outputs(1258) <= (inputs(118)) or (inputs(146));
    layer0_outputs(1259) <= (inputs(127)) or (inputs(87));
    layer0_outputs(1260) <= not(inputs(26)) or (inputs(81));
    layer0_outputs(1261) <= not(inputs(227)) or (inputs(99));
    layer0_outputs(1262) <= not((inputs(130)) or (inputs(214)));
    layer0_outputs(1263) <= not(inputs(85));
    layer0_outputs(1264) <= (inputs(9)) and (inputs(233));
    layer0_outputs(1265) <= inputs(97);
    layer0_outputs(1266) <= (inputs(12)) and (inputs(32));
    layer0_outputs(1267) <= (inputs(128)) and not (inputs(76));
    layer0_outputs(1268) <= (inputs(227)) or (inputs(217));
    layer0_outputs(1269) <= (inputs(122)) and not (inputs(1));
    layer0_outputs(1270) <= (inputs(241)) or (inputs(57));
    layer0_outputs(1271) <= '1';
    layer0_outputs(1272) <= '1';
    layer0_outputs(1273) <= (inputs(145)) and (inputs(4));
    layer0_outputs(1274) <= inputs(217);
    layer0_outputs(1275) <= (inputs(36)) and not (inputs(111));
    layer0_outputs(1276) <= '0';
    layer0_outputs(1277) <= '0';
    layer0_outputs(1278) <= not(inputs(179));
    layer0_outputs(1279) <= (inputs(34)) and not (inputs(237));
    layer0_outputs(1280) <= inputs(169);
    layer0_outputs(1281) <= not((inputs(37)) and (inputs(102)));
    layer0_outputs(1282) <= (inputs(191)) and (inputs(231));
    layer0_outputs(1283) <= not(inputs(104)) or (inputs(158));
    layer0_outputs(1284) <= (inputs(226)) or (inputs(193));
    layer0_outputs(1285) <= not(inputs(90));
    layer0_outputs(1286) <= inputs(138);
    layer0_outputs(1287) <= (inputs(145)) xor (inputs(0));
    layer0_outputs(1288) <= (inputs(175)) xor (inputs(156));
    layer0_outputs(1289) <= not(inputs(166));
    layer0_outputs(1290) <= '0';
    layer0_outputs(1291) <= not(inputs(38)) or (inputs(29));
    layer0_outputs(1292) <= not(inputs(72));
    layer0_outputs(1293) <= (inputs(15)) and (inputs(7));
    layer0_outputs(1294) <= not((inputs(214)) or (inputs(189)));
    layer0_outputs(1295) <= (inputs(233)) and not (inputs(0));
    layer0_outputs(1296) <= not(inputs(143)) or (inputs(251));
    layer0_outputs(1297) <= not(inputs(35));
    layer0_outputs(1298) <= inputs(122);
    layer0_outputs(1299) <= not(inputs(25));
    layer0_outputs(1300) <= inputs(99);
    layer0_outputs(1301) <= (inputs(196)) and not (inputs(249));
    layer0_outputs(1302) <= (inputs(80)) xor (inputs(11));
    layer0_outputs(1303) <= not((inputs(195)) or (inputs(140)));
    layer0_outputs(1304) <= not(inputs(114));
    layer0_outputs(1305) <= (inputs(212)) or (inputs(103));
    layer0_outputs(1306) <= not(inputs(187)) or (inputs(175));
    layer0_outputs(1307) <= not((inputs(28)) or (inputs(194)));
    layer0_outputs(1308) <= (inputs(239)) xor (inputs(63));
    layer0_outputs(1309) <= not(inputs(251));
    layer0_outputs(1310) <= '0';
    layer0_outputs(1311) <= not((inputs(252)) or (inputs(62)));
    layer0_outputs(1312) <= '0';
    layer0_outputs(1313) <= (inputs(166)) and not (inputs(69));
    layer0_outputs(1314) <= inputs(56);
    layer0_outputs(1315) <= inputs(8);
    layer0_outputs(1316) <= not((inputs(236)) or (inputs(137)));
    layer0_outputs(1317) <= not((inputs(62)) xor (inputs(234)));
    layer0_outputs(1318) <= (inputs(93)) or (inputs(0));
    layer0_outputs(1319) <= not((inputs(92)) and (inputs(14)));
    layer0_outputs(1320) <= not((inputs(43)) or (inputs(75)));
    layer0_outputs(1321) <= inputs(23);
    layer0_outputs(1322) <= inputs(139);
    layer0_outputs(1323) <= inputs(104);
    layer0_outputs(1324) <= (inputs(38)) and not (inputs(233));
    layer0_outputs(1325) <= inputs(44);
    layer0_outputs(1326) <= (inputs(135)) and not (inputs(177));
    layer0_outputs(1327) <= not(inputs(155)) or (inputs(214));
    layer0_outputs(1328) <= not((inputs(76)) or (inputs(120)));
    layer0_outputs(1329) <= '1';
    layer0_outputs(1330) <= '1';
    layer0_outputs(1331) <= not((inputs(139)) or (inputs(69)));
    layer0_outputs(1332) <= not(inputs(4)) or (inputs(214));
    layer0_outputs(1333) <= not((inputs(80)) xor (inputs(69)));
    layer0_outputs(1334) <= not(inputs(239));
    layer0_outputs(1335) <= (inputs(38)) or (inputs(160));
    layer0_outputs(1336) <= (inputs(253)) and not (inputs(196));
    layer0_outputs(1337) <= not(inputs(23));
    layer0_outputs(1338) <= inputs(24);
    layer0_outputs(1339) <= inputs(173);
    layer0_outputs(1340) <= (inputs(147)) and (inputs(144));
    layer0_outputs(1341) <= not(inputs(5)) or (inputs(194));
    layer0_outputs(1342) <= not(inputs(146)) or (inputs(116));
    layer0_outputs(1343) <= '0';
    layer0_outputs(1344) <= inputs(170);
    layer0_outputs(1345) <= not((inputs(87)) xor (inputs(227)));
    layer0_outputs(1346) <= inputs(154);
    layer0_outputs(1347) <= inputs(155);
    layer0_outputs(1348) <= (inputs(188)) and not (inputs(253));
    layer0_outputs(1349) <= inputs(150);
    layer0_outputs(1350) <= inputs(203);
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= '1';
    layer0_outputs(1353) <= inputs(42);
    layer0_outputs(1354) <= '0';
    layer0_outputs(1355) <= not((inputs(157)) or (inputs(69)));
    layer0_outputs(1356) <= not(inputs(92)) or (inputs(154));
    layer0_outputs(1357) <= not((inputs(220)) or (inputs(212)));
    layer0_outputs(1358) <= not(inputs(226)) or (inputs(102));
    layer0_outputs(1359) <= not(inputs(50)) or (inputs(207));
    layer0_outputs(1360) <= inputs(130);
    layer0_outputs(1361) <= inputs(5);
    layer0_outputs(1362) <= inputs(36);
    layer0_outputs(1363) <= inputs(119);
    layer0_outputs(1364) <= not(inputs(215));
    layer0_outputs(1365) <= (inputs(175)) and not (inputs(232));
    layer0_outputs(1366) <= (inputs(92)) or (inputs(66));
    layer0_outputs(1367) <= (inputs(16)) or (inputs(224));
    layer0_outputs(1368) <= not((inputs(212)) and (inputs(180)));
    layer0_outputs(1369) <= not(inputs(85));
    layer0_outputs(1370) <= (inputs(76)) or (inputs(48));
    layer0_outputs(1371) <= '1';
    layer0_outputs(1372) <= not(inputs(78));
    layer0_outputs(1373) <= inputs(204);
    layer0_outputs(1374) <= not(inputs(144));
    layer0_outputs(1375) <= inputs(254);
    layer0_outputs(1376) <= (inputs(200)) and (inputs(236));
    layer0_outputs(1377) <= not(inputs(129));
    layer0_outputs(1378) <= not(inputs(255)) or (inputs(214));
    layer0_outputs(1379) <= inputs(161);
    layer0_outputs(1380) <= not(inputs(125));
    layer0_outputs(1381) <= inputs(210);
    layer0_outputs(1382) <= inputs(24);
    layer0_outputs(1383) <= not(inputs(68));
    layer0_outputs(1384) <= '1';
    layer0_outputs(1385) <= not((inputs(124)) or (inputs(37)));
    layer0_outputs(1386) <= not((inputs(49)) or (inputs(125)));
    layer0_outputs(1387) <= '0';
    layer0_outputs(1388) <= not(inputs(128));
    layer0_outputs(1389) <= not(inputs(122));
    layer0_outputs(1390) <= inputs(143);
    layer0_outputs(1391) <= inputs(116);
    layer0_outputs(1392) <= (inputs(229)) or (inputs(4));
    layer0_outputs(1393) <= not((inputs(99)) or (inputs(139)));
    layer0_outputs(1394) <= not(inputs(37)) or (inputs(115));
    layer0_outputs(1395) <= inputs(199);
    layer0_outputs(1396) <= (inputs(196)) or (inputs(211));
    layer0_outputs(1397) <= not((inputs(7)) and (inputs(193)));
    layer0_outputs(1398) <= (inputs(39)) and not (inputs(187));
    layer0_outputs(1399) <= not(inputs(209));
    layer0_outputs(1400) <= '1';
    layer0_outputs(1401) <= not(inputs(167)) or (inputs(43));
    layer0_outputs(1402) <= '0';
    layer0_outputs(1403) <= not(inputs(72)) or (inputs(190));
    layer0_outputs(1404) <= not(inputs(229));
    layer0_outputs(1405) <= inputs(122);
    layer0_outputs(1406) <= (inputs(138)) or (inputs(177));
    layer0_outputs(1407) <= not((inputs(125)) or (inputs(188)));
    layer0_outputs(1408) <= not(inputs(26));
    layer0_outputs(1409) <= '1';
    layer0_outputs(1410) <= not(inputs(159));
    layer0_outputs(1411) <= (inputs(90)) and not (inputs(235));
    layer0_outputs(1412) <= inputs(99);
    layer0_outputs(1413) <= not(inputs(100));
    layer0_outputs(1414) <= not(inputs(102));
    layer0_outputs(1415) <= '0';
    layer0_outputs(1416) <= not(inputs(180));
    layer0_outputs(1417) <= not((inputs(204)) or (inputs(196)));
    layer0_outputs(1418) <= '1';
    layer0_outputs(1419) <= (inputs(213)) or (inputs(211));
    layer0_outputs(1420) <= not(inputs(126));
    layer0_outputs(1421) <= not((inputs(88)) or (inputs(104)));
    layer0_outputs(1422) <= (inputs(160)) or (inputs(173));
    layer0_outputs(1423) <= inputs(79);
    layer0_outputs(1424) <= not(inputs(254)) or (inputs(47));
    layer0_outputs(1425) <= not(inputs(53)) or (inputs(204));
    layer0_outputs(1426) <= inputs(120);
    layer0_outputs(1427) <= '1';
    layer0_outputs(1428) <= not(inputs(146));
    layer0_outputs(1429) <= (inputs(137)) and not (inputs(170));
    layer0_outputs(1430) <= (inputs(143)) or (inputs(68));
    layer0_outputs(1431) <= inputs(27);
    layer0_outputs(1432) <= not(inputs(103));
    layer0_outputs(1433) <= not(inputs(92));
    layer0_outputs(1434) <= not(inputs(159)) or (inputs(231));
    layer0_outputs(1435) <= not(inputs(84));
    layer0_outputs(1436) <= not(inputs(246));
    layer0_outputs(1437) <= '1';
    layer0_outputs(1438) <= not((inputs(50)) or (inputs(92)));
    layer0_outputs(1439) <= inputs(146);
    layer0_outputs(1440) <= not(inputs(119)) or (inputs(117));
    layer0_outputs(1441) <= not(inputs(177)) or (inputs(1));
    layer0_outputs(1442) <= not(inputs(37));
    layer0_outputs(1443) <= (inputs(128)) or (inputs(89));
    layer0_outputs(1444) <= inputs(59);
    layer0_outputs(1445) <= inputs(236);
    layer0_outputs(1446) <= '1';
    layer0_outputs(1447) <= not(inputs(189));
    layer0_outputs(1448) <= inputs(147);
    layer0_outputs(1449) <= (inputs(100)) and not (inputs(32));
    layer0_outputs(1450) <= (inputs(27)) xor (inputs(231));
    layer0_outputs(1451) <= not(inputs(20));
    layer0_outputs(1452) <= not(inputs(161)) or (inputs(101));
    layer0_outputs(1453) <= inputs(99);
    layer0_outputs(1454) <= not(inputs(50)) or (inputs(98));
    layer0_outputs(1455) <= not(inputs(15)) or (inputs(110));
    layer0_outputs(1456) <= (inputs(248)) and not (inputs(185));
    layer0_outputs(1457) <= not(inputs(135));
    layer0_outputs(1458) <= inputs(255);
    layer0_outputs(1459) <= inputs(151);
    layer0_outputs(1460) <= '0';
    layer0_outputs(1461) <= not(inputs(33)) or (inputs(98));
    layer0_outputs(1462) <= not((inputs(55)) and (inputs(60)));
    layer0_outputs(1463) <= '1';
    layer0_outputs(1464) <= not(inputs(215));
    layer0_outputs(1465) <= '1';
    layer0_outputs(1466) <= (inputs(101)) or (inputs(78));
    layer0_outputs(1467) <= not(inputs(0));
    layer0_outputs(1468) <= (inputs(242)) and not (inputs(66));
    layer0_outputs(1469) <= inputs(17);
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= inputs(82);
    layer0_outputs(1472) <= (inputs(202)) and (inputs(212));
    layer0_outputs(1473) <= '0';
    layer0_outputs(1474) <= '1';
    layer0_outputs(1475) <= not((inputs(82)) or (inputs(39)));
    layer0_outputs(1476) <= inputs(243);
    layer0_outputs(1477) <= not(inputs(135)) or (inputs(113));
    layer0_outputs(1478) <= inputs(107);
    layer0_outputs(1479) <= inputs(22);
    layer0_outputs(1480) <= not(inputs(95)) or (inputs(140));
    layer0_outputs(1481) <= inputs(199);
    layer0_outputs(1482) <= not((inputs(239)) or (inputs(162)));
    layer0_outputs(1483) <= (inputs(91)) or (inputs(83));
    layer0_outputs(1484) <= inputs(150);
    layer0_outputs(1485) <= not(inputs(65));
    layer0_outputs(1486) <= inputs(176);
    layer0_outputs(1487) <= (inputs(113)) and not (inputs(228));
    layer0_outputs(1488) <= not(inputs(26));
    layer0_outputs(1489) <= inputs(250);
    layer0_outputs(1490) <= not(inputs(188)) or (inputs(139));
    layer0_outputs(1491) <= inputs(231);
    layer0_outputs(1492) <= not(inputs(131));
    layer0_outputs(1493) <= '0';
    layer0_outputs(1494) <= inputs(119);
    layer0_outputs(1495) <= (inputs(39)) and not (inputs(108));
    layer0_outputs(1496) <= not((inputs(60)) and (inputs(55)));
    layer0_outputs(1497) <= not(inputs(10)) or (inputs(42));
    layer0_outputs(1498) <= not(inputs(120)) or (inputs(231));
    layer0_outputs(1499) <= (inputs(113)) or (inputs(84));
    layer0_outputs(1500) <= not(inputs(168)) or (inputs(67));
    layer0_outputs(1501) <= not(inputs(247));
    layer0_outputs(1502) <= not((inputs(203)) xor (inputs(249)));
    layer0_outputs(1503) <= inputs(40);
    layer0_outputs(1504) <= inputs(25);
    layer0_outputs(1505) <= not(inputs(77)) or (inputs(71));
    layer0_outputs(1506) <= inputs(83);
    layer0_outputs(1507) <= (inputs(11)) and not (inputs(219));
    layer0_outputs(1508) <= inputs(99);
    layer0_outputs(1509) <= (inputs(87)) and (inputs(126));
    layer0_outputs(1510) <= inputs(233);
    layer0_outputs(1511) <= (inputs(234)) and not (inputs(135));
    layer0_outputs(1512) <= not((inputs(206)) or (inputs(173)));
    layer0_outputs(1513) <= not((inputs(111)) or (inputs(219)));
    layer0_outputs(1514) <= '0';
    layer0_outputs(1515) <= not((inputs(59)) and (inputs(39)));
    layer0_outputs(1516) <= '0';
    layer0_outputs(1517) <= (inputs(49)) or (inputs(71));
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= (inputs(8)) and not (inputs(55));
    layer0_outputs(1520) <= inputs(67);
    layer0_outputs(1521) <= not((inputs(94)) or (inputs(93)));
    layer0_outputs(1522) <= not(inputs(178));
    layer0_outputs(1523) <= '1';
    layer0_outputs(1524) <= inputs(161);
    layer0_outputs(1525) <= '0';
    layer0_outputs(1526) <= not((inputs(65)) or (inputs(63)));
    layer0_outputs(1527) <= not(inputs(35));
    layer0_outputs(1528) <= not((inputs(235)) or (inputs(233)));
    layer0_outputs(1529) <= (inputs(15)) and not (inputs(147));
    layer0_outputs(1530) <= not((inputs(245)) or (inputs(221)));
    layer0_outputs(1531) <= not((inputs(229)) xor (inputs(7)));
    layer0_outputs(1532) <= not((inputs(203)) or (inputs(144)));
    layer0_outputs(1533) <= not(inputs(220));
    layer0_outputs(1534) <= (inputs(68)) or (inputs(45));
    layer0_outputs(1535) <= not(inputs(2)) or (inputs(145));
    layer0_outputs(1536) <= not(inputs(178));
    layer0_outputs(1537) <= not((inputs(161)) or (inputs(108)));
    layer0_outputs(1538) <= not((inputs(112)) or (inputs(255)));
    layer0_outputs(1539) <= not((inputs(173)) or (inputs(130)));
    layer0_outputs(1540) <= not((inputs(2)) or (inputs(21)));
    layer0_outputs(1541) <= not(inputs(141));
    layer0_outputs(1542) <= '1';
    layer0_outputs(1543) <= '1';
    layer0_outputs(1544) <= not(inputs(195));
    layer0_outputs(1545) <= not((inputs(251)) and (inputs(3)));
    layer0_outputs(1546) <= not(inputs(222)) or (inputs(34));
    layer0_outputs(1547) <= (inputs(173)) and not (inputs(178));
    layer0_outputs(1548) <= '1';
    layer0_outputs(1549) <= (inputs(211)) and not (inputs(116));
    layer0_outputs(1550) <= not(inputs(53));
    layer0_outputs(1551) <= (inputs(199)) and not (inputs(131));
    layer0_outputs(1552) <= not(inputs(171));
    layer0_outputs(1553) <= not(inputs(8));
    layer0_outputs(1554) <= (inputs(14)) or (inputs(95));
    layer0_outputs(1555) <= inputs(130);
    layer0_outputs(1556) <= inputs(142);
    layer0_outputs(1557) <= not(inputs(137));
    layer0_outputs(1558) <= '1';
    layer0_outputs(1559) <= (inputs(22)) or (inputs(217));
    layer0_outputs(1560) <= not(inputs(46));
    layer0_outputs(1561) <= (inputs(108)) and not (inputs(166));
    layer0_outputs(1562) <= not(inputs(189));
    layer0_outputs(1563) <= inputs(76);
    layer0_outputs(1564) <= '1';
    layer0_outputs(1565) <= (inputs(9)) or (inputs(93));
    layer0_outputs(1566) <= not((inputs(6)) or (inputs(124)));
    layer0_outputs(1567) <= (inputs(159)) or (inputs(212));
    layer0_outputs(1568) <= not(inputs(102));
    layer0_outputs(1569) <= not((inputs(221)) xor (inputs(153)));
    layer0_outputs(1570) <= not((inputs(227)) or (inputs(84)));
    layer0_outputs(1571) <= not((inputs(222)) or (inputs(152)));
    layer0_outputs(1572) <= (inputs(84)) and not (inputs(145));
    layer0_outputs(1573) <= inputs(178);
    layer0_outputs(1574) <= not(inputs(211));
    layer0_outputs(1575) <= inputs(89);
    layer0_outputs(1576) <= (inputs(12)) and (inputs(216));
    layer0_outputs(1577) <= '1';
    layer0_outputs(1578) <= not(inputs(110)) or (inputs(5));
    layer0_outputs(1579) <= '1';
    layer0_outputs(1580) <= inputs(7);
    layer0_outputs(1581) <= not(inputs(158)) or (inputs(172));
    layer0_outputs(1582) <= (inputs(237)) and not (inputs(53));
    layer0_outputs(1583) <= not(inputs(206));
    layer0_outputs(1584) <= (inputs(6)) and not (inputs(22));
    layer0_outputs(1585) <= (inputs(75)) and not (inputs(111));
    layer0_outputs(1586) <= (inputs(102)) and not (inputs(189));
    layer0_outputs(1587) <= inputs(146);
    layer0_outputs(1588) <= not(inputs(17)) or (inputs(62));
    layer0_outputs(1589) <= '0';
    layer0_outputs(1590) <= not((inputs(195)) or (inputs(226)));
    layer0_outputs(1591) <= inputs(228);
    layer0_outputs(1592) <= not((inputs(126)) or (inputs(111)));
    layer0_outputs(1593) <= '0';
    layer0_outputs(1594) <= inputs(22);
    layer0_outputs(1595) <= (inputs(176)) or (inputs(163));
    layer0_outputs(1596) <= '1';
    layer0_outputs(1597) <= not((inputs(109)) or (inputs(106)));
    layer0_outputs(1598) <= inputs(41);
    layer0_outputs(1599) <= (inputs(90)) and not (inputs(193));
    layer0_outputs(1600) <= (inputs(78)) and not (inputs(39));
    layer0_outputs(1601) <= not(inputs(235));
    layer0_outputs(1602) <= not(inputs(9)) or (inputs(100));
    layer0_outputs(1603) <= not(inputs(78));
    layer0_outputs(1604) <= not(inputs(174)) or (inputs(100));
    layer0_outputs(1605) <= (inputs(185)) and not (inputs(103));
    layer0_outputs(1606) <= (inputs(23)) and not (inputs(225));
    layer0_outputs(1607) <= not((inputs(54)) or (inputs(108)));
    layer0_outputs(1608) <= not(inputs(3));
    layer0_outputs(1609) <= not((inputs(139)) or (inputs(233)));
    layer0_outputs(1610) <= not((inputs(151)) or (inputs(111)));
    layer0_outputs(1611) <= not(inputs(54));
    layer0_outputs(1612) <= (inputs(61)) or (inputs(131));
    layer0_outputs(1613) <= not(inputs(203));
    layer0_outputs(1614) <= not((inputs(220)) xor (inputs(158)));
    layer0_outputs(1615) <= (inputs(108)) or (inputs(177));
    layer0_outputs(1616) <= (inputs(44)) and not (inputs(154));
    layer0_outputs(1617) <= not((inputs(73)) xor (inputs(183)));
    layer0_outputs(1618) <= '0';
    layer0_outputs(1619) <= '1';
    layer0_outputs(1620) <= not(inputs(24));
    layer0_outputs(1621) <= '1';
    layer0_outputs(1622) <= not(inputs(67)) or (inputs(38));
    layer0_outputs(1623) <= not((inputs(51)) or (inputs(92)));
    layer0_outputs(1624) <= not(inputs(119));
    layer0_outputs(1625) <= '0';
    layer0_outputs(1626) <= (inputs(240)) or (inputs(127));
    layer0_outputs(1627) <= (inputs(200)) and not (inputs(223));
    layer0_outputs(1628) <= (inputs(14)) and not (inputs(163));
    layer0_outputs(1629) <= inputs(157);
    layer0_outputs(1630) <= not((inputs(80)) and (inputs(255)));
    layer0_outputs(1631) <= '0';
    layer0_outputs(1632) <= (inputs(201)) and (inputs(76));
    layer0_outputs(1633) <= '0';
    layer0_outputs(1634) <= '1';
    layer0_outputs(1635) <= not((inputs(57)) and (inputs(121)));
    layer0_outputs(1636) <= not(inputs(14));
    layer0_outputs(1637) <= not((inputs(156)) or (inputs(47)));
    layer0_outputs(1638) <= not((inputs(248)) and (inputs(234)));
    layer0_outputs(1639) <= not(inputs(134)) or (inputs(222));
    layer0_outputs(1640) <= inputs(49);
    layer0_outputs(1641) <= not(inputs(116)) or (inputs(241));
    layer0_outputs(1642) <= '1';
    layer0_outputs(1643) <= (inputs(195)) and not (inputs(192));
    layer0_outputs(1644) <= not(inputs(224)) or (inputs(208));
    layer0_outputs(1645) <= '0';
    layer0_outputs(1646) <= not(inputs(118)) or (inputs(34));
    layer0_outputs(1647) <= not((inputs(105)) or (inputs(237)));
    layer0_outputs(1648) <= (inputs(9)) xor (inputs(127));
    layer0_outputs(1649) <= '1';
    layer0_outputs(1650) <= (inputs(130)) or (inputs(112));
    layer0_outputs(1651) <= (inputs(107)) or (inputs(122));
    layer0_outputs(1652) <= inputs(184);
    layer0_outputs(1653) <= not(inputs(156));
    layer0_outputs(1654) <= '1';
    layer0_outputs(1655) <= inputs(5);
    layer0_outputs(1656) <= inputs(115);
    layer0_outputs(1657) <= (inputs(72)) or (inputs(249));
    layer0_outputs(1658) <= not(inputs(45)) or (inputs(242));
    layer0_outputs(1659) <= inputs(23);
    layer0_outputs(1660) <= '0';
    layer0_outputs(1661) <= not(inputs(47)) or (inputs(36));
    layer0_outputs(1662) <= (inputs(76)) and (inputs(187));
    layer0_outputs(1663) <= not(inputs(116));
    layer0_outputs(1664) <= inputs(162);
    layer0_outputs(1665) <= not(inputs(255));
    layer0_outputs(1666) <= not((inputs(173)) or (inputs(85)));
    layer0_outputs(1667) <= (inputs(87)) and not (inputs(206));
    layer0_outputs(1668) <= (inputs(91)) or (inputs(28));
    layer0_outputs(1669) <= inputs(0);
    layer0_outputs(1670) <= not(inputs(63)) or (inputs(7));
    layer0_outputs(1671) <= not(inputs(204));
    layer0_outputs(1672) <= (inputs(3)) or (inputs(5));
    layer0_outputs(1673) <= (inputs(185)) and not (inputs(208));
    layer0_outputs(1674) <= '0';
    layer0_outputs(1675) <= inputs(68);
    layer0_outputs(1676) <= inputs(19);
    layer0_outputs(1677) <= inputs(234);
    layer0_outputs(1678) <= inputs(127);
    layer0_outputs(1679) <= inputs(18);
    layer0_outputs(1680) <= not(inputs(79));
    layer0_outputs(1681) <= not(inputs(22)) or (inputs(164));
    layer0_outputs(1682) <= (inputs(181)) and (inputs(182));
    layer0_outputs(1683) <= not(inputs(175));
    layer0_outputs(1684) <= not(inputs(86)) or (inputs(220));
    layer0_outputs(1685) <= '1';
    layer0_outputs(1686) <= not(inputs(24)) or (inputs(14));
    layer0_outputs(1687) <= (inputs(44)) and (inputs(27));
    layer0_outputs(1688) <= (inputs(188)) and not (inputs(179));
    layer0_outputs(1689) <= not((inputs(163)) xor (inputs(176)));
    layer0_outputs(1690) <= (inputs(69)) and not (inputs(174));
    layer0_outputs(1691) <= not(inputs(232));
    layer0_outputs(1692) <= '0';
    layer0_outputs(1693) <= inputs(54);
    layer0_outputs(1694) <= '1';
    layer0_outputs(1695) <= '1';
    layer0_outputs(1696) <= inputs(139);
    layer0_outputs(1697) <= not((inputs(205)) or (inputs(59)));
    layer0_outputs(1698) <= not(inputs(7));
    layer0_outputs(1699) <= (inputs(216)) and not (inputs(66));
    layer0_outputs(1700) <= inputs(100);
    layer0_outputs(1701) <= (inputs(83)) xor (inputs(97));
    layer0_outputs(1702) <= not(inputs(177));
    layer0_outputs(1703) <= '0';
    layer0_outputs(1704) <= (inputs(12)) and not (inputs(223));
    layer0_outputs(1705) <= not((inputs(224)) and (inputs(100)));
    layer0_outputs(1706) <= not(inputs(89));
    layer0_outputs(1707) <= not(inputs(242)) or (inputs(247));
    layer0_outputs(1708) <= (inputs(229)) and (inputs(173));
    layer0_outputs(1709) <= '0';
    layer0_outputs(1710) <= (inputs(196)) and not (inputs(191));
    layer0_outputs(1711) <= not((inputs(21)) xor (inputs(160)));
    layer0_outputs(1712) <= not((inputs(18)) and (inputs(11)));
    layer0_outputs(1713) <= (inputs(17)) and (inputs(99));
    layer0_outputs(1714) <= '1';
    layer0_outputs(1715) <= (inputs(6)) or (inputs(48));
    layer0_outputs(1716) <= not(inputs(97));
    layer0_outputs(1717) <= not(inputs(208)) or (inputs(54));
    layer0_outputs(1718) <= (inputs(148)) or (inputs(248));
    layer0_outputs(1719) <= (inputs(32)) and not (inputs(75));
    layer0_outputs(1720) <= (inputs(53)) or (inputs(203));
    layer0_outputs(1721) <= not(inputs(149));
    layer0_outputs(1722) <= not(inputs(10)) or (inputs(251));
    layer0_outputs(1723) <= (inputs(80)) or (inputs(222));
    layer0_outputs(1724) <= (inputs(31)) and (inputs(103));
    layer0_outputs(1725) <= not(inputs(132)) or (inputs(190));
    layer0_outputs(1726) <= not(inputs(46));
    layer0_outputs(1727) <= not(inputs(228));
    layer0_outputs(1728) <= (inputs(132)) or (inputs(192));
    layer0_outputs(1729) <= '1';
    layer0_outputs(1730) <= '0';
    layer0_outputs(1731) <= not(inputs(149));
    layer0_outputs(1732) <= not(inputs(18)) or (inputs(161));
    layer0_outputs(1733) <= not((inputs(175)) xor (inputs(148)));
    layer0_outputs(1734) <= not((inputs(169)) or (inputs(45)));
    layer0_outputs(1735) <= (inputs(65)) and (inputs(242));
    layer0_outputs(1736) <= not((inputs(22)) xor (inputs(95)));
    layer0_outputs(1737) <= not((inputs(176)) and (inputs(254)));
    layer0_outputs(1738) <= not(inputs(229));
    layer0_outputs(1739) <= not(inputs(137)) or (inputs(197));
    layer0_outputs(1740) <= not((inputs(222)) or (inputs(92)));
    layer0_outputs(1741) <= inputs(15);
    layer0_outputs(1742) <= (inputs(209)) and (inputs(240));
    layer0_outputs(1743) <= inputs(61);
    layer0_outputs(1744) <= '1';
    layer0_outputs(1745) <= not(inputs(115));
    layer0_outputs(1746) <= '0';
    layer0_outputs(1747) <= not(inputs(210));
    layer0_outputs(1748) <= '0';
    layer0_outputs(1749) <= (inputs(145)) and not (inputs(255));
    layer0_outputs(1750) <= not(inputs(219)) or (inputs(77));
    layer0_outputs(1751) <= not(inputs(146));
    layer0_outputs(1752) <= '1';
    layer0_outputs(1753) <= (inputs(62)) and not (inputs(216));
    layer0_outputs(1754) <= not(inputs(94));
    layer0_outputs(1755) <= not(inputs(69));
    layer0_outputs(1756) <= not((inputs(8)) and (inputs(151)));
    layer0_outputs(1757) <= (inputs(109)) or (inputs(139));
    layer0_outputs(1758) <= '0';
    layer0_outputs(1759) <= not((inputs(117)) and (inputs(198)));
    layer0_outputs(1760) <= not((inputs(179)) and (inputs(215)));
    layer0_outputs(1761) <= not(inputs(12));
    layer0_outputs(1762) <= not(inputs(84));
    layer0_outputs(1763) <= inputs(25);
    layer0_outputs(1764) <= not(inputs(207));
    layer0_outputs(1765) <= (inputs(84)) or (inputs(124));
    layer0_outputs(1766) <= '1';
    layer0_outputs(1767) <= inputs(36);
    layer0_outputs(1768) <= '1';
    layer0_outputs(1769) <= (inputs(235)) xor (inputs(108));
    layer0_outputs(1770) <= inputs(77);
    layer0_outputs(1771) <= inputs(179);
    layer0_outputs(1772) <= (inputs(150)) or (inputs(148));
    layer0_outputs(1773) <= inputs(119);
    layer0_outputs(1774) <= inputs(143);
    layer0_outputs(1775) <= (inputs(29)) or (inputs(251));
    layer0_outputs(1776) <= not((inputs(195)) or (inputs(177)));
    layer0_outputs(1777) <= not(inputs(44));
    layer0_outputs(1778) <= '1';
    layer0_outputs(1779) <= not(inputs(5));
    layer0_outputs(1780) <= not((inputs(245)) or (inputs(56)));
    layer0_outputs(1781) <= (inputs(131)) xor (inputs(85));
    layer0_outputs(1782) <= not((inputs(52)) and (inputs(155)));
    layer0_outputs(1783) <= inputs(154);
    layer0_outputs(1784) <= (inputs(70)) or (inputs(97));
    layer0_outputs(1785) <= not(inputs(110));
    layer0_outputs(1786) <= not(inputs(92));
    layer0_outputs(1787) <= not(inputs(159));
    layer0_outputs(1788) <= inputs(164);
    layer0_outputs(1789) <= not((inputs(227)) or (inputs(226)));
    layer0_outputs(1790) <= not((inputs(112)) and (inputs(40)));
    layer0_outputs(1791) <= (inputs(11)) and (inputs(237));
    layer0_outputs(1792) <= not(inputs(123)) or (inputs(193));
    layer0_outputs(1793) <= (inputs(34)) and not (inputs(212));
    layer0_outputs(1794) <= '1';
    layer0_outputs(1795) <= '1';
    layer0_outputs(1796) <= not(inputs(65));
    layer0_outputs(1797) <= '1';
    layer0_outputs(1798) <= not((inputs(113)) or (inputs(165)));
    layer0_outputs(1799) <= not((inputs(1)) and (inputs(151)));
    layer0_outputs(1800) <= not(inputs(50));
    layer0_outputs(1801) <= (inputs(189)) or (inputs(69));
    layer0_outputs(1802) <= not((inputs(180)) or (inputs(110)));
    layer0_outputs(1803) <= (inputs(238)) or (inputs(54));
    layer0_outputs(1804) <= not(inputs(78)) or (inputs(196));
    layer0_outputs(1805) <= (inputs(73)) or (inputs(176));
    layer0_outputs(1806) <= not(inputs(171)) or (inputs(163));
    layer0_outputs(1807) <= not(inputs(75));
    layer0_outputs(1808) <= '1';
    layer0_outputs(1809) <= (inputs(23)) and (inputs(152));
    layer0_outputs(1810) <= not(inputs(128));
    layer0_outputs(1811) <= inputs(92);
    layer0_outputs(1812) <= (inputs(70)) or (inputs(13));
    layer0_outputs(1813) <= not((inputs(104)) or (inputs(88)));
    layer0_outputs(1814) <= (inputs(83)) or (inputs(147));
    layer0_outputs(1815) <= not(inputs(17));
    layer0_outputs(1816) <= (inputs(215)) and not (inputs(61));
    layer0_outputs(1817) <= inputs(6);
    layer0_outputs(1818) <= (inputs(157)) or (inputs(98));
    layer0_outputs(1819) <= (inputs(162)) or (inputs(66));
    layer0_outputs(1820) <= not(inputs(235));
    layer0_outputs(1821) <= inputs(164);
    layer0_outputs(1822) <= not(inputs(181));
    layer0_outputs(1823) <= inputs(245);
    layer0_outputs(1824) <= not(inputs(174));
    layer0_outputs(1825) <= not(inputs(59));
    layer0_outputs(1826) <= '1';
    layer0_outputs(1827) <= not((inputs(224)) or (inputs(229)));
    layer0_outputs(1828) <= inputs(97);
    layer0_outputs(1829) <= not((inputs(254)) or (inputs(152)));
    layer0_outputs(1830) <= '0';
    layer0_outputs(1831) <= not((inputs(122)) or (inputs(14)));
    layer0_outputs(1832) <= inputs(225);
    layer0_outputs(1833) <= (inputs(67)) and not (inputs(173));
    layer0_outputs(1834) <= (inputs(192)) and not (inputs(248));
    layer0_outputs(1835) <= not((inputs(175)) or (inputs(218)));
    layer0_outputs(1836) <= not((inputs(240)) and (inputs(84)));
    layer0_outputs(1837) <= (inputs(214)) and not (inputs(137));
    layer0_outputs(1838) <= inputs(74);
    layer0_outputs(1839) <= not(inputs(103)) or (inputs(202));
    layer0_outputs(1840) <= not(inputs(26));
    layer0_outputs(1841) <= not(inputs(24));
    layer0_outputs(1842) <= (inputs(101)) or (inputs(187));
    layer0_outputs(1843) <= not(inputs(184));
    layer0_outputs(1844) <= (inputs(156)) and not (inputs(86));
    layer0_outputs(1845) <= not(inputs(120)) or (inputs(98));
    layer0_outputs(1846) <= inputs(175);
    layer0_outputs(1847) <= not(inputs(25));
    layer0_outputs(1848) <= (inputs(22)) or (inputs(116));
    layer0_outputs(1849) <= (inputs(94)) and not (inputs(152));
    layer0_outputs(1850) <= inputs(166);
    layer0_outputs(1851) <= (inputs(118)) or (inputs(69));
    layer0_outputs(1852) <= '0';
    layer0_outputs(1853) <= not((inputs(144)) and (inputs(245)));
    layer0_outputs(1854) <= '0';
    layer0_outputs(1855) <= not(inputs(174)) or (inputs(12));
    layer0_outputs(1856) <= '0';
    layer0_outputs(1857) <= not((inputs(179)) or (inputs(198)));
    layer0_outputs(1858) <= inputs(70);
    layer0_outputs(1859) <= inputs(2);
    layer0_outputs(1860) <= (inputs(163)) and not (inputs(207));
    layer0_outputs(1861) <= inputs(86);
    layer0_outputs(1862) <= (inputs(27)) and (inputs(252));
    layer0_outputs(1863) <= (inputs(133)) or (inputs(40));
    layer0_outputs(1864) <= not(inputs(150));
    layer0_outputs(1865) <= not(inputs(132)) or (inputs(6));
    layer0_outputs(1866) <= (inputs(33)) or (inputs(18));
    layer0_outputs(1867) <= (inputs(9)) or (inputs(6));
    layer0_outputs(1868) <= (inputs(83)) and not (inputs(134));
    layer0_outputs(1869) <= (inputs(61)) xor (inputs(180));
    layer0_outputs(1870) <= not((inputs(140)) or (inputs(159)));
    layer0_outputs(1871) <= (inputs(96)) and not (inputs(49));
    layer0_outputs(1872) <= not(inputs(213));
    layer0_outputs(1873) <= '0';
    layer0_outputs(1874) <= not((inputs(216)) or (inputs(103)));
    layer0_outputs(1875) <= '0';
    layer0_outputs(1876) <= not(inputs(74));
    layer0_outputs(1877) <= not((inputs(27)) or (inputs(79)));
    layer0_outputs(1878) <= not(inputs(183));
    layer0_outputs(1879) <= not(inputs(44));
    layer0_outputs(1880) <= (inputs(42)) and (inputs(40));
    layer0_outputs(1881) <= not(inputs(229));
    layer0_outputs(1882) <= not(inputs(89));
    layer0_outputs(1883) <= '0';
    layer0_outputs(1884) <= not(inputs(20));
    layer0_outputs(1885) <= not((inputs(77)) or (inputs(252)));
    layer0_outputs(1886) <= (inputs(221)) and (inputs(74));
    layer0_outputs(1887) <= '1';
    layer0_outputs(1888) <= inputs(231);
    layer0_outputs(1889) <= (inputs(172)) or (inputs(147));
    layer0_outputs(1890) <= (inputs(151)) xor (inputs(242));
    layer0_outputs(1891) <= not(inputs(209)) or (inputs(149));
    layer0_outputs(1892) <= not(inputs(190));
    layer0_outputs(1893) <= (inputs(146)) or (inputs(51));
    layer0_outputs(1894) <= (inputs(254)) and (inputs(63));
    layer0_outputs(1895) <= inputs(211);
    layer0_outputs(1896) <= (inputs(218)) or (inputs(162));
    layer0_outputs(1897) <= not(inputs(230));
    layer0_outputs(1898) <= (inputs(147)) or (inputs(127));
    layer0_outputs(1899) <= not(inputs(22)) or (inputs(97));
    layer0_outputs(1900) <= not(inputs(21)) or (inputs(129));
    layer0_outputs(1901) <= (inputs(105)) and not (inputs(253));
    layer0_outputs(1902) <= (inputs(223)) or (inputs(168));
    layer0_outputs(1903) <= (inputs(149)) and (inputs(185));
    layer0_outputs(1904) <= not(inputs(239));
    layer0_outputs(1905) <= inputs(170);
    layer0_outputs(1906) <= not(inputs(220));
    layer0_outputs(1907) <= '1';
    layer0_outputs(1908) <= (inputs(248)) or (inputs(33));
    layer0_outputs(1909) <= not((inputs(16)) or (inputs(4)));
    layer0_outputs(1910) <= not((inputs(143)) and (inputs(28)));
    layer0_outputs(1911) <= (inputs(127)) or (inputs(55));
    layer0_outputs(1912) <= (inputs(163)) and not (inputs(109));
    layer0_outputs(1913) <= (inputs(8)) xor (inputs(126));
    layer0_outputs(1914) <= '0';
    layer0_outputs(1915) <= not(inputs(135));
    layer0_outputs(1916) <= (inputs(58)) and not (inputs(63));
    layer0_outputs(1917) <= inputs(195);
    layer0_outputs(1918) <= not(inputs(70));
    layer0_outputs(1919) <= (inputs(11)) and (inputs(5));
    layer0_outputs(1920) <= (inputs(246)) and not (inputs(25));
    layer0_outputs(1921) <= not(inputs(172));
    layer0_outputs(1922) <= not(inputs(89));
    layer0_outputs(1923) <= inputs(84);
    layer0_outputs(1924) <= not((inputs(252)) or (inputs(234)));
    layer0_outputs(1925) <= (inputs(223)) or (inputs(5));
    layer0_outputs(1926) <= inputs(219);
    layer0_outputs(1927) <= (inputs(217)) or (inputs(219));
    layer0_outputs(1928) <= (inputs(71)) or (inputs(226));
    layer0_outputs(1929) <= (inputs(185)) and (inputs(172));
    layer0_outputs(1930) <= inputs(14);
    layer0_outputs(1931) <= not((inputs(170)) and (inputs(196)));
    layer0_outputs(1932) <= not(inputs(40));
    layer0_outputs(1933) <= (inputs(176)) or (inputs(143));
    layer0_outputs(1934) <= not(inputs(145));
    layer0_outputs(1935) <= (inputs(235)) or (inputs(219));
    layer0_outputs(1936) <= (inputs(60)) or (inputs(19));
    layer0_outputs(1937) <= inputs(238);
    layer0_outputs(1938) <= (inputs(217)) or (inputs(189));
    layer0_outputs(1939) <= '0';
    layer0_outputs(1940) <= not(inputs(160)) or (inputs(55));
    layer0_outputs(1941) <= (inputs(116)) or (inputs(147));
    layer0_outputs(1942) <= not(inputs(146)) or (inputs(223));
    layer0_outputs(1943) <= (inputs(145)) or (inputs(111));
    layer0_outputs(1944) <= not(inputs(208));
    layer0_outputs(1945) <= (inputs(110)) or (inputs(211));
    layer0_outputs(1946) <= not((inputs(68)) or (inputs(239)));
    layer0_outputs(1947) <= not(inputs(22)) or (inputs(28));
    layer0_outputs(1948) <= (inputs(165)) and not (inputs(221));
    layer0_outputs(1949) <= not(inputs(23));
    layer0_outputs(1950) <= inputs(56);
    layer0_outputs(1951) <= inputs(243);
    layer0_outputs(1952) <= '0';
    layer0_outputs(1953) <= not(inputs(105));
    layer0_outputs(1954) <= inputs(177);
    layer0_outputs(1955) <= not((inputs(78)) xor (inputs(44)));
    layer0_outputs(1956) <= inputs(58);
    layer0_outputs(1957) <= not((inputs(193)) or (inputs(120)));
    layer0_outputs(1958) <= not(inputs(177)) or (inputs(146));
    layer0_outputs(1959) <= '0';
    layer0_outputs(1960) <= (inputs(235)) and (inputs(91));
    layer0_outputs(1961) <= (inputs(120)) and not (inputs(254));
    layer0_outputs(1962) <= inputs(147);
    layer0_outputs(1963) <= not(inputs(119));
    layer0_outputs(1964) <= not((inputs(220)) or (inputs(144)));
    layer0_outputs(1965) <= not((inputs(93)) or (inputs(188)));
    layer0_outputs(1966) <= not((inputs(3)) xor (inputs(211)));
    layer0_outputs(1967) <= inputs(109);
    layer0_outputs(1968) <= '1';
    layer0_outputs(1969) <= not((inputs(21)) or (inputs(243)));
    layer0_outputs(1970) <= '1';
    layer0_outputs(1971) <= (inputs(32)) and not (inputs(30));
    layer0_outputs(1972) <= (inputs(162)) and not (inputs(135));
    layer0_outputs(1973) <= not(inputs(106)) or (inputs(179));
    layer0_outputs(1974) <= (inputs(2)) or (inputs(124));
    layer0_outputs(1975) <= '1';
    layer0_outputs(1976) <= inputs(167);
    layer0_outputs(1977) <= not(inputs(184));
    layer0_outputs(1978) <= '0';
    layer0_outputs(1979) <= not(inputs(197)) or (inputs(189));
    layer0_outputs(1980) <= inputs(155);
    layer0_outputs(1981) <= inputs(130);
    layer0_outputs(1982) <= (inputs(176)) and not (inputs(233));
    layer0_outputs(1983) <= not(inputs(60));
    layer0_outputs(1984) <= not(inputs(208)) or (inputs(27));
    layer0_outputs(1985) <= (inputs(55)) and not (inputs(107));
    layer0_outputs(1986) <= '1';
    layer0_outputs(1987) <= not(inputs(117)) or (inputs(41));
    layer0_outputs(1988) <= not(inputs(37));
    layer0_outputs(1989) <= not(inputs(177));
    layer0_outputs(1990) <= '1';
    layer0_outputs(1991) <= inputs(97);
    layer0_outputs(1992) <= (inputs(134)) and not (inputs(200));
    layer0_outputs(1993) <= (inputs(170)) and not (inputs(57));
    layer0_outputs(1994) <= inputs(204);
    layer0_outputs(1995) <= '0';
    layer0_outputs(1996) <= not(inputs(223)) or (inputs(126));
    layer0_outputs(1997) <= not(inputs(173));
    layer0_outputs(1998) <= (inputs(1)) or (inputs(218));
    layer0_outputs(1999) <= not((inputs(206)) or (inputs(251)));
    layer0_outputs(2000) <= inputs(74);
    layer0_outputs(2001) <= inputs(50);
    layer0_outputs(2002) <= inputs(10);
    layer0_outputs(2003) <= (inputs(182)) and not (inputs(132));
    layer0_outputs(2004) <= not(inputs(172));
    layer0_outputs(2005) <= (inputs(232)) and not (inputs(183));
    layer0_outputs(2006) <= (inputs(30)) or (inputs(60));
    layer0_outputs(2007) <= not((inputs(145)) or (inputs(69)));
    layer0_outputs(2008) <= not((inputs(44)) or (inputs(98)));
    layer0_outputs(2009) <= (inputs(220)) and not (inputs(127));
    layer0_outputs(2010) <= not(inputs(141));
    layer0_outputs(2011) <= (inputs(192)) or (inputs(212));
    layer0_outputs(2012) <= inputs(183);
    layer0_outputs(2013) <= not(inputs(106)) or (inputs(172));
    layer0_outputs(2014) <= not((inputs(207)) or (inputs(237)));
    layer0_outputs(2015) <= (inputs(58)) and (inputs(225));
    layer0_outputs(2016) <= not(inputs(220));
    layer0_outputs(2017) <= not(inputs(178)) or (inputs(236));
    layer0_outputs(2018) <= (inputs(50)) and (inputs(88));
    layer0_outputs(2019) <= inputs(77);
    layer0_outputs(2020) <= '0';
    layer0_outputs(2021) <= '0';
    layer0_outputs(2022) <= inputs(246);
    layer0_outputs(2023) <= not((inputs(3)) or (inputs(46)));
    layer0_outputs(2024) <= not(inputs(158)) or (inputs(77));
    layer0_outputs(2025) <= inputs(104);
    layer0_outputs(2026) <= inputs(134);
    layer0_outputs(2027) <= (inputs(70)) or (inputs(133));
    layer0_outputs(2028) <= not(inputs(115));
    layer0_outputs(2029) <= not(inputs(25));
    layer0_outputs(2030) <= not(inputs(117));
    layer0_outputs(2031) <= inputs(93);
    layer0_outputs(2032) <= (inputs(44)) or (inputs(205));
    layer0_outputs(2033) <= (inputs(108)) or (inputs(21));
    layer0_outputs(2034) <= (inputs(91)) or (inputs(111));
    layer0_outputs(2035) <= '1';
    layer0_outputs(2036) <= (inputs(65)) xor (inputs(216));
    layer0_outputs(2037) <= '0';
    layer0_outputs(2038) <= not(inputs(173)) or (inputs(253));
    layer0_outputs(2039) <= inputs(218);
    layer0_outputs(2040) <= not(inputs(217));
    layer0_outputs(2041) <= (inputs(205)) and not (inputs(51));
    layer0_outputs(2042) <= (inputs(75)) or (inputs(123));
    layer0_outputs(2043) <= not(inputs(20)) or (inputs(83));
    layer0_outputs(2044) <= (inputs(192)) or (inputs(232));
    layer0_outputs(2045) <= '1';
    layer0_outputs(2046) <= (inputs(251)) and (inputs(160));
    layer0_outputs(2047) <= not(inputs(87)) or (inputs(251));
    layer0_outputs(2048) <= (inputs(138)) or (inputs(107));
    layer0_outputs(2049) <= not(inputs(136)) or (inputs(138));
    layer0_outputs(2050) <= '0';
    layer0_outputs(2051) <= not(inputs(122)) or (inputs(11));
    layer0_outputs(2052) <= not(inputs(176));
    layer0_outputs(2053) <= (inputs(107)) or (inputs(47));
    layer0_outputs(2054) <= not(inputs(187)) or (inputs(251));
    layer0_outputs(2055) <= not(inputs(209));
    layer0_outputs(2056) <= inputs(41);
    layer0_outputs(2057) <= inputs(147);
    layer0_outputs(2058) <= inputs(92);
    layer0_outputs(2059) <= not(inputs(167)) or (inputs(186));
    layer0_outputs(2060) <= '1';
    layer0_outputs(2061) <= (inputs(54)) xor (inputs(2));
    layer0_outputs(2062) <= not((inputs(192)) or (inputs(229)));
    layer0_outputs(2063) <= (inputs(169)) or (inputs(16));
    layer0_outputs(2064) <= not(inputs(212)) or (inputs(135));
    layer0_outputs(2065) <= '0';
    layer0_outputs(2066) <= (inputs(158)) xor (inputs(222));
    layer0_outputs(2067) <= not(inputs(187));
    layer0_outputs(2068) <= '1';
    layer0_outputs(2069) <= not(inputs(100));
    layer0_outputs(2070) <= not(inputs(121));
    layer0_outputs(2071) <= (inputs(1)) or (inputs(190));
    layer0_outputs(2072) <= '1';
    layer0_outputs(2073) <= (inputs(150)) and not (inputs(254));
    layer0_outputs(2074) <= '0';
    layer0_outputs(2075) <= '0';
    layer0_outputs(2076) <= (inputs(31)) xor (inputs(2));
    layer0_outputs(2077) <= inputs(149);
    layer0_outputs(2078) <= (inputs(87)) xor (inputs(143));
    layer0_outputs(2079) <= not((inputs(127)) or (inputs(140)));
    layer0_outputs(2080) <= not((inputs(225)) or (inputs(45)));
    layer0_outputs(2081) <= (inputs(98)) and (inputs(57));
    layer0_outputs(2082) <= (inputs(251)) and not (inputs(114));
    layer0_outputs(2083) <= (inputs(62)) and not (inputs(238));
    layer0_outputs(2084) <= not((inputs(186)) or (inputs(142)));
    layer0_outputs(2085) <= inputs(248);
    layer0_outputs(2086) <= '1';
    layer0_outputs(2087) <= inputs(229);
    layer0_outputs(2088) <= '0';
    layer0_outputs(2089) <= not(inputs(129));
    layer0_outputs(2090) <= not(inputs(105));
    layer0_outputs(2091) <= '0';
    layer0_outputs(2092) <= '1';
    layer0_outputs(2093) <= inputs(21);
    layer0_outputs(2094) <= not((inputs(204)) or (inputs(223)));
    layer0_outputs(2095) <= (inputs(215)) and (inputs(8));
    layer0_outputs(2096) <= (inputs(110)) and not (inputs(14));
    layer0_outputs(2097) <= inputs(73);
    layer0_outputs(2098) <= (inputs(155)) or (inputs(68));
    layer0_outputs(2099) <= '1';
    layer0_outputs(2100) <= not((inputs(17)) and (inputs(23)));
    layer0_outputs(2101) <= not(inputs(20));
    layer0_outputs(2102) <= (inputs(40)) and not (inputs(164));
    layer0_outputs(2103) <= not(inputs(86));
    layer0_outputs(2104) <= not(inputs(32)) or (inputs(11));
    layer0_outputs(2105) <= inputs(174);
    layer0_outputs(2106) <= (inputs(60)) and not (inputs(240));
    layer0_outputs(2107) <= (inputs(218)) or (inputs(86));
    layer0_outputs(2108) <= (inputs(47)) or (inputs(46));
    layer0_outputs(2109) <= '1';
    layer0_outputs(2110) <= '0';
    layer0_outputs(2111) <= not(inputs(32)) or (inputs(153));
    layer0_outputs(2112) <= inputs(68);
    layer0_outputs(2113) <= inputs(91);
    layer0_outputs(2114) <= (inputs(136)) or (inputs(143));
    layer0_outputs(2115) <= inputs(97);
    layer0_outputs(2116) <= not(inputs(245));
    layer0_outputs(2117) <= inputs(139);
    layer0_outputs(2118) <= inputs(32);
    layer0_outputs(2119) <= inputs(157);
    layer0_outputs(2120) <= not((inputs(114)) xor (inputs(28)));
    layer0_outputs(2121) <= (inputs(170)) or (inputs(130));
    layer0_outputs(2122) <= not((inputs(247)) or (inputs(246)));
    layer0_outputs(2123) <= not(inputs(8)) or (inputs(13));
    layer0_outputs(2124) <= not(inputs(23));
    layer0_outputs(2125) <= not(inputs(181)) or (inputs(83));
    layer0_outputs(2126) <= (inputs(112)) or (inputs(99));
    layer0_outputs(2127) <= (inputs(113)) or (inputs(102));
    layer0_outputs(2128) <= not(inputs(202)) or (inputs(211));
    layer0_outputs(2129) <= '1';
    layer0_outputs(2130) <= not(inputs(176));
    layer0_outputs(2131) <= '1';
    layer0_outputs(2132) <= inputs(243);
    layer0_outputs(2133) <= not((inputs(56)) and (inputs(36)));
    layer0_outputs(2134) <= (inputs(149)) and not (inputs(104));
    layer0_outputs(2135) <= (inputs(69)) and not (inputs(2));
    layer0_outputs(2136) <= not(inputs(219));
    layer0_outputs(2137) <= '0';
    layer0_outputs(2138) <= '1';
    layer0_outputs(2139) <= not(inputs(93));
    layer0_outputs(2140) <= '0';
    layer0_outputs(2141) <= (inputs(128)) and not (inputs(205));
    layer0_outputs(2142) <= not(inputs(230)) or (inputs(63));
    layer0_outputs(2143) <= (inputs(170)) and not (inputs(9));
    layer0_outputs(2144) <= not(inputs(46));
    layer0_outputs(2145) <= not((inputs(80)) or (inputs(207)));
    layer0_outputs(2146) <= inputs(180);
    layer0_outputs(2147) <= not((inputs(71)) and (inputs(127)));
    layer0_outputs(2148) <= not((inputs(10)) xor (inputs(9)));
    layer0_outputs(2149) <= not(inputs(105));
    layer0_outputs(2150) <= inputs(211);
    layer0_outputs(2151) <= (inputs(31)) xor (inputs(232));
    layer0_outputs(2152) <= not(inputs(74));
    layer0_outputs(2153) <= not(inputs(213));
    layer0_outputs(2154) <= (inputs(44)) xor (inputs(75));
    layer0_outputs(2155) <= (inputs(95)) and (inputs(67));
    layer0_outputs(2156) <= (inputs(119)) xor (inputs(150));
    layer0_outputs(2157) <= not(inputs(230));
    layer0_outputs(2158) <= not(inputs(181)) or (inputs(110));
    layer0_outputs(2159) <= inputs(68);
    layer0_outputs(2160) <= not((inputs(115)) and (inputs(0)));
    layer0_outputs(2161) <= inputs(66);
    layer0_outputs(2162) <= not((inputs(246)) and (inputs(186)));
    layer0_outputs(2163) <= not(inputs(80));
    layer0_outputs(2164) <= not(inputs(210));
    layer0_outputs(2165) <= inputs(238);
    layer0_outputs(2166) <= inputs(135);
    layer0_outputs(2167) <= not(inputs(119));
    layer0_outputs(2168) <= (inputs(244)) or (inputs(41));
    layer0_outputs(2169) <= not(inputs(86));
    layer0_outputs(2170) <= (inputs(148)) or (inputs(158));
    layer0_outputs(2171) <= inputs(188);
    layer0_outputs(2172) <= inputs(83);
    layer0_outputs(2173) <= (inputs(149)) or (inputs(188));
    layer0_outputs(2174) <= not((inputs(149)) xor (inputs(149)));
    layer0_outputs(2175) <= not((inputs(208)) or (inputs(9)));
    layer0_outputs(2176) <= not(inputs(118)) or (inputs(223));
    layer0_outputs(2177) <= not(inputs(152));
    layer0_outputs(2178) <= (inputs(202)) and not (inputs(31));
    layer0_outputs(2179) <= inputs(77);
    layer0_outputs(2180) <= inputs(157);
    layer0_outputs(2181) <= (inputs(216)) and (inputs(217));
    layer0_outputs(2182) <= not(inputs(118)) or (inputs(191));
    layer0_outputs(2183) <= (inputs(208)) and (inputs(124));
    layer0_outputs(2184) <= not(inputs(92));
    layer0_outputs(2185) <= '0';
    layer0_outputs(2186) <= not(inputs(167));
    layer0_outputs(2187) <= inputs(158);
    layer0_outputs(2188) <= not((inputs(123)) xor (inputs(67)));
    layer0_outputs(2189) <= (inputs(242)) or (inputs(18));
    layer0_outputs(2190) <= inputs(159);
    layer0_outputs(2191) <= (inputs(176)) xor (inputs(10));
    layer0_outputs(2192) <= not((inputs(124)) or (inputs(202)));
    layer0_outputs(2193) <= inputs(228);
    layer0_outputs(2194) <= (inputs(145)) and not (inputs(77));
    layer0_outputs(2195) <= (inputs(85)) or (inputs(97));
    layer0_outputs(2196) <= inputs(76);
    layer0_outputs(2197) <= (inputs(5)) and (inputs(24));
    layer0_outputs(2198) <= not(inputs(77)) or (inputs(14));
    layer0_outputs(2199) <= not((inputs(1)) or (inputs(38)));
    layer0_outputs(2200) <= inputs(176);
    layer0_outputs(2201) <= not(inputs(239));
    layer0_outputs(2202) <= not((inputs(180)) xor (inputs(60)));
    layer0_outputs(2203) <= not((inputs(62)) or (inputs(45)));
    layer0_outputs(2204) <= not(inputs(241));
    layer0_outputs(2205) <= not((inputs(72)) and (inputs(200)));
    layer0_outputs(2206) <= not(inputs(8));
    layer0_outputs(2207) <= '0';
    layer0_outputs(2208) <= not(inputs(13));
    layer0_outputs(2209) <= inputs(247);
    layer0_outputs(2210) <= (inputs(222)) or (inputs(18));
    layer0_outputs(2211) <= inputs(153);
    layer0_outputs(2212) <= not((inputs(71)) and (inputs(36)));
    layer0_outputs(2213) <= not(inputs(44));
    layer0_outputs(2214) <= (inputs(146)) xor (inputs(226));
    layer0_outputs(2215) <= (inputs(120)) and not (inputs(140));
    layer0_outputs(2216) <= '0';
    layer0_outputs(2217) <= not(inputs(77)) or (inputs(105));
    layer0_outputs(2218) <= not(inputs(239)) or (inputs(12));
    layer0_outputs(2219) <= not((inputs(4)) or (inputs(16)));
    layer0_outputs(2220) <= not(inputs(221));
    layer0_outputs(2221) <= not(inputs(116));
    layer0_outputs(2222) <= not((inputs(81)) or (inputs(66)));
    layer0_outputs(2223) <= '1';
    layer0_outputs(2224) <= not(inputs(91));
    layer0_outputs(2225) <= (inputs(238)) and (inputs(240));
    layer0_outputs(2226) <= not(inputs(151));
    layer0_outputs(2227) <= not(inputs(214)) or (inputs(118));
    layer0_outputs(2228) <= (inputs(28)) or (inputs(19));
    layer0_outputs(2229) <= (inputs(210)) and not (inputs(120));
    layer0_outputs(2230) <= inputs(75);
    layer0_outputs(2231) <= '0';
    layer0_outputs(2232) <= (inputs(2)) or (inputs(25));
    layer0_outputs(2233) <= inputs(183);
    layer0_outputs(2234) <= (inputs(51)) and (inputs(239));
    layer0_outputs(2235) <= not(inputs(39)) or (inputs(155));
    layer0_outputs(2236) <= inputs(40);
    layer0_outputs(2237) <= not((inputs(19)) or (inputs(163)));
    layer0_outputs(2238) <= (inputs(231)) and not (inputs(52));
    layer0_outputs(2239) <= not((inputs(98)) xor (inputs(14)));
    layer0_outputs(2240) <= not(inputs(215)) or (inputs(136));
    layer0_outputs(2241) <= '1';
    layer0_outputs(2242) <= inputs(231);
    layer0_outputs(2243) <= '0';
    layer0_outputs(2244) <= not((inputs(48)) xor (inputs(172)));
    layer0_outputs(2245) <= not(inputs(155));
    layer0_outputs(2246) <= '1';
    layer0_outputs(2247) <= inputs(228);
    layer0_outputs(2248) <= inputs(166);
    layer0_outputs(2249) <= not(inputs(179)) or (inputs(31));
    layer0_outputs(2250) <= not(inputs(25));
    layer0_outputs(2251) <= inputs(94);
    layer0_outputs(2252) <= not((inputs(166)) or (inputs(134)));
    layer0_outputs(2253) <= (inputs(162)) and not (inputs(109));
    layer0_outputs(2254) <= not(inputs(183));
    layer0_outputs(2255) <= '1';
    layer0_outputs(2256) <= not(inputs(23)) or (inputs(207));
    layer0_outputs(2257) <= (inputs(108)) or (inputs(94));
    layer0_outputs(2258) <= inputs(59);
    layer0_outputs(2259) <= '1';
    layer0_outputs(2260) <= not((inputs(97)) or (inputs(188)));
    layer0_outputs(2261) <= '1';
    layer0_outputs(2262) <= inputs(239);
    layer0_outputs(2263) <= inputs(8);
    layer0_outputs(2264) <= (inputs(153)) and not (inputs(46));
    layer0_outputs(2265) <= not(inputs(227));
    layer0_outputs(2266) <= inputs(141);
    layer0_outputs(2267) <= not(inputs(153));
    layer0_outputs(2268) <= '0';
    layer0_outputs(2269) <= inputs(97);
    layer0_outputs(2270) <= (inputs(86)) and (inputs(10));
    layer0_outputs(2271) <= not((inputs(192)) or (inputs(237)));
    layer0_outputs(2272) <= not(inputs(164));
    layer0_outputs(2273) <= not((inputs(251)) or (inputs(64)));
    layer0_outputs(2274) <= not(inputs(108));
    layer0_outputs(2275) <= '0';
    layer0_outputs(2276) <= inputs(84);
    layer0_outputs(2277) <= (inputs(39)) or (inputs(0));
    layer0_outputs(2278) <= not(inputs(177));
    layer0_outputs(2279) <= not(inputs(211));
    layer0_outputs(2280) <= '0';
    layer0_outputs(2281) <= (inputs(195)) and not (inputs(31));
    layer0_outputs(2282) <= not(inputs(247));
    layer0_outputs(2283) <= not(inputs(16));
    layer0_outputs(2284) <= not(inputs(37));
    layer0_outputs(2285) <= (inputs(155)) and not (inputs(57));
    layer0_outputs(2286) <= inputs(168);
    layer0_outputs(2287) <= (inputs(106)) and not (inputs(113));
    layer0_outputs(2288) <= (inputs(225)) and not (inputs(59));
    layer0_outputs(2289) <= not(inputs(147));
    layer0_outputs(2290) <= '0';
    layer0_outputs(2291) <= not(inputs(157));
    layer0_outputs(2292) <= not((inputs(31)) xor (inputs(199)));
    layer0_outputs(2293) <= (inputs(49)) or (inputs(151));
    layer0_outputs(2294) <= (inputs(132)) and not (inputs(94));
    layer0_outputs(2295) <= not(inputs(84));
    layer0_outputs(2296) <= not(inputs(217)) or (inputs(85));
    layer0_outputs(2297) <= (inputs(71)) and not (inputs(222));
    layer0_outputs(2298) <= inputs(88);
    layer0_outputs(2299) <= not(inputs(244));
    layer0_outputs(2300) <= (inputs(64)) and not (inputs(77));
    layer0_outputs(2301) <= inputs(86);
    layer0_outputs(2302) <= '1';
    layer0_outputs(2303) <= '0';
    layer0_outputs(2304) <= not(inputs(76));
    layer0_outputs(2305) <= (inputs(85)) and not (inputs(6));
    layer0_outputs(2306) <= not(inputs(109)) or (inputs(135));
    layer0_outputs(2307) <= not((inputs(228)) or (inputs(161)));
    layer0_outputs(2308) <= (inputs(156)) or (inputs(227));
    layer0_outputs(2309) <= inputs(252);
    layer0_outputs(2310) <= inputs(224);
    layer0_outputs(2311) <= not(inputs(137)) or (inputs(230));
    layer0_outputs(2312) <= inputs(25);
    layer0_outputs(2313) <= not(inputs(94));
    layer0_outputs(2314) <= inputs(142);
    layer0_outputs(2315) <= (inputs(232)) and (inputs(165));
    layer0_outputs(2316) <= (inputs(153)) and (inputs(141));
    layer0_outputs(2317) <= inputs(136);
    layer0_outputs(2318) <= not((inputs(86)) or (inputs(210)));
    layer0_outputs(2319) <= not(inputs(89));
    layer0_outputs(2320) <= (inputs(100)) or (inputs(239));
    layer0_outputs(2321) <= inputs(107);
    layer0_outputs(2322) <= inputs(234);
    layer0_outputs(2323) <= (inputs(34)) and not (inputs(221));
    layer0_outputs(2324) <= inputs(147);
    layer0_outputs(2325) <= inputs(177);
    layer0_outputs(2326) <= inputs(98);
    layer0_outputs(2327) <= '0';
    layer0_outputs(2328) <= not(inputs(146));
    layer0_outputs(2329) <= (inputs(203)) and not (inputs(208));
    layer0_outputs(2330) <= not(inputs(90));
    layer0_outputs(2331) <= not(inputs(119));
    layer0_outputs(2332) <= not((inputs(0)) or (inputs(90)));
    layer0_outputs(2333) <= not(inputs(13));
    layer0_outputs(2334) <= (inputs(81)) and not (inputs(186));
    layer0_outputs(2335) <= (inputs(173)) and not (inputs(15));
    layer0_outputs(2336) <= not((inputs(184)) or (inputs(178)));
    layer0_outputs(2337) <= '0';
    layer0_outputs(2338) <= inputs(87);
    layer0_outputs(2339) <= (inputs(234)) and not (inputs(153));
    layer0_outputs(2340) <= not(inputs(242));
    layer0_outputs(2341) <= not(inputs(192));
    layer0_outputs(2342) <= inputs(247);
    layer0_outputs(2343) <= not((inputs(25)) xor (inputs(55)));
    layer0_outputs(2344) <= not(inputs(231));
    layer0_outputs(2345) <= not(inputs(36));
    layer0_outputs(2346) <= not(inputs(120));
    layer0_outputs(2347) <= not(inputs(220)) or (inputs(12));
    layer0_outputs(2348) <= '1';
    layer0_outputs(2349) <= inputs(212);
    layer0_outputs(2350) <= (inputs(25)) and not (inputs(237));
    layer0_outputs(2351) <= inputs(240);
    layer0_outputs(2352) <= not((inputs(253)) or (inputs(115)));
    layer0_outputs(2353) <= not(inputs(56)) or (inputs(82));
    layer0_outputs(2354) <= '0';
    layer0_outputs(2355) <= (inputs(249)) and (inputs(224));
    layer0_outputs(2356) <= inputs(8);
    layer0_outputs(2357) <= not(inputs(216)) or (inputs(181));
    layer0_outputs(2358) <= (inputs(11)) and not (inputs(4));
    layer0_outputs(2359) <= not(inputs(19));
    layer0_outputs(2360) <= '1';
    layer0_outputs(2361) <= not((inputs(2)) or (inputs(149)));
    layer0_outputs(2362) <= (inputs(131)) and (inputs(122));
    layer0_outputs(2363) <= not(inputs(72)) or (inputs(49));
    layer0_outputs(2364) <= not((inputs(94)) or (inputs(174)));
    layer0_outputs(2365) <= (inputs(1)) xor (inputs(120));
    layer0_outputs(2366) <= '1';
    layer0_outputs(2367) <= not(inputs(84)) or (inputs(0));
    layer0_outputs(2368) <= inputs(68);
    layer0_outputs(2369) <= '1';
    layer0_outputs(2370) <= '0';
    layer0_outputs(2371) <= not(inputs(104)) or (inputs(248));
    layer0_outputs(2372) <= inputs(168);
    layer0_outputs(2373) <= '1';
    layer0_outputs(2374) <= (inputs(124)) or (inputs(4));
    layer0_outputs(2375) <= inputs(59);
    layer0_outputs(2376) <= inputs(131);
    layer0_outputs(2377) <= (inputs(72)) and (inputs(132));
    layer0_outputs(2378) <= not(inputs(178)) or (inputs(97));
    layer0_outputs(2379) <= (inputs(106)) and not (inputs(164));
    layer0_outputs(2380) <= inputs(101);
    layer0_outputs(2381) <= not(inputs(130));
    layer0_outputs(2382) <= (inputs(101)) or (inputs(140));
    layer0_outputs(2383) <= not(inputs(165));
    layer0_outputs(2384) <= (inputs(166)) and not (inputs(230));
    layer0_outputs(2385) <= inputs(117);
    layer0_outputs(2386) <= not(inputs(68)) or (inputs(34));
    layer0_outputs(2387) <= (inputs(53)) and not (inputs(174));
    layer0_outputs(2388) <= '0';
    layer0_outputs(2389) <= not((inputs(252)) and (inputs(228)));
    layer0_outputs(2390) <= inputs(232);
    layer0_outputs(2391) <= (inputs(134)) and not (inputs(141));
    layer0_outputs(2392) <= not(inputs(12));
    layer0_outputs(2393) <= (inputs(181)) or (inputs(184));
    layer0_outputs(2394) <= (inputs(156)) and not (inputs(32));
    layer0_outputs(2395) <= not((inputs(0)) and (inputs(230)));
    layer0_outputs(2396) <= (inputs(203)) or (inputs(219));
    layer0_outputs(2397) <= (inputs(70)) and (inputs(174));
    layer0_outputs(2398) <= (inputs(91)) or (inputs(191));
    layer0_outputs(2399) <= not((inputs(48)) and (inputs(98)));
    layer0_outputs(2400) <= not(inputs(8)) or (inputs(159));
    layer0_outputs(2401) <= (inputs(20)) xor (inputs(38));
    layer0_outputs(2402) <= not(inputs(107));
    layer0_outputs(2403) <= not(inputs(163)) or (inputs(15));
    layer0_outputs(2404) <= not((inputs(61)) or (inputs(112)));
    layer0_outputs(2405) <= (inputs(217)) and not (inputs(62));
    layer0_outputs(2406) <= not(inputs(79)) or (inputs(4));
    layer0_outputs(2407) <= (inputs(161)) and not (inputs(58));
    layer0_outputs(2408) <= (inputs(148)) and not (inputs(220));
    layer0_outputs(2409) <= (inputs(200)) or (inputs(238));
    layer0_outputs(2410) <= not(inputs(195)) or (inputs(30));
    layer0_outputs(2411) <= not(inputs(101));
    layer0_outputs(2412) <= not((inputs(250)) or (inputs(66)));
    layer0_outputs(2413) <= '0';
    layer0_outputs(2414) <= inputs(164);
    layer0_outputs(2415) <= not(inputs(88)) or (inputs(192));
    layer0_outputs(2416) <= inputs(210);
    layer0_outputs(2417) <= (inputs(144)) and not (inputs(221));
    layer0_outputs(2418) <= not(inputs(41));
    layer0_outputs(2419) <= (inputs(118)) and (inputs(173));
    layer0_outputs(2420) <= inputs(194);
    layer0_outputs(2421) <= '1';
    layer0_outputs(2422) <= '1';
    layer0_outputs(2423) <= '0';
    layer0_outputs(2424) <= not(inputs(198)) or (inputs(93));
    layer0_outputs(2425) <= (inputs(155)) and (inputs(19));
    layer0_outputs(2426) <= not((inputs(44)) xor (inputs(164)));
    layer0_outputs(2427) <= not(inputs(106));
    layer0_outputs(2428) <= inputs(215);
    layer0_outputs(2429) <= not(inputs(74)) or (inputs(142));
    layer0_outputs(2430) <= (inputs(248)) and (inputs(54));
    layer0_outputs(2431) <= not(inputs(209)) or (inputs(134));
    layer0_outputs(2432) <= not(inputs(227)) or (inputs(165));
    layer0_outputs(2433) <= (inputs(232)) and not (inputs(168));
    layer0_outputs(2434) <= not(inputs(109));
    layer0_outputs(2435) <= not(inputs(212));
    layer0_outputs(2436) <= '0';
    layer0_outputs(2437) <= (inputs(45)) xor (inputs(47));
    layer0_outputs(2438) <= not((inputs(124)) or (inputs(154)));
    layer0_outputs(2439) <= not((inputs(36)) or (inputs(140)));
    layer0_outputs(2440) <= not((inputs(140)) or (inputs(253)));
    layer0_outputs(2441) <= (inputs(156)) or (inputs(18));
    layer0_outputs(2442) <= not(inputs(154));
    layer0_outputs(2443) <= (inputs(178)) and not (inputs(142));
    layer0_outputs(2444) <= not(inputs(202));
    layer0_outputs(2445) <= (inputs(223)) and not (inputs(96));
    layer0_outputs(2446) <= not((inputs(101)) or (inputs(118)));
    layer0_outputs(2447) <= not((inputs(208)) or (inputs(132)));
    layer0_outputs(2448) <= inputs(32);
    layer0_outputs(2449) <= not(inputs(153)) or (inputs(149));
    layer0_outputs(2450) <= (inputs(143)) and not (inputs(43));
    layer0_outputs(2451) <= not(inputs(167));
    layer0_outputs(2452) <= not(inputs(122)) or (inputs(225));
    layer0_outputs(2453) <= (inputs(126)) or (inputs(146));
    layer0_outputs(2454) <= not(inputs(217));
    layer0_outputs(2455) <= (inputs(110)) xor (inputs(106));
    layer0_outputs(2456) <= '0';
    layer0_outputs(2457) <= inputs(69);
    layer0_outputs(2458) <= inputs(31);
    layer0_outputs(2459) <= (inputs(0)) and (inputs(225));
    layer0_outputs(2460) <= not((inputs(75)) or (inputs(244)));
    layer0_outputs(2461) <= inputs(84);
    layer0_outputs(2462) <= not(inputs(80)) or (inputs(94));
    layer0_outputs(2463) <= not((inputs(239)) xor (inputs(150)));
    layer0_outputs(2464) <= not(inputs(1));
    layer0_outputs(2465) <= '1';
    layer0_outputs(2466) <= not(inputs(120));
    layer0_outputs(2467) <= (inputs(67)) and not (inputs(189));
    layer0_outputs(2468) <= not(inputs(60)) or (inputs(246));
    layer0_outputs(2469) <= not(inputs(71)) or (inputs(103));
    layer0_outputs(2470) <= (inputs(52)) or (inputs(55));
    layer0_outputs(2471) <= (inputs(6)) and (inputs(28));
    layer0_outputs(2472) <= not(inputs(180)) or (inputs(224));
    layer0_outputs(2473) <= not((inputs(236)) or (inputs(19)));
    layer0_outputs(2474) <= not(inputs(97)) or (inputs(205));
    layer0_outputs(2475) <= not(inputs(203));
    layer0_outputs(2476) <= '0';
    layer0_outputs(2477) <= inputs(99);
    layer0_outputs(2478) <= (inputs(120)) and not (inputs(100));
    layer0_outputs(2479) <= (inputs(80)) and not (inputs(65));
    layer0_outputs(2480) <= inputs(233);
    layer0_outputs(2481) <= '0';
    layer0_outputs(2482) <= (inputs(22)) and (inputs(10));
    layer0_outputs(2483) <= inputs(250);
    layer0_outputs(2484) <= not(inputs(57));
    layer0_outputs(2485) <= (inputs(92)) or (inputs(22));
    layer0_outputs(2486) <= '1';
    layer0_outputs(2487) <= (inputs(109)) and (inputs(30));
    layer0_outputs(2488) <= '1';
    layer0_outputs(2489) <= not((inputs(61)) or (inputs(32)));
    layer0_outputs(2490) <= not((inputs(59)) and (inputs(174)));
    layer0_outputs(2491) <= inputs(125);
    layer0_outputs(2492) <= (inputs(13)) and not (inputs(134));
    layer0_outputs(2493) <= not(inputs(243));
    layer0_outputs(2494) <= not(inputs(126));
    layer0_outputs(2495) <= (inputs(34)) and (inputs(248));
    layer0_outputs(2496) <= not(inputs(181));
    layer0_outputs(2497) <= inputs(233);
    layer0_outputs(2498) <= not(inputs(99));
    layer0_outputs(2499) <= '0';
    layer0_outputs(2500) <= inputs(120);
    layer0_outputs(2501) <= (inputs(78)) xor (inputs(78));
    layer0_outputs(2502) <= '0';
    layer0_outputs(2503) <= (inputs(177)) or (inputs(52));
    layer0_outputs(2504) <= '0';
    layer0_outputs(2505) <= (inputs(48)) or (inputs(163));
    layer0_outputs(2506) <= inputs(233);
    layer0_outputs(2507) <= '1';
    layer0_outputs(2508) <= inputs(22);
    layer0_outputs(2509) <= not(inputs(119));
    layer0_outputs(2510) <= (inputs(253)) and not (inputs(134));
    layer0_outputs(2511) <= '0';
    layer0_outputs(2512) <= '0';
    layer0_outputs(2513) <= '0';
    layer0_outputs(2514) <= '1';
    layer0_outputs(2515) <= inputs(31);
    layer0_outputs(2516) <= '1';
    layer0_outputs(2517) <= not(inputs(230));
    layer0_outputs(2518) <= (inputs(40)) and (inputs(225));
    layer0_outputs(2519) <= not(inputs(105));
    layer0_outputs(2520) <= inputs(67);
    layer0_outputs(2521) <= (inputs(213)) and (inputs(63));
    layer0_outputs(2522) <= not((inputs(178)) or (inputs(148)));
    layer0_outputs(2523) <= (inputs(236)) and not (inputs(155));
    layer0_outputs(2524) <= not(inputs(137));
    layer0_outputs(2525) <= '1';
    layer0_outputs(2526) <= not(inputs(224)) or (inputs(25));
    layer0_outputs(2527) <= not((inputs(139)) or (inputs(182)));
    layer0_outputs(2528) <= not(inputs(168)) or (inputs(247));
    layer0_outputs(2529) <= inputs(105);
    layer0_outputs(2530) <= not(inputs(221));
    layer0_outputs(2531) <= (inputs(1)) or (inputs(234));
    layer0_outputs(2532) <= (inputs(60)) or (inputs(64));
    layer0_outputs(2533) <= not(inputs(226));
    layer0_outputs(2534) <= '0';
    layer0_outputs(2535) <= (inputs(112)) and not (inputs(139));
    layer0_outputs(2536) <= inputs(122);
    layer0_outputs(2537) <= not((inputs(127)) or (inputs(45)));
    layer0_outputs(2538) <= not(inputs(118));
    layer0_outputs(2539) <= '1';
    layer0_outputs(2540) <= '0';
    layer0_outputs(2541) <= not((inputs(177)) or (inputs(255)));
    layer0_outputs(2542) <= (inputs(95)) or (inputs(238));
    layer0_outputs(2543) <= '1';
    layer0_outputs(2544) <= (inputs(24)) and (inputs(93));
    layer0_outputs(2545) <= not(inputs(177));
    layer0_outputs(2546) <= (inputs(223)) xor (inputs(12));
    layer0_outputs(2547) <= not((inputs(95)) or (inputs(48)));
    layer0_outputs(2548) <= inputs(102);
    layer0_outputs(2549) <= not((inputs(180)) and (inputs(180)));
    layer0_outputs(2550) <= not(inputs(148)) or (inputs(90));
    layer0_outputs(2551) <= inputs(86);
    layer0_outputs(2552) <= inputs(85);
    layer0_outputs(2553) <= not(inputs(128));
    layer0_outputs(2554) <= not(inputs(255)) or (inputs(189));
    layer0_outputs(2555) <= (inputs(77)) and not (inputs(150));
    layer0_outputs(2556) <= '1';
    layer0_outputs(2557) <= '1';
    layer0_outputs(2558) <= (inputs(125)) and (inputs(93));
    layer0_outputs(2559) <= '1';
    layer1_outputs(0) <= layer0_outputs(2213);
    layer1_outputs(1) <= (layer0_outputs(171)) and not (layer0_outputs(1503));
    layer1_outputs(2) <= not((layer0_outputs(2413)) xor (layer0_outputs(1089)));
    layer1_outputs(3) <= not(layer0_outputs(375));
    layer1_outputs(4) <= (layer0_outputs(2255)) or (layer0_outputs(2206));
    layer1_outputs(5) <= (layer0_outputs(1061)) and not (layer0_outputs(1370));
    layer1_outputs(6) <= not(layer0_outputs(1026));
    layer1_outputs(7) <= not(layer0_outputs(1830)) or (layer0_outputs(292));
    layer1_outputs(8) <= layer0_outputs(564);
    layer1_outputs(9) <= not(layer0_outputs(1746)) or (layer0_outputs(2484));
    layer1_outputs(10) <= layer0_outputs(676);
    layer1_outputs(11) <= (layer0_outputs(226)) and not (layer0_outputs(439));
    layer1_outputs(12) <= layer0_outputs(1139);
    layer1_outputs(13) <= not(layer0_outputs(2063));
    layer1_outputs(14) <= not(layer0_outputs(940)) or (layer0_outputs(1656));
    layer1_outputs(15) <= (layer0_outputs(284)) and not (layer0_outputs(331));
    layer1_outputs(16) <= not(layer0_outputs(1321));
    layer1_outputs(17) <= not(layer0_outputs(2416));
    layer1_outputs(18) <= '0';
    layer1_outputs(19) <= (layer0_outputs(2273)) or (layer0_outputs(1378));
    layer1_outputs(20) <= layer0_outputs(2375);
    layer1_outputs(21) <= layer0_outputs(973);
    layer1_outputs(22) <= (layer0_outputs(1397)) and not (layer0_outputs(325));
    layer1_outputs(23) <= '0';
    layer1_outputs(24) <= not(layer0_outputs(2323));
    layer1_outputs(25) <= not(layer0_outputs(1584));
    layer1_outputs(26) <= '0';
    layer1_outputs(27) <= not(layer0_outputs(2367)) or (layer0_outputs(299));
    layer1_outputs(28) <= (layer0_outputs(1011)) and not (layer0_outputs(951));
    layer1_outputs(29) <= '1';
    layer1_outputs(30) <= layer0_outputs(27);
    layer1_outputs(31) <= layer0_outputs(724);
    layer1_outputs(32) <= (layer0_outputs(582)) and (layer0_outputs(223));
    layer1_outputs(33) <= (layer0_outputs(1141)) and not (layer0_outputs(116));
    layer1_outputs(34) <= not((layer0_outputs(976)) or (layer0_outputs(364)));
    layer1_outputs(35) <= not((layer0_outputs(371)) or (layer0_outputs(575)));
    layer1_outputs(36) <= not((layer0_outputs(2281)) or (layer0_outputs(2335)));
    layer1_outputs(37) <= layer0_outputs(1547);
    layer1_outputs(38) <= not((layer0_outputs(2212)) and (layer0_outputs(1528)));
    layer1_outputs(39) <= not(layer0_outputs(2044));
    layer1_outputs(40) <= not(layer0_outputs(2445)) or (layer0_outputs(2493));
    layer1_outputs(41) <= (layer0_outputs(289)) and (layer0_outputs(1069));
    layer1_outputs(42) <= layer0_outputs(804);
    layer1_outputs(43) <= '1';
    layer1_outputs(44) <= (layer0_outputs(537)) and not (layer0_outputs(1669));
    layer1_outputs(45) <= (layer0_outputs(1045)) xor (layer0_outputs(2482));
    layer1_outputs(46) <= (layer0_outputs(706)) and (layer0_outputs(893));
    layer1_outputs(47) <= (layer0_outputs(880)) and not (layer0_outputs(1683));
    layer1_outputs(48) <= layer0_outputs(2342);
    layer1_outputs(49) <= (layer0_outputs(1691)) or (layer0_outputs(1411));
    layer1_outputs(50) <= not(layer0_outputs(953)) or (layer0_outputs(813));
    layer1_outputs(51) <= layer0_outputs(73);
    layer1_outputs(52) <= not((layer0_outputs(1555)) or (layer0_outputs(2552)));
    layer1_outputs(53) <= layer0_outputs(72);
    layer1_outputs(54) <= (layer0_outputs(742)) xor (layer0_outputs(1146));
    layer1_outputs(55) <= (layer0_outputs(20)) and (layer0_outputs(414));
    layer1_outputs(56) <= not(layer0_outputs(1221)) or (layer0_outputs(865));
    layer1_outputs(57) <= (layer0_outputs(19)) or (layer0_outputs(1300));
    layer1_outputs(58) <= (layer0_outputs(852)) and not (layer0_outputs(310));
    layer1_outputs(59) <= layer0_outputs(1322);
    layer1_outputs(60) <= '1';
    layer1_outputs(61) <= not((layer0_outputs(2039)) and (layer0_outputs(615)));
    layer1_outputs(62) <= not(layer0_outputs(2104)) or (layer0_outputs(558));
    layer1_outputs(63) <= not(layer0_outputs(2074)) or (layer0_outputs(801));
    layer1_outputs(64) <= not(layer0_outputs(146));
    layer1_outputs(65) <= layer0_outputs(287);
    layer1_outputs(66) <= (layer0_outputs(870)) or (layer0_outputs(915));
    layer1_outputs(67) <= '0';
    layer1_outputs(68) <= not(layer0_outputs(1646));
    layer1_outputs(69) <= (layer0_outputs(1706)) and (layer0_outputs(2271));
    layer1_outputs(70) <= not(layer0_outputs(1525)) or (layer0_outputs(378));
    layer1_outputs(71) <= (layer0_outputs(1348)) and not (layer0_outputs(1301));
    layer1_outputs(72) <= (layer0_outputs(2085)) and not (layer0_outputs(330));
    layer1_outputs(73) <= not((layer0_outputs(259)) or (layer0_outputs(2544)));
    layer1_outputs(74) <= not((layer0_outputs(610)) or (layer0_outputs(456)));
    layer1_outputs(75) <= layer0_outputs(585);
    layer1_outputs(76) <= not(layer0_outputs(2049)) or (layer0_outputs(2320));
    layer1_outputs(77) <= not((layer0_outputs(902)) and (layer0_outputs(1836)));
    layer1_outputs(78) <= (layer0_outputs(1958)) and not (layer0_outputs(2051));
    layer1_outputs(79) <= layer0_outputs(1926);
    layer1_outputs(80) <= (layer0_outputs(1353)) and not (layer0_outputs(1611));
    layer1_outputs(81) <= '1';
    layer1_outputs(82) <= (layer0_outputs(2154)) or (layer0_outputs(845));
    layer1_outputs(83) <= (layer0_outputs(96)) and not (layer0_outputs(2361));
    layer1_outputs(84) <= (layer0_outputs(35)) and not (layer0_outputs(113));
    layer1_outputs(85) <= (layer0_outputs(149)) and not (layer0_outputs(2105));
    layer1_outputs(86) <= not(layer0_outputs(1678)) or (layer0_outputs(969));
    layer1_outputs(87) <= layer0_outputs(815);
    layer1_outputs(88) <= (layer0_outputs(2235)) and (layer0_outputs(252));
    layer1_outputs(89) <= not(layer0_outputs(1804)) or (layer0_outputs(676));
    layer1_outputs(90) <= '1';
    layer1_outputs(91) <= not((layer0_outputs(1713)) or (layer0_outputs(1597)));
    layer1_outputs(92) <= layer0_outputs(1093);
    layer1_outputs(93) <= layer0_outputs(2011);
    layer1_outputs(94) <= not(layer0_outputs(13)) or (layer0_outputs(2184));
    layer1_outputs(95) <= not((layer0_outputs(1090)) or (layer0_outputs(2286)));
    layer1_outputs(96) <= (layer0_outputs(54)) and not (layer0_outputs(996));
    layer1_outputs(97) <= not((layer0_outputs(379)) and (layer0_outputs(2460)));
    layer1_outputs(98) <= not(layer0_outputs(1538)) or (layer0_outputs(430));
    layer1_outputs(99) <= layer0_outputs(2359);
    layer1_outputs(100) <= (layer0_outputs(1878)) and not (layer0_outputs(2276));
    layer1_outputs(101) <= not(layer0_outputs(965));
    layer1_outputs(102) <= not((layer0_outputs(1522)) and (layer0_outputs(1760)));
    layer1_outputs(103) <= not(layer0_outputs(1562)) or (layer0_outputs(51));
    layer1_outputs(104) <= not(layer0_outputs(824)) or (layer0_outputs(2262));
    layer1_outputs(105) <= layer0_outputs(1871);
    layer1_outputs(106) <= (layer0_outputs(666)) or (layer0_outputs(1967));
    layer1_outputs(107) <= layer0_outputs(383);
    layer1_outputs(108) <= (layer0_outputs(1286)) or (layer0_outputs(509));
    layer1_outputs(109) <= not((layer0_outputs(1782)) or (layer0_outputs(1704)));
    layer1_outputs(110) <= (layer0_outputs(570)) and not (layer0_outputs(1812));
    layer1_outputs(111) <= (layer0_outputs(448)) or (layer0_outputs(980));
    layer1_outputs(112) <= '1';
    layer1_outputs(113) <= not(layer0_outputs(1163));
    layer1_outputs(114) <= not((layer0_outputs(1399)) or (layer0_outputs(796)));
    layer1_outputs(115) <= (layer0_outputs(512)) and not (layer0_outputs(983));
    layer1_outputs(116) <= (layer0_outputs(1263)) and not (layer0_outputs(959));
    layer1_outputs(117) <= (layer0_outputs(2372)) or (layer0_outputs(1738));
    layer1_outputs(118) <= not(layer0_outputs(19));
    layer1_outputs(119) <= not(layer0_outputs(22));
    layer1_outputs(120) <= layer0_outputs(997);
    layer1_outputs(121) <= (layer0_outputs(1227)) and not (layer0_outputs(1104));
    layer1_outputs(122) <= not((layer0_outputs(2513)) or (layer0_outputs(668)));
    layer1_outputs(123) <= layer0_outputs(2498);
    layer1_outputs(124) <= layer0_outputs(1911);
    layer1_outputs(125) <= (layer0_outputs(370)) or (layer0_outputs(678));
    layer1_outputs(126) <= not(layer0_outputs(2387)) or (layer0_outputs(250));
    layer1_outputs(127) <= layer0_outputs(2471);
    layer1_outputs(128) <= not((layer0_outputs(204)) or (layer0_outputs(1929)));
    layer1_outputs(129) <= not(layer0_outputs(1957));
    layer1_outputs(130) <= '0';
    layer1_outputs(131) <= (layer0_outputs(1775)) and (layer0_outputs(164));
    layer1_outputs(132) <= not((layer0_outputs(1112)) or (layer0_outputs(486)));
    layer1_outputs(133) <= not((layer0_outputs(2546)) xor (layer0_outputs(1672)));
    layer1_outputs(134) <= layer0_outputs(1405);
    layer1_outputs(135) <= (layer0_outputs(73)) and not (layer0_outputs(2210));
    layer1_outputs(136) <= '1';
    layer1_outputs(137) <= (layer0_outputs(1884)) and not (layer0_outputs(1302));
    layer1_outputs(138) <= (layer0_outputs(1673)) or (layer0_outputs(595));
    layer1_outputs(139) <= not(layer0_outputs(71));
    layer1_outputs(140) <= (layer0_outputs(1992)) and not (layer0_outputs(1743));
    layer1_outputs(141) <= (layer0_outputs(1431)) and (layer0_outputs(1944));
    layer1_outputs(142) <= layer0_outputs(2519);
    layer1_outputs(143) <= (layer0_outputs(2144)) and (layer0_outputs(2386));
    layer1_outputs(144) <= '0';
    layer1_outputs(145) <= not(layer0_outputs(1420));
    layer1_outputs(146) <= (layer0_outputs(1684)) and not (layer0_outputs(891));
    layer1_outputs(147) <= not((layer0_outputs(1428)) and (layer0_outputs(723)));
    layer1_outputs(148) <= (layer0_outputs(503)) and not (layer0_outputs(1182));
    layer1_outputs(149) <= (layer0_outputs(285)) or (layer0_outputs(157));
    layer1_outputs(150) <= (layer0_outputs(495)) and not (layer0_outputs(1895));
    layer1_outputs(151) <= '0';
    layer1_outputs(152) <= (layer0_outputs(1513)) and not (layer0_outputs(2385));
    layer1_outputs(153) <= not((layer0_outputs(2145)) and (layer0_outputs(2412)));
    layer1_outputs(154) <= '1';
    layer1_outputs(155) <= not(layer0_outputs(2301));
    layer1_outputs(156) <= layer0_outputs(2078);
    layer1_outputs(157) <= not(layer0_outputs(96)) or (layer0_outputs(2291));
    layer1_outputs(158) <= (layer0_outputs(1554)) or (layer0_outputs(550));
    layer1_outputs(159) <= (layer0_outputs(2447)) and (layer0_outputs(2479));
    layer1_outputs(160) <= not(layer0_outputs(2552));
    layer1_outputs(161) <= '1';
    layer1_outputs(162) <= not(layer0_outputs(1806));
    layer1_outputs(163) <= (layer0_outputs(2350)) or (layer0_outputs(2128));
    layer1_outputs(164) <= not(layer0_outputs(1840)) or (layer0_outputs(2076));
    layer1_outputs(165) <= (layer0_outputs(146)) and (layer0_outputs(1073));
    layer1_outputs(166) <= not(layer0_outputs(1133)) or (layer0_outputs(230));
    layer1_outputs(167) <= layer0_outputs(1712);
    layer1_outputs(168) <= not(layer0_outputs(2099)) or (layer0_outputs(571));
    layer1_outputs(169) <= (layer0_outputs(857)) or (layer0_outputs(1324));
    layer1_outputs(170) <= not((layer0_outputs(18)) and (layer0_outputs(581)));
    layer1_outputs(171) <= not((layer0_outputs(1860)) or (layer0_outputs(1783)));
    layer1_outputs(172) <= layer0_outputs(1666);
    layer1_outputs(173) <= '1';
    layer1_outputs(174) <= not(layer0_outputs(1717));
    layer1_outputs(175) <= not(layer0_outputs(751));
    layer1_outputs(176) <= (layer0_outputs(2027)) and (layer0_outputs(1383));
    layer1_outputs(177) <= not(layer0_outputs(2340)) or (layer0_outputs(118));
    layer1_outputs(178) <= (layer0_outputs(1715)) and not (layer0_outputs(1464));
    layer1_outputs(179) <= not(layer0_outputs(1737)) or (layer0_outputs(193));
    layer1_outputs(180) <= (layer0_outputs(547)) and (layer0_outputs(1353));
    layer1_outputs(181) <= layer0_outputs(392);
    layer1_outputs(182) <= not(layer0_outputs(29));
    layer1_outputs(183) <= '1';
    layer1_outputs(184) <= layer0_outputs(875);
    layer1_outputs(185) <= not(layer0_outputs(1864));
    layer1_outputs(186) <= '0';
    layer1_outputs(187) <= not(layer0_outputs(703)) or (layer0_outputs(1833));
    layer1_outputs(188) <= (layer0_outputs(685)) or (layer0_outputs(1326));
    layer1_outputs(189) <= not(layer0_outputs(1927)) or (layer0_outputs(91));
    layer1_outputs(190) <= not((layer0_outputs(2242)) and (layer0_outputs(2330)));
    layer1_outputs(191) <= (layer0_outputs(874)) or (layer0_outputs(320));
    layer1_outputs(192) <= (layer0_outputs(1896)) or (layer0_outputs(2457));
    layer1_outputs(193) <= not(layer0_outputs(2291));
    layer1_outputs(194) <= '0';
    layer1_outputs(195) <= not((layer0_outputs(252)) or (layer0_outputs(729)));
    layer1_outputs(196) <= not(layer0_outputs(2284));
    layer1_outputs(197) <= '0';
    layer1_outputs(198) <= not(layer0_outputs(544)) or (layer0_outputs(617));
    layer1_outputs(199) <= layer0_outputs(1012);
    layer1_outputs(200) <= layer0_outputs(145);
    layer1_outputs(201) <= not(layer0_outputs(498)) or (layer0_outputs(2452));
    layer1_outputs(202) <= not(layer0_outputs(1363)) or (layer0_outputs(1365));
    layer1_outputs(203) <= not(layer0_outputs(1655)) or (layer0_outputs(1492));
    layer1_outputs(204) <= not((layer0_outputs(592)) and (layer0_outputs(527)));
    layer1_outputs(205) <= not(layer0_outputs(2411));
    layer1_outputs(206) <= layer0_outputs(934);
    layer1_outputs(207) <= not(layer0_outputs(2516));
    layer1_outputs(208) <= '0';
    layer1_outputs(209) <= layer0_outputs(1401);
    layer1_outputs(210) <= not(layer0_outputs(1695)) or (layer0_outputs(2147));
    layer1_outputs(211) <= not((layer0_outputs(1619)) or (layer0_outputs(580)));
    layer1_outputs(212) <= not(layer0_outputs(1608)) or (layer0_outputs(541));
    layer1_outputs(213) <= not(layer0_outputs(928));
    layer1_outputs(214) <= layer0_outputs(1789);
    layer1_outputs(215) <= (layer0_outputs(2134)) xor (layer0_outputs(1265));
    layer1_outputs(216) <= (layer0_outputs(664)) and (layer0_outputs(1866));
    layer1_outputs(217) <= (layer0_outputs(399)) and not (layer0_outputs(1255));
    layer1_outputs(218) <= not(layer0_outputs(2043));
    layer1_outputs(219) <= (layer0_outputs(2025)) and not (layer0_outputs(1128));
    layer1_outputs(220) <= '0';
    layer1_outputs(221) <= not(layer0_outputs(1580)) or (layer0_outputs(1287));
    layer1_outputs(222) <= not(layer0_outputs(2498));
    layer1_outputs(223) <= layer0_outputs(47);
    layer1_outputs(224) <= layer0_outputs(1643);
    layer1_outputs(225) <= (layer0_outputs(83)) and not (layer0_outputs(1005));
    layer1_outputs(226) <= not((layer0_outputs(1661)) and (layer0_outputs(381)));
    layer1_outputs(227) <= '0';
    layer1_outputs(228) <= layer0_outputs(315);
    layer1_outputs(229) <= not(layer0_outputs(560)) or (layer0_outputs(522));
    layer1_outputs(230) <= (layer0_outputs(2186)) and not (layer0_outputs(1319));
    layer1_outputs(231) <= layer0_outputs(610);
    layer1_outputs(232) <= not(layer0_outputs(788)) or (layer0_outputs(844));
    layer1_outputs(233) <= not(layer0_outputs(730));
    layer1_outputs(234) <= '0';
    layer1_outputs(235) <= not((layer0_outputs(614)) or (layer0_outputs(2133)));
    layer1_outputs(236) <= layer0_outputs(1700);
    layer1_outputs(237) <= (layer0_outputs(487)) and not (layer0_outputs(108));
    layer1_outputs(238) <= not(layer0_outputs(1533));
    layer1_outputs(239) <= '1';
    layer1_outputs(240) <= '1';
    layer1_outputs(241) <= '1';
    layer1_outputs(242) <= (layer0_outputs(468)) and not (layer0_outputs(957));
    layer1_outputs(243) <= (layer0_outputs(1239)) xor (layer0_outputs(1708));
    layer1_outputs(244) <= '0';
    layer1_outputs(245) <= not(layer0_outputs(2110)) or (layer0_outputs(788));
    layer1_outputs(246) <= '0';
    layer1_outputs(247) <= not(layer0_outputs(194));
    layer1_outputs(248) <= not((layer0_outputs(2538)) xor (layer0_outputs(1650)));
    layer1_outputs(249) <= layer0_outputs(1610);
    layer1_outputs(250) <= not(layer0_outputs(2215));
    layer1_outputs(251) <= not((layer0_outputs(741)) and (layer0_outputs(1293)));
    layer1_outputs(252) <= not(layer0_outputs(1125));
    layer1_outputs(253) <= not(layer0_outputs(427)) or (layer0_outputs(307));
    layer1_outputs(254) <= layer0_outputs(1144);
    layer1_outputs(255) <= not(layer0_outputs(1952));
    layer1_outputs(256) <= not(layer0_outputs(2125));
    layer1_outputs(257) <= not(layer0_outputs(1008));
    layer1_outputs(258) <= not((layer0_outputs(191)) or (layer0_outputs(184)));
    layer1_outputs(259) <= (layer0_outputs(1155)) and not (layer0_outputs(2166));
    layer1_outputs(260) <= (layer0_outputs(766)) or (layer0_outputs(1742));
    layer1_outputs(261) <= layer0_outputs(1068);
    layer1_outputs(262) <= not(layer0_outputs(2371));
    layer1_outputs(263) <= layer0_outputs(1280);
    layer1_outputs(264) <= (layer0_outputs(1110)) and (layer0_outputs(1961));
    layer1_outputs(265) <= layer0_outputs(2400);
    layer1_outputs(266) <= (layer0_outputs(2180)) and not (layer0_outputs(2165));
    layer1_outputs(267) <= layer0_outputs(1735);
    layer1_outputs(268) <= '0';
    layer1_outputs(269) <= '0';
    layer1_outputs(270) <= (layer0_outputs(1763)) and not (layer0_outputs(2515));
    layer1_outputs(271) <= (layer0_outputs(136)) and not (layer0_outputs(1505));
    layer1_outputs(272) <= not(layer0_outputs(515)) or (layer0_outputs(1252));
    layer1_outputs(273) <= (layer0_outputs(1948)) xor (layer0_outputs(2017));
    layer1_outputs(274) <= not(layer0_outputs(1956)) or (layer0_outputs(134));
    layer1_outputs(275) <= (layer0_outputs(237)) and (layer0_outputs(2026));
    layer1_outputs(276) <= not(layer0_outputs(1118));
    layer1_outputs(277) <= not(layer0_outputs(1757));
    layer1_outputs(278) <= not(layer0_outputs(2054));
    layer1_outputs(279) <= not((layer0_outputs(1636)) xor (layer0_outputs(2091)));
    layer1_outputs(280) <= '1';
    layer1_outputs(281) <= not((layer0_outputs(2136)) and (layer0_outputs(2444)));
    layer1_outputs(282) <= (layer0_outputs(1348)) and not (layer0_outputs(461));
    layer1_outputs(283) <= not((layer0_outputs(1451)) and (layer0_outputs(611)));
    layer1_outputs(284) <= layer0_outputs(464);
    layer1_outputs(285) <= not(layer0_outputs(2405));
    layer1_outputs(286) <= (layer0_outputs(792)) and not (layer0_outputs(1876));
    layer1_outputs(287) <= (layer0_outputs(1714)) and not (layer0_outputs(1667));
    layer1_outputs(288) <= not(layer0_outputs(530));
    layer1_outputs(289) <= layer0_outputs(2266);
    layer1_outputs(290) <= (layer0_outputs(64)) and not (layer0_outputs(742));
    layer1_outputs(291) <= not(layer0_outputs(1819));
    layer1_outputs(292) <= layer0_outputs(1499);
    layer1_outputs(293) <= not(layer0_outputs(1733));
    layer1_outputs(294) <= layer0_outputs(222);
    layer1_outputs(295) <= '0';
    layer1_outputs(296) <= not((layer0_outputs(2392)) and (layer0_outputs(1210)));
    layer1_outputs(297) <= (layer0_outputs(430)) and (layer0_outputs(2222));
    layer1_outputs(298) <= '1';
    layer1_outputs(299) <= not(layer0_outputs(1022)) or (layer0_outputs(2047));
    layer1_outputs(300) <= not((layer0_outputs(684)) or (layer0_outputs(1728)));
    layer1_outputs(301) <= (layer0_outputs(794)) and not (layer0_outputs(2288));
    layer1_outputs(302) <= '0';
    layer1_outputs(303) <= layer0_outputs(2175);
    layer1_outputs(304) <= '1';
    layer1_outputs(305) <= layer0_outputs(2331);
    layer1_outputs(306) <= not(layer0_outputs(1623)) or (layer0_outputs(1018));
    layer1_outputs(307) <= (layer0_outputs(1460)) and not (layer0_outputs(1893));
    layer1_outputs(308) <= not(layer0_outputs(2358));
    layer1_outputs(309) <= not(layer0_outputs(1299));
    layer1_outputs(310) <= not(layer0_outputs(504));
    layer1_outputs(311) <= not(layer0_outputs(2354)) or (layer0_outputs(583));
    layer1_outputs(312) <= layer0_outputs(558);
    layer1_outputs(313) <= not((layer0_outputs(2430)) or (layer0_outputs(2532)));
    layer1_outputs(314) <= not((layer0_outputs(688)) and (layer0_outputs(277)));
    layer1_outputs(315) <= '1';
    layer1_outputs(316) <= not(layer0_outputs(1090));
    layer1_outputs(317) <= layer0_outputs(632);
    layer1_outputs(318) <= '1';
    layer1_outputs(319) <= '1';
    layer1_outputs(320) <= '0';
    layer1_outputs(321) <= (layer0_outputs(1896)) and (layer0_outputs(698));
    layer1_outputs(322) <= not((layer0_outputs(59)) or (layer0_outputs(2456)));
    layer1_outputs(323) <= '1';
    layer1_outputs(324) <= '1';
    layer1_outputs(325) <= not((layer0_outputs(1477)) and (layer0_outputs(2360)));
    layer1_outputs(326) <= not((layer0_outputs(821)) or (layer0_outputs(138)));
    layer1_outputs(327) <= (layer0_outputs(2038)) and (layer0_outputs(1320));
    layer1_outputs(328) <= (layer0_outputs(376)) xor (layer0_outputs(500));
    layer1_outputs(329) <= not((layer0_outputs(677)) and (layer0_outputs(30)));
    layer1_outputs(330) <= not(layer0_outputs(2379));
    layer1_outputs(331) <= layer0_outputs(722);
    layer1_outputs(332) <= not((layer0_outputs(1712)) or (layer0_outputs(1596)));
    layer1_outputs(333) <= '1';
    layer1_outputs(334) <= not(layer0_outputs(140)) or (layer0_outputs(517));
    layer1_outputs(335) <= (layer0_outputs(1688)) or (layer0_outputs(408));
    layer1_outputs(336) <= not((layer0_outputs(1251)) or (layer0_outputs(381)));
    layer1_outputs(337) <= not(layer0_outputs(2216)) or (layer0_outputs(692));
    layer1_outputs(338) <= not(layer0_outputs(82));
    layer1_outputs(339) <= layer0_outputs(90);
    layer1_outputs(340) <= layer0_outputs(1861);
    layer1_outputs(341) <= '1';
    layer1_outputs(342) <= '0';
    layer1_outputs(343) <= not((layer0_outputs(947)) or (layer0_outputs(1457)));
    layer1_outputs(344) <= not((layer0_outputs(614)) or (layer0_outputs(1572)));
    layer1_outputs(345) <= (layer0_outputs(1250)) and (layer0_outputs(1435));
    layer1_outputs(346) <= (layer0_outputs(785)) and not (layer0_outputs(368));
    layer1_outputs(347) <= layer0_outputs(2381);
    layer1_outputs(348) <= layer0_outputs(2330);
    layer1_outputs(349) <= (layer0_outputs(700)) or (layer0_outputs(797));
    layer1_outputs(350) <= (layer0_outputs(766)) and not (layer0_outputs(71));
    layer1_outputs(351) <= not(layer0_outputs(2472));
    layer1_outputs(352) <= not(layer0_outputs(2324));
    layer1_outputs(353) <= (layer0_outputs(1038)) or (layer0_outputs(1559));
    layer1_outputs(354) <= layer0_outputs(458);
    layer1_outputs(355) <= layer0_outputs(1827);
    layer1_outputs(356) <= '0';
    layer1_outputs(357) <= (layer0_outputs(1932)) or (layer0_outputs(1800));
    layer1_outputs(358) <= '1';
    layer1_outputs(359) <= '0';
    layer1_outputs(360) <= '1';
    layer1_outputs(361) <= not(layer0_outputs(42));
    layer1_outputs(362) <= (layer0_outputs(453)) and not (layer0_outputs(1306));
    layer1_outputs(363) <= '0';
    layer1_outputs(364) <= not(layer0_outputs(326));
    layer1_outputs(365) <= '0';
    layer1_outputs(366) <= not(layer0_outputs(1571)) or (layer0_outputs(740));
    layer1_outputs(367) <= layer0_outputs(479);
    layer1_outputs(368) <= '0';
    layer1_outputs(369) <= not(layer0_outputs(526)) or (layer0_outputs(2197));
    layer1_outputs(370) <= not(layer0_outputs(1094)) or (layer0_outputs(2376));
    layer1_outputs(371) <= (layer0_outputs(1285)) and not (layer0_outputs(571));
    layer1_outputs(372) <= not(layer0_outputs(447)) or (layer0_outputs(2274));
    layer1_outputs(373) <= layer0_outputs(1835);
    layer1_outputs(374) <= layer0_outputs(510);
    layer1_outputs(375) <= (layer0_outputs(208)) and (layer0_outputs(1764));
    layer1_outputs(376) <= (layer0_outputs(1681)) or (layer0_outputs(202));
    layer1_outputs(377) <= (layer0_outputs(221)) and (layer0_outputs(44));
    layer1_outputs(378) <= (layer0_outputs(636)) and not (layer0_outputs(1088));
    layer1_outputs(379) <= layer0_outputs(1366);
    layer1_outputs(380) <= not((layer0_outputs(426)) or (layer0_outputs(1168)));
    layer1_outputs(381) <= layer0_outputs(2344);
    layer1_outputs(382) <= (layer0_outputs(1320)) and not (layer0_outputs(1598));
    layer1_outputs(383) <= (layer0_outputs(738)) and not (layer0_outputs(2337));
    layer1_outputs(384) <= not((layer0_outputs(2433)) and (layer0_outputs(1289)));
    layer1_outputs(385) <= not(layer0_outputs(2013)) or (layer0_outputs(804));
    layer1_outputs(386) <= (layer0_outputs(1363)) or (layer0_outputs(800));
    layer1_outputs(387) <= layer0_outputs(407);
    layer1_outputs(388) <= layer0_outputs(249);
    layer1_outputs(389) <= not((layer0_outputs(1356)) and (layer0_outputs(641)));
    layer1_outputs(390) <= layer0_outputs(854);
    layer1_outputs(391) <= layer0_outputs(1955);
    layer1_outputs(392) <= not((layer0_outputs(1274)) and (layer0_outputs(843)));
    layer1_outputs(393) <= not((layer0_outputs(1387)) or (layer0_outputs(2062)));
    layer1_outputs(394) <= not(layer0_outputs(1092));
    layer1_outputs(395) <= not((layer0_outputs(559)) and (layer0_outputs(1191)));
    layer1_outputs(396) <= layer0_outputs(283);
    layer1_outputs(397) <= not(layer0_outputs(2401));
    layer1_outputs(398) <= layer0_outputs(1546);
    layer1_outputs(399) <= (layer0_outputs(1872)) and (layer0_outputs(403));
    layer1_outputs(400) <= '0';
    layer1_outputs(401) <= '1';
    layer1_outputs(402) <= (layer0_outputs(1561)) and not (layer0_outputs(182));
    layer1_outputs(403) <= '0';
    layer1_outputs(404) <= not((layer0_outputs(1006)) or (layer0_outputs(2005)));
    layer1_outputs(405) <= (layer0_outputs(1759)) and (layer0_outputs(851));
    layer1_outputs(406) <= (layer0_outputs(65)) and (layer0_outputs(2402));
    layer1_outputs(407) <= (layer0_outputs(1864)) and (layer0_outputs(2446));
    layer1_outputs(408) <= not((layer0_outputs(661)) and (layer0_outputs(2042)));
    layer1_outputs(409) <= layer0_outputs(916);
    layer1_outputs(410) <= layer0_outputs(2191);
    layer1_outputs(411) <= layer0_outputs(474);
    layer1_outputs(412) <= (layer0_outputs(1512)) and not (layer0_outputs(2171));
    layer1_outputs(413) <= layer0_outputs(326);
    layer1_outputs(414) <= layer0_outputs(478);
    layer1_outputs(415) <= (layer0_outputs(1309)) and not (layer0_outputs(411));
    layer1_outputs(416) <= not(layer0_outputs(762));
    layer1_outputs(417) <= layer0_outputs(1132);
    layer1_outputs(418) <= (layer0_outputs(1868)) or (layer0_outputs(2292));
    layer1_outputs(419) <= (layer0_outputs(1882)) and not (layer0_outputs(871));
    layer1_outputs(420) <= (layer0_outputs(2500)) and (layer0_outputs(1608));
    layer1_outputs(421) <= layer0_outputs(1032);
    layer1_outputs(422) <= '1';
    layer1_outputs(423) <= '0';
    layer1_outputs(424) <= (layer0_outputs(696)) and (layer0_outputs(1118));
    layer1_outputs(425) <= layer0_outputs(1739);
    layer1_outputs(426) <= '1';
    layer1_outputs(427) <= not(layer0_outputs(520)) or (layer0_outputs(2233));
    layer1_outputs(428) <= layer0_outputs(85);
    layer1_outputs(429) <= not(layer0_outputs(1006)) or (layer0_outputs(2526));
    layer1_outputs(430) <= '1';
    layer1_outputs(431) <= (layer0_outputs(535)) and not (layer0_outputs(2533));
    layer1_outputs(432) <= not(layer0_outputs(828));
    layer1_outputs(433) <= (layer0_outputs(969)) and not (layer0_outputs(2181));
    layer1_outputs(434) <= not((layer0_outputs(1244)) and (layer0_outputs(1834)));
    layer1_outputs(435) <= not((layer0_outputs(1108)) and (layer0_outputs(199)));
    layer1_outputs(436) <= not(layer0_outputs(2233));
    layer1_outputs(437) <= (layer0_outputs(12)) or (layer0_outputs(247));
    layer1_outputs(438) <= '0';
    layer1_outputs(439) <= not(layer0_outputs(2117));
    layer1_outputs(440) <= '0';
    layer1_outputs(441) <= not(layer0_outputs(1381));
    layer1_outputs(442) <= not((layer0_outputs(1156)) or (layer0_outputs(351)));
    layer1_outputs(443) <= '0';
    layer1_outputs(444) <= not(layer0_outputs(1236));
    layer1_outputs(445) <= (layer0_outputs(552)) and not (layer0_outputs(1291));
    layer1_outputs(446) <= (layer0_outputs(74)) and not (layer0_outputs(1370));
    layer1_outputs(447) <= not(layer0_outputs(485)) or (layer0_outputs(1447));
    layer1_outputs(448) <= not((layer0_outputs(1407)) and (layer0_outputs(1604)));
    layer1_outputs(449) <= (layer0_outputs(1705)) xor (layer0_outputs(546));
    layer1_outputs(450) <= not((layer0_outputs(831)) or (layer0_outputs(2104)));
    layer1_outputs(451) <= not(layer0_outputs(422)) or (layer0_outputs(888));
    layer1_outputs(452) <= not(layer0_outputs(745)) or (layer0_outputs(1737));
    layer1_outputs(453) <= (layer0_outputs(2244)) or (layer0_outputs(1804));
    layer1_outputs(454) <= '1';
    layer1_outputs(455) <= (layer0_outputs(1234)) and (layer0_outputs(2286));
    layer1_outputs(456) <= '0';
    layer1_outputs(457) <= (layer0_outputs(1589)) and not (layer0_outputs(2160));
    layer1_outputs(458) <= (layer0_outputs(40)) or (layer0_outputs(333));
    layer1_outputs(459) <= layer0_outputs(516);
    layer1_outputs(460) <= not((layer0_outputs(1955)) or (layer0_outputs(1526)));
    layer1_outputs(461) <= (layer0_outputs(1918)) and (layer0_outputs(1357));
    layer1_outputs(462) <= layer0_outputs(1825);
    layer1_outputs(463) <= '1';
    layer1_outputs(464) <= (layer0_outputs(1490)) and (layer0_outputs(1186));
    layer1_outputs(465) <= not((layer0_outputs(1204)) and (layer0_outputs(294)));
    layer1_outputs(466) <= (layer0_outputs(1718)) or (layer0_outputs(1854));
    layer1_outputs(467) <= not(layer0_outputs(2138)) or (layer0_outputs(204));
    layer1_outputs(468) <= layer0_outputs(1225);
    layer1_outputs(469) <= (layer0_outputs(633)) and not (layer0_outputs(1445));
    layer1_outputs(470) <= (layer0_outputs(2179)) and not (layer0_outputs(194));
    layer1_outputs(471) <= not(layer0_outputs(415));
    layer1_outputs(472) <= (layer0_outputs(2006)) or (layer0_outputs(805));
    layer1_outputs(473) <= '1';
    layer1_outputs(474) <= (layer0_outputs(1867)) and (layer0_outputs(1262));
    layer1_outputs(475) <= (layer0_outputs(717)) and (layer0_outputs(1380));
    layer1_outputs(476) <= (layer0_outputs(884)) or (layer0_outputs(1461));
    layer1_outputs(477) <= (layer0_outputs(2468)) and not (layer0_outputs(1606));
    layer1_outputs(478) <= (layer0_outputs(108)) and (layer0_outputs(997));
    layer1_outputs(479) <= not(layer0_outputs(1710));
    layer1_outputs(480) <= '1';
    layer1_outputs(481) <= (layer0_outputs(2003)) and not (layer0_outputs(147));
    layer1_outputs(482) <= not((layer0_outputs(473)) xor (layer0_outputs(1759)));
    layer1_outputs(483) <= (layer0_outputs(2380)) or (layer0_outputs(1009));
    layer1_outputs(484) <= not(layer0_outputs(1066)) or (layer0_outputs(2549));
    layer1_outputs(485) <= (layer0_outputs(569)) and not (layer0_outputs(110));
    layer1_outputs(486) <= '0';
    layer1_outputs(487) <= not(layer0_outputs(2036)) or (layer0_outputs(2056));
    layer1_outputs(488) <= (layer0_outputs(1898)) and not (layer0_outputs(489));
    layer1_outputs(489) <= not((layer0_outputs(664)) and (layer0_outputs(2558)));
    layer1_outputs(490) <= (layer0_outputs(1654)) and not (layer0_outputs(1810));
    layer1_outputs(491) <= not(layer0_outputs(1279));
    layer1_outputs(492) <= not((layer0_outputs(233)) and (layer0_outputs(1741)));
    layer1_outputs(493) <= layer0_outputs(1097);
    layer1_outputs(494) <= '0';
    layer1_outputs(495) <= (layer0_outputs(2263)) or (layer0_outputs(335));
    layer1_outputs(496) <= not(layer0_outputs(526)) or (layer0_outputs(2274));
    layer1_outputs(497) <= (layer0_outputs(1083)) and not (layer0_outputs(1667));
    layer1_outputs(498) <= '0';
    layer1_outputs(499) <= layer0_outputs(1765);
    layer1_outputs(500) <= not(layer0_outputs(1798)) or (layer0_outputs(2114));
    layer1_outputs(501) <= not(layer0_outputs(1687));
    layer1_outputs(502) <= layer0_outputs(791);
    layer1_outputs(503) <= not(layer0_outputs(720)) or (layer0_outputs(877));
    layer1_outputs(504) <= layer0_outputs(1275);
    layer1_outputs(505) <= not(layer0_outputs(253)) or (layer0_outputs(1037));
    layer1_outputs(506) <= (layer0_outputs(2178)) and not (layer0_outputs(1429));
    layer1_outputs(507) <= not(layer0_outputs(1066));
    layer1_outputs(508) <= not(layer0_outputs(479)) or (layer0_outputs(529));
    layer1_outputs(509) <= not((layer0_outputs(76)) or (layer0_outputs(377)));
    layer1_outputs(510) <= layer0_outputs(578);
    layer1_outputs(511) <= layer0_outputs(1261);
    layer1_outputs(512) <= '1';
    layer1_outputs(513) <= not((layer0_outputs(1998)) or (layer0_outputs(1373)));
    layer1_outputs(514) <= not(layer0_outputs(2158));
    layer1_outputs(515) <= not((layer0_outputs(774)) or (layer0_outputs(2114)));
    layer1_outputs(516) <= '0';
    layer1_outputs(517) <= not((layer0_outputs(268)) and (layer0_outputs(955)));
    layer1_outputs(518) <= layer0_outputs(254);
    layer1_outputs(519) <= not(layer0_outputs(2454)) or (layer0_outputs(1576));
    layer1_outputs(520) <= '1';
    layer1_outputs(521) <= layer0_outputs(990);
    layer1_outputs(522) <= not(layer0_outputs(2482)) or (layer0_outputs(1439));
    layer1_outputs(523) <= (layer0_outputs(1892)) and not (layer0_outputs(388));
    layer1_outputs(524) <= not((layer0_outputs(820)) and (layer0_outputs(1088)));
    layer1_outputs(525) <= not(layer0_outputs(986));
    layer1_outputs(526) <= not((layer0_outputs(2095)) or (layer0_outputs(1155)));
    layer1_outputs(527) <= not(layer0_outputs(1497)) or (layer0_outputs(2132));
    layer1_outputs(528) <= layer0_outputs(267);
    layer1_outputs(529) <= not((layer0_outputs(384)) and (layer0_outputs(1000)));
    layer1_outputs(530) <= (layer0_outputs(2295)) or (layer0_outputs(899));
    layer1_outputs(531) <= not((layer0_outputs(674)) or (layer0_outputs(1209)));
    layer1_outputs(532) <= layer0_outputs(2224);
    layer1_outputs(533) <= not((layer0_outputs(389)) and (layer0_outputs(609)));
    layer1_outputs(534) <= not(layer0_outputs(465)) or (layer0_outputs(1963));
    layer1_outputs(535) <= not((layer0_outputs(1623)) or (layer0_outputs(1983)));
    layer1_outputs(536) <= layer0_outputs(1772);
    layer1_outputs(537) <= not(layer0_outputs(760)) or (layer0_outputs(89));
    layer1_outputs(538) <= '1';
    layer1_outputs(539) <= not((layer0_outputs(238)) and (layer0_outputs(489)));
    layer1_outputs(540) <= not(layer0_outputs(1994)) or (layer0_outputs(2040));
    layer1_outputs(541) <= not(layer0_outputs(1433));
    layer1_outputs(542) <= '1';
    layer1_outputs(543) <= not(layer0_outputs(2105));
    layer1_outputs(544) <= (layer0_outputs(2109)) and not (layer0_outputs(264));
    layer1_outputs(545) <= '0';
    layer1_outputs(546) <= not((layer0_outputs(703)) and (layer0_outputs(1494)));
    layer1_outputs(547) <= (layer0_outputs(1204)) and not (layer0_outputs(2287));
    layer1_outputs(548) <= (layer0_outputs(629)) or (layer0_outputs(1496));
    layer1_outputs(549) <= not(layer0_outputs(105)) or (layer0_outputs(590));
    layer1_outputs(550) <= not(layer0_outputs(390));
    layer1_outputs(551) <= (layer0_outputs(1442)) and not (layer0_outputs(699));
    layer1_outputs(552) <= not(layer0_outputs(1686));
    layer1_outputs(553) <= not(layer0_outputs(877)) or (layer0_outputs(465));
    layer1_outputs(554) <= not(layer0_outputs(1143));
    layer1_outputs(555) <= not((layer0_outputs(399)) and (layer0_outputs(1655)));
    layer1_outputs(556) <= not(layer0_outputs(1772));
    layer1_outputs(557) <= not(layer0_outputs(1492));
    layer1_outputs(558) <= not((layer0_outputs(1349)) or (layer0_outputs(303)));
    layer1_outputs(559) <= (layer0_outputs(1885)) and (layer0_outputs(1219));
    layer1_outputs(560) <= layer0_outputs(756);
    layer1_outputs(561) <= not(layer0_outputs(309));
    layer1_outputs(562) <= (layer0_outputs(687)) and not (layer0_outputs(1496));
    layer1_outputs(563) <= not((layer0_outputs(103)) and (layer0_outputs(1078)));
    layer1_outputs(564) <= (layer0_outputs(2090)) or (layer0_outputs(160));
    layer1_outputs(565) <= '0';
    layer1_outputs(566) <= (layer0_outputs(1277)) and not (layer0_outputs(2488));
    layer1_outputs(567) <= not(layer0_outputs(696)) or (layer0_outputs(596));
    layer1_outputs(568) <= not(layer0_outputs(2259)) or (layer0_outputs(1185));
    layer1_outputs(569) <= layer0_outputs(1468);
    layer1_outputs(570) <= (layer0_outputs(597)) and not (layer0_outputs(774));
    layer1_outputs(571) <= not((layer0_outputs(1950)) xor (layer0_outputs(127)));
    layer1_outputs(572) <= not((layer0_outputs(1375)) or (layer0_outputs(1326)));
    layer1_outputs(573) <= not(layer0_outputs(2475)) or (layer0_outputs(2001));
    layer1_outputs(574) <= not(layer0_outputs(1602)) or (layer0_outputs(2374));
    layer1_outputs(575) <= (layer0_outputs(2304)) and (layer0_outputs(978));
    layer1_outputs(576) <= (layer0_outputs(1914)) or (layer0_outputs(1177));
    layer1_outputs(577) <= not((layer0_outputs(476)) and (layer0_outputs(2188)));
    layer1_outputs(578) <= (layer0_outputs(1045)) and not (layer0_outputs(2118));
    layer1_outputs(579) <= not(layer0_outputs(2014)) or (layer0_outputs(2234));
    layer1_outputs(580) <= (layer0_outputs(1983)) and not (layer0_outputs(1960));
    layer1_outputs(581) <= layer0_outputs(2491);
    layer1_outputs(582) <= layer0_outputs(2124);
    layer1_outputs(583) <= '1';
    layer1_outputs(584) <= not(layer0_outputs(1404));
    layer1_outputs(585) <= (layer0_outputs(2415)) and (layer0_outputs(691));
    layer1_outputs(586) <= (layer0_outputs(2003)) and not (layer0_outputs(923));
    layer1_outputs(587) <= (layer0_outputs(622)) or (layer0_outputs(1926));
    layer1_outputs(588) <= (layer0_outputs(1190)) and not (layer0_outputs(1902));
    layer1_outputs(589) <= not(layer0_outputs(1023)) or (layer0_outputs(1026));
    layer1_outputs(590) <= '0';
    layer1_outputs(591) <= not(layer0_outputs(1079));
    layer1_outputs(592) <= layer0_outputs(2188);
    layer1_outputs(593) <= (layer0_outputs(1041)) and not (layer0_outputs(1036));
    layer1_outputs(594) <= layer0_outputs(519);
    layer1_outputs(595) <= layer0_outputs(2307);
    layer1_outputs(596) <= (layer0_outputs(416)) and not (layer0_outputs(1933));
    layer1_outputs(597) <= '0';
    layer1_outputs(598) <= '1';
    layer1_outputs(599) <= not(layer0_outputs(239));
    layer1_outputs(600) <= not((layer0_outputs(1650)) or (layer0_outputs(2451)));
    layer1_outputs(601) <= not(layer0_outputs(606));
    layer1_outputs(602) <= (layer0_outputs(429)) and not (layer0_outputs(395));
    layer1_outputs(603) <= not(layer0_outputs(2192)) or (layer0_outputs(266));
    layer1_outputs(604) <= '0';
    layer1_outputs(605) <= not(layer0_outputs(133));
    layer1_outputs(606) <= (layer0_outputs(219)) and not (layer0_outputs(1109));
    layer1_outputs(607) <= (layer0_outputs(106)) and (layer0_outputs(1959));
    layer1_outputs(608) <= (layer0_outputs(2193)) and (layer0_outputs(1605));
    layer1_outputs(609) <= not(layer0_outputs(1777)) or (layer0_outputs(697));
    layer1_outputs(610) <= (layer0_outputs(1641)) and not (layer0_outputs(2417));
    layer1_outputs(611) <= not((layer0_outputs(931)) or (layer0_outputs(366)));
    layer1_outputs(612) <= not((layer0_outputs(2094)) and (layer0_outputs(462)));
    layer1_outputs(613) <= (layer0_outputs(1022)) and (layer0_outputs(542));
    layer1_outputs(614) <= not(layer0_outputs(1273));
    layer1_outputs(615) <= layer0_outputs(1323);
    layer1_outputs(616) <= not(layer0_outputs(1099));
    layer1_outputs(617) <= layer0_outputs(655);
    layer1_outputs(618) <= not((layer0_outputs(1345)) or (layer0_outputs(2399)));
    layer1_outputs(619) <= (layer0_outputs(2148)) xor (layer0_outputs(121));
    layer1_outputs(620) <= not(layer0_outputs(1782));
    layer1_outputs(621) <= layer0_outputs(2306);
    layer1_outputs(622) <= not((layer0_outputs(35)) and (layer0_outputs(299)));
    layer1_outputs(623) <= '0';
    layer1_outputs(624) <= not(layer0_outputs(314));
    layer1_outputs(625) <= not(layer0_outputs(2237));
    layer1_outputs(626) <= (layer0_outputs(644)) and not (layer0_outputs(1425));
    layer1_outputs(627) <= '0';
    layer1_outputs(628) <= not(layer0_outputs(1462));
    layer1_outputs(629) <= not((layer0_outputs(2066)) or (layer0_outputs(209)));
    layer1_outputs(630) <= (layer0_outputs(198)) and not (layer0_outputs(2557));
    layer1_outputs(631) <= '1';
    layer1_outputs(632) <= (layer0_outputs(394)) or (layer0_outputs(2048));
    layer1_outputs(633) <= not(layer0_outputs(752));
    layer1_outputs(634) <= not((layer0_outputs(1126)) or (layer0_outputs(403)));
    layer1_outputs(635) <= (layer0_outputs(1874)) and not (layer0_outputs(2469));
    layer1_outputs(636) <= (layer0_outputs(1203)) and (layer0_outputs(1028));
    layer1_outputs(637) <= layer0_outputs(1025);
    layer1_outputs(638) <= not(layer0_outputs(2310));
    layer1_outputs(639) <= '0';
    layer1_outputs(640) <= not(layer0_outputs(91)) or (layer0_outputs(2057));
    layer1_outputs(641) <= layer0_outputs(1084);
    layer1_outputs(642) <= layer0_outputs(1557);
    layer1_outputs(643) <= (layer0_outputs(1036)) or (layer0_outputs(906));
    layer1_outputs(644) <= (layer0_outputs(2554)) and (layer0_outputs(2112));
    layer1_outputs(645) <= (layer0_outputs(1987)) and not (layer0_outputs(1484));
    layer1_outputs(646) <= (layer0_outputs(2139)) and not (layer0_outputs(782));
    layer1_outputs(647) <= layer0_outputs(1084);
    layer1_outputs(648) <= (layer0_outputs(1769)) or (layer0_outputs(1511));
    layer1_outputs(649) <= '1';
    layer1_outputs(650) <= layer0_outputs(129);
    layer1_outputs(651) <= layer0_outputs(1832);
    layer1_outputs(652) <= not((layer0_outputs(1493)) xor (layer0_outputs(1494)));
    layer1_outputs(653) <= not(layer0_outputs(86)) or (layer0_outputs(67));
    layer1_outputs(654) <= not((layer0_outputs(2409)) or (layer0_outputs(1419)));
    layer1_outputs(655) <= not((layer0_outputs(1120)) or (layer0_outputs(1846)));
    layer1_outputs(656) <= '1';
    layer1_outputs(657) <= '1';
    layer1_outputs(658) <= not(layer0_outputs(70)) or (layer0_outputs(770));
    layer1_outputs(659) <= not(layer0_outputs(1304)) or (layer0_outputs(1015));
    layer1_outputs(660) <= (layer0_outputs(977)) and not (layer0_outputs(2012));
    layer1_outputs(661) <= layer0_outputs(860);
    layer1_outputs(662) <= layer0_outputs(1360);
    layer1_outputs(663) <= (layer0_outputs(1890)) or (layer0_outputs(365));
    layer1_outputs(664) <= not(layer0_outputs(2496));
    layer1_outputs(665) <= not(layer0_outputs(1559)) or (layer0_outputs(1632));
    layer1_outputs(666) <= not(layer0_outputs(2492)) or (layer0_outputs(1705));
    layer1_outputs(667) <= layer0_outputs(135);
    layer1_outputs(668) <= not((layer0_outputs(2428)) or (layer0_outputs(1481)));
    layer1_outputs(669) <= not((layer0_outputs(2492)) and (layer0_outputs(580)));
    layer1_outputs(670) <= layer0_outputs(2087);
    layer1_outputs(671) <= (layer0_outputs(987)) and not (layer0_outputs(1273));
    layer1_outputs(672) <= not((layer0_outputs(357)) or (layer0_outputs(461)));
    layer1_outputs(673) <= not(layer0_outputs(822)) or (layer0_outputs(1100));
    layer1_outputs(674) <= layer0_outputs(920);
    layer1_outputs(675) <= not(layer0_outputs(822)) or (layer0_outputs(652));
    layer1_outputs(676) <= not(layer0_outputs(418));
    layer1_outputs(677) <= '1';
    layer1_outputs(678) <= not(layer0_outputs(1389));
    layer1_outputs(679) <= (layer0_outputs(1158)) and not (layer0_outputs(496));
    layer1_outputs(680) <= (layer0_outputs(853)) and (layer0_outputs(985));
    layer1_outputs(681) <= not((layer0_outputs(2249)) or (layer0_outputs(579)));
    layer1_outputs(682) <= not(layer0_outputs(2494));
    layer1_outputs(683) <= not((layer0_outputs(328)) or (layer0_outputs(1803)));
    layer1_outputs(684) <= layer0_outputs(61);
    layer1_outputs(685) <= not((layer0_outputs(2073)) and (layer0_outputs(1292)));
    layer1_outputs(686) <= not(layer0_outputs(1573)) or (layer0_outputs(1709));
    layer1_outputs(687) <= not((layer0_outputs(2124)) and (layer0_outputs(875)));
    layer1_outputs(688) <= not((layer0_outputs(301)) xor (layer0_outputs(1749)));
    layer1_outputs(689) <= not((layer0_outputs(1242)) and (layer0_outputs(1451)));
    layer1_outputs(690) <= (layer0_outputs(1726)) and not (layer0_outputs(2179));
    layer1_outputs(691) <= not(layer0_outputs(2529));
    layer1_outputs(692) <= not((layer0_outputs(1930)) and (layer0_outputs(812)));
    layer1_outputs(693) <= not((layer0_outputs(2346)) xor (layer0_outputs(189)));
    layer1_outputs(694) <= (layer0_outputs(1580)) or (layer0_outputs(819));
    layer1_outputs(695) <= not((layer0_outputs(216)) xor (layer0_outputs(169)));
    layer1_outputs(696) <= not(layer0_outputs(2443));
    layer1_outputs(697) <= not(layer0_outputs(42));
    layer1_outputs(698) <= layer0_outputs(2517);
    layer1_outputs(699) <= not(layer0_outputs(2429)) or (layer0_outputs(616));
    layer1_outputs(700) <= not(layer0_outputs(1421)) or (layer0_outputs(1742));
    layer1_outputs(701) <= layer0_outputs(1124);
    layer1_outputs(702) <= not(layer0_outputs(805)) or (layer0_outputs(270));
    layer1_outputs(703) <= not(layer0_outputs(1339));
    layer1_outputs(704) <= not((layer0_outputs(2378)) and (layer0_outputs(686)));
    layer1_outputs(705) <= not(layer0_outputs(1530)) or (layer0_outputs(14));
    layer1_outputs(706) <= not(layer0_outputs(23)) or (layer0_outputs(1573));
    layer1_outputs(707) <= (layer0_outputs(563)) and not (layer0_outputs(411));
    layer1_outputs(708) <= (layer0_outputs(651)) or (layer0_outputs(51));
    layer1_outputs(709) <= (layer0_outputs(2307)) and not (layer0_outputs(2225));
    layer1_outputs(710) <= '1';
    layer1_outputs(711) <= not(layer0_outputs(2494)) or (layer0_outputs(1202));
    layer1_outputs(712) <= (layer0_outputs(1276)) and not (layer0_outputs(289));
    layer1_outputs(713) <= not((layer0_outputs(1062)) or (layer0_outputs(650)));
    layer1_outputs(714) <= not(layer0_outputs(287));
    layer1_outputs(715) <= (layer0_outputs(1181)) or (layer0_outputs(1344));
    layer1_outputs(716) <= (layer0_outputs(2469)) and not (layer0_outputs(112));
    layer1_outputs(717) <= not(layer0_outputs(2039)) or (layer0_outputs(1057));
    layer1_outputs(718) <= not(layer0_outputs(539));
    layer1_outputs(719) <= '1';
    layer1_outputs(720) <= not(layer0_outputs(2241));
    layer1_outputs(721) <= not((layer0_outputs(999)) and (layer0_outputs(716)));
    layer1_outputs(722) <= (layer0_outputs(1367)) and not (layer0_outputs(2006));
    layer1_outputs(723) <= '0';
    layer1_outputs(724) <= (layer0_outputs(2158)) or (layer0_outputs(2190));
    layer1_outputs(725) <= (layer0_outputs(2547)) and (layer0_outputs(881));
    layer1_outputs(726) <= not(layer0_outputs(835));
    layer1_outputs(727) <= (layer0_outputs(578)) or (layer0_outputs(1419));
    layer1_outputs(728) <= (layer0_outputs(648)) and not (layer0_outputs(987));
    layer1_outputs(729) <= not(layer0_outputs(501)) or (layer0_outputs(186));
    layer1_outputs(730) <= layer0_outputs(2248);
    layer1_outputs(731) <= '1';
    layer1_outputs(732) <= '1';
    layer1_outputs(733) <= '0';
    layer1_outputs(734) <= '0';
    layer1_outputs(735) <= not(layer0_outputs(1725));
    layer1_outputs(736) <= '0';
    layer1_outputs(737) <= layer0_outputs(949);
    layer1_outputs(738) <= '1';
    layer1_outputs(739) <= not(layer0_outputs(1303)) or (layer0_outputs(1216));
    layer1_outputs(740) <= layer0_outputs(598);
    layer1_outputs(741) <= layer0_outputs(2199);
    layer1_outputs(742) <= (layer0_outputs(781)) and not (layer0_outputs(1948));
    layer1_outputs(743) <= (layer0_outputs(369)) and not (layer0_outputs(1674));
    layer1_outputs(744) <= (layer0_outputs(1411)) and not (layer0_outputs(1229));
    layer1_outputs(745) <= not(layer0_outputs(2294));
    layer1_outputs(746) <= (layer0_outputs(1071)) and not (layer0_outputs(1640));
    layer1_outputs(747) <= layer0_outputs(879);
    layer1_outputs(748) <= layer0_outputs(1824);
    layer1_outputs(749) <= not((layer0_outputs(2315)) or (layer0_outputs(1876)));
    layer1_outputs(750) <= not((layer0_outputs(625)) and (layer0_outputs(1233)));
    layer1_outputs(751) <= (layer0_outputs(1198)) and not (layer0_outputs(834));
    layer1_outputs(752) <= layer0_outputs(626);
    layer1_outputs(753) <= (layer0_outputs(1931)) and (layer0_outputs(2532));
    layer1_outputs(754) <= (layer0_outputs(1877)) and not (layer0_outputs(1444));
    layer1_outputs(755) <= not(layer0_outputs(841));
    layer1_outputs(756) <= not((layer0_outputs(2219)) and (layer0_outputs(2537)));
    layer1_outputs(757) <= not((layer0_outputs(136)) and (layer0_outputs(2228)));
    layer1_outputs(758) <= (layer0_outputs(1436)) or (layer0_outputs(182));
    layer1_outputs(759) <= not((layer0_outputs(760)) xor (layer0_outputs(434)));
    layer1_outputs(760) <= layer0_outputs(1828);
    layer1_outputs(761) <= (layer0_outputs(2404)) and (layer0_outputs(2272));
    layer1_outputs(762) <= not(layer0_outputs(1501));
    layer1_outputs(763) <= (layer0_outputs(577)) or (layer0_outputs(1014));
    layer1_outputs(764) <= layer0_outputs(1147);
    layer1_outputs(765) <= '0';
    layer1_outputs(766) <= (layer0_outputs(1159)) and (layer0_outputs(2419));
    layer1_outputs(767) <= not(layer0_outputs(1569));
    layer1_outputs(768) <= not((layer0_outputs(1385)) or (layer0_outputs(1422)));
    layer1_outputs(769) <= (layer0_outputs(165)) and not (layer0_outputs(268));
    layer1_outputs(770) <= '0';
    layer1_outputs(771) <= not((layer0_outputs(783)) and (layer0_outputs(2432)));
    layer1_outputs(772) <= (layer0_outputs(2079)) and not (layer0_outputs(1915));
    layer1_outputs(773) <= not((layer0_outputs(1187)) and (layer0_outputs(2275)));
    layer1_outputs(774) <= (layer0_outputs(1708)) and not (layer0_outputs(1604));
    layer1_outputs(775) <= not((layer0_outputs(1565)) or (layer0_outputs(1382)));
    layer1_outputs(776) <= '1';
    layer1_outputs(777) <= '0';
    layer1_outputs(778) <= layer0_outputs(1393);
    layer1_outputs(779) <= layer0_outputs(1527);
    layer1_outputs(780) <= not((layer0_outputs(1174)) or (layer0_outputs(849)));
    layer1_outputs(781) <= not((layer0_outputs(1800)) and (layer0_outputs(2201)));
    layer1_outputs(782) <= not(layer0_outputs(794)) or (layer0_outputs(2396));
    layer1_outputs(783) <= layer0_outputs(2164);
    layer1_outputs(784) <= layer0_outputs(860);
    layer1_outputs(785) <= layer0_outputs(1821);
    layer1_outputs(786) <= (layer0_outputs(859)) and not (layer0_outputs(1391));
    layer1_outputs(787) <= (layer0_outputs(1905)) or (layer0_outputs(2214));
    layer1_outputs(788) <= not(layer0_outputs(244));
    layer1_outputs(789) <= '1';
    layer1_outputs(790) <= (layer0_outputs(1568)) and not (layer0_outputs(410));
    layer1_outputs(791) <= layer0_outputs(257);
    layer1_outputs(792) <= not((layer0_outputs(1639)) or (layer0_outputs(949)));
    layer1_outputs(793) <= not((layer0_outputs(2108)) or (layer0_outputs(1991)));
    layer1_outputs(794) <= not((layer0_outputs(573)) or (layer0_outputs(1070)));
    layer1_outputs(795) <= (layer0_outputs(810)) and not (layer0_outputs(425));
    layer1_outputs(796) <= not(layer0_outputs(1431)) or (layer0_outputs(1126));
    layer1_outputs(797) <= (layer0_outputs(2343)) and not (layer0_outputs(226));
    layer1_outputs(798) <= '1';
    layer1_outputs(799) <= not(layer0_outputs(348)) or (layer0_outputs(1884));
    layer1_outputs(800) <= '0';
    layer1_outputs(801) <= not((layer0_outputs(806)) or (layer0_outputs(1915)));
    layer1_outputs(802) <= not(layer0_outputs(1566)) or (layer0_outputs(1998));
    layer1_outputs(803) <= not(layer0_outputs(167)) or (layer0_outputs(304));
    layer1_outputs(804) <= not(layer0_outputs(1346));
    layer1_outputs(805) <= (layer0_outputs(353)) and not (layer0_outputs(40));
    layer1_outputs(806) <= not(layer0_outputs(280)) or (layer0_outputs(744));
    layer1_outputs(807) <= '1';
    layer1_outputs(808) <= (layer0_outputs(282)) and (layer0_outputs(211));
    layer1_outputs(809) <= (layer0_outputs(1741)) or (layer0_outputs(1178));
    layer1_outputs(810) <= '1';
    layer1_outputs(811) <= not(layer0_outputs(1436));
    layer1_outputs(812) <= not((layer0_outputs(1278)) and (layer0_outputs(2313)));
    layer1_outputs(813) <= not(layer0_outputs(878)) or (layer0_outputs(2431));
    layer1_outputs(814) <= not((layer0_outputs(972)) or (layer0_outputs(2000)));
    layer1_outputs(815) <= not(layer0_outputs(587)) or (layer0_outputs(1898));
    layer1_outputs(816) <= (layer0_outputs(337)) and not (layer0_outputs(768));
    layer1_outputs(817) <= not(layer0_outputs(1335));
    layer1_outputs(818) <= not(layer0_outputs(327));
    layer1_outputs(819) <= (layer0_outputs(1839)) or (layer0_outputs(2219));
    layer1_outputs(820) <= not((layer0_outputs(699)) and (layer0_outputs(689)));
    layer1_outputs(821) <= not((layer0_outputs(1238)) or (layer0_outputs(1435)));
    layer1_outputs(822) <= not(layer0_outputs(512)) or (layer0_outputs(312));
    layer1_outputs(823) <= not((layer0_outputs(984)) and (layer0_outputs(1377)));
    layer1_outputs(824) <= not(layer0_outputs(2412));
    layer1_outputs(825) <= not(layer0_outputs(1091)) or (layer0_outputs(1364));
    layer1_outputs(826) <= (layer0_outputs(675)) and not (layer0_outputs(1448));
    layer1_outputs(827) <= layer0_outputs(1522);
    layer1_outputs(828) <= (layer0_outputs(190)) or (layer0_outputs(2523));
    layer1_outputs(829) <= not(layer0_outputs(1456));
    layer1_outputs(830) <= not((layer0_outputs(191)) and (layer0_outputs(1201)));
    layer1_outputs(831) <= (layer0_outputs(2386)) and not (layer0_outputs(95));
    layer1_outputs(832) <= (layer0_outputs(2135)) and (layer0_outputs(2541));
    layer1_outputs(833) <= layer0_outputs(1615);
    layer1_outputs(834) <= layer0_outputs(826);
    layer1_outputs(835) <= not((layer0_outputs(1440)) and (layer0_outputs(1801)));
    layer1_outputs(836) <= layer0_outputs(649);
    layer1_outputs(837) <= not(layer0_outputs(1961));
    layer1_outputs(838) <= (layer0_outputs(779)) or (layer0_outputs(2371));
    layer1_outputs(839) <= '1';
    layer1_outputs(840) <= (layer0_outputs(1783)) or (layer0_outputs(2253));
    layer1_outputs(841) <= not(layer0_outputs(1479));
    layer1_outputs(842) <= not(layer0_outputs(334)) or (layer0_outputs(1423));
    layer1_outputs(843) <= '0';
    layer1_outputs(844) <= (layer0_outputs(1035)) or (layer0_outputs(1220));
    layer1_outputs(845) <= layer0_outputs(212);
    layer1_outputs(846) <= not(layer0_outputs(1054));
    layer1_outputs(847) <= (layer0_outputs(1027)) and not (layer0_outputs(1923));
    layer1_outputs(848) <= '0';
    layer1_outputs(849) <= (layer0_outputs(2245)) and not (layer0_outputs(1498));
    layer1_outputs(850) <= '1';
    layer1_outputs(851) <= (layer0_outputs(672)) or (layer0_outputs(1426));
    layer1_outputs(852) <= '1';
    layer1_outputs(853) <= layer0_outputs(1201);
    layer1_outputs(854) <= not((layer0_outputs(823)) and (layer0_outputs(210)));
    layer1_outputs(855) <= not(layer0_outputs(167));
    layer1_outputs(856) <= (layer0_outputs(179)) and (layer0_outputs(455));
    layer1_outputs(857) <= not(layer0_outputs(524));
    layer1_outputs(858) <= not(layer0_outputs(1974)) or (layer0_outputs(2029));
    layer1_outputs(859) <= not((layer0_outputs(1664)) and (layer0_outputs(1713)));
    layer1_outputs(860) <= not((layer0_outputs(1108)) xor (layer0_outputs(424)));
    layer1_outputs(861) <= not(layer0_outputs(2317));
    layer1_outputs(862) <= layer0_outputs(1278);
    layer1_outputs(863) <= (layer0_outputs(1578)) and (layer0_outputs(743));
    layer1_outputs(864) <= layer0_outputs(2442);
    layer1_outputs(865) <= not(layer0_outputs(1280));
    layer1_outputs(866) <= layer0_outputs(784);
    layer1_outputs(867) <= layer0_outputs(2062);
    layer1_outputs(868) <= (layer0_outputs(1040)) and (layer0_outputs(1086));
    layer1_outputs(869) <= layer0_outputs(741);
    layer1_outputs(870) <= not(layer0_outputs(1309));
    layer1_outputs(871) <= not(layer0_outputs(298));
    layer1_outputs(872) <= not((layer0_outputs(1784)) or (layer0_outputs(2357)));
    layer1_outputs(873) <= (layer0_outputs(2)) and not (layer0_outputs(2349));
    layer1_outputs(874) <= layer0_outputs(1567);
    layer1_outputs(875) <= '0';
    layer1_outputs(876) <= not((layer0_outputs(1916)) or (layer0_outputs(1887)));
    layer1_outputs(877) <= not((layer0_outputs(2168)) and (layer0_outputs(671)));
    layer1_outputs(878) <= not(layer0_outputs(528)) or (layer0_outputs(322));
    layer1_outputs(879) <= not((layer0_outputs(1934)) and (layer0_outputs(2030)));
    layer1_outputs(880) <= layer0_outputs(1164);
    layer1_outputs(881) <= not(layer0_outputs(6));
    layer1_outputs(882) <= layer0_outputs(1261);
    layer1_outputs(883) <= (layer0_outputs(1038)) and not (layer0_outputs(2026));
    layer1_outputs(884) <= (layer0_outputs(389)) and (layer0_outputs(10));
    layer1_outputs(885) <= layer0_outputs(1599);
    layer1_outputs(886) <= not((layer0_outputs(2192)) or (layer0_outputs(1778)));
    layer1_outputs(887) <= not(layer0_outputs(2025)) or (layer0_outputs(1929));
    layer1_outputs(888) <= layer0_outputs(909);
    layer1_outputs(889) <= not(layer0_outputs(515)) or (layer0_outputs(484));
    layer1_outputs(890) <= layer0_outputs(459);
    layer1_outputs(891) <= not(layer0_outputs(2232));
    layer1_outputs(892) <= '0';
    layer1_outputs(893) <= not((layer0_outputs(320)) xor (layer0_outputs(579)));
    layer1_outputs(894) <= (layer0_outputs(166)) and not (layer0_outputs(1471));
    layer1_outputs(895) <= layer0_outputs(2553);
    layer1_outputs(896) <= '0';
    layer1_outputs(897) <= layer0_outputs(995);
    layer1_outputs(898) <= (layer0_outputs(1880)) and (layer0_outputs(1721));
    layer1_outputs(899) <= layer0_outputs(359);
    layer1_outputs(900) <= not(layer0_outputs(858)) or (layer0_outputs(2126));
    layer1_outputs(901) <= not(layer0_outputs(1878));
    layer1_outputs(902) <= (layer0_outputs(1238)) and (layer0_outputs(2139));
    layer1_outputs(903) <= (layer0_outputs(2472)) and not (layer0_outputs(933));
    layer1_outputs(904) <= not(layer0_outputs(228));
    layer1_outputs(905) <= (layer0_outputs(2546)) and (layer0_outputs(2047));
    layer1_outputs(906) <= not((layer0_outputs(1211)) or (layer0_outputs(1994)));
    layer1_outputs(907) <= (layer0_outputs(141)) and not (layer0_outputs(946));
    layer1_outputs(908) <= (layer0_outputs(1619)) and not (layer0_outputs(1553));
    layer1_outputs(909) <= (layer0_outputs(1035)) and (layer0_outputs(2202));
    layer1_outputs(910) <= (layer0_outputs(1564)) xor (layer0_outputs(895));
    layer1_outputs(911) <= (layer0_outputs(1111)) or (layer0_outputs(266));
    layer1_outputs(912) <= layer0_outputs(2024);
    layer1_outputs(913) <= not(layer0_outputs(2041)) or (layer0_outputs(650));
    layer1_outputs(914) <= (layer0_outputs(1521)) and not (layer0_outputs(1390));
    layer1_outputs(915) <= not(layer0_outputs(1663));
    layer1_outputs(916) <= not(layer0_outputs(425)) or (layer0_outputs(2155));
    layer1_outputs(917) <= not(layer0_outputs(2404));
    layer1_outputs(918) <= not((layer0_outputs(534)) or (layer0_outputs(2151)));
    layer1_outputs(919) <= '1';
    layer1_outputs(920) <= layer0_outputs(33);
    layer1_outputs(921) <= '1';
    layer1_outputs(922) <= not(layer0_outputs(1274));
    layer1_outputs(923) <= not(layer0_outputs(43));
    layer1_outputs(924) <= not(layer0_outputs(1421));
    layer1_outputs(925) <= not(layer0_outputs(661)) or (layer0_outputs(132));
    layer1_outputs(926) <= layer0_outputs(118);
    layer1_outputs(927) <= (layer0_outputs(293)) and not (layer0_outputs(1813));
    layer1_outputs(928) <= not(layer0_outputs(1936));
    layer1_outputs(929) <= not((layer0_outputs(975)) or (layer0_outputs(1362)));
    layer1_outputs(930) <= not(layer0_outputs(737));
    layer1_outputs(931) <= (layer0_outputs(1670)) and not (layer0_outputs(1671));
    layer1_outputs(932) <= not(layer0_outputs(2439)) or (layer0_outputs(1223));
    layer1_outputs(933) <= not(layer0_outputs(2512));
    layer1_outputs(934) <= '1';
    layer1_outputs(935) <= '1';
    layer1_outputs(936) <= not(layer0_outputs(1809));
    layer1_outputs(937) <= (layer0_outputs(2107)) and (layer0_outputs(2187));
    layer1_outputs(938) <= not(layer0_outputs(195));
    layer1_outputs(939) <= (layer0_outputs(2493)) and not (layer0_outputs(1117));
    layer1_outputs(940) <= (layer0_outputs(905)) or (layer0_outputs(1368));
    layer1_outputs(941) <= (layer0_outputs(1398)) and not (layer0_outputs(1807));
    layer1_outputs(942) <= layer0_outputs(2345);
    layer1_outputs(943) <= not(layer0_outputs(1453));
    layer1_outputs(944) <= layer0_outputs(2102);
    layer1_outputs(945) <= not(layer0_outputs(2249)) or (layer0_outputs(2059));
    layer1_outputs(946) <= not((layer0_outputs(317)) or (layer0_outputs(1845)));
    layer1_outputs(947) <= (layer0_outputs(778)) or (layer0_outputs(1050));
    layer1_outputs(948) <= '0';
    layer1_outputs(949) <= not((layer0_outputs(138)) xor (layer0_outputs(2551)));
    layer1_outputs(950) <= (layer0_outputs(333)) and (layer0_outputs(786));
    layer1_outputs(951) <= '0';
    layer1_outputs(952) <= (layer0_outputs(1844)) or (layer0_outputs(1993));
    layer1_outputs(953) <= layer0_outputs(651);
    layer1_outputs(954) <= not(layer0_outputs(1137));
    layer1_outputs(955) <= '0';
    layer1_outputs(956) <= '0';
    layer1_outputs(957) <= (layer0_outputs(1174)) and not (layer0_outputs(985));
    layer1_outputs(958) <= layer0_outputs(2040);
    layer1_outputs(959) <= not((layer0_outputs(355)) or (layer0_outputs(2530)));
    layer1_outputs(960) <= not((layer0_outputs(1186)) xor (layer0_outputs(1871)));
    layer1_outputs(961) <= not((layer0_outputs(1723)) or (layer0_outputs(2443)));
    layer1_outputs(962) <= layer0_outputs(197);
    layer1_outputs(963) <= (layer0_outputs(1552)) and (layer0_outputs(1528));
    layer1_outputs(964) <= not(layer0_outputs(2526)) or (layer0_outputs(605));
    layer1_outputs(965) <= not(layer0_outputs(2500));
    layer1_outputs(966) <= (layer0_outputs(324)) and not (layer0_outputs(878));
    layer1_outputs(967) <= not((layer0_outputs(1128)) or (layer0_outputs(1551)));
    layer1_outputs(968) <= (layer0_outputs(2028)) and not (layer0_outputs(157));
    layer1_outputs(969) <= not((layer0_outputs(1446)) or (layer0_outputs(148)));
    layer1_outputs(970) <= layer0_outputs(2453);
    layer1_outputs(971) <= layer0_outputs(634);
    layer1_outputs(972) <= '1';
    layer1_outputs(973) <= '0';
    layer1_outputs(974) <= not((layer0_outputs(1552)) or (layer0_outputs(807)));
    layer1_outputs(975) <= layer0_outputs(144);
    layer1_outputs(976) <= (layer0_outputs(2164)) or (layer0_outputs(1455));
    layer1_outputs(977) <= (layer0_outputs(211)) and not (layer0_outputs(1239));
    layer1_outputs(978) <= layer0_outputs(808);
    layer1_outputs(979) <= (layer0_outputs(563)) and not (layer0_outputs(1946));
    layer1_outputs(980) <= '0';
    layer1_outputs(981) <= not(layer0_outputs(2542));
    layer1_outputs(982) <= not(layer0_outputs(688)) or (layer0_outputs(274));
    layer1_outputs(983) <= layer0_outputs(557);
    layer1_outputs(984) <= '0';
    layer1_outputs(985) <= '1';
    layer1_outputs(986) <= not(layer0_outputs(1595)) or (layer0_outputs(600));
    layer1_outputs(987) <= not(layer0_outputs(551)) or (layer0_outputs(24));
    layer1_outputs(988) <= layer0_outputs(637);
    layer1_outputs(989) <= not(layer0_outputs(2449)) or (layer0_outputs(590));
    layer1_outputs(990) <= (layer0_outputs(1318)) or (layer0_outputs(45));
    layer1_outputs(991) <= '0';
    layer1_outputs(992) <= (layer0_outputs(842)) and (layer0_outputs(1458));
    layer1_outputs(993) <= (layer0_outputs(1369)) xor (layer0_outputs(695));
    layer1_outputs(994) <= not(layer0_outputs(2356));
    layer1_outputs(995) <= (layer0_outputs(1543)) or (layer0_outputs(31));
    layer1_outputs(996) <= not((layer0_outputs(514)) or (layer0_outputs(2211)));
    layer1_outputs(997) <= not((layer0_outputs(2338)) or (layer0_outputs(543)));
    layer1_outputs(998) <= not((layer0_outputs(1698)) and (layer0_outputs(944)));
    layer1_outputs(999) <= not(layer0_outputs(452));
    layer1_outputs(1000) <= (layer0_outputs(1509)) and (layer0_outputs(719));
    layer1_outputs(1001) <= not(layer0_outputs(1984));
    layer1_outputs(1002) <= (layer0_outputs(2346)) or (layer0_outputs(776));
    layer1_outputs(1003) <= (layer0_outputs(260)) and (layer0_outputs(943));
    layer1_outputs(1004) <= not(layer0_outputs(119));
    layer1_outputs(1005) <= not(layer0_outputs(358)) or (layer0_outputs(163));
    layer1_outputs(1006) <= layer0_outputs(1077);
    layer1_outputs(1007) <= layer0_outputs(233);
    layer1_outputs(1008) <= not(layer0_outputs(192));
    layer1_outputs(1009) <= '1';
    layer1_outputs(1010) <= '1';
    layer1_outputs(1011) <= (layer0_outputs(2479)) and (layer0_outputs(618));
    layer1_outputs(1012) <= (layer0_outputs(1734)) and not (layer0_outputs(642));
    layer1_outputs(1013) <= layer0_outputs(962);
    layer1_outputs(1014) <= (layer0_outputs(335)) and (layer0_outputs(1571));
    layer1_outputs(1015) <= not((layer0_outputs(440)) and (layer0_outputs(1386)));
    layer1_outputs(1016) <= (layer0_outputs(1886)) and not (layer0_outputs(435));
    layer1_outputs(1017) <= '1';
    layer1_outputs(1018) <= not(layer0_outputs(2487)) or (layer0_outputs(1717));
    layer1_outputs(1019) <= '1';
    layer1_outputs(1020) <= not(layer0_outputs(843));
    layer1_outputs(1021) <= not(layer0_outputs(2115));
    layer1_outputs(1022) <= not(layer0_outputs(919)) or (layer0_outputs(988));
    layer1_outputs(1023) <= '1';
    layer1_outputs(1024) <= '1';
    layer1_outputs(1025) <= (layer0_outputs(2506)) or (layer0_outputs(1944));
    layer1_outputs(1026) <= layer0_outputs(362);
    layer1_outputs(1027) <= layer0_outputs(525);
    layer1_outputs(1028) <= not(layer0_outputs(2538)) or (layer0_outputs(360));
    layer1_outputs(1029) <= not(layer0_outputs(354)) or (layer0_outputs(2256));
    layer1_outputs(1030) <= (layer0_outputs(998)) and not (layer0_outputs(178));
    layer1_outputs(1031) <= not((layer0_outputs(989)) or (layer0_outputs(1180)));
    layer1_outputs(1032) <= layer0_outputs(107);
    layer1_outputs(1033) <= layer0_outputs(1592);
    layer1_outputs(1034) <= '0';
    layer1_outputs(1035) <= not(layer0_outputs(343)) or (layer0_outputs(2141));
    layer1_outputs(1036) <= not((layer0_outputs(556)) and (layer0_outputs(48)));
    layer1_outputs(1037) <= '1';
    layer1_outputs(1038) <= '1';
    layer1_outputs(1039) <= (layer0_outputs(2033)) or (layer0_outputs(1613));
    layer1_outputs(1040) <= (layer0_outputs(492)) or (layer0_outputs(1230));
    layer1_outputs(1041) <= not((layer0_outputs(1173)) or (layer0_outputs(1064)));
    layer1_outputs(1042) <= not((layer0_outputs(1105)) and (layer0_outputs(1019)));
    layer1_outputs(1043) <= (layer0_outputs(721)) and not (layer0_outputs(847));
    layer1_outputs(1044) <= not(layer0_outputs(584)) or (layer0_outputs(837));
    layer1_outputs(1045) <= not((layer0_outputs(1410)) or (layer0_outputs(1182)));
    layer1_outputs(1046) <= not(layer0_outputs(459)) or (layer0_outputs(567));
    layer1_outputs(1047) <= (layer0_outputs(1485)) and not (layer0_outputs(2044));
    layer1_outputs(1048) <= (layer0_outputs(188)) and not (layer0_outputs(2441));
    layer1_outputs(1049) <= (layer0_outputs(2106)) and (layer0_outputs(749));
    layer1_outputs(1050) <= (layer0_outputs(1217)) and not (layer0_outputs(2141));
    layer1_outputs(1051) <= not(layer0_outputs(311));
    layer1_outputs(1052) <= '1';
    layer1_outputs(1053) <= not((layer0_outputs(1701)) and (layer0_outputs(198)));
    layer1_outputs(1054) <= '1';
    layer1_outputs(1055) <= (layer0_outputs(666)) and not (layer0_outputs(2521));
    layer1_outputs(1056) <= layer0_outputs(595);
    layer1_outputs(1057) <= not(layer0_outputs(2435)) or (layer0_outputs(910));
    layer1_outputs(1058) <= '0';
    layer1_outputs(1059) <= (layer0_outputs(1626)) and (layer0_outputs(175));
    layer1_outputs(1060) <= (layer0_outputs(1802)) and not (layer0_outputs(244));
    layer1_outputs(1061) <= not(layer0_outputs(340));
    layer1_outputs(1062) <= not(layer0_outputs(393)) or (layer0_outputs(109));
    layer1_outputs(1063) <= (layer0_outputs(1083)) and not (layer0_outputs(814));
    layer1_outputs(1064) <= '0';
    layer1_outputs(1065) <= layer0_outputs(2322);
    layer1_outputs(1066) <= not((layer0_outputs(549)) and (layer0_outputs(1033)));
    layer1_outputs(1067) <= '0';
    layer1_outputs(1068) <= not((layer0_outputs(1020)) xor (layer0_outputs(2529)));
    layer1_outputs(1069) <= not(layer0_outputs(592)) or (layer0_outputs(2172));
    layer1_outputs(1070) <= '1';
    layer1_outputs(1071) <= layer0_outputs(731);
    layer1_outputs(1072) <= (layer0_outputs(1806)) xor (layer0_outputs(75));
    layer1_outputs(1073) <= '1';
    layer1_outputs(1074) <= layer0_outputs(1091);
    layer1_outputs(1075) <= not(layer0_outputs(1242)) or (layer0_outputs(50));
    layer1_outputs(1076) <= not((layer0_outputs(1199)) or (layer0_outputs(2157)));
    layer1_outputs(1077) <= (layer0_outputs(235)) and not (layer0_outputs(2440));
    layer1_outputs(1078) <= '1';
    layer1_outputs(1079) <= not(layer0_outputs(728));
    layer1_outputs(1080) <= '0';
    layer1_outputs(1081) <= layer0_outputs(203);
    layer1_outputs(1082) <= not(layer0_outputs(99));
    layer1_outputs(1083) <= not(layer0_outputs(1980));
    layer1_outputs(1084) <= (layer0_outputs(1184)) or (layer0_outputs(1540));
    layer1_outputs(1085) <= (layer0_outputs(382)) and not (layer0_outputs(1478));
    layer1_outputs(1086) <= not(layer0_outputs(1814));
    layer1_outputs(1087) <= (layer0_outputs(1408)) and (layer0_outputs(1506));
    layer1_outputs(1088) <= not(layer0_outputs(895));
    layer1_outputs(1089) <= not(layer0_outputs(2266));
    layer1_outputs(1090) <= '0';
    layer1_outputs(1091) <= not(layer0_outputs(195));
    layer1_outputs(1092) <= (layer0_outputs(423)) and not (layer0_outputs(2373));
    layer1_outputs(1093) <= (layer0_outputs(2513)) or (layer0_outputs(2257));
    layer1_outputs(1094) <= not((layer0_outputs(393)) and (layer0_outputs(321)));
    layer1_outputs(1095) <= not((layer0_outputs(1811)) or (layer0_outputs(917)));
    layer1_outputs(1096) <= not(layer0_outputs(241)) or (layer0_outputs(2159));
    layer1_outputs(1097) <= layer0_outputs(1917);
    layer1_outputs(1098) <= (layer0_outputs(1336)) and not (layer0_outputs(65));
    layer1_outputs(1099) <= layer0_outputs(232);
    layer1_outputs(1100) <= layer0_outputs(681);
    layer1_outputs(1101) <= not(layer0_outputs(752)) or (layer0_outputs(682));
    layer1_outputs(1102) <= layer0_outputs(683);
    layer1_outputs(1103) <= '1';
    layer1_outputs(1104) <= not((layer0_outputs(2432)) or (layer0_outputs(2162)));
    layer1_outputs(1105) <= not((layer0_outputs(544)) or (layer0_outputs(2303)));
    layer1_outputs(1106) <= not((layer0_outputs(156)) or (layer0_outputs(313)));
    layer1_outputs(1107) <= not(layer0_outputs(1594));
    layer1_outputs(1108) <= (layer0_outputs(620)) and not (layer0_outputs(596));
    layer1_outputs(1109) <= (layer0_outputs(1364)) and (layer0_outputs(0));
    layer1_outputs(1110) <= not(layer0_outputs(594));
    layer1_outputs(1111) <= '1';
    layer1_outputs(1112) <= (layer0_outputs(1936)) and not (layer0_outputs(129));
    layer1_outputs(1113) <= not((layer0_outputs(1417)) or (layer0_outputs(933)));
    layer1_outputs(1114) <= layer0_outputs(1985);
    layer1_outputs(1115) <= not(layer0_outputs(2125));
    layer1_outputs(1116) <= not(layer0_outputs(1482)) or (layer0_outputs(633));
    layer1_outputs(1117) <= not(layer0_outputs(2254));
    layer1_outputs(1118) <= not((layer0_outputs(539)) and (layer0_outputs(2237)));
    layer1_outputs(1119) <= '0';
    layer1_outputs(1120) <= not(layer0_outputs(2462));
    layer1_outputs(1121) <= not(layer0_outputs(1145));
    layer1_outputs(1122) <= layer0_outputs(2177);
    layer1_outputs(1123) <= not(layer0_outputs(1823)) or (layer0_outputs(1670));
    layer1_outputs(1124) <= layer0_outputs(954);
    layer1_outputs(1125) <= not(layer0_outputs(1486));
    layer1_outputs(1126) <= not(layer0_outputs(702));
    layer1_outputs(1127) <= not(layer0_outputs(2487)) or (layer0_outputs(1745));
    layer1_outputs(1128) <= not((layer0_outputs(1824)) or (layer0_outputs(1076)));
    layer1_outputs(1129) <= not(layer0_outputs(968));
    layer1_outputs(1130) <= not(layer0_outputs(81)) or (layer0_outputs(904));
    layer1_outputs(1131) <= not(layer0_outputs(1096)) or (layer0_outputs(1917));
    layer1_outputs(1132) <= layer0_outputs(174);
    layer1_outputs(1133) <= layer0_outputs(901);
    layer1_outputs(1134) <= (layer0_outputs(966)) or (layer0_outputs(230));
    layer1_outputs(1135) <= not(layer0_outputs(2208)) or (layer0_outputs(1243));
    layer1_outputs(1136) <= not(layer0_outputs(2375));
    layer1_outputs(1137) <= (layer0_outputs(6)) and not (layer0_outputs(36));
    layer1_outputs(1138) <= (layer0_outputs(61)) or (layer0_outputs(799));
    layer1_outputs(1139) <= (layer0_outputs(1234)) or (layer0_outputs(2024));
    layer1_outputs(1140) <= layer0_outputs(2548);
    layer1_outputs(1141) <= (layer0_outputs(2092)) or (layer0_outputs(716));
    layer1_outputs(1142) <= not(layer0_outputs(2342));
    layer1_outputs(1143) <= layer0_outputs(960);
    layer1_outputs(1144) <= (layer0_outputs(1257)) and (layer0_outputs(1850));
    layer1_outputs(1145) <= '0';
    layer1_outputs(1146) <= layer0_outputs(68);
    layer1_outputs(1147) <= (layer0_outputs(36)) and not (layer0_outputs(2507));
    layer1_outputs(1148) <= not(layer0_outputs(220));
    layer1_outputs(1149) <= not(layer0_outputs(90)) or (layer0_outputs(2173));
    layer1_outputs(1150) <= (layer0_outputs(953)) and not (layer0_outputs(533));
    layer1_outputs(1151) <= '1';
    layer1_outputs(1152) <= not(layer0_outputs(1842));
    layer1_outputs(1153) <= not(layer0_outputs(293));
    layer1_outputs(1154) <= not(layer0_outputs(665));
    layer1_outputs(1155) <= (layer0_outputs(747)) and not (layer0_outputs(888));
    layer1_outputs(1156) <= (layer0_outputs(1138)) and (layer0_outputs(1731));
    layer1_outputs(1157) <= not(layer0_outputs(1873)) or (layer0_outputs(2009));
    layer1_outputs(1158) <= not(layer0_outputs(1136)) or (layer0_outputs(1425));
    layer1_outputs(1159) <= layer0_outputs(1535);
    layer1_outputs(1160) <= not(layer0_outputs(1541)) or (layer0_outputs(1774));
    layer1_outputs(1161) <= not(layer0_outputs(419)) or (layer0_outputs(1203));
    layer1_outputs(1162) <= not(layer0_outputs(1867)) or (layer0_outputs(1807));
    layer1_outputs(1163) <= not((layer0_outputs(152)) or (layer0_outputs(739)));
    layer1_outputs(1164) <= '0';
    layer1_outputs(1165) <= not(layer0_outputs(1644));
    layer1_outputs(1166) <= '0';
    layer1_outputs(1167) <= not(layer0_outputs(1258));
    layer1_outputs(1168) <= not(layer0_outputs(1260)) or (layer0_outputs(1859));
    layer1_outputs(1169) <= not(layer0_outputs(2434)) or (layer0_outputs(1154));
    layer1_outputs(1170) <= (layer0_outputs(458)) and (layer0_outputs(890));
    layer1_outputs(1171) <= not(layer0_outputs(2253)) or (layer0_outputs(249));
    layer1_outputs(1172) <= not((layer0_outputs(2021)) xor (layer0_outputs(2312)));
    layer1_outputs(1173) <= layer0_outputs(874);
    layer1_outputs(1174) <= '0';
    layer1_outputs(1175) <= layer0_outputs(963);
    layer1_outputs(1176) <= not(layer0_outputs(2558));
    layer1_outputs(1177) <= not(layer0_outputs(1865));
    layer1_outputs(1178) <= not(layer0_outputs(79));
    layer1_outputs(1179) <= not(layer0_outputs(2222));
    layer1_outputs(1180) <= not(layer0_outputs(102));
    layer1_outputs(1181) <= not((layer0_outputs(530)) and (layer0_outputs(1438)));
    layer1_outputs(1182) <= not(layer0_outputs(1590));
    layer1_outputs(1183) <= '0';
    layer1_outputs(1184) <= not((layer0_outputs(2271)) and (layer0_outputs(1462)));
    layer1_outputs(1185) <= layer0_outputs(34);
    layer1_outputs(1186) <= not((layer0_outputs(273)) or (layer0_outputs(937)));
    layer1_outputs(1187) <= layer0_outputs(1012);
    layer1_outputs(1188) <= not(layer0_outputs(1445));
    layer1_outputs(1189) <= (layer0_outputs(251)) or (layer0_outputs(2126));
    layer1_outputs(1190) <= not((layer0_outputs(1700)) or (layer0_outputs(2394)));
    layer1_outputs(1191) <= not(layer0_outputs(993)) or (layer0_outputs(238));
    layer1_outputs(1192) <= not(layer0_outputs(1879));
    layer1_outputs(1193) <= layer0_outputs(2267);
    layer1_outputs(1194) <= (layer0_outputs(265)) and (layer0_outputs(2177));
    layer1_outputs(1195) <= layer0_outputs(1315);
    layer1_outputs(1196) <= '0';
    layer1_outputs(1197) <= not(layer0_outputs(2489)) or (layer0_outputs(709));
    layer1_outputs(1198) <= not(layer0_outputs(468));
    layer1_outputs(1199) <= not(layer0_outputs(1087)) or (layer0_outputs(1542));
    layer1_outputs(1200) <= '1';
    layer1_outputs(1201) <= (layer0_outputs(1590)) and not (layer0_outputs(1297));
    layer1_outputs(1202) <= (layer0_outputs(37)) and (layer0_outputs(1754));
    layer1_outputs(1203) <= layer0_outputs(402);
    layer1_outputs(1204) <= layer0_outputs(961);
    layer1_outputs(1205) <= not(layer0_outputs(1191)) or (layer0_outputs(845));
    layer1_outputs(1206) <= not(layer0_outputs(477)) or (layer0_outputs(1143));
    layer1_outputs(1207) <= '1';
    layer1_outputs(1208) <= '1';
    layer1_outputs(1209) <= layer0_outputs(536);
    layer1_outputs(1210) <= layer0_outputs(1912);
    layer1_outputs(1211) <= (layer0_outputs(839)) and not (layer0_outputs(1797));
    layer1_outputs(1212) <= not((layer0_outputs(1010)) and (layer0_outputs(1755)));
    layer1_outputs(1213) <= '0';
    layer1_outputs(1214) <= not(layer0_outputs(499));
    layer1_outputs(1215) <= layer0_outputs(2194);
    layer1_outputs(1216) <= not(layer0_outputs(1666));
    layer1_outputs(1217) <= layer0_outputs(2478);
    layer1_outputs(1218) <= not((layer0_outputs(469)) or (layer0_outputs(1903)));
    layer1_outputs(1219) <= '0';
    layer1_outputs(1220) <= not((layer0_outputs(409)) or (layer0_outputs(2142)));
    layer1_outputs(1221) <= (layer0_outputs(332)) and not (layer0_outputs(1565));
    layer1_outputs(1222) <= layer0_outputs(125);
    layer1_outputs(1223) <= layer0_outputs(612);
    layer1_outputs(1224) <= not(layer0_outputs(1281));
    layer1_outputs(1225) <= not((layer0_outputs(2057)) or (layer0_outputs(386)));
    layer1_outputs(1226) <= not((layer0_outputs(1957)) and (layer0_outputs(1495)));
    layer1_outputs(1227) <= layer0_outputs(965);
    layer1_outputs(1228) <= not(layer0_outputs(516)) or (layer0_outputs(731));
    layer1_outputs(1229) <= (layer0_outputs(2442)) and not (layer0_outputs(722));
    layer1_outputs(1230) <= layer0_outputs(1351);
    layer1_outputs(1231) <= not(layer0_outputs(1482));
    layer1_outputs(1232) <= not((layer0_outputs(2067)) and (layer0_outputs(401)));
    layer1_outputs(1233) <= not(layer0_outputs(205));
    layer1_outputs(1234) <= (layer0_outputs(291)) xor (layer0_outputs(1722));
    layer1_outputs(1235) <= not((layer0_outputs(768)) and (layer0_outputs(816)));
    layer1_outputs(1236) <= (layer0_outputs(656)) and (layer0_outputs(1498));
    layer1_outputs(1237) <= not(layer0_outputs(1603)) or (layer0_outputs(2329));
    layer1_outputs(1238) <= not((layer0_outputs(566)) and (layer0_outputs(216)));
    layer1_outputs(1239) <= layer0_outputs(1403);
    layer1_outputs(1240) <= not((layer0_outputs(732)) and (layer0_outputs(112)));
    layer1_outputs(1241) <= (layer0_outputs(1058)) and (layer0_outputs(2327));
    layer1_outputs(1242) <= not(layer0_outputs(1907));
    layer1_outputs(1243) <= (layer0_outputs(1881)) and not (layer0_outputs(1560));
    layer1_outputs(1244) <= not(layer0_outputs(690));
    layer1_outputs(1245) <= not(layer0_outputs(1627)) or (layer0_outputs(718));
    layer1_outputs(1246) <= '1';
    layer1_outputs(1247) <= not(layer0_outputs(1432));
    layer1_outputs(1248) <= (layer0_outputs(1159)) and (layer0_outputs(2511));
    layer1_outputs(1249) <= '0';
    layer1_outputs(1250) <= not(layer0_outputs(1872)) or (layer0_outputs(57));
    layer1_outputs(1251) <= layer0_outputs(2002);
    layer1_outputs(1252) <= layer0_outputs(2022);
    layer1_outputs(1253) <= not(layer0_outputs(466)) or (layer0_outputs(1669));
    layer1_outputs(1254) <= '1';
    layer1_outputs(1255) <= not((layer0_outputs(2055)) and (layer0_outputs(1949)));
    layer1_outputs(1256) <= layer0_outputs(2189);
    layer1_outputs(1257) <= not((layer0_outputs(1146)) and (layer0_outputs(1834)));
    layer1_outputs(1258) <= not(layer0_outputs(2351));
    layer1_outputs(1259) <= layer0_outputs(2322);
    layer1_outputs(1260) <= not((layer0_outputs(227)) or (layer0_outputs(1338)));
    layer1_outputs(1261) <= '1';
    layer1_outputs(1262) <= '0';
    layer1_outputs(1263) <= '1';
    layer1_outputs(1264) <= (layer0_outputs(771)) or (layer0_outputs(1025));
    layer1_outputs(1265) <= layer0_outputs(889);
    layer1_outputs(1266) <= layer0_outputs(398);
    layer1_outputs(1267) <= not(layer0_outputs(1009)) or (layer0_outputs(1982));
    layer1_outputs(1268) <= layer0_outputs(2517);
    layer1_outputs(1269) <= (layer0_outputs(891)) and not (layer0_outputs(717));
    layer1_outputs(1270) <= not((layer0_outputs(1770)) and (layer0_outputs(698)));
    layer1_outputs(1271) <= layer0_outputs(2187);
    layer1_outputs(1272) <= not((layer0_outputs(1935)) and (layer0_outputs(2504)));
    layer1_outputs(1273) <= not(layer0_outputs(344));
    layer1_outputs(1274) <= not((layer0_outputs(2023)) and (layer0_outputs(1949)));
    layer1_outputs(1275) <= (layer0_outputs(820)) and not (layer0_outputs(1725));
    layer1_outputs(1276) <= not(layer0_outputs(1847));
    layer1_outputs(1277) <= (layer0_outputs(533)) or (layer0_outputs(2369));
    layer1_outputs(1278) <= not((layer0_outputs(1925)) or (layer0_outputs(589)));
    layer1_outputs(1279) <= (layer0_outputs(1106)) and (layer0_outputs(521));
    layer1_outputs(1280) <= layer0_outputs(1399);
    layer1_outputs(1281) <= not((layer0_outputs(684)) or (layer0_outputs(1591)));
    layer1_outputs(1282) <= not(layer0_outputs(206)) or (layer0_outputs(2087));
    layer1_outputs(1283) <= layer0_outputs(1209);
    layer1_outputs(1284) <= not(layer0_outputs(336));
    layer1_outputs(1285) <= (layer0_outputs(1013)) and not (layer0_outputs(2070));
    layer1_outputs(1286) <= (layer0_outputs(432)) and not (layer0_outputs(1019));
    layer1_outputs(1287) <= (layer0_outputs(1962)) and not (layer0_outputs(1452));
    layer1_outputs(1288) <= not((layer0_outputs(2297)) and (layer0_outputs(2031)));
    layer1_outputs(1289) <= (layer0_outputs(1973)) and not (layer0_outputs(2321));
    layer1_outputs(1290) <= (layer0_outputs(1093)) and not (layer0_outputs(142));
    layer1_outputs(1291) <= not(layer0_outputs(861)) or (layer0_outputs(1457));
    layer1_outputs(1292) <= not((layer0_outputs(2017)) and (layer0_outputs(1067)));
    layer1_outputs(1293) <= '1';
    layer1_outputs(1294) <= '0';
    layer1_outputs(1295) <= not((layer0_outputs(715)) and (layer0_outputs(2145)));
    layer1_outputs(1296) <= not(layer0_outputs(2122)) or (layer0_outputs(1001));
    layer1_outputs(1297) <= '1';
    layer1_outputs(1298) <= (layer0_outputs(1434)) and not (layer0_outputs(46));
    layer1_outputs(1299) <= (layer0_outputs(409)) and not (layer0_outputs(745));
    layer1_outputs(1300) <= layer0_outputs(150);
    layer1_outputs(1301) <= not((layer0_outputs(127)) and (layer0_outputs(1977)));
    layer1_outputs(1302) <= layer0_outputs(970);
    layer1_outputs(1303) <= not((layer0_outputs(1466)) or (layer0_outputs(1818)));
    layer1_outputs(1304) <= '0';
    layer1_outputs(1305) <= not(layer0_outputs(1361)) or (layer0_outputs(2326));
    layer1_outputs(1306) <= not((layer0_outputs(1075)) and (layer0_outputs(1820)));
    layer1_outputs(1307) <= not(layer0_outputs(511));
    layer1_outputs(1308) <= '0';
    layer1_outputs(1309) <= (layer0_outputs(1269)) xor (layer0_outputs(2464));
    layer1_outputs(1310) <= '1';
    layer1_outputs(1311) <= '0';
    layer1_outputs(1312) <= (layer0_outputs(1808)) or (layer0_outputs(599));
    layer1_outputs(1313) <= not(layer0_outputs(795));
    layer1_outputs(1314) <= layer0_outputs(1690);
    layer1_outputs(1315) <= (layer0_outputs(657)) or (layer0_outputs(603));
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= '1';
    layer1_outputs(1318) <= not(layer0_outputs(952));
    layer1_outputs(1319) <= (layer0_outputs(1304)) and not (layer0_outputs(1481));
    layer1_outputs(1320) <= '1';
    layer1_outputs(1321) <= not(layer0_outputs(1857));
    layer1_outputs(1322) <= not(layer0_outputs(1651));
    layer1_outputs(1323) <= '1';
    layer1_outputs(1324) <= not((layer0_outputs(421)) or (layer0_outputs(2433)));
    layer1_outputs(1325) <= (layer0_outputs(602)) and not (layer0_outputs(221));
    layer1_outputs(1326) <= layer0_outputs(1938);
    layer1_outputs(1327) <= (layer0_outputs(1972)) and (layer0_outputs(2293));
    layer1_outputs(1328) <= layer0_outputs(840);
    layer1_outputs(1329) <= layer0_outputs(824);
    layer1_outputs(1330) <= not(layer0_outputs(1945)) or (layer0_outputs(2211));
    layer1_outputs(1331) <= not(layer0_outputs(302)) or (layer0_outputs(2185));
    layer1_outputs(1332) <= layer0_outputs(2319);
    layer1_outputs(1333) <= layer0_outputs(1449);
    layer1_outputs(1334) <= (layer0_outputs(1664)) xor (layer0_outputs(279));
    layer1_outputs(1335) <= (layer0_outputs(2555)) or (layer0_outputs(1240));
    layer1_outputs(1336) <= (layer0_outputs(1210)) or (layer0_outputs(292));
    layer1_outputs(1337) <= not(layer0_outputs(1396));
    layer1_outputs(1338) <= '0';
    layer1_outputs(1339) <= not(layer0_outputs(77)) or (layer0_outputs(463));
    layer1_outputs(1340) <= '0';
    layer1_outputs(1341) <= (layer0_outputs(1751)) and (layer0_outputs(1781));
    layer1_outputs(1342) <= (layer0_outputs(1882)) or (layer0_outputs(1329));
    layer1_outputs(1343) <= not(layer0_outputs(827));
    layer1_outputs(1344) <= (layer0_outputs(2176)) xor (layer0_outputs(2408));
    layer1_outputs(1345) <= '1';
    layer1_outputs(1346) <= not(layer0_outputs(2519));
    layer1_outputs(1347) <= layer0_outputs(2406);
    layer1_outputs(1348) <= layer0_outputs(602);
    layer1_outputs(1349) <= not((layer0_outputs(935)) and (layer0_outputs(2130)));
    layer1_outputs(1350) <= not((layer0_outputs(915)) or (layer0_outputs(642)));
    layer1_outputs(1351) <= layer0_outputs(375);
    layer1_outputs(1352) <= not(layer0_outputs(2505));
    layer1_outputs(1353) <= not(layer0_outputs(325)) or (layer0_outputs(1852));
    layer1_outputs(1354) <= layer0_outputs(1873);
    layer1_outputs(1355) <= '1';
    layer1_outputs(1356) <= layer0_outputs(1953);
    layer1_outputs(1357) <= (layer0_outputs(1964)) and not (layer0_outputs(1723));
    layer1_outputs(1358) <= not(layer0_outputs(1152)) or (layer0_outputs(356));
    layer1_outputs(1359) <= not((layer0_outputs(13)) and (layer0_outputs(2508)));
    layer1_outputs(1360) <= layer0_outputs(264);
    layer1_outputs(1361) <= (layer0_outputs(1386)) xor (layer0_outputs(1679));
    layer1_outputs(1362) <= layer0_outputs(597);
    layer1_outputs(1363) <= not(layer0_outputs(856));
    layer1_outputs(1364) <= layer0_outputs(176);
    layer1_outputs(1365) <= not((layer0_outputs(1053)) and (layer0_outputs(898)));
    layer1_outputs(1366) <= '0';
    layer1_outputs(1367) <= (layer0_outputs(2515)) and not (layer0_outputs(1514));
    layer1_outputs(1368) <= layer0_outputs(2445);
    layer1_outputs(1369) <= not((layer0_outputs(1398)) and (layer0_outputs(520)));
    layer1_outputs(1370) <= layer0_outputs(549);
    layer1_outputs(1371) <= layer0_outputs(2491);
    layer1_outputs(1372) <= '0';
    layer1_outputs(1373) <= (layer0_outputs(2191)) and (layer0_outputs(12));
    layer1_outputs(1374) <= (layer0_outputs(2352)) and (layer0_outputs(1530));
    layer1_outputs(1375) <= '1';
    layer1_outputs(1376) <= not((layer0_outputs(838)) or (layer0_outputs(352)));
    layer1_outputs(1377) <= (layer0_outputs(2523)) and not (layer0_outputs(59));
    layer1_outputs(1378) <= layer0_outputs(1488);
    layer1_outputs(1379) <= (layer0_outputs(162)) xor (layer0_outputs(192));
    layer1_outputs(1380) <= not(layer0_outputs(2471));
    layer1_outputs(1381) <= not(layer0_outputs(57));
    layer1_outputs(1382) <= not(layer0_outputs(1785));
    layer1_outputs(1383) <= not((layer0_outputs(1105)) and (layer0_outputs(2455)));
    layer1_outputs(1384) <= not(layer0_outputs(863));
    layer1_outputs(1385) <= not(layer0_outputs(1065));
    layer1_outputs(1386) <= layer0_outputs(187);
    layer1_outputs(1387) <= not(layer0_outputs(1692)) or (layer0_outputs(449));
    layer1_outputs(1388) <= (layer0_outputs(1231)) and (layer0_outputs(361));
    layer1_outputs(1389) <= '1';
    layer1_outputs(1390) <= (layer0_outputs(1976)) and not (layer0_outputs(921));
    layer1_outputs(1391) <= not((layer0_outputs(2203)) and (layer0_outputs(806)));
    layer1_outputs(1392) <= (layer0_outputs(1196)) and (layer0_outputs(2356));
    layer1_outputs(1393) <= (layer0_outputs(2476)) and (layer0_outputs(1077));
    layer1_outputs(1394) <= '0';
    layer1_outputs(1395) <= not(layer0_outputs(2143));
    layer1_outputs(1396) <= '0';
    layer1_outputs(1397) <= layer0_outputs(1526);
    layer1_outputs(1398) <= layer0_outputs(1179);
    layer1_outputs(1399) <= '0';
    layer1_outputs(1400) <= not((layer0_outputs(884)) and (layer0_outputs(1040)));
    layer1_outputs(1401) <= '0';
    layer1_outputs(1402) <= not((layer0_outputs(1910)) or (layer0_outputs(2559)));
    layer1_outputs(1403) <= '1';
    layer1_outputs(1404) <= not((layer0_outputs(2238)) or (layer0_outputs(683)));
    layer1_outputs(1405) <= (layer0_outputs(1111)) and not (layer0_outputs(863));
    layer1_outputs(1406) <= layer0_outputs(2184);
    layer1_outputs(1407) <= layer0_outputs(85);
    layer1_outputs(1408) <= not(layer0_outputs(83));
    layer1_outputs(1409) <= (layer0_outputs(1647)) and (layer0_outputs(2096));
    layer1_outputs(1410) <= not(layer0_outputs(1614));
    layer1_outputs(1411) <= not(layer0_outputs(503)) or (layer0_outputs(2186));
    layer1_outputs(1412) <= (layer0_outputs(1696)) and (layer0_outputs(1682));
    layer1_outputs(1413) <= not(layer0_outputs(2189));
    layer1_outputs(1414) <= layer0_outputs(783);
    layer1_outputs(1415) <= not(layer0_outputs(78));
    layer1_outputs(1416) <= not(layer0_outputs(826)) or (layer0_outputs(2410));
    layer1_outputs(1417) <= (layer0_outputs(1453)) and (layer0_outputs(1199));
    layer1_outputs(1418) <= (layer0_outputs(673)) and not (layer0_outputs(88));
    layer1_outputs(1419) <= (layer0_outputs(2528)) and (layer0_outputs(2065));
    layer1_outputs(1420) <= not(layer0_outputs(2149));
    layer1_outputs(1421) <= not(layer0_outputs(1063));
    layer1_outputs(1422) <= (layer0_outputs(2463)) and not (layer0_outputs(130));
    layer1_outputs(1423) <= (layer0_outputs(450)) and not (layer0_outputs(41));
    layer1_outputs(1424) <= (layer0_outputs(2165)) and not (layer0_outputs(1272));
    layer1_outputs(1425) <= not(layer0_outputs(241));
    layer1_outputs(1426) <= layer0_outputs(1129);
    layer1_outputs(1427) <= not((layer0_outputs(1969)) or (layer0_outputs(2368)));
    layer1_outputs(1428) <= '1';
    layer1_outputs(1429) <= not((layer0_outputs(199)) or (layer0_outputs(941)));
    layer1_outputs(1430) <= (layer0_outputs(1237)) and (layer0_outputs(811));
    layer1_outputs(1431) <= layer0_outputs(2071);
    layer1_outputs(1432) <= (layer0_outputs(452)) and (layer0_outputs(311));
    layer1_outputs(1433) <= layer0_outputs(787);
    layer1_outputs(1434) <= (layer0_outputs(1173)) and not (layer0_outputs(34));
    layer1_outputs(1435) <= (layer0_outputs(1121)) or (layer0_outputs(800));
    layer1_outputs(1436) <= (layer0_outputs(439)) or (layer0_outputs(2205));
    layer1_outputs(1437) <= not(layer0_outputs(638)) or (layer0_outputs(1594));
    layer1_outputs(1438) <= not(layer0_outputs(2206));
    layer1_outputs(1439) <= not(layer0_outputs(560));
    layer1_outputs(1440) <= layer0_outputs(844);
    layer1_outputs(1441) <= '0';
    layer1_outputs(1442) <= not(layer0_outputs(653)) or (layer0_outputs(131));
    layer1_outputs(1443) <= not(layer0_outputs(2098));
    layer1_outputs(1444) <= not(layer0_outputs(1275)) or (layer0_outputs(1418));
    layer1_outputs(1445) <= layer0_outputs(511);
    layer1_outputs(1446) <= (layer0_outputs(1524)) or (layer0_outputs(1176));
    layer1_outputs(1447) <= not(layer0_outputs(1013));
    layer1_outputs(1448) <= layer0_outputs(672);
    layer1_outputs(1449) <= (layer0_outputs(1024)) and not (layer0_outputs(2550));
    layer1_outputs(1450) <= '0';
    layer1_outputs(1451) <= (layer0_outputs(1480)) and (layer0_outputs(2217));
    layer1_outputs(1452) <= not((layer0_outputs(2326)) and (layer0_outputs(1624)));
    layer1_outputs(1453) <= not(layer0_outputs(445));
    layer1_outputs(1454) <= (layer0_outputs(896)) and (layer0_outputs(76));
    layer1_outputs(1455) <= not((layer0_outputs(939)) and (layer0_outputs(442)));
    layer1_outputs(1456) <= '1';
    layer1_outputs(1457) <= layer0_outputs(1652);
    layer1_outputs(1458) <= layer0_outputs(2005);
    layer1_outputs(1459) <= layer0_outputs(2295);
    layer1_outputs(1460) <= '0';
    layer1_outputs(1461) <= not(layer0_outputs(1771));
    layer1_outputs(1462) <= not(layer0_outputs(1401)) or (layer0_outputs(1732));
    layer1_outputs(1463) <= not(layer0_outputs(1153)) or (layer0_outputs(133));
    layer1_outputs(1464) <= (layer0_outputs(1361)) and (layer0_outputs(729));
    layer1_outputs(1465) <= layer0_outputs(790);
    layer1_outputs(1466) <= not((layer0_outputs(1883)) or (layer0_outputs(882)));
    layer1_outputs(1467) <= not(layer0_outputs(373));
    layer1_outputs(1468) <= layer0_outputs(1101);
    layer1_outputs(1469) <= layer0_outputs(1404);
    layer1_outputs(1470) <= '1';
    layer1_outputs(1471) <= not(layer0_outputs(807));
    layer1_outputs(1472) <= layer0_outputs(32);
    layer1_outputs(1473) <= not(layer0_outputs(2444)) or (layer0_outputs(599));
    layer1_outputs(1474) <= not(layer0_outputs(829));
    layer1_outputs(1475) <= layer0_outputs(1691);
    layer1_outputs(1476) <= (layer0_outputs(853)) and not (layer0_outputs(1463));
    layer1_outputs(1477) <= layer0_outputs(2119);
    layer1_outputs(1478) <= not((layer0_outputs(1962)) or (layer0_outputs(747)));
    layer1_outputs(1479) <= not(layer0_outputs(1638));
    layer1_outputs(1480) <= not(layer0_outputs(631));
    layer1_outputs(1481) <= not((layer0_outputs(1376)) or (layer0_outputs(784)));
    layer1_outputs(1482) <= not(layer0_outputs(2398));
    layer1_outputs(1483) <= not(layer0_outputs(2034));
    layer1_outputs(1484) <= not(layer0_outputs(2414));
    layer1_outputs(1485) <= layer0_outputs(149);
    layer1_outputs(1486) <= (layer0_outputs(445)) and not (layer0_outputs(364));
    layer1_outputs(1487) <= not((layer0_outputs(2140)) xor (layer0_outputs(1766)));
    layer1_outputs(1488) <= '1';
    layer1_outputs(1489) <= '1';
    layer1_outputs(1490) <= not(layer0_outputs(1575)) or (layer0_outputs(529));
    layer1_outputs(1491) <= '1';
    layer1_outputs(1492) <= (layer0_outputs(973)) and not (layer0_outputs(553));
    layer1_outputs(1493) <= (layer0_outputs(1358)) and not (layer0_outputs(87));
    layer1_outputs(1494) <= '0';
    layer1_outputs(1495) <= '0';
    layer1_outputs(1496) <= not((layer0_outputs(2019)) or (layer0_outputs(387)));
    layer1_outputs(1497) <= not(layer0_outputs(1405)) or (layer0_outputs(591));
    layer1_outputs(1498) <= not((layer0_outputs(1426)) and (layer0_outputs(2147)));
    layer1_outputs(1499) <= not(layer0_outputs(1727));
    layer1_outputs(1500) <= (layer0_outputs(355)) and not (layer0_outputs(2278));
    layer1_outputs(1501) <= layer0_outputs(1899);
    layer1_outputs(1502) <= (layer0_outputs(2212)) and (layer0_outputs(1002));
    layer1_outputs(1503) <= not(layer0_outputs(407)) or (layer0_outputs(536));
    layer1_outputs(1504) <= (layer0_outputs(2135)) or (layer0_outputs(1303));
    layer1_outputs(1505) <= not(layer0_outputs(1347));
    layer1_outputs(1506) <= not(layer0_outputs(925)) or (layer0_outputs(1337));
    layer1_outputs(1507) <= not((layer0_outputs(1916)) and (layer0_outputs(1183)));
    layer1_outputs(1508) <= not(layer0_outputs(2167));
    layer1_outputs(1509) <= not(layer0_outputs(2536));
    layer1_outputs(1510) <= not(layer0_outputs(1706));
    layer1_outputs(1511) <= layer0_outputs(360);
    layer1_outputs(1512) <= (layer0_outputs(1841)) and not (layer0_outputs(1924));
    layer1_outputs(1513) <= '0';
    layer1_outputs(1514) <= not(layer0_outputs(2269));
    layer1_outputs(1515) <= not((layer0_outputs(1175)) xor (layer0_outputs(219)));
    layer1_outputs(1516) <= not(layer0_outputs(1049)) or (layer0_outputs(1226));
    layer1_outputs(1517) <= '1';
    layer1_outputs(1518) <= (layer0_outputs(637)) and (layer0_outputs(200));
    layer1_outputs(1519) <= not((layer0_outputs(471)) and (layer0_outputs(2347)));
    layer1_outputs(1520) <= (layer0_outputs(1788)) or (layer0_outputs(319));
    layer1_outputs(1521) <= layer0_outputs(1781);
    layer1_outputs(1522) <= not(layer0_outputs(1702));
    layer1_outputs(1523) <= '0';
    layer1_outputs(1524) <= '1';
    layer1_outputs(1525) <= (layer0_outputs(380)) and not (layer0_outputs(846));
    layer1_outputs(1526) <= (layer0_outputs(306)) and not (layer0_outputs(2154));
    layer1_outputs(1527) <= layer0_outputs(854);
    layer1_outputs(1528) <= not(layer0_outputs(708)) or (layer0_outputs(1798));
    layer1_outputs(1529) <= not(layer0_outputs(1556)) or (layer0_outputs(2223));
    layer1_outputs(1530) <= (layer0_outputs(2317)) or (layer0_outputs(1330));
    layer1_outputs(1531) <= (layer0_outputs(522)) and not (layer0_outputs(1110));
    layer1_outputs(1532) <= not(layer0_outputs(302));
    layer1_outputs(1533) <= not((layer0_outputs(1301)) and (layer0_outputs(164)));
    layer1_outputs(1534) <= '0';
    layer1_outputs(1535) <= not(layer0_outputs(1095)) or (layer0_outputs(1837));
    layer1_outputs(1536) <= not(layer0_outputs(1395));
    layer1_outputs(1537) <= not(layer0_outputs(798));
    layer1_outputs(1538) <= (layer0_outputs(903)) or (layer0_outputs(1651));
    layer1_outputs(1539) <= '1';
    layer1_outputs(1540) <= not(layer0_outputs(1680)) or (layer0_outputs(1715));
    layer1_outputs(1541) <= layer0_outputs(253);
    layer1_outputs(1542) <= not(layer0_outputs(179));
    layer1_outputs(1543) <= not((layer0_outputs(1635)) and (layer0_outputs(275)));
    layer1_outputs(1544) <= not(layer0_outputs(174));
    layer1_outputs(1545) <= not(layer0_outputs(746));
    layer1_outputs(1546) <= not((layer0_outputs(1010)) or (layer0_outputs(796)));
    layer1_outputs(1547) <= (layer0_outputs(2273)) or (layer0_outputs(1030));
    layer1_outputs(1548) <= not((layer0_outputs(818)) and (layer0_outputs(1057)));
    layer1_outputs(1549) <= not(layer0_outputs(1217)) or (layer0_outputs(31));
    layer1_outputs(1550) <= layer0_outputs(2466);
    layer1_outputs(1551) <= '0';
    layer1_outputs(1552) <= not(layer0_outputs(350)) or (layer0_outputs(137));
    layer1_outputs(1553) <= (layer0_outputs(290)) and (layer0_outputs(2088));
    layer1_outputs(1554) <= '0';
    layer1_outputs(1555) <= not((layer0_outputs(451)) or (layer0_outputs(866)));
    layer1_outputs(1556) <= not((layer0_outputs(622)) or (layer0_outputs(2278)));
    layer1_outputs(1557) <= not(layer0_outputs(2216)) or (layer0_outputs(961));
    layer1_outputs(1558) <= (layer0_outputs(2426)) and (layer0_outputs(1968));
    layer1_outputs(1559) <= '1';
    layer1_outputs(1560) <= (layer0_outputs(2116)) and not (layer0_outputs(971));
    layer1_outputs(1561) <= layer0_outputs(1885);
    layer1_outputs(1562) <= (layer0_outputs(154)) and (layer0_outputs(1505));
    layer1_outputs(1563) <= layer0_outputs(63);
    layer1_outputs(1564) <= not(layer0_outputs(1585));
    layer1_outputs(1565) <= not((layer0_outputs(1537)) and (layer0_outputs(2289)));
    layer1_outputs(1566) <= (layer0_outputs(1125)) and not (layer0_outputs(1403));
    layer1_outputs(1567) <= not(layer0_outputs(1900));
    layer1_outputs(1568) <= not(layer0_outputs(1801));
    layer1_outputs(1569) <= '0';
    layer1_outputs(1570) <= (layer0_outputs(1544)) and not (layer0_outputs(373));
    layer1_outputs(1571) <= not(layer0_outputs(1825));
    layer1_outputs(1572) <= (layer0_outputs(2069)) and not (layer0_outputs(630));
    layer1_outputs(1573) <= not((layer0_outputs(1922)) or (layer0_outputs(1967)));
    layer1_outputs(1574) <= (layer0_outputs(418)) and not (layer0_outputs(890));
    layer1_outputs(1575) <= not(layer0_outputs(1511)) or (layer0_outputs(263));
    layer1_outputs(1576) <= (layer0_outputs(1985)) and (layer0_outputs(655));
    layer1_outputs(1577) <= '0';
    layer1_outputs(1578) <= (layer0_outputs(2301)) or (layer0_outputs(2085));
    layer1_outputs(1579) <= not(layer0_outputs(2007));
    layer1_outputs(1580) <= not(layer0_outputs(28));
    layer1_outputs(1581) <= (layer0_outputs(1483)) or (layer0_outputs(574));
    layer1_outputs(1582) <= not(layer0_outputs(1172)) or (layer0_outputs(2209));
    layer1_outputs(1583) <= (layer0_outputs(100)) xor (layer0_outputs(834));
    layer1_outputs(1584) <= not(layer0_outputs(1063));
    layer1_outputs(1585) <= '1';
    layer1_outputs(1586) <= not((layer0_outputs(2089)) and (layer0_outputs(55)));
    layer1_outputs(1587) <= (layer0_outputs(1475)) and not (layer0_outputs(1609));
    layer1_outputs(1588) <= (layer0_outputs(1626)) or (layer0_outputs(653));
    layer1_outputs(1589) <= (layer0_outputs(224)) or (layer0_outputs(95));
    layer1_outputs(1590) <= (layer0_outputs(1044)) and (layer0_outputs(1773));
    layer1_outputs(1591) <= not((layer0_outputs(1156)) or (layer0_outputs(876)));
    layer1_outputs(1592) <= not(layer0_outputs(2285));
    layer1_outputs(1593) <= not(layer0_outputs(1152)) or (layer0_outputs(1770));
    layer1_outputs(1594) <= '1';
    layer1_outputs(1595) <= not(layer0_outputs(347)) or (layer0_outputs(1841));
    layer1_outputs(1596) <= not(layer0_outputs(2209));
    layer1_outputs(1597) <= '1';
    layer1_outputs(1598) <= not(layer0_outputs(1786));
    layer1_outputs(1599) <= layer0_outputs(2343);
    layer1_outputs(1600) <= (layer0_outputs(67)) or (layer0_outputs(554));
    layer1_outputs(1601) <= '0';
    layer1_outputs(1602) <= (layer0_outputs(1167)) and not (layer0_outputs(247));
    layer1_outputs(1603) <= '0';
    layer1_outputs(1604) <= not(layer0_outputs(2176)) or (layer0_outputs(1656));
    layer1_outputs(1605) <= '1';
    layer1_outputs(1606) <= not(layer0_outputs(1739));
    layer1_outputs(1607) <= (layer0_outputs(1265)) and not (layer0_outputs(2123));
    layer1_outputs(1608) <= layer0_outputs(1860);
    layer1_outputs(1609) <= '0';
    layer1_outputs(1610) <= not(layer0_outputs(258));
    layer1_outputs(1611) <= '0';
    layer1_outputs(1612) <= layer0_outputs(402);
    layer1_outputs(1613) <= (layer0_outputs(120)) or (layer0_outputs(2106));
    layer1_outputs(1614) <= (layer0_outputs(345)) and not (layer0_outputs(1380));
    layer1_outputs(1615) <= layer0_outputs(2082);
    layer1_outputs(1616) <= (layer0_outputs(718)) or (layer0_outputs(2335));
    layer1_outputs(1617) <= (layer0_outputs(870)) and not (layer0_outputs(1625));
    layer1_outputs(1618) <= (layer0_outputs(2541)) and not (layer0_outputs(2521));
    layer1_outputs(1619) <= layer0_outputs(2364);
    layer1_outputs(1620) <= not(layer0_outputs(317)) or (layer0_outputs(2339));
    layer1_outputs(1621) <= (layer0_outputs(1856)) and not (layer0_outputs(1887));
    layer1_outputs(1622) <= (layer0_outputs(2283)) and not (layer0_outputs(1820));
    layer1_outputs(1623) <= (layer0_outputs(864)) and not (layer0_outputs(2315));
    layer1_outputs(1624) <= (layer0_outputs(54)) or (layer0_outputs(1510));
    layer1_outputs(1625) <= '0';
    layer1_outputs(1626) <= (layer0_outputs(555)) and not (layer0_outputs(384));
    layer1_outputs(1627) <= not(layer0_outputs(1246)) or (layer0_outputs(2031));
    layer1_outputs(1628) <= (layer0_outputs(177)) and not (layer0_outputs(2052));
    layer1_outputs(1629) <= layer0_outputs(1255);
    layer1_outputs(1630) <= (layer0_outputs(2549)) xor (layer0_outputs(2228));
    layer1_outputs(1631) <= layer0_outputs(1413);
    layer1_outputs(1632) <= '1';
    layer1_outputs(1633) <= layer0_outputs(1943);
    layer1_outputs(1634) <= '0';
    layer1_outputs(1635) <= '1';
    layer1_outputs(1636) <= not((layer0_outputs(631)) or (layer0_outputs(679)));
    layer1_outputs(1637) <= (layer0_outputs(2524)) and not (layer0_outputs(2328));
    layer1_outputs(1638) <= '0';
    layer1_outputs(1639) <= layer0_outputs(2022);
    layer1_outputs(1640) <= not(layer0_outputs(867));
    layer1_outputs(1641) <= layer0_outputs(924);
    layer1_outputs(1642) <= not(layer0_outputs(710)) or (layer0_outputs(483));
    layer1_outputs(1643) <= layer0_outputs(1491);
    layer1_outputs(1644) <= not(layer0_outputs(793)) or (layer0_outputs(1854));
    layer1_outputs(1645) <= not(layer0_outputs(1406));
    layer1_outputs(1646) <= (layer0_outputs(704)) and (layer0_outputs(2008));
    layer1_outputs(1647) <= (layer0_outputs(1784)) or (layer0_outputs(1540));
    layer1_outputs(1648) <= not(layer0_outputs(892));
    layer1_outputs(1649) <= layer0_outputs(736);
    layer1_outputs(1650) <= layer0_outputs(1047);
    layer1_outputs(1651) <= layer0_outputs(2333);
    layer1_outputs(1652) <= not(layer0_outputs(925)) or (layer0_outputs(2019));
    layer1_outputs(1653) <= not(layer0_outputs(2243)) or (layer0_outputs(188));
    layer1_outputs(1654) <= not((layer0_outputs(491)) or (layer0_outputs(2336)));
    layer1_outputs(1655) <= not(layer0_outputs(1113));
    layer1_outputs(1656) <= (layer0_outputs(2344)) and not (layer0_outputs(0));
    layer1_outputs(1657) <= not(layer0_outputs(499));
    layer1_outputs(1658) <= '1';
    layer1_outputs(1659) <= not(layer0_outputs(1828));
    layer1_outputs(1660) <= not(layer0_outputs(1560));
    layer1_outputs(1661) <= (layer0_outputs(1459)) and (layer0_outputs(582));
    layer1_outputs(1662) <= not((layer0_outputs(2251)) or (layer0_outputs(1869)));
    layer1_outputs(1663) <= layer0_outputs(567);
    layer1_outputs(1664) <= not((layer0_outputs(2217)) and (layer0_outputs(2133)));
    layer1_outputs(1665) <= layer0_outputs(2250);
    layer1_outputs(1666) <= (layer0_outputs(1794)) or (layer0_outputs(2505));
    layer1_outputs(1667) <= layer0_outputs(1620);
    layer1_outputs(1668) <= (layer0_outputs(1286)) and not (layer0_outputs(505));
    layer1_outputs(1669) <= not(layer0_outputs(1707));
    layer1_outputs(1670) <= not(layer0_outputs(498));
    layer1_outputs(1671) <= (layer0_outputs(300)) or (layer0_outputs(52));
    layer1_outputs(1672) <= not(layer0_outputs(695)) or (layer0_outputs(1041));
    layer1_outputs(1673) <= '0';
    layer1_outputs(1674) <= layer0_outputs(2205);
    layer1_outputs(1675) <= (layer0_outputs(658)) and not (layer0_outputs(1237));
    layer1_outputs(1676) <= layer0_outputs(2390);
    layer1_outputs(1677) <= layer0_outputs(132);
    layer1_outputs(1678) <= '0';
    layer1_outputs(1679) <= '0';
    layer1_outputs(1680) <= not(layer0_outputs(47));
    layer1_outputs(1681) <= not((layer0_outputs(2458)) and (layer0_outputs(850)));
    layer1_outputs(1682) <= not(layer0_outputs(1919)) or (layer0_outputs(1677));
    layer1_outputs(1683) <= not((layer0_outputs(606)) and (layer0_outputs(1087)));
    layer1_outputs(1684) <= '0';
    layer1_outputs(1685) <= (layer0_outputs(638)) xor (layer0_outputs(86));
    layer1_outputs(1686) <= layer0_outputs(2260);
    layer1_outputs(1687) <= not(layer0_outputs(2157));
    layer1_outputs(1688) <= not(layer0_outputs(2250));
    layer1_outputs(1689) <= not(layer0_outputs(2051));
    layer1_outputs(1690) <= layer0_outputs(992);
    layer1_outputs(1691) <= (layer0_outputs(334)) and not (layer0_outputs(2119));
    layer1_outputs(1692) <= not((layer0_outputs(1253)) or (layer0_outputs(1208)));
    layer1_outputs(1693) <= not((layer0_outputs(1618)) and (layer0_outputs(2438)));
    layer1_outputs(1694) <= layer0_outputs(1247);
    layer1_outputs(1695) <= not(layer0_outputs(1073)) or (layer0_outputs(920));
    layer1_outputs(1696) <= not(layer0_outputs(1995)) or (layer0_outputs(1564));
    layer1_outputs(1697) <= (layer0_outputs(349)) and not (layer0_outputs(1855));
    layer1_outputs(1698) <= not(layer0_outputs(1113)) or (layer0_outputs(310));
    layer1_outputs(1699) <= not(layer0_outputs(2393)) or (layer0_outputs(792));
    layer1_outputs(1700) <= '0';
    layer1_outputs(1701) <= '1';
    layer1_outputs(1702) <= not(layer0_outputs(2284)) or (layer0_outputs(87));
    layer1_outputs(1703) <= '0';
    layer1_outputs(1704) <= not(layer0_outputs(372)) or (layer0_outputs(1471));
    layer1_outputs(1705) <= layer0_outputs(847);
    layer1_outputs(1706) <= not(layer0_outputs(538)) or (layer0_outputs(1709));
    layer1_outputs(1707) <= not(layer0_outputs(128)) or (layer0_outputs(670));
    layer1_outputs(1708) <= layer0_outputs(861);
    layer1_outputs(1709) <= not((layer0_outputs(2402)) or (layer0_outputs(837)));
    layer1_outputs(1710) <= not(layer0_outputs(2194)) or (layer0_outputs(1314));
    layer1_outputs(1711) <= (layer0_outputs(586)) and not (layer0_outputs(1803));
    layer1_outputs(1712) <= (layer0_outputs(927)) and not (layer0_outputs(2163));
    layer1_outputs(1713) <= '0';
    layer1_outputs(1714) <= (layer0_outputs(968)) and not (layer0_outputs(574));
    layer1_outputs(1715) <= (layer0_outputs(1097)) and not (layer0_outputs(2341));
    layer1_outputs(1716) <= (layer0_outputs(46)) and (layer0_outputs(1693));
    layer1_outputs(1717) <= not(layer0_outputs(1213)) or (layer0_outputs(2090));
    layer1_outputs(1718) <= not((layer0_outputs(1428)) and (layer0_outputs(39)));
    layer1_outputs(1719) <= not((layer0_outputs(2297)) and (layer0_outputs(257)));
    layer1_outputs(1720) <= not(layer0_outputs(2461));
    layer1_outputs(1721) <= not(layer0_outputs(1504));
    layer1_outputs(1722) <= not(layer0_outputs(478)) or (layer0_outputs(872));
    layer1_outputs(1723) <= (layer0_outputs(669)) and not (layer0_outputs(475));
    layer1_outputs(1724) <= not((layer0_outputs(942)) and (layer0_outputs(1251)));
    layer1_outputs(1725) <= not(layer0_outputs(871)) or (layer0_outputs(1332));
    layer1_outputs(1726) <= not(layer0_outputs(583));
    layer1_outputs(1727) <= layer0_outputs(1918);
    layer1_outputs(1728) <= '1';
    layer1_outputs(1729) <= (layer0_outputs(173)) and (layer0_outputs(2103));
    layer1_outputs(1730) <= layer0_outputs(246);
    layer1_outputs(1731) <= (layer0_outputs(1995)) and (layer0_outputs(2518));
    layer1_outputs(1732) <= not(layer0_outputs(1908)) or (layer0_outputs(1951));
    layer1_outputs(1733) <= layer0_outputs(281);
    layer1_outputs(1734) <= layer0_outputs(2089);
    layer1_outputs(1735) <= layer0_outputs(938);
    layer1_outputs(1736) <= (layer0_outputs(1978)) and not (layer0_outputs(1214));
    layer1_outputs(1737) <= layer0_outputs(1002);
    layer1_outputs(1738) <= '0';
    layer1_outputs(1739) <= (layer0_outputs(1279)) and (layer0_outputs(663));
    layer1_outputs(1740) <= not(layer0_outputs(2504)) or (layer0_outputs(2460));
    layer1_outputs(1741) <= not(layer0_outputs(1357));
    layer1_outputs(1742) <= not(layer0_outputs(1814));
    layer1_outputs(1743) <= (layer0_outputs(2509)) and not (layer0_outputs(611));
    layer1_outputs(1744) <= '0';
    layer1_outputs(1745) <= not(layer0_outputs(93));
    layer1_outputs(1746) <= not((layer0_outputs(1064)) and (layer0_outputs(1161)));
    layer1_outputs(1747) <= not((layer0_outputs(1579)) or (layer0_outputs(1271)));
    layer1_outputs(1748) <= layer0_outputs(2503);
    layer1_outputs(1749) <= '1';
    layer1_outputs(1750) <= not((layer0_outputs(405)) or (layer0_outputs(2355)));
    layer1_outputs(1751) <= '1';
    layer1_outputs(1752) <= (layer0_outputs(2130)) and not (layer0_outputs(608));
    layer1_outputs(1753) <= not((layer0_outputs(1913)) and (layer0_outputs(2064)));
    layer1_outputs(1754) <= not(layer0_outputs(2203)) or (layer0_outputs(220));
    layer1_outputs(1755) <= '1';
    layer1_outputs(1756) <= not(layer0_outputs(2484)) or (layer0_outputs(789));
    layer1_outputs(1757) <= layer0_outputs(1786);
    layer1_outputs(1758) <= layer0_outputs(2156);
    layer1_outputs(1759) <= not(layer0_outputs(2254)) or (layer0_outputs(2332));
    layer1_outputs(1760) <= not(layer0_outputs(645)) or (layer0_outputs(285));
    layer1_outputs(1761) <= not(layer0_outputs(2415));
    layer1_outputs(1762) <= not(layer0_outputs(1971)) or (layer0_outputs(1333));
    layer1_outputs(1763) <= '1';
    layer1_outputs(1764) <= (layer0_outputs(855)) and not (layer0_outputs(1472));
    layer1_outputs(1765) <= (layer0_outputs(1605)) and not (layer0_outputs(288));
    layer1_outputs(1766) <= not(layer0_outputs(262)) or (layer0_outputs(368));
    layer1_outputs(1767) <= (layer0_outputs(1333)) and (layer0_outputs(531));
    layer1_outputs(1768) <= not(layer0_outputs(1149)) or (layer0_outputs(1507));
    layer1_outputs(1769) <= layer0_outputs(2341);
    layer1_outputs(1770) <= not(layer0_outputs(569)) or (layer0_outputs(840));
    layer1_outputs(1771) <= layer0_outputs(1900);
    layer1_outputs(1772) <= not(layer0_outputs(647));
    layer1_outputs(1773) <= not(layer0_outputs(1031));
    layer1_outputs(1774) <= '1';
    layer1_outputs(1775) <= not((layer0_outputs(2182)) or (layer0_outputs(385)));
    layer1_outputs(1776) <= '1';
    layer1_outputs(1777) <= '0';
    layer1_outputs(1778) <= '1';
    layer1_outputs(1779) <= layer0_outputs(1432);
    layer1_outputs(1780) <= not((layer0_outputs(1757)) and (layer0_outputs(316)));
    layer1_outputs(1781) <= '0';
    layer1_outputs(1782) <= '0';
    layer1_outputs(1783) <= '0';
    layer1_outputs(1784) <= (layer0_outputs(2053)) and not (layer0_outputs(444));
    layer1_outputs(1785) <= not(layer0_outputs(2016));
    layer1_outputs(1786) <= not(layer0_outputs(2434)) or (layer0_outputs(2015));
    layer1_outputs(1787) <= not(layer0_outputs(212));
    layer1_outputs(1788) <= layer0_outputs(1591);
    layer1_outputs(1789) <= not(layer0_outputs(1965));
    layer1_outputs(1790) <= not(layer0_outputs(977)) or (layer0_outputs(53));
    layer1_outputs(1791) <= not(layer0_outputs(715)) or (layer0_outputs(283));
    layer1_outputs(1792) <= (layer0_outputs(37)) and (layer0_outputs(1888));
    layer1_outputs(1793) <= not(layer0_outputs(815));
    layer1_outputs(1794) <= '1';
    layer1_outputs(1795) <= not(layer0_outputs(1124));
    layer1_outputs(1796) <= not(layer0_outputs(1840));
    layer1_outputs(1797) <= not(layer0_outputs(2298)) or (layer0_outputs(1588));
    layer1_outputs(1798) <= not(layer0_outputs(1029));
    layer1_outputs(1799) <= not(layer0_outputs(168)) or (layer0_outputs(1160));
    layer1_outputs(1800) <= (layer0_outputs(1065)) and not (layer0_outputs(1859));
    layer1_outputs(1801) <= (layer0_outputs(1999)) xor (layer0_outputs(2146));
    layer1_outputs(1802) <= not(layer0_outputs(2103)) or (layer0_outputs(2270));
    layer1_outputs(1803) <= (layer0_outputs(1847)) and (layer0_outputs(391));
    layer1_outputs(1804) <= (layer0_outputs(8)) and not (layer0_outputs(2080));
    layer1_outputs(1805) <= layer0_outputs(773);
    layer1_outputs(1806) <= not(layer0_outputs(2480));
    layer1_outputs(1807) <= (layer0_outputs(2068)) and not (layer0_outputs(234));
    layer1_outputs(1808) <= not((layer0_outputs(1750)) and (layer0_outputs(1443)));
    layer1_outputs(1809) <= (layer0_outputs(910)) or (layer0_outputs(2196));
    layer1_outputs(1810) <= not(layer0_outputs(553));
    layer1_outputs(1811) <= not((layer0_outputs(612)) and (layer0_outputs(577)));
    layer1_outputs(1812) <= (layer0_outputs(2411)) and (layer0_outputs(1897));
    layer1_outputs(1813) <= (layer0_outputs(2300)) and not (layer0_outputs(356));
    layer1_outputs(1814) <= '1';
    layer1_outputs(1815) <= not((layer0_outputs(122)) and (layer0_outputs(1791)));
    layer1_outputs(1816) <= (layer0_outputs(497)) and not (layer0_outputs(2041));
    layer1_outputs(1817) <= (layer0_outputs(446)) xor (layer0_outputs(2308));
    layer1_outputs(1818) <= (layer0_outputs(1740)) or (layer0_outputs(2377));
    layer1_outputs(1819) <= '0';
    layer1_outputs(1820) <= not((layer0_outputs(654)) and (layer0_outputs(756)));
    layer1_outputs(1821) <= not((layer0_outputs(1441)) and (layer0_outputs(2522)));
    layer1_outputs(1822) <= '0';
    layer1_outputs(1823) <= (layer0_outputs(1747)) and not (layer0_outputs(346));
    layer1_outputs(1824) <= not(layer0_outputs(464));
    layer1_outputs(1825) <= (layer0_outputs(453)) and (layer0_outputs(1977));
    layer1_outputs(1826) <= not((layer0_outputs(450)) or (layer0_outputs(1815)));
    layer1_outputs(1827) <= '1';
    layer1_outputs(1828) <= (layer0_outputs(1561)) or (layer0_outputs(1731));
    layer1_outputs(1829) <= not((layer0_outputs(1849)) and (layer0_outputs(152)));
    layer1_outputs(1830) <= (layer0_outputs(1098)) and (layer0_outputs(1991));
    layer1_outputs(1831) <= '1';
    layer1_outputs(1832) <= (layer0_outputs(248)) and not (layer0_outputs(1694));
    layer1_outputs(1833) <= (layer0_outputs(205)) or (layer0_outputs(743));
    layer1_outputs(1834) <= (layer0_outputs(919)) or (layer0_outputs(2384));
    layer1_outputs(1835) <= (layer0_outputs(780)) and not (layer0_outputs(532));
    layer1_outputs(1836) <= not((layer0_outputs(1637)) and (layer0_outputs(1648)));
    layer1_outputs(1837) <= '0';
    layer1_outputs(1838) <= layer0_outputs(75);
    layer1_outputs(1839) <= '1';
    layer1_outputs(1840) <= not(layer0_outputs(1394));
    layer1_outputs(1841) <= not(layer0_outputs(267));
    layer1_outputs(1842) <= (layer0_outputs(467)) and (layer0_outputs(21));
    layer1_outputs(1843) <= not((layer0_outputs(573)) or (layer0_outputs(2382)));
    layer1_outputs(1844) <= '0';
    layer1_outputs(1845) <= '1';
    layer1_outputs(1846) <= '1';
    layer1_outputs(1847) <= not((layer0_outputs(1440)) or (layer0_outputs(242)));
    layer1_outputs(1848) <= not(layer0_outputs(1220)) or (layer0_outputs(2121));
    layer1_outputs(1849) <= layer0_outputs(410);
    layer1_outputs(1850) <= '0';
    layer1_outputs(1851) <= not((layer0_outputs(1236)) or (layer0_outputs(2013)));
    layer1_outputs(1852) <= not(layer0_outputs(2027)) or (layer0_outputs(1668));
    layer1_outputs(1853) <= not((layer0_outputs(1660)) and (layer0_outputs(1589)));
    layer1_outputs(1854) <= not(layer0_outputs(1235)) or (layer0_outputs(1037));
    layer1_outputs(1855) <= not(layer0_outputs(1072));
    layer1_outputs(1856) <= layer0_outputs(1976);
    layer1_outputs(1857) <= not(layer0_outputs(2313));
    layer1_outputs(1858) <= not(layer0_outputs(2431)) or (layer0_outputs(98));
    layer1_outputs(1859) <= not((layer0_outputs(2070)) or (layer0_outputs(1267)));
    layer1_outputs(1860) <= layer0_outputs(911);
    layer1_outputs(1861) <= not((layer0_outputs(1797)) or (layer0_outputs(1583)));
    layer1_outputs(1862) <= not((layer0_outputs(144)) and (layer0_outputs(2470)));
    layer1_outputs(1863) <= layer0_outputs(608);
    layer1_outputs(1864) <= (layer0_outputs(1075)) and not (layer0_outputs(243));
    layer1_outputs(1865) <= not(layer0_outputs(1889)) or (layer0_outputs(2198));
    layer1_outputs(1866) <= layer0_outputs(2069);
    layer1_outputs(1867) <= not(layer0_outputs(2331));
    layer1_outputs(1868) <= (layer0_outputs(1226)) or (layer0_outputs(322));
    layer1_outputs(1869) <= not(layer0_outputs(524));
    layer1_outputs(1870) <= '1';
    layer1_outputs(1871) <= layer0_outputs(125);
    layer1_outputs(1872) <= not(layer0_outputs(2277));
    layer1_outputs(1873) <= '1';
    layer1_outputs(1874) <= '0';
    layer1_outputs(1875) <= '1';
    layer1_outputs(1876) <= layer0_outputs(1296);
    layer1_outputs(1877) <= layer0_outputs(2270);
    layer1_outputs(1878) <= '0';
    layer1_outputs(1879) <= (layer0_outputs(1593)) or (layer0_outputs(2453));
    layer1_outputs(1880) <= not((layer0_outputs(1641)) and (layer0_outputs(272)));
    layer1_outputs(1881) <= not(layer0_outputs(1502)) or (layer0_outputs(448));
    layer1_outputs(1882) <= '1';
    layer1_outputs(1883) <= (layer0_outputs(115)) and not (layer0_outputs(408));
    layer1_outputs(1884) <= (layer0_outputs(1582)) and not (layer0_outputs(1400));
    layer1_outputs(1885) <= '1';
    layer1_outputs(1886) <= (layer0_outputs(1935)) and (layer0_outputs(1384));
    layer1_outputs(1887) <= (layer0_outputs(284)) and not (layer0_outputs(1148));
    layer1_outputs(1888) <= not(layer0_outputs(1074)) or (layer0_outputs(1130));
    layer1_outputs(1889) <= not((layer0_outputs(348)) or (layer0_outputs(2117)));
    layer1_outputs(1890) <= '0';
    layer1_outputs(1891) <= not(layer0_outputs(1755)) or (layer0_outputs(2520));
    layer1_outputs(1892) <= layer0_outputs(1805);
    layer1_outputs(1893) <= not(layer0_outputs(477));
    layer1_outputs(1894) <= layer0_outputs(162);
    layer1_outputs(1895) <= not(layer0_outputs(2131)) or (layer0_outputs(1517));
    layer1_outputs(1896) <= not((layer0_outputs(278)) and (layer0_outputs(978)));
    layer1_outputs(1897) <= not((layer0_outputs(1424)) or (layer0_outputs(1756)));
    layer1_outputs(1898) <= not(layer0_outputs(1520));
    layer1_outputs(1899) <= (layer0_outputs(2496)) and (layer0_outputs(1776));
    layer1_outputs(1900) <= (layer0_outputs(388)) and not (layer0_outputs(1799));
    layer1_outputs(1901) <= '1';
    layer1_outputs(1902) <= not(layer0_outputs(1535));
    layer1_outputs(1903) <= (layer0_outputs(1975)) or (layer0_outputs(1463));
    layer1_outputs(1904) <= layer0_outputs(2245);
    layer1_outputs(1905) <= (layer0_outputs(1355)) and not (layer0_outputs(2150));
    layer1_outputs(1906) <= '1';
    layer1_outputs(1907) <= not(layer0_outputs(705)) or (layer0_outputs(723));
    layer1_outputs(1908) <= layer0_outputs(2150);
    layer1_outputs(1909) <= not(layer0_outputs(1851)) or (layer0_outputs(879));
    layer1_outputs(1910) <= not(layer0_outputs(2536));
    layer1_outputs(1911) <= not((layer0_outputs(150)) or (layer0_outputs(1449)));
    layer1_outputs(1912) <= not(layer0_outputs(280));
    layer1_outputs(1913) <= layer0_outputs(1595);
    layer1_outputs(1914) <= layer0_outputs(1277);
    layer1_outputs(1915) <= layer0_outputs(1620);
    layer1_outputs(1916) <= (layer0_outputs(1853)) and not (layer0_outputs(1305));
    layer1_outputs(1917) <= (layer0_outputs(1574)) and not (layer0_outputs(764));
    layer1_outputs(1918) <= not((layer0_outputs(1581)) or (layer0_outputs(548)));
    layer1_outputs(1919) <= (layer0_outputs(1115)) and not (layer0_outputs(865));
    layer1_outputs(1920) <= layer0_outputs(307);
    layer1_outputs(1921) <= not(layer0_outputs(1148)) or (layer0_outputs(500));
    layer1_outputs(1922) <= '0';
    layer1_outputs(1923) <= not((layer0_outputs(883)) and (layer0_outputs(346)));
    layer1_outputs(1924) <= layer0_outputs(916);
    layer1_outputs(1925) <= (layer0_outputs(1780)) and not (layer0_outputs(272));
    layer1_outputs(1926) <= not(layer0_outputs(1665)) or (layer0_outputs(591));
    layer1_outputs(1927) <= (layer0_outputs(1531)) and (layer0_outputs(228));
    layer1_outputs(1928) <= '0';
    layer1_outputs(1929) <= not(layer0_outputs(2351));
    layer1_outputs(1930) <= layer0_outputs(912);
    layer1_outputs(1931) <= not((layer0_outputs(406)) or (layer0_outputs(99)));
    layer1_outputs(1932) <= not((layer0_outputs(1429)) or (layer0_outputs(2318)));
    layer1_outputs(1933) <= not(layer0_outputs(1114)) or (layer0_outputs(1532));
    layer1_outputs(1934) <= (layer0_outputs(130)) or (layer0_outputs(1550));
    layer1_outputs(1935) <= layer0_outputs(1116);
    layer1_outputs(1936) <= not((layer0_outputs(2405)) or (layer0_outputs(2533)));
    layer1_outputs(1937) <= not(layer0_outputs(1295)) or (layer0_outputs(1366));
    layer1_outputs(1938) <= not((layer0_outputs(1323)) or (layer0_outputs(1402)));
    layer1_outputs(1939) <= layer0_outputs(864);
    layer1_outputs(1940) <= layer0_outputs(2256);
    layer1_outputs(1941) <= (layer0_outputs(1379)) and (layer0_outputs(901));
    layer1_outputs(1942) <= not((layer0_outputs(370)) or (layer0_outputs(2287)));
    layer1_outputs(1943) <= '0';
    layer1_outputs(1944) <= (layer0_outputs(2425)) and (layer0_outputs(1787));
    layer1_outputs(1945) <= not(layer0_outputs(2391)) or (layer0_outputs(1082));
    layer1_outputs(1946) <= '1';
    layer1_outputs(1947) <= (layer0_outputs(1004)) and not (layer0_outputs(1649));
    layer1_outputs(1948) <= (layer0_outputs(1162)) and not (layer0_outputs(2542));
    layer1_outputs(1949) <= '1';
    layer1_outputs(1950) <= (layer0_outputs(687)) and not (layer0_outputs(1206));
    layer1_outputs(1951) <= layer0_outputs(701);
    layer1_outputs(1952) <= layer0_outputs(1106);
    layer1_outputs(1953) <= not(layer0_outputs(1909));
    layer1_outputs(1954) <= '0';
    layer1_outputs(1955) <= not((layer0_outputs(227)) or (layer0_outputs(886)));
    layer1_outputs(1956) <= not(layer0_outputs(1388));
    layer1_outputs(1957) <= (layer0_outputs(1563)) and (layer0_outputs(2149));
    layer1_outputs(1958) <= layer0_outputs(1294);
    layer1_outputs(1959) <= layer0_outputs(1413);
    layer1_outputs(1960) <= layer0_outputs(1142);
    layer1_outputs(1961) <= not(layer0_outputs(1920)) or (layer0_outputs(1452));
    layer1_outputs(1962) <= not(layer0_outputs(1051)) or (layer0_outputs(1094));
    layer1_outputs(1963) <= not(layer0_outputs(1456));
    layer1_outputs(1964) <= not(layer0_outputs(707)) or (layer0_outputs(727));
    layer1_outputs(1965) <= (layer0_outputs(643)) and (layer0_outputs(1053));
    layer1_outputs(1966) <= (layer0_outputs(1684)) and (layer0_outputs(11));
    layer1_outputs(1967) <= (layer0_outputs(710)) xor (layer0_outputs(1642));
    layer1_outputs(1968) <= '1';
    layer1_outputs(1969) <= not(layer0_outputs(2389));
    layer1_outputs(1970) <= (layer0_outputs(825)) and not (layer0_outputs(397));
    layer1_outputs(1971) <= not((layer0_outputs(534)) and (layer0_outputs(634)));
    layer1_outputs(1972) <= not(layer0_outputs(2055));
    layer1_outputs(1973) <= not((layer0_outputs(2459)) or (layer0_outputs(2098)));
    layer1_outputs(1974) <= (layer0_outputs(1966)) and (layer0_outputs(124));
    layer1_outputs(1975) <= not(layer0_outputs(996));
    layer1_outputs(1976) <= layer0_outputs(1895);
    layer1_outputs(1977) <= (layer0_outputs(1001)) and not (layer0_outputs(314));
    layer1_outputs(1978) <= (layer0_outputs(2202)) and not (layer0_outputs(1819));
    layer1_outputs(1979) <= not(layer0_outputs(2195));
    layer1_outputs(1980) <= layer0_outputs(1325);
    layer1_outputs(1981) <= (layer0_outputs(1024)) and not (layer0_outputs(2210));
    layer1_outputs(1982) <= (layer0_outputs(2473)) and (layer0_outputs(1175));
    layer1_outputs(1983) <= '0';
    layer1_outputs(1984) <= layer0_outputs(734);
    layer1_outputs(1985) <= (layer0_outputs(1848)) or (layer0_outputs(1600));
    layer1_outputs(1986) <= not(layer0_outputs(1448));
    layer1_outputs(1987) <= layer0_outputs(297);
    layer1_outputs(1988) <= not(layer0_outputs(324));
    layer1_outputs(1989) <= (layer0_outputs(2466)) or (layer0_outputs(1215));
    layer1_outputs(1990) <= '0';
    layer1_outputs(1991) <= '1';
    layer1_outputs(1992) <= not((layer0_outputs(1541)) xor (layer0_outputs(1007)));
    layer1_outputs(1993) <= not(layer0_outputs(1115));
    layer1_outputs(1994) <= not(layer0_outputs(2318)) or (layer0_outputs(2156));
    layer1_outputs(1995) <= layer0_outputs(1469);
    layer1_outputs(1996) <= not(layer0_outputs(1954));
    layer1_outputs(1997) <= not((layer0_outputs(586)) xor (layer0_outputs(1099)));
    layer1_outputs(1998) <= '1';
    layer1_outputs(1999) <= not((layer0_outputs(2524)) and (layer0_outputs(1104)));
    layer1_outputs(2000) <= not(layer0_outputs(1225));
    layer1_outputs(2001) <= not(layer0_outputs(173)) or (layer0_outputs(2190));
    layer1_outputs(2002) <= not(layer0_outputs(236));
    layer1_outputs(2003) <= not(layer0_outputs(363)) or (layer0_outputs(518));
    layer1_outputs(2004) <= layer0_outputs(1515);
    layer1_outputs(2005) <= not(layer0_outputs(1822)) or (layer0_outputs(1728));
    layer1_outputs(2006) <= layer0_outputs(271);
    layer1_outputs(2007) <= '1';
    layer1_outputs(2008) <= '0';
    layer1_outputs(2009) <= not(layer0_outputs(817));
    layer1_outputs(2010) <= '0';
    layer1_outputs(2011) <= layer0_outputs(1702);
    layer1_outputs(2012) <= not((layer0_outputs(1200)) or (layer0_outputs(1416)));
    layer1_outputs(2013) <= not((layer0_outputs(1444)) or (layer0_outputs(1659)));
    layer1_outputs(2014) <= (layer0_outputs(493)) and not (layer0_outputs(1696));
    layer1_outputs(2015) <= not((layer0_outputs(243)) or (layer0_outputs(2325)));
    layer1_outputs(2016) <= '1';
    layer1_outputs(2017) <= not((layer0_outputs(32)) and (layer0_outputs(84)));
    layer1_outputs(2018) <= '0';
    layer1_outputs(2019) <= not(layer0_outputs(1796)) or (layer0_outputs(208));
    layer1_outputs(2020) <= not((layer0_outputs(1244)) or (layer0_outputs(1947)));
    layer1_outputs(2021) <= (layer0_outputs(201)) and not (layer0_outputs(323));
    layer1_outputs(2022) <= (layer0_outputs(206)) and not (layer0_outputs(1736));
    layer1_outputs(2023) <= layer0_outputs(1305);
    layer1_outputs(2024) <= (layer0_outputs(2294)) and not (layer0_outputs(2544));
    layer1_outputs(2025) <= not((layer0_outputs(2465)) and (layer0_outputs(2316)));
    layer1_outputs(2026) <= (layer0_outputs(2101)) and not (layer0_outputs(2372));
    layer1_outputs(2027) <= (layer0_outputs(2452)) and not (layer0_outputs(290));
    layer1_outputs(2028) <= not(layer0_outputs(2122)) or (layer0_outputs(1102));
    layer1_outputs(2029) <= '0';
    layer1_outputs(2030) <= not(layer0_outputs(1350));
    layer1_outputs(2031) <= (layer0_outputs(2160)) and not (layer0_outputs(1892));
    layer1_outputs(2032) <= (layer0_outputs(1536)) and not (layer0_outputs(581));
    layer1_outputs(2033) <= (layer0_outputs(2094)) and not (layer0_outputs(1248));
    layer1_outputs(2034) <= not(layer0_outputs(1381));
    layer1_outputs(2035) <= not(layer0_outputs(1229));
    layer1_outputs(2036) <= (layer0_outputs(1643)) and not (layer0_outputs(111));
    layer1_outputs(2037) <= not((layer0_outputs(2449)) and (layer0_outputs(2414)));
    layer1_outputs(2038) <= not((layer0_outputs(508)) or (layer0_outputs(623)));
    layer1_outputs(2039) <= (layer0_outputs(880)) and (layer0_outputs(2302));
    layer1_outputs(2040) <= not(layer0_outputs(903)) or (layer0_outputs(104));
    layer1_outputs(2041) <= '1';
    layer1_outputs(2042) <= (layer0_outputs(894)) and not (layer0_outputs(604));
    layer1_outputs(2043) <= layer0_outputs(754);
    layer1_outputs(2044) <= layer0_outputs(1407);
    layer1_outputs(2045) <= (layer0_outputs(990)) xor (layer0_outputs(1474));
    layer1_outputs(2046) <= not(layer0_outputs(1519));
    layer1_outputs(2047) <= (layer0_outputs(80)) and not (layer0_outputs(680));
    layer1_outputs(2048) <= '0';
    layer1_outputs(2049) <= (layer0_outputs(931)) and not (layer0_outputs(2299));
    layer1_outputs(2050) <= '1';
    layer1_outputs(2051) <= not(layer0_outputs(197));
    layer1_outputs(2052) <= layer0_outputs(270);
    layer1_outputs(2053) <= layer0_outputs(701);
    layer1_outputs(2054) <= not((layer0_outputs(876)) and (layer0_outputs(619)));
    layer1_outputs(2055) <= (layer0_outputs(470)) and (layer0_outputs(2076));
    layer1_outputs(2056) <= (layer0_outputs(154)) and not (layer0_outputs(309));
    layer1_outputs(2057) <= not(layer0_outputs(1958));
    layer1_outputs(2058) <= not(layer0_outputs(1316));
    layer1_outputs(2059) <= '1';
    layer1_outputs(2060) <= not(layer0_outputs(131));
    layer1_outputs(2061) <= not((layer0_outputs(2416)) or (layer0_outputs(342)));
    layer1_outputs(2062) <= not((layer0_outputs(2239)) and (layer0_outputs(620)));
    layer1_outputs(2063) <= layer0_outputs(1388);
    layer1_outputs(2064) <= (layer0_outputs(2537)) or (layer0_outputs(791));
    layer1_outputs(2065) <= (layer0_outputs(158)) and not (layer0_outputs(8));
    layer1_outputs(2066) <= not(layer0_outputs(994));
    layer1_outputs(2067) <= (layer0_outputs(767)) or (layer0_outputs(1288));
    layer1_outputs(2068) <= '0';
    layer1_outputs(2069) <= (layer0_outputs(1931)) or (layer0_outputs(2255));
    layer1_outputs(2070) <= layer0_outputs(17);
    layer1_outputs(2071) <= not(layer0_outputs(1689));
    layer1_outputs(2072) <= (layer0_outputs(1861)) and not (layer0_outputs(413));
    layer1_outputs(2073) <= not(layer0_outputs(1831));
    layer1_outputs(2074) <= layer0_outputs(1821);
    layer1_outputs(2075) <= not(layer0_outputs(1214)) or (layer0_outputs(1135));
    layer1_outputs(2076) <= not(layer0_outputs(1447));
    layer1_outputs(2077) <= (layer0_outputs(751)) or (layer0_outputs(1127));
    layer1_outputs(2078) <= '0';
    layer1_outputs(2079) <= (layer0_outputs(2232)) or (layer0_outputs(1607));
    layer1_outputs(2080) <= not((layer0_outputs(2056)) or (layer0_outputs(2551)));
    layer1_outputs(2081) <= not((layer0_outputs(1198)) and (layer0_outputs(980)));
    layer1_outputs(2082) <= (layer0_outputs(1382)) and not (layer0_outputs(1439));
    layer1_outputs(2083) <= layer0_outputs(535);
    layer1_outputs(2084) <= layer0_outputs(1107);
    layer1_outputs(2085) <= layer0_outputs(659);
    layer1_outputs(2086) <= not(layer0_outputs(1243));
    layer1_outputs(2087) <= not(layer0_outputs(2450)) or (layer0_outputs(64));
    layer1_outputs(2088) <= '0';
    layer1_outputs(2089) <= not(layer0_outputs(705)) or (layer0_outputs(799));
    layer1_outputs(2090) <= not(layer0_outputs(1412));
    layer1_outputs(2091) <= (layer0_outputs(1321)) and (layer0_outputs(2014));
    layer1_outputs(2092) <= not(layer0_outputs(186));
    layer1_outputs(2093) <= not(layer0_outputs(278));
    layer1_outputs(2094) <= (layer0_outputs(2264)) or (layer0_outputs(848));
    layer1_outputs(2095) <= '1';
    layer1_outputs(2096) <= (layer0_outputs(1060)) or (layer0_outputs(1119));
    layer1_outputs(2097) <= not((layer0_outputs(613)) and (layer0_outputs(1950)));
    layer1_outputs(2098) <= (layer0_outputs(1459)) or (layer0_outputs(2497));
    layer1_outputs(2099) <= '1';
    layer1_outputs(2100) <= (layer0_outputs(2214)) and not (layer0_outputs(1660));
    layer1_outputs(2101) <= not(layer0_outputs(158));
    layer1_outputs(2102) <= (layer0_outputs(1965)) and not (layer0_outputs(1610));
    layer1_outputs(2103) <= not(layer0_outputs(1687));
    layer1_outputs(2104) <= (layer0_outputs(1454)) and (layer0_outputs(2276));
    layer1_outputs(2105) <= not((layer0_outputs(480)) and (layer0_outputs(518)));
    layer1_outputs(2106) <= (layer0_outputs(139)) and not (layer0_outputs(971));
    layer1_outputs(2107) <= (layer0_outputs(2525)) and (layer0_outputs(734));
    layer1_outputs(2108) <= not(layer0_outputs(1602)) or (layer0_outputs(813));
    layer1_outputs(2109) <= layer0_outputs(2314);
    layer1_outputs(2110) <= not(layer0_outputs(724)) or (layer0_outputs(2258));
    layer1_outputs(2111) <= '0';
    layer1_outputs(2112) <= (layer0_outputs(1369)) and not (layer0_outputs(575));
    layer1_outputs(2113) <= not(layer0_outputs(2282)) or (layer0_outputs(1527));
    layer1_outputs(2114) <= (layer0_outputs(2220)) and not (layer0_outputs(2328));
    layer1_outputs(2115) <= not(layer0_outputs(1744)) or (layer0_outputs(229));
    layer1_outputs(2116) <= (layer0_outputs(2437)) and (layer0_outputs(1544));
    layer1_outputs(2117) <= layer0_outputs(922);
    layer1_outputs(2118) <= layer0_outputs(361);
    layer1_outputs(2119) <= not(layer0_outputs(2152)) or (layer0_outputs(1316));
    layer1_outputs(2120) <= layer0_outputs(1450);
    layer1_outputs(2121) <= '0';
    layer1_outputs(2122) <= (layer0_outputs(1632)) or (layer0_outputs(1908));
    layer1_outputs(2123) <= (layer0_outputs(584)) and (layer0_outputs(321));
    layer1_outputs(2124) <= layer0_outputs(475);
    layer1_outputs(2125) <= (layer0_outputs(1578)) and not (layer0_outputs(1763));
    layer1_outputs(2126) <= not(layer0_outputs(1988));
    layer1_outputs(2127) <= '0';
    layer1_outputs(2128) <= not(layer0_outputs(2075)) or (layer0_outputs(885));
    layer1_outputs(2129) <= layer0_outputs(1652);
    layer1_outputs(2130) <= not(layer0_outputs(1508)) or (layer0_outputs(1534));
    layer1_outputs(2131) <= not(layer0_outputs(927));
    layer1_outputs(2132) <= layer0_outputs(1933);
    layer1_outputs(2133) <= not(layer0_outputs(1254));
    layer1_outputs(2134) <= layer0_outputs(28);
    layer1_outputs(2135) <= '0';
    layer1_outputs(2136) <= not(layer0_outputs(1843));
    layer1_outputs(2137) <= (layer0_outputs(2173)) and not (layer0_outputs(1344));
    layer1_outputs(2138) <= layer0_outputs(2418);
    layer1_outputs(2139) <= '0';
    layer1_outputs(2140) <= not((layer0_outputs(1080)) or (layer0_outputs(134)));
    layer1_outputs(2141) <= not((layer0_outputs(1844)) xor (layer0_outputs(942)));
    layer1_outputs(2142) <= not(layer0_outputs(704));
    layer1_outputs(2143) <= (layer0_outputs(2429)) and not (layer0_outputs(1534));
    layer1_outputs(2144) <= layer0_outputs(2400);
    layer1_outputs(2145) <= layer0_outputs(769);
    layer1_outputs(2146) <= not(layer0_outputs(1241));
    layer1_outputs(2147) <= not(layer0_outputs(1659)) or (layer0_outputs(692));
    layer1_outputs(2148) <= layer0_outputs(1047);
    layer1_outputs(2149) <= (layer0_outputs(1292)) or (layer0_outputs(1120));
    layer1_outputs(2150) <= layer0_outputs(58);
    layer1_outputs(2151) <= (layer0_outputs(1285)) and not (layer0_outputs(668));
    layer1_outputs(2152) <= not(layer0_outputs(1307)) or (layer0_outputs(1575));
    layer1_outputs(2153) <= not(layer0_outputs(2485));
    layer1_outputs(2154) <= not(layer0_outputs(433)) or (layer0_outputs(1042));
    layer1_outputs(2155) <= not(layer0_outputs(737)) or (layer0_outputs(2247));
    layer1_outputs(2156) <= layer0_outputs(2290);
    layer1_outputs(2157) <= not(layer0_outputs(2257)) or (layer0_outputs(2108));
    layer1_outputs(2158) <= '1';
    layer1_outputs(2159) <= '0';
    layer1_outputs(2160) <= not((layer0_outputs(419)) and (layer0_outputs(2388)));
    layer1_outputs(2161) <= layer0_outputs(1420);
    layer1_outputs(2162) <= not((layer0_outputs(629)) xor (layer0_outputs(1479)));
    layer1_outputs(2163) <= not((layer0_outputs(460)) or (layer0_outputs(856)));
    layer1_outputs(2164) <= '1';
    layer1_outputs(2165) <= layer0_outputs(467);
    layer1_outputs(2166) <= not(layer0_outputs(1880)) or (layer0_outputs(2240));
    layer1_outputs(2167) <= '1';
    layer1_outputs(2168) <= not(layer0_outputs(1945));
    layer1_outputs(2169) <= not(layer0_outputs(1568));
    layer1_outputs(2170) <= (layer0_outputs(1947)) and not (layer0_outputs(2148));
    layer1_outputs(2171) <= (layer0_outputs(964)) and not (layer0_outputs(1914));
    layer1_outputs(2172) <= not(layer0_outputs(1858));
    layer1_outputs(2173) <= not((layer0_outputs(119)) and (layer0_outputs(2547)));
    layer1_outputs(2174) <= layer0_outputs(185);
    layer1_outputs(2175) <= (layer0_outputs(1337)) and (layer0_outputs(2378));
    layer1_outputs(2176) <= not(layer0_outputs(1816));
    layer1_outputs(2177) <= '0';
    layer1_outputs(2178) <= not(layer0_outputs(2230));
    layer1_outputs(2179) <= (layer0_outputs(1899)) and (layer0_outputs(2199));
    layer1_outputs(2180) <= not(layer0_outputs(2080)) or (layer0_outputs(214));
    layer1_outputs(2181) <= not(layer0_outputs(2522));
    layer1_outputs(2182) <= (layer0_outputs(765)) and not (layer0_outputs(1921));
    layer1_outputs(2183) <= (layer0_outputs(1996)) or (layer0_outputs(1752));
    layer1_outputs(2184) <= layer0_outputs(58);
    layer1_outputs(2185) <= '0';
    layer1_outputs(2186) <= (layer0_outputs(519)) and not (layer0_outputs(331));
    layer1_outputs(2187) <= '1';
    layer1_outputs(2188) <= not(layer0_outputs(1764)) or (layer0_outputs(1392));
    layer1_outputs(2189) <= not(layer0_outputs(1178)) or (layer0_outputs(2427));
    layer1_outputs(2190) <= layer0_outputs(2084);
    layer1_outputs(2191) <= not((layer0_outputs(1446)) and (layer0_outputs(1963)));
    layer1_outputs(2192) <= not(layer0_outputs(1487)) or (layer0_outputs(938));
    layer1_outputs(2193) <= not(layer0_outputs(1092));
    layer1_outputs(2194) <= '0';
    layer1_outputs(2195) <= (layer0_outputs(2038)) and not (layer0_outputs(1032));
    layer1_outputs(2196) <= not((layer0_outputs(1495)) or (layer0_outputs(323)));
    layer1_outputs(2197) <= (layer0_outputs(2501)) and not (layer0_outputs(103));
    layer1_outputs(2198) <= layer0_outputs(662);
    layer1_outputs(2199) <= (layer0_outputs(618)) and (layer0_outputs(2010));
    layer1_outputs(2200) <= (layer0_outputs(78)) and not (layer0_outputs(1167));
    layer1_outputs(2201) <= not(layer0_outputs(1973));
    layer1_outputs(2202) <= '0';
    layer1_outputs(2203) <= not(layer0_outputs(1583)) or (layer0_outputs(377));
    layer1_outputs(2204) <= (layer0_outputs(29)) or (layer0_outputs(1761));
    layer1_outputs(2205) <= (layer0_outputs(1123)) and not (layer0_outputs(2531));
    layer1_outputs(2206) <= (layer0_outputs(1508)) and not (layer0_outputs(276));
    layer1_outputs(2207) <= (layer0_outputs(1416)) or (layer0_outputs(759));
    layer1_outputs(2208) <= not((layer0_outputs(1212)) xor (layer0_outputs(1538)));
    layer1_outputs(2209) <= not(layer0_outputs(2311)) or (layer0_outputs(1727));
    layer1_outputs(2210) <= (layer0_outputs(2555)) and (layer0_outputs(2042));
    layer1_outputs(2211) <= layer0_outputs(1349);
    layer1_outputs(2212) <= not((layer0_outputs(2305)) or (layer0_outputs(454)));
    layer1_outputs(2213) <= (layer0_outputs(491)) or (layer0_outputs(483));
    layer1_outputs(2214) <= not(layer0_outputs(2010));
    layer1_outputs(2215) <= layer0_outputs(1928);
    layer1_outputs(2216) <= not(layer0_outputs(143)) or (layer0_outputs(545));
    layer1_outputs(2217) <= (layer0_outputs(1213)) and not (layer0_outputs(338));
    layer1_outputs(2218) <= '0';
    layer1_outputs(2219) <= not(layer0_outputs(374)) or (layer0_outputs(1183));
    layer1_outputs(2220) <= (layer0_outputs(1838)) and not (layer0_outputs(1932));
    layer1_outputs(2221) <= '0';
    layer1_outputs(2222) <= not((layer0_outputs(1576)) or (layer0_outputs(1612)));
    layer1_outputs(2223) <= not(layer0_outputs(2420)) or (layer0_outputs(25));
    layer1_outputs(2224) <= '0';
    layer1_outputs(2225) <= layer0_outputs(2072);
    layer1_outputs(2226) <= layer0_outputs(2325);
    layer1_outputs(2227) <= layer0_outputs(1488);
    layer1_outputs(2228) <= not(layer0_outputs(2309));
    layer1_outputs(2229) <= (layer0_outputs(1671)) and not (layer0_outputs(744));
    layer1_outputs(2230) <= layer0_outputs(660);
    layer1_outputs(2231) <= not(layer0_outputs(964));
    layer1_outputs(2232) <= not(layer0_outputs(1283));
    layer1_outputs(2233) <= not(layer0_outputs(151)) or (layer0_outputs(1960));
    layer1_outputs(2234) <= not(layer0_outputs(1587));
    layer1_outputs(2235) <= not(layer0_outputs(400));
    layer1_outputs(2236) <= (layer0_outputs(312)) and not (layer0_outputs(936));
    layer1_outputs(2237) <= (layer0_outputs(624)) or (layer0_outputs(1845));
    layer1_outputs(2238) <= not(layer0_outputs(1675));
    layer1_outputs(2239) <= '0';
    layer1_outputs(2240) <= (layer0_outputs(2376)) or (layer0_outputs(929));
    layer1_outputs(2241) <= layer0_outputs(1719);
    layer1_outputs(2242) <= not(layer0_outputs(1109)) or (layer0_outputs(641));
    layer1_outputs(2243) <= not((layer0_outputs(1548)) and (layer0_outputs(1477)));
    layer1_outputs(2244) <= '0';
    layer1_outputs(2245) <= not(layer0_outputs(2396)) or (layer0_outputs(862));
    layer1_outputs(2246) <= (layer0_outputs(193)) and not (layer0_outputs(750));
    layer1_outputs(2247) <= layer0_outputs(1938);
    layer1_outputs(2248) <= (layer0_outputs(1295)) or (layer0_outputs(2198));
    layer1_outputs(2249) <= '1';
    layer1_outputs(2250) <= not((layer0_outputs(1997)) and (layer0_outputs(92)));
    layer1_outputs(2251) <= layer0_outputs(1338);
    layer1_outputs(2252) <= (layer0_outputs(1629)) and not (layer0_outputs(1704));
    layer1_outputs(2253) <= (layer0_outputs(1837)) and not (layer0_outputs(2365));
    layer1_outputs(2254) <= not((layer0_outputs(1790)) and (layer0_outputs(848)));
    layer1_outputs(2255) <= (layer0_outputs(1832)) and (layer0_outputs(1582));
    layer1_outputs(2256) <= not(layer0_outputs(680)) or (layer0_outputs(1499));
    layer1_outputs(2257) <= not((layer0_outputs(671)) or (layer0_outputs(1185)));
    layer1_outputs(2258) <= not(layer0_outputs(1189)) or (layer0_outputs(183));
    layer1_outputs(2259) <= '1';
    layer1_outputs(2260) <= not(layer0_outputs(1701));
    layer1_outputs(2261) <= (layer0_outputs(1749)) and not (layer0_outputs(107));
    layer1_outputs(2262) <= not(layer0_outputs(2195));
    layer1_outputs(2263) <= not(layer0_outputs(576)) or (layer0_outputs(178));
    layer1_outputs(2264) <= '1';
    layer1_outputs(2265) <= not(layer0_outputs(1372));
    layer1_outputs(2266) <= '0';
    layer1_outputs(2267) <= (layer0_outputs(94)) or (layer0_outputs(2323));
    layer1_outputs(2268) <= layer0_outputs(1284);
    layer1_outputs(2269) <= (layer0_outputs(1475)) and not (layer0_outputs(733));
    layer1_outputs(2270) <= not(layer0_outputs(1268));
    layer1_outputs(2271) <= (layer0_outputs(600)) and not (layer0_outputs(1672));
    layer1_outputs(2272) <= not(layer0_outputs(1512));
    layer1_outputs(2273) <= '0';
    layer1_outputs(2274) <= not((layer0_outputs(1606)) or (layer0_outputs(989)));
    layer1_outputs(2275) <= not(layer0_outputs(2398));
    layer1_outputs(2276) <= not(layer0_outputs(201));
    layer1_outputs(2277) <= layer0_outputs(1922);
    layer1_outputs(2278) <= not(layer0_outputs(892));
    layer1_outputs(2279) <= not(layer0_outputs(2269));
    layer1_outputs(2280) <= not(layer0_outputs(2034));
    layer1_outputs(2281) <= layer0_outputs(970);
    layer1_outputs(2282) <= '1';
    layer1_outputs(2283) <= not(layer0_outputs(623));
    layer1_outputs(2284) <= (layer0_outputs(2020)) and not (layer0_outputs(2246));
    layer1_outputs(2285) <= not((layer0_outputs(1777)) and (layer0_outputs(1341)));
    layer1_outputs(2286) <= '1';
    layer1_outputs(2287) <= '0';
    layer1_outputs(2288) <= (layer0_outputs(442)) and (layer0_outputs(2430));
    layer1_outputs(2289) <= layer0_outputs(2483);
    layer1_outputs(2290) <= '0';
    layer1_outputs(2291) <= (layer0_outputs(213)) and not (layer0_outputs(329));
    layer1_outputs(2292) <= not(layer0_outputs(1414)) or (layer0_outputs(217));
    layer1_outputs(2293) <= layer0_outputs(256);
    layer1_outputs(2294) <= layer0_outputs(1818);
    layer1_outputs(2295) <= (layer0_outputs(2049)) and not (layer0_outputs(2128));
    layer1_outputs(2296) <= layer0_outputs(1170);
    layer1_outputs(2297) <= layer0_outputs(1051);
    layer1_outputs(2298) <= (layer0_outputs(225)) and (layer0_outputs(2032));
    layer1_outputs(2299) <= not((layer0_outputs(689)) or (layer0_outputs(62)));
    layer1_outputs(2300) <= '0';
    layer1_outputs(2301) <= (layer0_outputs(2144)) and not (layer0_outputs(1005));
    layer1_outputs(2302) <= (layer0_outputs(913)) or (layer0_outputs(1839));
    layer1_outputs(2303) <= (layer0_outputs(406)) and not (layer0_outputs(1245));
    layer1_outputs(2304) <= not(layer0_outputs(1253)) or (layer0_outputs(2151));
    layer1_outputs(2305) <= not(layer0_outputs(437)) or (layer0_outputs(187));
    layer1_outputs(2306) <= not(layer0_outputs(725));
    layer1_outputs(2307) <= not(layer0_outputs(706)) or (layer0_outputs(795));
    layer1_outputs(2308) <= (layer0_outputs(245)) and (layer0_outputs(260));
    layer1_outputs(2309) <= not(layer0_outputs(2213));
    layer1_outputs(2310) <= not((layer0_outputs(2111)) and (layer0_outputs(1472)));
    layer1_outputs(2311) <= not(layer0_outputs(1410));
    layer1_outputs(2312) <= layer0_outputs(640);
    layer1_outputs(2313) <= layer0_outputs(2172);
    layer1_outputs(2314) <= (layer0_outputs(2428)) and not (layer0_outputs(1014));
    layer1_outputs(2315) <= (layer0_outputs(1318)) and (layer0_outputs(2397));
    layer1_outputs(2316) <= not((layer0_outputs(2545)) xor (layer0_outputs(1240)));
    layer1_outputs(2317) <= not((layer0_outputs(2483)) or (layer0_outputs(1317)));
    layer1_outputs(2318) <= (layer0_outputs(1823)) and not (layer0_outputs(2000));
    layer1_outputs(2319) <= not(layer0_outputs(1027));
    layer1_outputs(2320) <= not(layer0_outputs(240));
    layer1_outputs(2321) <= layer0_outputs(1788);
    layer1_outputs(2322) <= not((layer0_outputs(1663)) and (layer0_outputs(378)));
    layer1_outputs(2323) <= (layer0_outputs(1649)) or (layer0_outputs(667));
    layer1_outputs(2324) <= layer0_outputs(1796);
    layer1_outputs(2325) <= (layer0_outputs(952)) and not (layer0_outputs(1720));
    layer1_outputs(2326) <= (layer0_outputs(438)) and (layer0_outputs(1870));
    layer1_outputs(2327) <= not(layer0_outputs(218)) or (layer0_outputs(2161));
    layer1_outputs(2328) <= layer0_outputs(2097);
    layer1_outputs(2329) <= not(layer0_outputs(2394));
    layer1_outputs(2330) <= (layer0_outputs(568)) and not (layer0_outputs(1221));
    layer1_outputs(2331) <= not((layer0_outputs(562)) or (layer0_outputs(2163)));
    layer1_outputs(2332) <= layer0_outputs(995);
    layer1_outputs(2333) <= not((layer0_outputs(523)) xor (layer0_outputs(1748)));
    layer1_outputs(2334) <= not((layer0_outputs(1130)) or (layer0_outputs(392)));
    layer1_outputs(2335) <= not(layer0_outputs(2252));
    layer1_outputs(2336) <= (layer0_outputs(2512)) and not (layer0_outputs(2422));
    layer1_outputs(2337) <= '1';
    layer1_outputs(2338) <= not((layer0_outputs(537)) and (layer0_outputs(1657)));
    layer1_outputs(2339) <= (layer0_outputs(1342)) or (layer0_outputs(2004));
    layer1_outputs(2340) <= '0';
    layer1_outputs(2341) <= not(layer0_outputs(254));
    layer1_outputs(2342) <= '1';
    layer1_outputs(2343) <= not(layer0_outputs(1205)) or (layer0_outputs(2340));
    layer1_outputs(2344) <= (layer0_outputs(785)) and (layer0_outputs(231));
    layer1_outputs(2345) <= not((layer0_outputs(639)) and (layer0_outputs(2279)));
    layer1_outputs(2346) <= not(layer0_outputs(1));
    layer1_outputs(2347) <= '1';
    layer1_outputs(2348) <= not((layer0_outputs(755)) and (layer0_outputs(1858)));
    layer1_outputs(2349) <= not(layer0_outputs(564));
    layer1_outputs(2350) <= not((layer0_outputs(1586)) and (layer0_outputs(974)));
    layer1_outputs(2351) <= '1';
    layer1_outputs(2352) <= (layer0_outputs(1169)) and not (layer0_outputs(97));
    layer1_outputs(2353) <= layer0_outputs(396);
    layer1_outputs(2354) <= not((layer0_outputs(1441)) and (layer0_outputs(1942)));
    layer1_outputs(2355) <= layer0_outputs(2403);
    layer1_outputs(2356) <= layer0_outputs(2409);
    layer1_outputs(2357) <= not(layer0_outputs(1132));
    layer1_outputs(2358) <= '0';
    layer1_outputs(2359) <= layer0_outputs(1732);
    layer1_outputs(2360) <= not((layer0_outputs(1621)) and (layer0_outputs(2262)));
    layer1_outputs(2361) <= (layer0_outputs(363)) and not (layer0_outputs(1283));
    layer1_outputs(2362) <= (layer0_outputs(2383)) and not (layer0_outputs(2077));
    layer1_outputs(2363) <= not(layer0_outputs(2169)) or (layer0_outputs(1360));
    layer1_outputs(2364) <= layer0_outputs(2146);
    layer1_outputs(2365) <= '1';
    layer1_outputs(2366) <= '0';
    layer1_outputs(2367) <= '0';
    layer1_outputs(2368) <= (layer0_outputs(2030)) and not (layer0_outputs(2420));
    layer1_outputs(2369) <= not(layer0_outputs(750));
    layer1_outputs(2370) <= not((layer0_outputs(1312)) and (layer0_outputs(697)));
    layer1_outputs(2371) <= not((layer0_outputs(673)) and (layer0_outputs(235)));
    layer1_outputs(2372) <= (layer0_outputs(887)) and (layer0_outputs(2478));
    layer1_outputs(2373) <= (layer0_outputs(1601)) and not (layer0_outputs(1350));
    layer1_outputs(2374) <= (layer0_outputs(2153)) and not (layer0_outputs(1048));
    layer1_outputs(2375) <= not((layer0_outputs(1930)) and (layer0_outputs(1098)));
    layer1_outputs(2376) <= not(layer0_outputs(1810)) or (layer0_outputs(354));
    layer1_outputs(2377) <= (layer0_outputs(769)) or (layer0_outputs(632));
    layer1_outputs(2378) <= not(layer0_outputs(66)) or (layer0_outputs(101));
    layer1_outputs(2379) <= '1';
    layer1_outputs(2380) <= layer0_outputs(443);
    layer1_outputs(2381) <= layer0_outputs(2379);
    layer1_outputs(2382) <= '1';
    layer1_outputs(2383) <= not((layer0_outputs(161)) and (layer0_outputs(2407)));
    layer1_outputs(2384) <= not((layer0_outputs(932)) and (layer0_outputs(627)));
    layer1_outputs(2385) <= not(layer0_outputs(1497)) or (layer0_outputs(2215));
    layer1_outputs(2386) <= not((layer0_outputs(256)) or (layer0_outputs(1028)));
    layer1_outputs(2387) <= layer0_outputs(2464);
    layer1_outputs(2388) <= not((layer0_outputs(1112)) or (layer0_outputs(2520)));
    layer1_outputs(2389) <= not((layer0_outputs(1868)) and (layer0_outputs(1219)));
    layer1_outputs(2390) <= (layer0_outputs(2029)) or (layer0_outputs(318));
    layer1_outputs(2391) <= layer0_outputs(1753);
    layer1_outputs(2392) <= '1';
    layer1_outputs(2393) <= layer0_outputs(2193);
    layer1_outputs(2394) <= not(layer0_outputs(855));
    layer1_outputs(2395) <= '1';
    layer1_outputs(2396) <= layer0_outputs(1059);
    layer1_outputs(2397) <= not(layer0_outputs(473));
    layer1_outputs(2398) <= '0';
    layer1_outputs(2399) <= (layer0_outputs(15)) and not (layer0_outputs(135));
    layer1_outputs(2400) <= not(layer0_outputs(1711)) or (layer0_outputs(196));
    layer1_outputs(2401) <= layer0_outputs(1222);
    layer1_outputs(2402) <= (layer0_outputs(2508)) and not (layer0_outputs(1016));
    layer1_outputs(2403) <= (layer0_outputs(867)) and (layer0_outputs(998));
    layer1_outputs(2404) <= layer0_outputs(2023);
    layer1_outputs(2405) <= not(layer0_outputs(2531));
    layer1_outputs(2406) <= '0';
    layer1_outputs(2407) <= layer0_outputs(1789);
    layer1_outputs(2408) <= not((layer0_outputs(1760)) and (layer0_outputs(2200)));
    layer1_outputs(2409) <= layer0_outputs(225);
    layer1_outputs(2410) <= layer0_outputs(1817);
    layer1_outputs(2411) <= not((layer0_outputs(2334)) and (layer0_outputs(177)));
    layer1_outputs(2412) <= '0';
    layer1_outputs(2413) <= (layer0_outputs(2100)) and not (layer0_outputs(2021));
    layer1_outputs(2414) <= layer0_outputs(1767);
    layer1_outputs(2415) <= (layer0_outputs(288)) or (layer0_outputs(897));
    layer1_outputs(2416) <= layer0_outputs(1802);
    layer1_outputs(2417) <= not((layer0_outputs(97)) or (layer0_outputs(1981)));
    layer1_outputs(2418) <= (layer0_outputs(1765)) or (layer0_outputs(2071));
    layer1_outputs(2419) <= not(layer0_outputs(259)) or (layer0_outputs(1912));
    layer1_outputs(2420) <= not((layer0_outputs(1454)) and (layer0_outputs(2435)));
    layer1_outputs(2421) <= '1';
    layer1_outputs(2422) <= (layer0_outputs(831)) and not (layer0_outputs(1989));
    layer1_outputs(2423) <= not(layer0_outputs(986));
    layer1_outputs(2424) <= (layer0_outputs(412)) and not (layer0_outputs(767));
    layer1_outputs(2425) <= layer0_outputs(1391);
    layer1_outputs(2426) <= not(layer0_outputs(1780));
    layer1_outputs(2427) <= not(layer0_outputs(2535)) or (layer0_outputs(1937));
    layer1_outputs(2428) <= layer0_outputs(48);
    layer1_outputs(2429) <= (layer0_outputs(514)) or (layer0_outputs(2456));
    layer1_outputs(2430) <= (layer0_outputs(1140)) and (layer0_outputs(1761));
    layer1_outputs(2431) <= not(layer0_outputs(1374));
    layer1_outputs(2432) <= not(layer0_outputs(281));
    layer1_outputs(2433) <= (layer0_outputs(295)) or (layer0_outputs(2349));
    layer1_outputs(2434) <= '1';
    layer1_outputs(2435) <= '0';
    layer1_outputs(2436) <= (layer0_outputs(709)) and (layer0_outputs(455));
    layer1_outputs(2437) <= layer0_outputs(1393);
    layer1_outputs(2438) <= (layer0_outputs(589)) and not (layer0_outputs(184));
    layer1_outputs(2439) <= layer0_outputs(400);
    layer1_outputs(2440) <= '1';
    layer1_outputs(2441) <= (layer0_outputs(2463)) and (layer0_outputs(2311));
    layer1_outputs(2442) <= layer0_outputs(506);
    layer1_outputs(2443) <= not(layer0_outputs(988));
    layer1_outputs(2444) <= not(layer0_outputs(1150));
    layer1_outputs(2445) <= not(layer0_outputs(1972)) or (layer0_outputs(981));
    layer1_outputs(2446) <= layer0_outputs(628);
    layer1_outputs(2447) <= (layer0_outputs(2380)) and (layer0_outputs(739));
    layer1_outputs(2448) <= (layer0_outputs(1331)) and not (layer0_outputs(2413));
    layer1_outputs(2449) <= not(layer0_outputs(2333));
    layer1_outputs(2450) <= not(layer0_outputs(5));
    layer1_outputs(2451) <= (layer0_outputs(1862)) or (layer0_outputs(1298));
    layer1_outputs(2452) <= not(layer0_outputs(2227));
    layer1_outputs(2453) <= not(layer0_outputs(2074)) or (layer0_outputs(17));
    layer1_outputs(2454) <= layer0_outputs(550);
    layer1_outputs(2455) <= '0';
    layer1_outputs(2456) <= (layer0_outputs(1176)) and not (layer0_outputs(2320));
    layer1_outputs(2457) <= '1';
    layer1_outputs(2458) <= (layer0_outputs(1587)) and not (layer0_outputs(339));
    layer1_outputs(2459) <= '1';
    layer1_outputs(2460) <= '1';
    layer1_outputs(2461) <= '0';
    layer1_outputs(2462) <= (layer0_outputs(236)) or (layer0_outputs(639));
    layer1_outputs(2463) <= not(layer0_outputs(2367));
    layer1_outputs(2464) <= '0';
    layer1_outputs(2465) <= not((layer0_outputs(2451)) and (layer0_outputs(1826)));
    layer1_outputs(2466) <= not(layer0_outputs(1524));
    layer1_outputs(2467) <= (layer0_outputs(2275)) and not (layer0_outputs(1332));
    layer1_outputs(2468) <= (layer0_outputs(1721)) and not (layer0_outputs(1722));
    layer1_outputs(2469) <= (layer0_outputs(123)) and (layer0_outputs(2296));
    layer1_outputs(2470) <= not(layer0_outputs(914)) or (layer0_outputs(250));
    layer1_outputs(2471) <= (layer0_outputs(155)) or (layer0_outputs(1553));
    layer1_outputs(2472) <= (layer0_outputs(1137)) and not (layer0_outputs(2352));
    layer1_outputs(2473) <= layer0_outputs(1181);
    layer1_outputs(2474) <= (layer0_outputs(62)) or (layer0_outputs(541));
    layer1_outputs(2475) <= layer0_outputs(1202);
    layer1_outputs(2476) <= not((layer0_outputs(2113)) or (layer0_outputs(301)));
    layer1_outputs(2477) <= layer0_outputs(352);
    layer1_outputs(2478) <= (layer0_outputs(1622)) and not (layer0_outputs(142));
    layer1_outputs(2479) <= not((layer0_outputs(1616)) xor (layer0_outputs(682)));
    layer1_outputs(2480) <= (layer0_outputs(1343)) or (layer0_outputs(1851));
    layer1_outputs(2481) <= (layer0_outputs(2277)) and not (layer0_outputs(1870));
    layer1_outputs(2482) <= not((layer0_outputs(1529)) xor (layer0_outputs(1134)));
    layer1_outputs(2483) <= not(layer0_outputs(1850));
    layer1_outputs(2484) <= not(layer0_outputs(415)) or (layer0_outputs(508));
    layer1_outputs(2485) <= layer0_outputs(809);
    layer1_outputs(2486) <= not((layer0_outputs(2381)) xor (layer0_outputs(532)));
    layer1_outputs(2487) <= layer0_outputs(2265);
    layer1_outputs(2488) <= '0';
    layer1_outputs(2489) <= not(layer0_outputs(1647));
    layer1_outputs(2490) <= not((layer0_outputs(2477)) or (layer0_outputs(397)));
    layer1_outputs(2491) <= not(layer0_outputs(833)) or (layer0_outputs(2229));
    layer1_outputs(2492) <= (layer0_outputs(401)) and (layer0_outputs(922));
    layer1_outputs(2493) <= (layer0_outputs(426)) and not (layer0_outputs(68));
    layer1_outputs(2494) <= not(layer0_outputs(1979)) or (layer0_outputs(1853));
    layer1_outputs(2495) <= '1';
    layer1_outputs(2496) <= (layer0_outputs(2288)) and not (layer0_outputs(802));
    layer1_outputs(2497) <= not(layer0_outputs(1383)) or (layer0_outputs(1771));
    layer1_outputs(2498) <= not(layer0_outputs(2127));
    layer1_outputs(2499) <= (layer0_outputs(565)) or (layer0_outputs(1909));
    layer1_outputs(2500) <= layer0_outputs(463);
    layer1_outputs(2501) <= not((layer0_outputs(1062)) and (layer0_outputs(1153)));
    layer1_outputs(2502) <= (layer0_outputs(1284)) or (layer0_outputs(251));
    layer1_outputs(2503) <= (layer0_outputs(2410)) and (layer0_outputs(1218));
    layer1_outputs(2504) <= layer0_outputs(21);
    layer1_outputs(2505) <= (layer0_outputs(56)) or (layer0_outputs(1718));
    layer1_outputs(2506) <= (layer0_outputs(2252)) and not (layer0_outputs(929));
    layer1_outputs(2507) <= '1';
    layer1_outputs(2508) <= '1';
    layer1_outputs(2509) <= not(layer0_outputs(1866)) or (layer0_outputs(1636));
    layer1_outputs(2510) <= (layer0_outputs(487)) and not (layer0_outputs(306));
    layer1_outputs(2511) <= (layer0_outputs(1180)) xor (layer0_outputs(1607));
    layer1_outputs(2512) <= (layer0_outputs(1396)) and (layer0_outputs(670));
    layer1_outputs(2513) <= layer0_outputs(643);
    layer1_outputs(2514) <= (layer0_outputs(1308)) xor (layer0_outputs(1720));
    layer1_outputs(2515) <= not(layer0_outputs(1613)) or (layer0_outputs(1169));
    layer1_outputs(2516) <= '1';
    layer1_outputs(2517) <= (layer0_outputs(1054)) and (layer0_outputs(2527));
    layer1_outputs(2518) <= not(layer0_outputs(917));
    layer1_outputs(2519) <= not(layer0_outputs(261));
    layer1_outputs(2520) <= (layer0_outputs(1311)) and (layer0_outputs(730));
    layer1_outputs(2521) <= '0';
    layer1_outputs(2522) <= not(layer0_outputs(776)) or (layer0_outputs(480));
    layer1_outputs(2523) <= (layer0_outputs(1531)) and not (layer0_outputs(1371));
    layer1_outputs(2524) <= not(layer0_outputs(2226));
    layer1_outputs(2525) <= not((layer0_outputs(2086)) or (layer0_outputs(1216)));
    layer1_outputs(2526) <= '0';
    layer1_outputs(2527) <= (layer0_outputs(1776)) and not (layer0_outputs(1389));
    layer1_outputs(2528) <= '0';
    layer1_outputs(2529) <= (layer0_outputs(109)) or (layer0_outputs(56));
    layer1_outputs(2530) <= '0';
    layer1_outputs(2531) <= (layer0_outputs(1046)) or (layer0_outputs(2174));
    layer1_outputs(2532) <= '1';
    layer1_outputs(2533) <= not(layer0_outputs(1177));
    layer1_outputs(2534) <= layer0_outputs(1937);
    layer1_outputs(2535) <= layer0_outputs(1964);
    layer1_outputs(2536) <= '0';
    layer1_outputs(2537) <= (layer0_outputs(2221)) and (layer0_outputs(436));
    layer1_outputs(2538) <= '0';
    layer1_outputs(2539) <= layer0_outputs(759);
    layer1_outputs(2540) <= not(layer0_outputs(1424)) or (layer0_outputs(1160));
    layer1_outputs(2541) <= (layer0_outputs(1476)) and not (layer0_outputs(1754));
    layer1_outputs(2542) <= (layer0_outputs(441)) and not (layer0_outputs(1208));
    layer1_outputs(2543) <= not(layer0_outputs(1711));
    layer1_outputs(2544) <= (layer0_outputs(1257)) and not (layer0_outputs(738));
    layer1_outputs(2545) <= (layer0_outputs(282)) and not (layer0_outputs(1102));
    layer1_outputs(2546) <= not(layer0_outputs(1194));
    layer1_outputs(2547) <= layer0_outputs(1747);
    layer1_outputs(2548) <= '1';
    layer1_outputs(2549) <= not(layer0_outputs(2321));
    layer1_outputs(2550) <= not(layer0_outputs(180));
    layer1_outputs(2551) <= (layer0_outputs(2332)) and not (layer0_outputs(838));
    layer1_outputs(2552) <= '1';
    layer1_outputs(2553) <= '0';
    layer1_outputs(2554) <= not(layer0_outputs(1355));
    layer1_outputs(2555) <= '1';
    layer1_outputs(2556) <= '0';
    layer1_outputs(2557) <= (layer0_outputs(2178)) or (layer0_outputs(1624));
    layer1_outputs(2558) <= '0';
    layer1_outputs(2559) <= (layer0_outputs(69)) and (layer0_outputs(113));
    layer2_outputs(0) <= '0';
    layer2_outputs(1) <= '1';
    layer2_outputs(2) <= (layer1_outputs(1821)) and not (layer1_outputs(1842));
    layer2_outputs(3) <= (layer1_outputs(570)) xor (layer1_outputs(1298));
    layer2_outputs(4) <= layer1_outputs(1774);
    layer2_outputs(5) <= not(layer1_outputs(2326));
    layer2_outputs(6) <= (layer1_outputs(1397)) and not (layer1_outputs(499));
    layer2_outputs(7) <= not(layer1_outputs(579)) or (layer1_outputs(115));
    layer2_outputs(8) <= layer1_outputs(1250);
    layer2_outputs(9) <= not((layer1_outputs(1466)) or (layer1_outputs(2083)));
    layer2_outputs(10) <= (layer1_outputs(1698)) and not (layer1_outputs(1859));
    layer2_outputs(11) <= layer1_outputs(1721);
    layer2_outputs(12) <= (layer1_outputs(1498)) or (layer1_outputs(222));
    layer2_outputs(13) <= layer1_outputs(237);
    layer2_outputs(14) <= (layer1_outputs(2507)) and (layer1_outputs(1609));
    layer2_outputs(15) <= layer1_outputs(2084);
    layer2_outputs(16) <= not(layer1_outputs(864)) or (layer1_outputs(131));
    layer2_outputs(17) <= not(layer1_outputs(1817)) or (layer1_outputs(1418));
    layer2_outputs(18) <= layer1_outputs(167);
    layer2_outputs(19) <= not((layer1_outputs(2519)) or (layer1_outputs(1321)));
    layer2_outputs(20) <= not(layer1_outputs(1825));
    layer2_outputs(21) <= not(layer1_outputs(1601)) or (layer1_outputs(1057));
    layer2_outputs(22) <= not(layer1_outputs(2186)) or (layer1_outputs(1858));
    layer2_outputs(23) <= layer1_outputs(676);
    layer2_outputs(24) <= not(layer1_outputs(1897));
    layer2_outputs(25) <= layer1_outputs(885);
    layer2_outputs(26) <= not(layer1_outputs(1019)) or (layer1_outputs(2302));
    layer2_outputs(27) <= not(layer1_outputs(2221)) or (layer1_outputs(612));
    layer2_outputs(28) <= not((layer1_outputs(782)) and (layer1_outputs(663)));
    layer2_outputs(29) <= (layer1_outputs(1989)) and not (layer1_outputs(350));
    layer2_outputs(30) <= not(layer1_outputs(1043));
    layer2_outputs(31) <= (layer1_outputs(2053)) or (layer1_outputs(2261));
    layer2_outputs(32) <= '1';
    layer2_outputs(33) <= not(layer1_outputs(2449));
    layer2_outputs(34) <= not(layer1_outputs(887));
    layer2_outputs(35) <= '0';
    layer2_outputs(36) <= not(layer1_outputs(313));
    layer2_outputs(37) <= not((layer1_outputs(2164)) or (layer1_outputs(40)));
    layer2_outputs(38) <= layer1_outputs(2009);
    layer2_outputs(39) <= layer1_outputs(1084);
    layer2_outputs(40) <= (layer1_outputs(1836)) or (layer1_outputs(358));
    layer2_outputs(41) <= '0';
    layer2_outputs(42) <= layer1_outputs(2381);
    layer2_outputs(43) <= not(layer1_outputs(1831)) or (layer1_outputs(553));
    layer2_outputs(44) <= not(layer1_outputs(2031));
    layer2_outputs(45) <= (layer1_outputs(374)) and not (layer1_outputs(1933));
    layer2_outputs(46) <= not((layer1_outputs(650)) or (layer1_outputs(2378)));
    layer2_outputs(47) <= '1';
    layer2_outputs(48) <= not((layer1_outputs(1193)) and (layer1_outputs(1227)));
    layer2_outputs(49) <= layer1_outputs(1919);
    layer2_outputs(50) <= layer1_outputs(198);
    layer2_outputs(51) <= layer1_outputs(789);
    layer2_outputs(52) <= (layer1_outputs(1036)) and not (layer1_outputs(143));
    layer2_outputs(53) <= '1';
    layer2_outputs(54) <= layer1_outputs(91);
    layer2_outputs(55) <= layer1_outputs(884);
    layer2_outputs(56) <= not(layer1_outputs(1951));
    layer2_outputs(57) <= not(layer1_outputs(2041)) or (layer1_outputs(975));
    layer2_outputs(58) <= '1';
    layer2_outputs(59) <= not(layer1_outputs(1710));
    layer2_outputs(60) <= not(layer1_outputs(1041));
    layer2_outputs(61) <= (layer1_outputs(468)) and not (layer1_outputs(1373));
    layer2_outputs(62) <= not((layer1_outputs(254)) or (layer1_outputs(246)));
    layer2_outputs(63) <= layer1_outputs(1433);
    layer2_outputs(64) <= not(layer1_outputs(1719));
    layer2_outputs(65) <= '1';
    layer2_outputs(66) <= layer1_outputs(2293);
    layer2_outputs(67) <= not(layer1_outputs(2201));
    layer2_outputs(68) <= not(layer1_outputs(1362));
    layer2_outputs(69) <= '1';
    layer2_outputs(70) <= not((layer1_outputs(1291)) or (layer1_outputs(1126)));
    layer2_outputs(71) <= not(layer1_outputs(890)) or (layer1_outputs(2315));
    layer2_outputs(72) <= not(layer1_outputs(2062)) or (layer1_outputs(1946));
    layer2_outputs(73) <= not(layer1_outputs(797));
    layer2_outputs(74) <= '1';
    layer2_outputs(75) <= (layer1_outputs(2060)) and (layer1_outputs(1459));
    layer2_outputs(76) <= '0';
    layer2_outputs(77) <= not((layer1_outputs(1451)) and (layer1_outputs(1361)));
    layer2_outputs(78) <= '1';
    layer2_outputs(79) <= '1';
    layer2_outputs(80) <= not(layer1_outputs(1545));
    layer2_outputs(81) <= (layer1_outputs(1253)) and not (layer1_outputs(312));
    layer2_outputs(82) <= not((layer1_outputs(961)) or (layer1_outputs(2206)));
    layer2_outputs(83) <= not(layer1_outputs(2235)) or (layer1_outputs(1522));
    layer2_outputs(84) <= not(layer1_outputs(245));
    layer2_outputs(85) <= not((layer1_outputs(2343)) and (layer1_outputs(188)));
    layer2_outputs(86) <= not(layer1_outputs(472)) or (layer1_outputs(849));
    layer2_outputs(87) <= not(layer1_outputs(1640)) or (layer1_outputs(1980));
    layer2_outputs(88) <= not(layer1_outputs(385));
    layer2_outputs(89) <= layer1_outputs(1650);
    layer2_outputs(90) <= layer1_outputs(1138);
    layer2_outputs(91) <= not(layer1_outputs(17)) or (layer1_outputs(2020));
    layer2_outputs(92) <= layer1_outputs(1581);
    layer2_outputs(93) <= (layer1_outputs(1344)) or (layer1_outputs(1818));
    layer2_outputs(94) <= not((layer1_outputs(1173)) and (layer1_outputs(1646)));
    layer2_outputs(95) <= not((layer1_outputs(2338)) xor (layer1_outputs(333)));
    layer2_outputs(96) <= not(layer1_outputs(1979));
    layer2_outputs(97) <= not(layer1_outputs(1333)) or (layer1_outputs(2017));
    layer2_outputs(98) <= not(layer1_outputs(205));
    layer2_outputs(99) <= layer1_outputs(2150);
    layer2_outputs(100) <= (layer1_outputs(1479)) and not (layer1_outputs(129));
    layer2_outputs(101) <= not((layer1_outputs(170)) and (layer1_outputs(1357)));
    layer2_outputs(102) <= layer1_outputs(2342);
    layer2_outputs(103) <= '0';
    layer2_outputs(104) <= not((layer1_outputs(2346)) or (layer1_outputs(1862)));
    layer2_outputs(105) <= layer1_outputs(180);
    layer2_outputs(106) <= '0';
    layer2_outputs(107) <= layer1_outputs(1976);
    layer2_outputs(108) <= not((layer1_outputs(465)) and (layer1_outputs(209)));
    layer2_outputs(109) <= layer1_outputs(1790);
    layer2_outputs(110) <= not(layer1_outputs(1392)) or (layer1_outputs(324));
    layer2_outputs(111) <= not(layer1_outputs(282));
    layer2_outputs(112) <= not((layer1_outputs(279)) or (layer1_outputs(1353)));
    layer2_outputs(113) <= (layer1_outputs(232)) or (layer1_outputs(1424));
    layer2_outputs(114) <= (layer1_outputs(1956)) or (layer1_outputs(625));
    layer2_outputs(115) <= (layer1_outputs(1645)) and not (layer1_outputs(2259));
    layer2_outputs(116) <= layer1_outputs(1938);
    layer2_outputs(117) <= not(layer1_outputs(1567)) or (layer1_outputs(1463));
    layer2_outputs(118) <= '0';
    layer2_outputs(119) <= not(layer1_outputs(2006)) or (layer1_outputs(1275));
    layer2_outputs(120) <= not(layer1_outputs(416));
    layer2_outputs(121) <= '1';
    layer2_outputs(122) <= not(layer1_outputs(2222)) or (layer1_outputs(648));
    layer2_outputs(123) <= not(layer1_outputs(2238));
    layer2_outputs(124) <= not(layer1_outputs(2369));
    layer2_outputs(125) <= not(layer1_outputs(1053)) or (layer1_outputs(1578));
    layer2_outputs(126) <= not(layer1_outputs(179)) or (layer1_outputs(1713));
    layer2_outputs(127) <= (layer1_outputs(2257)) or (layer1_outputs(1938));
    layer2_outputs(128) <= not((layer1_outputs(1237)) or (layer1_outputs(1749)));
    layer2_outputs(129) <= layer1_outputs(296);
    layer2_outputs(130) <= '0';
    layer2_outputs(131) <= (layer1_outputs(1288)) and not (layer1_outputs(1008));
    layer2_outputs(132) <= not(layer1_outputs(2371));
    layer2_outputs(133) <= not(layer1_outputs(147));
    layer2_outputs(134) <= (layer1_outputs(194)) and not (layer1_outputs(2413));
    layer2_outputs(135) <= layer1_outputs(1289);
    layer2_outputs(136) <= layer1_outputs(1981);
    layer2_outputs(137) <= layer1_outputs(314);
    layer2_outputs(138) <= (layer1_outputs(1933)) or (layer1_outputs(124));
    layer2_outputs(139) <= layer1_outputs(1125);
    layer2_outputs(140) <= not((layer1_outputs(1509)) xor (layer1_outputs(1611)));
    layer2_outputs(141) <= '0';
    layer2_outputs(142) <= not(layer1_outputs(1025)) or (layer1_outputs(1658));
    layer2_outputs(143) <= '1';
    layer2_outputs(144) <= '0';
    layer2_outputs(145) <= (layer1_outputs(1339)) and not (layer1_outputs(0));
    layer2_outputs(146) <= not(layer1_outputs(1746)) or (layer1_outputs(2475));
    layer2_outputs(147) <= '1';
    layer2_outputs(148) <= not(layer1_outputs(2488)) or (layer1_outputs(731));
    layer2_outputs(149) <= layer1_outputs(1580);
    layer2_outputs(150) <= (layer1_outputs(1411)) and not (layer1_outputs(2325));
    layer2_outputs(151) <= layer1_outputs(2125);
    layer2_outputs(152) <= not((layer1_outputs(431)) or (layer1_outputs(294)));
    layer2_outputs(153) <= not(layer1_outputs(958));
    layer2_outputs(154) <= layer1_outputs(1015);
    layer2_outputs(155) <= '0';
    layer2_outputs(156) <= layer1_outputs(1315);
    layer2_outputs(157) <= layer1_outputs(361);
    layer2_outputs(158) <= (layer1_outputs(1018)) and not (layer1_outputs(116));
    layer2_outputs(159) <= layer1_outputs(1949);
    layer2_outputs(160) <= not(layer1_outputs(1458));
    layer2_outputs(161) <= (layer1_outputs(169)) or (layer1_outputs(1902));
    layer2_outputs(162) <= (layer1_outputs(215)) or (layer1_outputs(1647));
    layer2_outputs(163) <= layer1_outputs(1776);
    layer2_outputs(164) <= (layer1_outputs(152)) and not (layer1_outputs(2341));
    layer2_outputs(165) <= (layer1_outputs(483)) and (layer1_outputs(1062));
    layer2_outputs(166) <= layer1_outputs(1374);
    layer2_outputs(167) <= not(layer1_outputs(1686)) or (layer1_outputs(1760));
    layer2_outputs(168) <= (layer1_outputs(2251)) and not (layer1_outputs(462));
    layer2_outputs(169) <= layer1_outputs(1166);
    layer2_outputs(170) <= not(layer1_outputs(1102));
    layer2_outputs(171) <= not(layer1_outputs(1384));
    layer2_outputs(172) <= not((layer1_outputs(2202)) or (layer1_outputs(13)));
    layer2_outputs(173) <= (layer1_outputs(2095)) and not (layer1_outputs(1329));
    layer2_outputs(174) <= not((layer1_outputs(1797)) and (layer1_outputs(2551)));
    layer2_outputs(175) <= (layer1_outputs(307)) and (layer1_outputs(1978));
    layer2_outputs(176) <= not(layer1_outputs(1985));
    layer2_outputs(177) <= layer1_outputs(1500);
    layer2_outputs(178) <= not((layer1_outputs(1369)) or (layer1_outputs(335)));
    layer2_outputs(179) <= not((layer1_outputs(2178)) and (layer1_outputs(2331)));
    layer2_outputs(180) <= layer1_outputs(1421);
    layer2_outputs(181) <= layer1_outputs(1286);
    layer2_outputs(182) <= layer1_outputs(2338);
    layer2_outputs(183) <= (layer1_outputs(2268)) and (layer1_outputs(1123));
    layer2_outputs(184) <= '1';
    layer2_outputs(185) <= not((layer1_outputs(919)) and (layer1_outputs(140)));
    layer2_outputs(186) <= (layer1_outputs(1671)) and (layer1_outputs(1773));
    layer2_outputs(187) <= not(layer1_outputs(216)) or (layer1_outputs(1503));
    layer2_outputs(188) <= '1';
    layer2_outputs(189) <= not(layer1_outputs(2489));
    layer2_outputs(190) <= not((layer1_outputs(1086)) or (layer1_outputs(11)));
    layer2_outputs(191) <= layer1_outputs(747);
    layer2_outputs(192) <= not((layer1_outputs(2105)) or (layer1_outputs(429)));
    layer2_outputs(193) <= not((layer1_outputs(1203)) and (layer1_outputs(885)));
    layer2_outputs(194) <= layer1_outputs(1379);
    layer2_outputs(195) <= layer1_outputs(832);
    layer2_outputs(196) <= (layer1_outputs(189)) and not (layer1_outputs(1724));
    layer2_outputs(197) <= layer1_outputs(2184);
    layer2_outputs(198) <= not(layer1_outputs(2243));
    layer2_outputs(199) <= (layer1_outputs(1356)) and not (layer1_outputs(835));
    layer2_outputs(200) <= not(layer1_outputs(2211));
    layer2_outputs(201) <= layer1_outputs(2547);
    layer2_outputs(202) <= (layer1_outputs(614)) and not (layer1_outputs(2290));
    layer2_outputs(203) <= not(layer1_outputs(305));
    layer2_outputs(204) <= not(layer1_outputs(1252));
    layer2_outputs(205) <= layer1_outputs(1074);
    layer2_outputs(206) <= not(layer1_outputs(1356));
    layer2_outputs(207) <= (layer1_outputs(1804)) or (layer1_outputs(354));
    layer2_outputs(208) <= layer1_outputs(836);
    layer2_outputs(209) <= not(layer1_outputs(989));
    layer2_outputs(210) <= not((layer1_outputs(1875)) or (layer1_outputs(2088)));
    layer2_outputs(211) <= (layer1_outputs(575)) and not (layer1_outputs(2133));
    layer2_outputs(212) <= not(layer1_outputs(766)) or (layer1_outputs(607));
    layer2_outputs(213) <= (layer1_outputs(2415)) and (layer1_outputs(548));
    layer2_outputs(214) <= not(layer1_outputs(1028)) or (layer1_outputs(1798));
    layer2_outputs(215) <= layer1_outputs(151);
    layer2_outputs(216) <= not(layer1_outputs(1368)) or (layer1_outputs(1082));
    layer2_outputs(217) <= layer1_outputs(2424);
    layer2_outputs(218) <= not(layer1_outputs(1738)) or (layer1_outputs(1230));
    layer2_outputs(219) <= '0';
    layer2_outputs(220) <= layer1_outputs(859);
    layer2_outputs(221) <= '0';
    layer2_outputs(222) <= not((layer1_outputs(1030)) and (layer1_outputs(1185)));
    layer2_outputs(223) <= (layer1_outputs(1517)) and not (layer1_outputs(1334));
    layer2_outputs(224) <= layer1_outputs(2025);
    layer2_outputs(225) <= not((layer1_outputs(10)) and (layer1_outputs(948)));
    layer2_outputs(226) <= not(layer1_outputs(2270));
    layer2_outputs(227) <= not(layer1_outputs(1129));
    layer2_outputs(228) <= (layer1_outputs(31)) and (layer1_outputs(1614));
    layer2_outputs(229) <= (layer1_outputs(617)) and (layer1_outputs(1399));
    layer2_outputs(230) <= not(layer1_outputs(36));
    layer2_outputs(231) <= layer1_outputs(1455);
    layer2_outputs(232) <= not(layer1_outputs(1329)) or (layer1_outputs(491));
    layer2_outputs(233) <= (layer1_outputs(1695)) and not (layer1_outputs(815));
    layer2_outputs(234) <= (layer1_outputs(109)) and not (layer1_outputs(311));
    layer2_outputs(235) <= not(layer1_outputs(364)) or (layer1_outputs(1760));
    layer2_outputs(236) <= layer1_outputs(1961);
    layer2_outputs(237) <= (layer1_outputs(2337)) or (layer1_outputs(988));
    layer2_outputs(238) <= not(layer1_outputs(501)) or (layer1_outputs(165));
    layer2_outputs(239) <= not((layer1_outputs(2434)) or (layer1_outputs(1712)));
    layer2_outputs(240) <= layer1_outputs(1805);
    layer2_outputs(241) <= (layer1_outputs(223)) xor (layer1_outputs(1081));
    layer2_outputs(242) <= (layer1_outputs(1894)) and (layer1_outputs(273));
    layer2_outputs(243) <= not(layer1_outputs(1791)) or (layer1_outputs(1307));
    layer2_outputs(244) <= (layer1_outputs(34)) xor (layer1_outputs(1095));
    layer2_outputs(245) <= (layer1_outputs(2152)) and not (layer1_outputs(81));
    layer2_outputs(246) <= not(layer1_outputs(281));
    layer2_outputs(247) <= (layer1_outputs(1934)) or (layer1_outputs(1117));
    layer2_outputs(248) <= not(layer1_outputs(2153));
    layer2_outputs(249) <= (layer1_outputs(1265)) and not (layer1_outputs(2364));
    layer2_outputs(250) <= (layer1_outputs(2339)) and not (layer1_outputs(19));
    layer2_outputs(251) <= not(layer1_outputs(2491));
    layer2_outputs(252) <= not(layer1_outputs(2116)) or (layer1_outputs(1188));
    layer2_outputs(253) <= not((layer1_outputs(2285)) or (layer1_outputs(820)));
    layer2_outputs(254) <= not(layer1_outputs(515)) or (layer1_outputs(405));
    layer2_outputs(255) <= (layer1_outputs(2192)) and (layer1_outputs(408));
    layer2_outputs(256) <= not((layer1_outputs(2112)) and (layer1_outputs(160)));
    layer2_outputs(257) <= (layer1_outputs(1371)) or (layer1_outputs(940));
    layer2_outputs(258) <= '0';
    layer2_outputs(259) <= not(layer1_outputs(1685));
    layer2_outputs(260) <= '1';
    layer2_outputs(261) <= (layer1_outputs(666)) and not (layer1_outputs(1592));
    layer2_outputs(262) <= not(layer1_outputs(1428));
    layer2_outputs(263) <= not((layer1_outputs(283)) and (layer1_outputs(1860)));
    layer2_outputs(264) <= not(layer1_outputs(2311)) or (layer1_outputs(1053));
    layer2_outputs(265) <= (layer1_outputs(1874)) and not (layer1_outputs(1010));
    layer2_outputs(266) <= (layer1_outputs(2081)) or (layer1_outputs(1941));
    layer2_outputs(267) <= '0';
    layer2_outputs(268) <= (layer1_outputs(77)) and not (layer1_outputs(931));
    layer2_outputs(269) <= not(layer1_outputs(201));
    layer2_outputs(270) <= (layer1_outputs(891)) and not (layer1_outputs(2315));
    layer2_outputs(271) <= not(layer1_outputs(27));
    layer2_outputs(272) <= not(layer1_outputs(1872)) or (layer1_outputs(1909));
    layer2_outputs(273) <= not(layer1_outputs(1107)) or (layer1_outputs(567));
    layer2_outputs(274) <= '0';
    layer2_outputs(275) <= layer1_outputs(2008);
    layer2_outputs(276) <= (layer1_outputs(1695)) and (layer1_outputs(1521));
    layer2_outputs(277) <= not(layer1_outputs(576));
    layer2_outputs(278) <= not(layer1_outputs(1758));
    layer2_outputs(279) <= not(layer1_outputs(488));
    layer2_outputs(280) <= '1';
    layer2_outputs(281) <= '1';
    layer2_outputs(282) <= not(layer1_outputs(615)) or (layer1_outputs(2448));
    layer2_outputs(283) <= (layer1_outputs(928)) and not (layer1_outputs(2510));
    layer2_outputs(284) <= not(layer1_outputs(790));
    layer2_outputs(285) <= not(layer1_outputs(1386)) or (layer1_outputs(1801));
    layer2_outputs(286) <= not(layer1_outputs(1767));
    layer2_outputs(287) <= not(layer1_outputs(1167)) or (layer1_outputs(570));
    layer2_outputs(288) <= (layer1_outputs(1398)) and (layer1_outputs(1291));
    layer2_outputs(289) <= layer1_outputs(1216);
    layer2_outputs(290) <= layer1_outputs(1746);
    layer2_outputs(291) <= (layer1_outputs(2094)) or (layer1_outputs(844));
    layer2_outputs(292) <= layer1_outputs(1415);
    layer2_outputs(293) <= not(layer1_outputs(907)) or (layer1_outputs(705));
    layer2_outputs(294) <= layer1_outputs(414);
    layer2_outputs(295) <= layer1_outputs(691);
    layer2_outputs(296) <= (layer1_outputs(1568)) and not (layer1_outputs(2514));
    layer2_outputs(297) <= layer1_outputs(149);
    layer2_outputs(298) <= not(layer1_outputs(926));
    layer2_outputs(299) <= not(layer1_outputs(1332)) or (layer1_outputs(1420));
    layer2_outputs(300) <= not(layer1_outputs(1493));
    layer2_outputs(301) <= (layer1_outputs(1925)) and not (layer1_outputs(303));
    layer2_outputs(302) <= not((layer1_outputs(1482)) and (layer1_outputs(1887)));
    layer2_outputs(303) <= layer1_outputs(854);
    layer2_outputs(304) <= not((layer1_outputs(55)) or (layer1_outputs(821)));
    layer2_outputs(305) <= (layer1_outputs(2105)) and (layer1_outputs(1414));
    layer2_outputs(306) <= not(layer1_outputs(1133));
    layer2_outputs(307) <= not(layer1_outputs(1929));
    layer2_outputs(308) <= layer1_outputs(678);
    layer2_outputs(309) <= (layer1_outputs(2051)) and not (layer1_outputs(538));
    layer2_outputs(310) <= not((layer1_outputs(2067)) or (layer1_outputs(193)));
    layer2_outputs(311) <= (layer1_outputs(1050)) and not (layer1_outputs(563));
    layer2_outputs(312) <= layer1_outputs(581);
    layer2_outputs(313) <= not((layer1_outputs(1725)) and (layer1_outputs(2452)));
    layer2_outputs(314) <= not((layer1_outputs(514)) or (layer1_outputs(874)));
    layer2_outputs(315) <= layer1_outputs(2432);
    layer2_outputs(316) <= not(layer1_outputs(667));
    layer2_outputs(317) <= layer1_outputs(2429);
    layer2_outputs(318) <= (layer1_outputs(457)) and not (layer1_outputs(1415));
    layer2_outputs(319) <= not(layer1_outputs(336));
    layer2_outputs(320) <= not((layer1_outputs(749)) and (layer1_outputs(1628)));
    layer2_outputs(321) <= not(layer1_outputs(1714));
    layer2_outputs(322) <= not(layer1_outputs(1283));
    layer2_outputs(323) <= not(layer1_outputs(1236)) or (layer1_outputs(1151));
    layer2_outputs(324) <= not((layer1_outputs(512)) and (layer1_outputs(216)));
    layer2_outputs(325) <= layer1_outputs(1100);
    layer2_outputs(326) <= (layer1_outputs(2134)) and not (layer1_outputs(1005));
    layer2_outputs(327) <= not((layer1_outputs(2084)) or (layer1_outputs(2321)));
    layer2_outputs(328) <= (layer1_outputs(1104)) and not (layer1_outputs(538));
    layer2_outputs(329) <= not((layer1_outputs(2466)) and (layer1_outputs(2161)));
    layer2_outputs(330) <= layer1_outputs(860);
    layer2_outputs(331) <= '1';
    layer2_outputs(332) <= (layer1_outputs(146)) xor (layer1_outputs(2238));
    layer2_outputs(333) <= layer1_outputs(1233);
    layer2_outputs(334) <= '1';
    layer2_outputs(335) <= not(layer1_outputs(818));
    layer2_outputs(336) <= not(layer1_outputs(2296));
    layer2_outputs(337) <= (layer1_outputs(2148)) and not (layer1_outputs(162));
    layer2_outputs(338) <= (layer1_outputs(1409)) and not (layer1_outputs(1807));
    layer2_outputs(339) <= '0';
    layer2_outputs(340) <= layer1_outputs(412);
    layer2_outputs(341) <= '0';
    layer2_outputs(342) <= not(layer1_outputs(1314)) or (layer1_outputs(567));
    layer2_outputs(343) <= (layer1_outputs(2226)) and (layer1_outputs(2286));
    layer2_outputs(344) <= layer1_outputs(1793);
    layer2_outputs(345) <= '1';
    layer2_outputs(346) <= (layer1_outputs(1993)) and not (layer1_outputs(1663));
    layer2_outputs(347) <= (layer1_outputs(2067)) and not (layer1_outputs(1223));
    layer2_outputs(348) <= (layer1_outputs(649)) and (layer1_outputs(2056));
    layer2_outputs(349) <= not((layer1_outputs(1431)) and (layer1_outputs(1814)));
    layer2_outputs(350) <= not(layer1_outputs(1448));
    layer2_outputs(351) <= not(layer1_outputs(2054)) or (layer1_outputs(2380));
    layer2_outputs(352) <= not(layer1_outputs(2285));
    layer2_outputs(353) <= layer1_outputs(796);
    layer2_outputs(354) <= not((layer1_outputs(1790)) and (layer1_outputs(1449)));
    layer2_outputs(355) <= (layer1_outputs(1612)) and not (layer1_outputs(1434));
    layer2_outputs(356) <= (layer1_outputs(1954)) or (layer1_outputs(1132));
    layer2_outputs(357) <= not(layer1_outputs(1742));
    layer2_outputs(358) <= '1';
    layer2_outputs(359) <= (layer1_outputs(2131)) and not (layer1_outputs(664));
    layer2_outputs(360) <= '0';
    layer2_outputs(361) <= layer1_outputs(1764);
    layer2_outputs(362) <= not(layer1_outputs(1743));
    layer2_outputs(363) <= (layer1_outputs(2511)) and not (layer1_outputs(1989));
    layer2_outputs(364) <= (layer1_outputs(703)) or (layer1_outputs(665));
    layer2_outputs(365) <= not(layer1_outputs(1178));
    layer2_outputs(366) <= not(layer1_outputs(2336));
    layer2_outputs(367) <= (layer1_outputs(2060)) or (layer1_outputs(1485));
    layer2_outputs(368) <= not(layer1_outputs(993));
    layer2_outputs(369) <= layer1_outputs(2383);
    layer2_outputs(370) <= not(layer1_outputs(1386));
    layer2_outputs(371) <= (layer1_outputs(2204)) and not (layer1_outputs(2451));
    layer2_outputs(372) <= '0';
    layer2_outputs(373) <= '1';
    layer2_outputs(374) <= layer1_outputs(592);
    layer2_outputs(375) <= layer1_outputs(2413);
    layer2_outputs(376) <= not(layer1_outputs(580));
    layer2_outputs(377) <= (layer1_outputs(1550)) and not (layer1_outputs(199));
    layer2_outputs(378) <= not(layer1_outputs(1096));
    layer2_outputs(379) <= '1';
    layer2_outputs(380) <= not(layer1_outputs(1637)) or (layer1_outputs(2140));
    layer2_outputs(381) <= '0';
    layer2_outputs(382) <= not(layer1_outputs(1428));
    layer2_outputs(383) <= layer1_outputs(2372);
    layer2_outputs(384) <= not((layer1_outputs(1216)) or (layer1_outputs(114)));
    layer2_outputs(385) <= layer1_outputs(802);
    layer2_outputs(386) <= (layer1_outputs(212)) and (layer1_outputs(658));
    layer2_outputs(387) <= not(layer1_outputs(655)) or (layer1_outputs(408));
    layer2_outputs(388) <= not(layer1_outputs(664));
    layer2_outputs(389) <= (layer1_outputs(2061)) and (layer1_outputs(424));
    layer2_outputs(390) <= not(layer1_outputs(1090)) or (layer1_outputs(915));
    layer2_outputs(391) <= not(layer1_outputs(1214));
    layer2_outputs(392) <= layer1_outputs(829);
    layer2_outputs(393) <= not((layer1_outputs(756)) or (layer1_outputs(1079)));
    layer2_outputs(394) <= not(layer1_outputs(1059)) or (layer1_outputs(2423));
    layer2_outputs(395) <= not(layer1_outputs(1720));
    layer2_outputs(396) <= (layer1_outputs(52)) xor (layer1_outputs(81));
    layer2_outputs(397) <= (layer1_outputs(1894)) and not (layer1_outputs(960));
    layer2_outputs(398) <= (layer1_outputs(653)) and (layer1_outputs(1303));
    layer2_outputs(399) <= not((layer1_outputs(2021)) xor (layer1_outputs(1949)));
    layer2_outputs(400) <= not((layer1_outputs(2389)) and (layer1_outputs(2191)));
    layer2_outputs(401) <= not((layer1_outputs(1014)) or (layer1_outputs(916)));
    layer2_outputs(402) <= not(layer1_outputs(355));
    layer2_outputs(403) <= layer1_outputs(642);
    layer2_outputs(404) <= not((layer1_outputs(1673)) xor (layer1_outputs(297)));
    layer2_outputs(405) <= layer1_outputs(2015);
    layer2_outputs(406) <= (layer1_outputs(1562)) or (layer1_outputs(29));
    layer2_outputs(407) <= not(layer1_outputs(532));
    layer2_outputs(408) <= (layer1_outputs(946)) or (layer1_outputs(1627));
    layer2_outputs(409) <= not(layer1_outputs(1685));
    layer2_outputs(410) <= not(layer1_outputs(1014));
    layer2_outputs(411) <= layer1_outputs(634);
    layer2_outputs(412) <= not((layer1_outputs(1231)) or (layer1_outputs(2522)));
    layer2_outputs(413) <= not(layer1_outputs(1852));
    layer2_outputs(414) <= '0';
    layer2_outputs(415) <= (layer1_outputs(1636)) or (layer1_outputs(6));
    layer2_outputs(416) <= not(layer1_outputs(591)) or (layer1_outputs(764));
    layer2_outputs(417) <= not((layer1_outputs(44)) or (layer1_outputs(2556)));
    layer2_outputs(418) <= (layer1_outputs(1097)) and not (layer1_outputs(636));
    layer2_outputs(419) <= (layer1_outputs(1844)) and (layer1_outputs(470));
    layer2_outputs(420) <= not(layer1_outputs(2171));
    layer2_outputs(421) <= not(layer1_outputs(1161));
    layer2_outputs(422) <= layer1_outputs(2349);
    layer2_outputs(423) <= (layer1_outputs(242)) xor (layer1_outputs(1049));
    layer2_outputs(424) <= '0';
    layer2_outputs(425) <= not((layer1_outputs(220)) xor (layer1_outputs(1058)));
    layer2_outputs(426) <= (layer1_outputs(750)) and not (layer1_outputs(2535));
    layer2_outputs(427) <= layer1_outputs(532);
    layer2_outputs(428) <= (layer1_outputs(1844)) and not (layer1_outputs(2175));
    layer2_outputs(429) <= layer1_outputs(987);
    layer2_outputs(430) <= (layer1_outputs(1631)) and not (layer1_outputs(1314));
    layer2_outputs(431) <= not((layer1_outputs(1903)) or (layer1_outputs(1794)));
    layer2_outputs(432) <= not(layer1_outputs(316));
    layer2_outputs(433) <= (layer1_outputs(114)) or (layer1_outputs(586));
    layer2_outputs(434) <= not(layer1_outputs(1244)) or (layer1_outputs(1683));
    layer2_outputs(435) <= (layer1_outputs(2267)) or (layer1_outputs(868));
    layer2_outputs(436) <= layer1_outputs(549);
    layer2_outputs(437) <= layer1_outputs(1133);
    layer2_outputs(438) <= (layer1_outputs(197)) and (layer1_outputs(1967));
    layer2_outputs(439) <= '0';
    layer2_outputs(440) <= '0';
    layer2_outputs(441) <= not(layer1_outputs(335));
    layer2_outputs(442) <= '0';
    layer2_outputs(443) <= not((layer1_outputs(772)) or (layer1_outputs(1143)));
    layer2_outputs(444) <= (layer1_outputs(1174)) and not (layer1_outputs(705));
    layer2_outputs(445) <= not((layer1_outputs(208)) or (layer1_outputs(997)));
    layer2_outputs(446) <= not(layer1_outputs(80)) or (layer1_outputs(980));
    layer2_outputs(447) <= layer1_outputs(568);
    layer2_outputs(448) <= layer1_outputs(1336);
    layer2_outputs(449) <= '0';
    layer2_outputs(450) <= not(layer1_outputs(2361));
    layer2_outputs(451) <= not(layer1_outputs(587)) or (layer1_outputs(683));
    layer2_outputs(452) <= layer1_outputs(1339);
    layer2_outputs(453) <= layer1_outputs(644);
    layer2_outputs(454) <= '1';
    layer2_outputs(455) <= (layer1_outputs(2068)) and (layer1_outputs(2308));
    layer2_outputs(456) <= not(layer1_outputs(1340)) or (layer1_outputs(2522));
    layer2_outputs(457) <= layer1_outputs(1556);
    layer2_outputs(458) <= '1';
    layer2_outputs(459) <= layer1_outputs(920);
    layer2_outputs(460) <= not((layer1_outputs(298)) or (layer1_outputs(1038)));
    layer2_outputs(461) <= '0';
    layer2_outputs(462) <= (layer1_outputs(158)) and (layer1_outputs(1484));
    layer2_outputs(463) <= not(layer1_outputs(287));
    layer2_outputs(464) <= not((layer1_outputs(1432)) or (layer1_outputs(2498)));
    layer2_outputs(465) <= (layer1_outputs(223)) and (layer1_outputs(2304));
    layer2_outputs(466) <= not((layer1_outputs(2108)) and (layer1_outputs(2555)));
    layer2_outputs(467) <= (layer1_outputs(2200)) or (layer1_outputs(750));
    layer2_outputs(468) <= layer1_outputs(1770);
    layer2_outputs(469) <= layer1_outputs(1630);
    layer2_outputs(470) <= (layer1_outputs(1044)) and not (layer1_outputs(1627));
    layer2_outputs(471) <= (layer1_outputs(1272)) or (layer1_outputs(2351));
    layer2_outputs(472) <= (layer1_outputs(2260)) and not (layer1_outputs(494));
    layer2_outputs(473) <= not(layer1_outputs(833));
    layer2_outputs(474) <= (layer1_outputs(239)) or (layer1_outputs(2516));
    layer2_outputs(475) <= not(layer1_outputs(1233)) or (layer1_outputs(1112));
    layer2_outputs(476) <= layer1_outputs(934);
    layer2_outputs(477) <= (layer1_outputs(993)) and (layer1_outputs(1400));
    layer2_outputs(478) <= not(layer1_outputs(409));
    layer2_outputs(479) <= not(layer1_outputs(1769));
    layer2_outputs(480) <= not(layer1_outputs(1279));
    layer2_outputs(481) <= not(layer1_outputs(1162));
    layer2_outputs(482) <= not(layer1_outputs(861));
    layer2_outputs(483) <= layer1_outputs(2476);
    layer2_outputs(484) <= (layer1_outputs(1077)) and (layer1_outputs(1308));
    layer2_outputs(485) <= not(layer1_outputs(2020)) or (layer1_outputs(982));
    layer2_outputs(486) <= '0';
    layer2_outputs(487) <= not(layer1_outputs(1074)) or (layer1_outputs(1957));
    layer2_outputs(488) <= layer1_outputs(1347);
    layer2_outputs(489) <= not(layer1_outputs(156));
    layer2_outputs(490) <= not(layer1_outputs(1652));
    layer2_outputs(491) <= layer1_outputs(529);
    layer2_outputs(492) <= not((layer1_outputs(2155)) or (layer1_outputs(2515)));
    layer2_outputs(493) <= layer1_outputs(1954);
    layer2_outputs(494) <= layer1_outputs(1997);
    layer2_outputs(495) <= (layer1_outputs(812)) xor (layer1_outputs(1531));
    layer2_outputs(496) <= not(layer1_outputs(963));
    layer2_outputs(497) <= not((layer1_outputs(1968)) xor (layer1_outputs(1378)));
    layer2_outputs(498) <= (layer1_outputs(1945)) and not (layer1_outputs(1182));
    layer2_outputs(499) <= '1';
    layer2_outputs(500) <= (layer1_outputs(1213)) and not (layer1_outputs(318));
    layer2_outputs(501) <= (layer1_outputs(219)) and not (layer1_outputs(95));
    layer2_outputs(502) <= not(layer1_outputs(2013));
    layer2_outputs(503) <= layer1_outputs(1088);
    layer2_outputs(504) <= (layer1_outputs(2057)) or (layer1_outputs(1221));
    layer2_outputs(505) <= '0';
    layer2_outputs(506) <= (layer1_outputs(741)) and not (layer1_outputs(66));
    layer2_outputs(507) <= not(layer1_outputs(2376));
    layer2_outputs(508) <= '0';
    layer2_outputs(509) <= not(layer1_outputs(1160));
    layer2_outputs(510) <= '1';
    layer2_outputs(511) <= layer1_outputs(557);
    layer2_outputs(512) <= layer1_outputs(761);
    layer2_outputs(513) <= not(layer1_outputs(1359));
    layer2_outputs(514) <= not(layer1_outputs(691));
    layer2_outputs(515) <= not((layer1_outputs(137)) and (layer1_outputs(22)));
    layer2_outputs(516) <= not((layer1_outputs(882)) and (layer1_outputs(2475)));
    layer2_outputs(517) <= not(layer1_outputs(597));
    layer2_outputs(518) <= not(layer1_outputs(582)) or (layer1_outputs(1879));
    layer2_outputs(519) <= layer1_outputs(850);
    layer2_outputs(520) <= not(layer1_outputs(676)) or (layer1_outputs(461));
    layer2_outputs(521) <= layer1_outputs(1370);
    layer2_outputs(522) <= layer1_outputs(559);
    layer2_outputs(523) <= (layer1_outputs(389)) and (layer1_outputs(1615));
    layer2_outputs(524) <= not(layer1_outputs(2032)) or (layer1_outputs(378));
    layer2_outputs(525) <= not(layer1_outputs(2097));
    layer2_outputs(526) <= (layer1_outputs(742)) and (layer1_outputs(2387));
    layer2_outputs(527) <= not(layer1_outputs(2162));
    layer2_outputs(528) <= layer1_outputs(2096);
    layer2_outputs(529) <= layer1_outputs(1679);
    layer2_outputs(530) <= not(layer1_outputs(455));
    layer2_outputs(531) <= (layer1_outputs(76)) and (layer1_outputs(511));
    layer2_outputs(532) <= not(layer1_outputs(842));
    layer2_outputs(533) <= not(layer1_outputs(1518));
    layer2_outputs(534) <= '0';
    layer2_outputs(535) <= not(layer1_outputs(1408));
    layer2_outputs(536) <= not(layer1_outputs(2090)) or (layer1_outputs(507));
    layer2_outputs(537) <= (layer1_outputs(1526)) or (layer1_outputs(582));
    layer2_outputs(538) <= layer1_outputs(96);
    layer2_outputs(539) <= not(layer1_outputs(751));
    layer2_outputs(540) <= layer1_outputs(2107);
    layer2_outputs(541) <= not(layer1_outputs(1303));
    layer2_outputs(542) <= layer1_outputs(346);
    layer2_outputs(543) <= not(layer1_outputs(1351));
    layer2_outputs(544) <= not((layer1_outputs(737)) and (layer1_outputs(2293)));
    layer2_outputs(545) <= (layer1_outputs(2431)) or (layer1_outputs(2321));
    layer2_outputs(546) <= not(layer1_outputs(1400)) or (layer1_outputs(896));
    layer2_outputs(547) <= (layer1_outputs(9)) or (layer1_outputs(123));
    layer2_outputs(548) <= not(layer1_outputs(2388));
    layer2_outputs(549) <= (layer1_outputs(624)) or (layer1_outputs(772));
    layer2_outputs(550) <= '1';
    layer2_outputs(551) <= layer1_outputs(1526);
    layer2_outputs(552) <= layer1_outputs(500);
    layer2_outputs(553) <= not((layer1_outputs(1108)) and (layer1_outputs(21)));
    layer2_outputs(554) <= not(layer1_outputs(207)) or (layer1_outputs(2248));
    layer2_outputs(555) <= not(layer1_outputs(2518)) or (layer1_outputs(1659));
    layer2_outputs(556) <= (layer1_outputs(2136)) and (layer1_outputs(2120));
    layer2_outputs(557) <= (layer1_outputs(1470)) or (layer1_outputs(2343));
    layer2_outputs(558) <= '0';
    layer2_outputs(559) <= not(layer1_outputs(2106));
    layer2_outputs(560) <= (layer1_outputs(427)) and not (layer1_outputs(1957));
    layer2_outputs(561) <= (layer1_outputs(313)) and (layer1_outputs(940));
    layer2_outputs(562) <= layer1_outputs(1425);
    layer2_outputs(563) <= (layer1_outputs(12)) or (layer1_outputs(2307));
    layer2_outputs(564) <= not(layer1_outputs(2058)) or (layer1_outputs(2336));
    layer2_outputs(565) <= '0';
    layer2_outputs(566) <= (layer1_outputs(140)) and not (layer1_outputs(495));
    layer2_outputs(567) <= (layer1_outputs(643)) and (layer1_outputs(1302));
    layer2_outputs(568) <= not(layer1_outputs(1829));
    layer2_outputs(569) <= not(layer1_outputs(1690));
    layer2_outputs(570) <= not((layer1_outputs(183)) xor (layer1_outputs(2279)));
    layer2_outputs(571) <= not((layer1_outputs(1797)) or (layer1_outputs(89)));
    layer2_outputs(572) <= (layer1_outputs(765)) and not (layer1_outputs(1257));
    layer2_outputs(573) <= not(layer1_outputs(24)) or (layer1_outputs(1915));
    layer2_outputs(574) <= not((layer1_outputs(1982)) and (layer1_outputs(1152)));
    layer2_outputs(575) <= '0';
    layer2_outputs(576) <= layer1_outputs(1889);
    layer2_outputs(577) <= (layer1_outputs(498)) xor (layer1_outputs(873));
    layer2_outputs(578) <= (layer1_outputs(997)) or (layer1_outputs(1824));
    layer2_outputs(579) <= not(layer1_outputs(2410)) or (layer1_outputs(1779));
    layer2_outputs(580) <= not(layer1_outputs(142));
    layer2_outputs(581) <= not((layer1_outputs(1702)) or (layer1_outputs(385)));
    layer2_outputs(582) <= not(layer1_outputs(2440)) or (layer1_outputs(2189));
    layer2_outputs(583) <= layer1_outputs(879);
    layer2_outputs(584) <= (layer1_outputs(976)) and not (layer1_outputs(141));
    layer2_outputs(585) <= not(layer1_outputs(1951));
    layer2_outputs(586) <= (layer1_outputs(1324)) and not (layer1_outputs(383));
    layer2_outputs(587) <= (layer1_outputs(2404)) and not (layer1_outputs(1834));
    layer2_outputs(588) <= (layer1_outputs(102)) xor (layer1_outputs(126));
    layer2_outputs(589) <= (layer1_outputs(505)) and not (layer1_outputs(1215));
    layer2_outputs(590) <= not(layer1_outputs(1160));
    layer2_outputs(591) <= not((layer1_outputs(559)) xor (layer1_outputs(1762)));
    layer2_outputs(592) <= layer1_outputs(2120);
    layer2_outputs(593) <= '1';
    layer2_outputs(594) <= (layer1_outputs(2130)) and not (layer1_outputs(1322));
    layer2_outputs(595) <= not(layer1_outputs(2458));
    layer2_outputs(596) <= (layer1_outputs(1307)) and not (layer1_outputs(2311));
    layer2_outputs(597) <= layer1_outputs(2093);
    layer2_outputs(598) <= layer1_outputs(74);
    layer2_outputs(599) <= (layer1_outputs(478)) and (layer1_outputs(2373));
    layer2_outputs(600) <= (layer1_outputs(2432)) or (layer1_outputs(588));
    layer2_outputs(601) <= not(layer1_outputs(2085));
    layer2_outputs(602) <= not((layer1_outputs(603)) xor (layer1_outputs(522)));
    layer2_outputs(603) <= not((layer1_outputs(94)) and (layer1_outputs(1165)));
    layer2_outputs(604) <= (layer1_outputs(1669)) and not (layer1_outputs(272));
    layer2_outputs(605) <= (layer1_outputs(166)) and not (layer1_outputs(584));
    layer2_outputs(606) <= (layer1_outputs(843)) and not (layer1_outputs(934));
    layer2_outputs(607) <= layer1_outputs(987);
    layer2_outputs(608) <= (layer1_outputs(2119)) and not (layer1_outputs(1379));
    layer2_outputs(609) <= (layer1_outputs(660)) or (layer1_outputs(2218));
    layer2_outputs(610) <= (layer1_outputs(686)) and not (layer1_outputs(293));
    layer2_outputs(611) <= layer1_outputs(1869);
    layer2_outputs(612) <= not(layer1_outputs(1184));
    layer2_outputs(613) <= layer1_outputs(2501);
    layer2_outputs(614) <= '1';
    layer2_outputs(615) <= layer1_outputs(791);
    layer2_outputs(616) <= (layer1_outputs(1226)) xor (layer1_outputs(1987));
    layer2_outputs(617) <= layer1_outputs(1792);
    layer2_outputs(618) <= layer1_outputs(1758);
    layer2_outputs(619) <= layer1_outputs(122);
    layer2_outputs(620) <= not(layer1_outputs(2083));
    layer2_outputs(621) <= (layer1_outputs(89)) and not (layer1_outputs(1149));
    layer2_outputs(622) <= not(layer1_outputs(2423));
    layer2_outputs(623) <= layer1_outputs(256);
    layer2_outputs(624) <= not(layer1_outputs(1189));
    layer2_outputs(625) <= not(layer1_outputs(459));
    layer2_outputs(626) <= not((layer1_outputs(2003)) or (layer1_outputs(1066)));
    layer2_outputs(627) <= layer1_outputs(1769);
    layer2_outputs(628) <= not(layer1_outputs(817));
    layer2_outputs(629) <= '0';
    layer2_outputs(630) <= '1';
    layer2_outputs(631) <= layer1_outputs(1864);
    layer2_outputs(632) <= not(layer1_outputs(747));
    layer2_outputs(633) <= not(layer1_outputs(830));
    layer2_outputs(634) <= not(layer1_outputs(3)) or (layer1_outputs(1935));
    layer2_outputs(635) <= (layer1_outputs(894)) and (layer1_outputs(808));
    layer2_outputs(636) <= (layer1_outputs(834)) and not (layer1_outputs(558));
    layer2_outputs(637) <= '1';
    layer2_outputs(638) <= layer1_outputs(2492);
    layer2_outputs(639) <= not((layer1_outputs(2190)) and (layer1_outputs(2157)));
    layer2_outputs(640) <= not(layer1_outputs(2296));
    layer2_outputs(641) <= '0';
    layer2_outputs(642) <= not(layer1_outputs(1667));
    layer2_outputs(643) <= (layer1_outputs(1007)) and not (layer1_outputs(2126));
    layer2_outputs(644) <= '1';
    layer2_outputs(645) <= not(layer1_outputs(951));
    layer2_outputs(646) <= not(layer1_outputs(1092)) or (layer1_outputs(2527));
    layer2_outputs(647) <= (layer1_outputs(2351)) and (layer1_outputs(68));
    layer2_outputs(648) <= not(layer1_outputs(1856));
    layer2_outputs(649) <= not(layer1_outputs(2371));
    layer2_outputs(650) <= (layer1_outputs(244)) and not (layer1_outputs(677));
    layer2_outputs(651) <= (layer1_outputs(1552)) and not (layer1_outputs(2549));
    layer2_outputs(652) <= not(layer1_outputs(577));
    layer2_outputs(653) <= (layer1_outputs(1227)) and (layer1_outputs(1707));
    layer2_outputs(654) <= not((layer1_outputs(2034)) xor (layer1_outputs(40)));
    layer2_outputs(655) <= (layer1_outputs(231)) and not (layer1_outputs(1732));
    layer2_outputs(656) <= not(layer1_outputs(953));
    layer2_outputs(657) <= not((layer1_outputs(2045)) or (layer1_outputs(1387)));
    layer2_outputs(658) <= layer1_outputs(2233);
    layer2_outputs(659) <= not(layer1_outputs(861));
    layer2_outputs(660) <= layer1_outputs(2416);
    layer2_outputs(661) <= (layer1_outputs(780)) and not (layer1_outputs(2214));
    layer2_outputs(662) <= not(layer1_outputs(544));
    layer2_outputs(663) <= not((layer1_outputs(1849)) and (layer1_outputs(1683)));
    layer2_outputs(664) <= (layer1_outputs(267)) and not (layer1_outputs(1336));
    layer2_outputs(665) <= (layer1_outputs(1338)) and not (layer1_outputs(2117));
    layer2_outputs(666) <= not(layer1_outputs(2360)) or (layer1_outputs(1381));
    layer2_outputs(667) <= layer1_outputs(1097);
    layer2_outputs(668) <= layer1_outputs(92);
    layer2_outputs(669) <= (layer1_outputs(1843)) and not (layer1_outputs(154));
    layer2_outputs(670) <= (layer1_outputs(786)) or (layer1_outputs(2115));
    layer2_outputs(671) <= not(layer1_outputs(1039));
    layer2_outputs(672) <= (layer1_outputs(351)) and not (layer1_outputs(2173));
    layer2_outputs(673) <= layer1_outputs(697);
    layer2_outputs(674) <= '1';
    layer2_outputs(675) <= layer1_outputs(979);
    layer2_outputs(676) <= layer1_outputs(1042);
    layer2_outputs(677) <= not(layer1_outputs(1880));
    layer2_outputs(678) <= (layer1_outputs(890)) and (layer1_outputs(1335));
    layer2_outputs(679) <= '1';
    layer2_outputs(680) <= '1';
    layer2_outputs(681) <= not(layer1_outputs(1106)) or (layer1_outputs(696));
    layer2_outputs(682) <= (layer1_outputs(1125)) and (layer1_outputs(290));
    layer2_outputs(683) <= layer1_outputs(1884);
    layer2_outputs(684) <= '1';
    layer2_outputs(685) <= not(layer1_outputs(1995)) or (layer1_outputs(1191));
    layer2_outputs(686) <= not(layer1_outputs(1071)) or (layer1_outputs(1362));
    layer2_outputs(687) <= layer1_outputs(1691);
    layer2_outputs(688) <= (layer1_outputs(770)) or (layer1_outputs(1146));
    layer2_outputs(689) <= not((layer1_outputs(310)) and (layer1_outputs(1081)));
    layer2_outputs(690) <= not(layer1_outputs(1318)) or (layer1_outputs(524));
    layer2_outputs(691) <= not(layer1_outputs(1337));
    layer2_outputs(692) <= '1';
    layer2_outputs(693) <= (layer1_outputs(1022)) and not (layer1_outputs(1058));
    layer2_outputs(694) <= layer1_outputs(2414);
    layer2_outputs(695) <= not((layer1_outputs(2456)) and (layer1_outputs(2521)));
    layer2_outputs(696) <= layer1_outputs(857);
    layer2_outputs(697) <= '1';
    layer2_outputs(698) <= not(layer1_outputs(2355)) or (layer1_outputs(1353));
    layer2_outputs(699) <= '0';
    layer2_outputs(700) <= (layer1_outputs(1033)) and not (layer1_outputs(1465));
    layer2_outputs(701) <= layer1_outputs(970);
    layer2_outputs(702) <= not(layer1_outputs(2300));
    layer2_outputs(703) <= (layer1_outputs(1549)) and not (layer1_outputs(1711));
    layer2_outputs(704) <= '0';
    layer2_outputs(705) <= not(layer1_outputs(317)) or (layer1_outputs(945));
    layer2_outputs(706) <= not(layer1_outputs(196));
    layer2_outputs(707) <= layer1_outputs(1737);
    layer2_outputs(708) <= not((layer1_outputs(851)) and (layer1_outputs(243)));
    layer2_outputs(709) <= (layer1_outputs(361)) and (layer1_outputs(1122));
    layer2_outputs(710) <= not((layer1_outputs(1651)) or (layer1_outputs(2323)));
    layer2_outputs(711) <= layer1_outputs(2074);
    layer2_outputs(712) <= (layer1_outputs(1388)) and not (layer1_outputs(391));
    layer2_outputs(713) <= (layer1_outputs(2363)) or (layer1_outputs(469));
    layer2_outputs(714) <= (layer1_outputs(1277)) or (layer1_outputs(306));
    layer2_outputs(715) <= layer1_outputs(2280);
    layer2_outputs(716) <= not((layer1_outputs(823)) xor (layer1_outputs(760)));
    layer2_outputs(717) <= '1';
    layer2_outputs(718) <= layer1_outputs(1878);
    layer2_outputs(719) <= layer1_outputs(1222);
    layer2_outputs(720) <= not(layer1_outputs(2182)) or (layer1_outputs(1278));
    layer2_outputs(721) <= (layer1_outputs(1916)) and (layer1_outputs(214));
    layer2_outputs(722) <= not(layer1_outputs(1218)) or (layer1_outputs(2500));
    layer2_outputs(723) <= not(layer1_outputs(58)) or (layer1_outputs(2433));
    layer2_outputs(724) <= not((layer1_outputs(2340)) and (layer1_outputs(2528)));
    layer2_outputs(725) <= (layer1_outputs(120)) and (layer1_outputs(2145));
    layer2_outputs(726) <= '0';
    layer2_outputs(727) <= layer1_outputs(1481);
    layer2_outputs(728) <= not((layer1_outputs(2357)) and (layer1_outputs(71)));
    layer2_outputs(729) <= layer1_outputs(1730);
    layer2_outputs(730) <= layer1_outputs(1341);
    layer2_outputs(731) <= (layer1_outputs(1675)) or (layer1_outputs(439));
    layer2_outputs(732) <= layer1_outputs(1430);
    layer2_outputs(733) <= (layer1_outputs(2109)) or (layer1_outputs(900));
    layer2_outputs(734) <= not((layer1_outputs(1723)) or (layer1_outputs(2479)));
    layer2_outputs(735) <= '1';
    layer2_outputs(736) <= not(layer1_outputs(52));
    layer2_outputs(737) <= layer1_outputs(300);
    layer2_outputs(738) <= (layer1_outputs(2277)) and not (layer1_outputs(1047));
    layer2_outputs(739) <= not((layer1_outputs(1026)) or (layer1_outputs(2471)));
    layer2_outputs(740) <= (layer1_outputs(1345)) and (layer1_outputs(2228));
    layer2_outputs(741) <= (layer1_outputs(1040)) or (layer1_outputs(654));
    layer2_outputs(742) <= '1';
    layer2_outputs(743) <= layer1_outputs(1986);
    layer2_outputs(744) <= not(layer1_outputs(1717)) or (layer1_outputs(128));
    layer2_outputs(745) <= (layer1_outputs(726)) or (layer1_outputs(28));
    layer2_outputs(746) <= not(layer1_outputs(880));
    layer2_outputs(747) <= not(layer1_outputs(420));
    layer2_outputs(748) <= layer1_outputs(1442);
    layer2_outputs(749) <= not((layer1_outputs(1435)) or (layer1_outputs(2330)));
    layer2_outputs(750) <= (layer1_outputs(2247)) and (layer1_outputs(762));
    layer2_outputs(751) <= (layer1_outputs(964)) and not (layer1_outputs(428));
    layer2_outputs(752) <= not(layer1_outputs(395)) or (layer1_outputs(840));
    layer2_outputs(753) <= layer1_outputs(1586);
    layer2_outputs(754) <= layer1_outputs(2497);
    layer2_outputs(755) <= not(layer1_outputs(2186));
    layer2_outputs(756) <= not(layer1_outputs(338)) or (layer1_outputs(1344));
    layer2_outputs(757) <= '1';
    layer2_outputs(758) <= not((layer1_outputs(474)) or (layer1_outputs(369)));
    layer2_outputs(759) <= layer1_outputs(59);
    layer2_outputs(760) <= layer1_outputs(2389);
    layer2_outputs(761) <= (layer1_outputs(2137)) xor (layer1_outputs(1453));
    layer2_outputs(762) <= layer1_outputs(1977);
    layer2_outputs(763) <= (layer1_outputs(621)) and (layer1_outputs(601));
    layer2_outputs(764) <= (layer1_outputs(2127)) and not (layer1_outputs(1632));
    layer2_outputs(765) <= layer1_outputs(1210);
    layer2_outputs(766) <= not(layer1_outputs(628));
    layer2_outputs(767) <= layer1_outputs(419);
    layer2_outputs(768) <= '0';
    layer2_outputs(769) <= layer1_outputs(1720);
    layer2_outputs(770) <= not(layer1_outputs(1926));
    layer2_outputs(771) <= not(layer1_outputs(1304)) or (layer1_outputs(1559));
    layer2_outputs(772) <= layer1_outputs(2397);
    layer2_outputs(773) <= (layer1_outputs(1098)) and not (layer1_outputs(2215));
    layer2_outputs(774) <= (layer1_outputs(215)) and not (layer1_outputs(985));
    layer2_outputs(775) <= not((layer1_outputs(827)) and (layer1_outputs(15)));
    layer2_outputs(776) <= (layer1_outputs(1049)) and (layer1_outputs(733));
    layer2_outputs(777) <= (layer1_outputs(62)) and (layer1_outputs(933));
    layer2_outputs(778) <= not(layer1_outputs(637));
    layer2_outputs(779) <= not(layer1_outputs(1259));
    layer2_outputs(780) <= not((layer1_outputs(1625)) and (layer1_outputs(368)));
    layer2_outputs(781) <= layer1_outputs(1891);
    layer2_outputs(782) <= not(layer1_outputs(381));
    layer2_outputs(783) <= not(layer1_outputs(2362));
    layer2_outputs(784) <= (layer1_outputs(969)) and (layer1_outputs(400));
    layer2_outputs(785) <= not(layer1_outputs(555));
    layer2_outputs(786) <= not(layer1_outputs(969)) or (layer1_outputs(1728));
    layer2_outputs(787) <= (layer1_outputs(167)) and not (layer1_outputs(1455));
    layer2_outputs(788) <= not((layer1_outputs(44)) or (layer1_outputs(1452)));
    layer2_outputs(789) <= (layer1_outputs(2499)) xor (layer1_outputs(541));
    layer2_outputs(790) <= layer1_outputs(226);
    layer2_outputs(791) <= '1';
    layer2_outputs(792) <= (layer1_outputs(256)) and (layer1_outputs(801));
    layer2_outputs(793) <= (layer1_outputs(2256)) and not (layer1_outputs(2417));
    layer2_outputs(794) <= not(layer1_outputs(2547)) or (layer1_outputs(1688));
    layer2_outputs(795) <= not(layer1_outputs(1623));
    layer2_outputs(796) <= not(layer1_outputs(1224)) or (layer1_outputs(1506));
    layer2_outputs(797) <= (layer1_outputs(1310)) xor (layer1_outputs(407));
    layer2_outputs(798) <= layer1_outputs(1828);
    layer2_outputs(799) <= not((layer1_outputs(1156)) and (layer1_outputs(1266)));
    layer2_outputs(800) <= not((layer1_outputs(857)) and (layer1_outputs(912)));
    layer2_outputs(801) <= (layer1_outputs(1606)) and (layer1_outputs(2218));
    layer2_outputs(802) <= not(layer1_outputs(2474));
    layer2_outputs(803) <= layer1_outputs(458);
    layer2_outputs(804) <= not(layer1_outputs(902));
    layer2_outputs(805) <= not((layer1_outputs(1963)) or (layer1_outputs(999)));
    layer2_outputs(806) <= layer1_outputs(1350);
    layer2_outputs(807) <= not(layer1_outputs(1560));
    layer2_outputs(808) <= (layer1_outputs(98)) and not (layer1_outputs(709));
    layer2_outputs(809) <= (layer1_outputs(1646)) or (layer1_outputs(1713));
    layer2_outputs(810) <= not(layer1_outputs(316));
    layer2_outputs(811) <= layer1_outputs(1729);
    layer2_outputs(812) <= layer1_outputs(1795);
    layer2_outputs(813) <= (layer1_outputs(560)) and not (layer1_outputs(295));
    layer2_outputs(814) <= not(layer1_outputs(111)) or (layer1_outputs(717));
    layer2_outputs(815) <= (layer1_outputs(1727)) and not (layer1_outputs(2502));
    layer2_outputs(816) <= '0';
    layer2_outputs(817) <= (layer1_outputs(1891)) or (layer1_outputs(1385));
    layer2_outputs(818) <= not(layer1_outputs(1804));
    layer2_outputs(819) <= layer1_outputs(1556);
    layer2_outputs(820) <= not(layer1_outputs(759));
    layer2_outputs(821) <= (layer1_outputs(276)) and (layer1_outputs(1328));
    layer2_outputs(822) <= not(layer1_outputs(873));
    layer2_outputs(823) <= not(layer1_outputs(421));
    layer2_outputs(824) <= not(layer1_outputs(1881)) or (layer1_outputs(1564));
    layer2_outputs(825) <= not((layer1_outputs(474)) or (layer1_outputs(572)));
    layer2_outputs(826) <= layer1_outputs(2291);
    layer2_outputs(827) <= not(layer1_outputs(1942));
    layer2_outputs(828) <= layer1_outputs(1791);
    layer2_outputs(829) <= not(layer1_outputs(375));
    layer2_outputs(830) <= not(layer1_outputs(1979));
    layer2_outputs(831) <= (layer1_outputs(856)) and (layer1_outputs(2546));
    layer2_outputs(832) <= '1';
    layer2_outputs(833) <= layer1_outputs(233);
    layer2_outputs(834) <= layer1_outputs(2445);
    layer2_outputs(835) <= (layer1_outputs(55)) and (layer1_outputs(1871));
    layer2_outputs(836) <= layer1_outputs(1300);
    layer2_outputs(837) <= layer1_outputs(36);
    layer2_outputs(838) <= '0';
    layer2_outputs(839) <= not(layer1_outputs(2241));
    layer2_outputs(840) <= not((layer1_outputs(392)) and (layer1_outputs(531)));
    layer2_outputs(841) <= (layer1_outputs(840)) and not (layer1_outputs(1971));
    layer2_outputs(842) <= layer1_outputs(2386);
    layer2_outputs(843) <= not(layer1_outputs(952));
    layer2_outputs(844) <= (layer1_outputs(546)) or (layer1_outputs(1378));
    layer2_outputs(845) <= not(layer1_outputs(713));
    layer2_outputs(846) <= '1';
    layer2_outputs(847) <= layer1_outputs(963);
    layer2_outputs(848) <= '0';
    layer2_outputs(849) <= layer1_outputs(1433);
    layer2_outputs(850) <= '0';
    layer2_outputs(851) <= not(layer1_outputs(2500)) or (layer1_outputs(1035));
    layer2_outputs(852) <= '1';
    layer2_outputs(853) <= layer1_outputs(190);
    layer2_outputs(854) <= not((layer1_outputs(2166)) or (layer1_outputs(1228)));
    layer2_outputs(855) <= (layer1_outputs(1278)) and not (layer1_outputs(192));
    layer2_outputs(856) <= not(layer1_outputs(1704));
    layer2_outputs(857) <= (layer1_outputs(1302)) and (layer1_outputs(961));
    layer2_outputs(858) <= (layer1_outputs(292)) or (layer1_outputs(823));
    layer2_outputs(859) <= not((layer1_outputs(1718)) or (layer1_outputs(1137)));
    layer2_outputs(860) <= (layer1_outputs(2065)) and not (layer1_outputs(638));
    layer2_outputs(861) <= (layer1_outputs(300)) and not (layer1_outputs(349));
    layer2_outputs(862) <= not(layer1_outputs(325)) or (layer1_outputs(1118));
    layer2_outputs(863) <= not(layer1_outputs(2442)) or (layer1_outputs(2309));
    layer2_outputs(864) <= not((layer1_outputs(2044)) or (layer1_outputs(707)));
    layer2_outputs(865) <= not(layer1_outputs(1482));
    layer2_outputs(866) <= layer1_outputs(2381);
    layer2_outputs(867) <= not(layer1_outputs(2390));
    layer2_outputs(868) <= (layer1_outputs(2526)) and not (layer1_outputs(731));
    layer2_outputs(869) <= not(layer1_outputs(2265));
    layer2_outputs(870) <= '0';
    layer2_outputs(871) <= '0';
    layer2_outputs(872) <= not(layer1_outputs(501)) or (layer1_outputs(1571));
    layer2_outputs(873) <= (layer1_outputs(2495)) and (layer1_outputs(2437));
    layer2_outputs(874) <= (layer1_outputs(1765)) and (layer1_outputs(1111));
    layer2_outputs(875) <= not((layer1_outputs(593)) and (layer1_outputs(454)));
    layer2_outputs(876) <= not(layer1_outputs(2102));
    layer2_outputs(877) <= (layer1_outputs(895)) xor (layer1_outputs(2024));
    layer2_outputs(878) <= not((layer1_outputs(518)) and (layer1_outputs(217)));
    layer2_outputs(879) <= '1';
    layer2_outputs(880) <= (layer1_outputs(1570)) and not (layer1_outputs(2512));
    layer2_outputs(881) <= not((layer1_outputs(1969)) xor (layer1_outputs(763)));
    layer2_outputs(882) <= not((layer1_outputs(2463)) and (layer1_outputs(1993)));
    layer2_outputs(883) <= (layer1_outputs(698)) and not (layer1_outputs(1996));
    layer2_outputs(884) <= layer1_outputs(1446);
    layer2_outputs(885) <= not(layer1_outputs(1808));
    layer2_outputs(886) <= (layer1_outputs(261)) and (layer1_outputs(2200));
    layer2_outputs(887) <= (layer1_outputs(695)) and (layer1_outputs(2295));
    layer2_outputs(888) <= (layer1_outputs(2099)) xor (layer1_outputs(2467));
    layer2_outputs(889) <= (layer1_outputs(255)) xor (layer1_outputs(352));
    layer2_outputs(890) <= '0';
    layer2_outputs(891) <= not((layer1_outputs(336)) or (layer1_outputs(1830)));
    layer2_outputs(892) <= '0';
    layer2_outputs(893) <= not(layer1_outputs(1472)) or (layer1_outputs(1457));
    layer2_outputs(894) <= not(layer1_outputs(1947)) or (layer1_outputs(1597));
    layer2_outputs(895) <= '0';
    layer2_outputs(896) <= layer1_outputs(1295);
    layer2_outputs(897) <= '1';
    layer2_outputs(898) <= not(layer1_outputs(1706)) or (layer1_outputs(27));
    layer2_outputs(899) <= '0';
    layer2_outputs(900) <= not(layer1_outputs(953)) or (layer1_outputs(1460));
    layer2_outputs(901) <= not(layer1_outputs(374));
    layer2_outputs(902) <= not(layer1_outputs(2349));
    layer2_outputs(903) <= not(layer1_outputs(17));
    layer2_outputs(904) <= (layer1_outputs(2035)) and not (layer1_outputs(225));
    layer2_outputs(905) <= not(layer1_outputs(1772));
    layer2_outputs(906) <= not(layer1_outputs(534));
    layer2_outputs(907) <= not((layer1_outputs(449)) and (layer1_outputs(1085)));
    layer2_outputs(908) <= (layer1_outputs(1888)) and not (layer1_outputs(1237));
    layer2_outputs(909) <= '0';
    layer2_outputs(910) <= not(layer1_outputs(32));
    layer2_outputs(911) <= layer1_outputs(1370);
    layer2_outputs(912) <= not((layer1_outputs(1987)) and (layer1_outputs(1876)));
    layer2_outputs(913) <= not(layer1_outputs(373)) or (layer1_outputs(648));
    layer2_outputs(914) <= not(layer1_outputs(2348));
    layer2_outputs(915) <= layer1_outputs(22);
    layer2_outputs(916) <= not((layer1_outputs(1946)) xor (layer1_outputs(2168)));
    layer2_outputs(917) <= not(layer1_outputs(1667));
    layer2_outputs(918) <= not(layer1_outputs(1206));
    layer2_outputs(919) <= not(layer1_outputs(1785)) or (layer1_outputs(2503));
    layer2_outputs(920) <= (layer1_outputs(1441)) and not (layer1_outputs(1317));
    layer2_outputs(921) <= (layer1_outputs(166)) and (layer1_outputs(1501));
    layer2_outputs(922) <= '1';
    layer2_outputs(923) <= not(layer1_outputs(2189));
    layer2_outputs(924) <= layer1_outputs(584);
    layer2_outputs(925) <= not(layer1_outputs(71));
    layer2_outputs(926) <= not((layer1_outputs(2534)) or (layer1_outputs(1859)));
    layer2_outputs(927) <= (layer1_outputs(1124)) and not (layer1_outputs(1786));
    layer2_outputs(928) <= layer1_outputs(1622);
    layer2_outputs(929) <= '1';
    layer2_outputs(930) <= '0';
    layer2_outputs(931) <= (layer1_outputs(1365)) and (layer1_outputs(1910));
    layer2_outputs(932) <= not((layer1_outputs(2151)) or (layer1_outputs(397)));
    layer2_outputs(933) <= (layer1_outputs(955)) and not (layer1_outputs(2541));
    layer2_outputs(934) <= layer1_outputs(1741);
    layer2_outputs(935) <= layer1_outputs(2345);
    layer2_outputs(936) <= not(layer1_outputs(895)) or (layer1_outputs(2366));
    layer2_outputs(937) <= layer1_outputs(1789);
    layer2_outputs(938) <= not((layer1_outputs(688)) and (layer1_outputs(2335)));
    layer2_outputs(939) <= '1';
    layer2_outputs(940) <= (layer1_outputs(1070)) and (layer1_outputs(518));
    layer2_outputs(941) <= not(layer1_outputs(370));
    layer2_outputs(942) <= '1';
    layer2_outputs(943) <= layer1_outputs(2451);
    layer2_outputs(944) <= not((layer1_outputs(2004)) and (layer1_outputs(2089)));
    layer2_outputs(945) <= (layer1_outputs(1129)) and not (layer1_outputs(41));
    layer2_outputs(946) <= not(layer1_outputs(2450));
    layer2_outputs(947) <= not(layer1_outputs(1260));
    layer2_outputs(948) <= (layer1_outputs(2242)) and not (layer1_outputs(1112));
    layer2_outputs(949) <= not((layer1_outputs(2016)) or (layer1_outputs(323)));
    layer2_outputs(950) <= not(layer1_outputs(762));
    layer2_outputs(951) <= layer1_outputs(2539);
    layer2_outputs(952) <= layer1_outputs(673);
    layer2_outputs(953) <= layer1_outputs(756);
    layer2_outputs(954) <= not(layer1_outputs(1288));
    layer2_outputs(955) <= not((layer1_outputs(1155)) or (layer1_outputs(1901)));
    layer2_outputs(956) <= not(layer1_outputs(1251));
    layer2_outputs(957) <= not((layer1_outputs(2327)) or (layer1_outputs(2176)));
    layer2_outputs(958) <= '1';
    layer2_outputs(959) <= not(layer1_outputs(425));
    layer2_outputs(960) <= '1';
    layer2_outputs(961) <= not(layer1_outputs(1567));
    layer2_outputs(962) <= layer1_outputs(2540);
    layer2_outputs(963) <= not(layer1_outputs(2097));
    layer2_outputs(964) <= not(layer1_outputs(2542));
    layer2_outputs(965) <= not(layer1_outputs(450)) or (layer1_outputs(1558));
    layer2_outputs(966) <= (layer1_outputs(1710)) and not (layer1_outputs(2024));
    layer2_outputs(967) <= layer1_outputs(1174);
    layer2_outputs(968) <= (layer1_outputs(1564)) and not (layer1_outputs(2245));
    layer2_outputs(969) <= layer1_outputs(775);
    layer2_outputs(970) <= '0';
    layer2_outputs(971) <= (layer1_outputs(444)) or (layer1_outputs(1406));
    layer2_outputs(972) <= not(layer1_outputs(1309));
    layer2_outputs(973) <= '1';
    layer2_outputs(974) <= '0';
    layer2_outputs(975) <= not(layer1_outputs(1159));
    layer2_outputs(976) <= not(layer1_outputs(1469));
    layer2_outputs(977) <= '0';
    layer2_outputs(978) <= '0';
    layer2_outputs(979) <= (layer1_outputs(1343)) and not (layer1_outputs(403));
    layer2_outputs(980) <= layer1_outputs(444);
    layer2_outputs(981) <= not(layer1_outputs(2233)) or (layer1_outputs(1608));
    layer2_outputs(982) <= (layer1_outputs(2352)) and not (layer1_outputs(2152));
    layer2_outputs(983) <= '0';
    layer2_outputs(984) <= (layer1_outputs(411)) or (layer1_outputs(2519));
    layer2_outputs(985) <= not(layer1_outputs(681));
    layer2_outputs(986) <= '1';
    layer2_outputs(987) <= (layer1_outputs(2147)) and not (layer1_outputs(506));
    layer2_outputs(988) <= (layer1_outputs(2422)) and (layer1_outputs(1940));
    layer2_outputs(989) <= not(layer1_outputs(1080));
    layer2_outputs(990) <= layer1_outputs(421);
    layer2_outputs(991) <= not((layer1_outputs(1527)) or (layer1_outputs(510)));
    layer2_outputs(992) <= (layer1_outputs(2049)) or (layer1_outputs(625));
    layer2_outputs(993) <= not(layer1_outputs(2402)) or (layer1_outputs(1464));
    layer2_outputs(994) <= layer1_outputs(1600);
    layer2_outputs(995) <= '1';
    layer2_outputs(996) <= layer1_outputs(867);
    layer2_outputs(997) <= not(layer1_outputs(16));
    layer2_outputs(998) <= layer1_outputs(2219);
    layer2_outputs(999) <= not((layer1_outputs(1190)) and (layer1_outputs(1596)));
    layer2_outputs(1000) <= '1';
    layer2_outputs(1001) <= not(layer1_outputs(1656)) or (layer1_outputs(1599));
    layer2_outputs(1002) <= not((layer1_outputs(8)) or (layer1_outputs(2553)));
    layer2_outputs(1003) <= (layer1_outputs(2181)) and (layer1_outputs(31));
    layer2_outputs(1004) <= layer1_outputs(1863);
    layer2_outputs(1005) <= layer1_outputs(844);
    layer2_outputs(1006) <= '0';
    layer2_outputs(1007) <= '1';
    layer2_outputs(1008) <= (layer1_outputs(1703)) or (layer1_outputs(155));
    layer2_outputs(1009) <= not(layer1_outputs(1061));
    layer2_outputs(1010) <= not(layer1_outputs(2504));
    layer2_outputs(1011) <= layer1_outputs(2470);
    layer2_outputs(1012) <= (layer1_outputs(1846)) and (layer1_outputs(1741));
    layer2_outputs(1013) <= '0';
    layer2_outputs(1014) <= '1';
    layer2_outputs(1015) <= not((layer1_outputs(237)) or (layer1_outputs(1784)));
    layer2_outputs(1016) <= (layer1_outputs(792)) xor (layer1_outputs(545));
    layer2_outputs(1017) <= layer1_outputs(769);
    layer2_outputs(1018) <= layer1_outputs(1860);
    layer2_outputs(1019) <= (layer1_outputs(1253)) and not (layer1_outputs(465));
    layer2_outputs(1020) <= not(layer1_outputs(982)) or (layer1_outputs(1116));
    layer2_outputs(1021) <= (layer1_outputs(1500)) and (layer1_outputs(2048));
    layer2_outputs(1022) <= layer1_outputs(2513);
    layer2_outputs(1023) <= not(layer1_outputs(1273)) or (layer1_outputs(1640));
    layer2_outputs(1024) <= (layer1_outputs(189)) and not (layer1_outputs(706));
    layer2_outputs(1025) <= (layer1_outputs(1566)) and not (layer1_outputs(1694));
    layer2_outputs(1026) <= '1';
    layer2_outputs(1027) <= (layer1_outputs(176)) and not (layer1_outputs(922));
    layer2_outputs(1028) <= (layer1_outputs(1316)) and not (layer1_outputs(2262));
    layer2_outputs(1029) <= '0';
    layer2_outputs(1030) <= not(layer1_outputs(1272));
    layer2_outputs(1031) <= layer1_outputs(2468);
    layer2_outputs(1032) <= layer1_outputs(262);
    layer2_outputs(1033) <= '0';
    layer2_outputs(1034) <= not(layer1_outputs(2362));
    layer2_outputs(1035) <= '1';
    layer2_outputs(1036) <= layer1_outputs(629);
    layer2_outputs(1037) <= not(layer1_outputs(1921)) or (layer1_outputs(1477));
    layer2_outputs(1038) <= layer1_outputs(329);
    layer2_outputs(1039) <= not(layer1_outputs(1065)) or (layer1_outputs(399));
    layer2_outputs(1040) <= not((layer1_outputs(2094)) and (layer1_outputs(327)));
    layer2_outputs(1041) <= not(layer1_outputs(2080)) or (layer1_outputs(1248));
    layer2_outputs(1042) <= (layer1_outputs(379)) and (layer1_outputs(2440));
    layer2_outputs(1043) <= layer1_outputs(1621);
    layer2_outputs(1044) <= not(layer1_outputs(424)) or (layer1_outputs(2220));
    layer2_outputs(1045) <= (layer1_outputs(1543)) or (layer1_outputs(2468));
    layer2_outputs(1046) <= (layer1_outputs(2317)) xor (layer1_outputs(1645));
    layer2_outputs(1047) <= '0';
    layer2_outputs(1048) <= (layer1_outputs(1850)) and not (layer1_outputs(1653));
    layer2_outputs(1049) <= not(layer1_outputs(1493)) or (layer1_outputs(285));
    layer2_outputs(1050) <= layer1_outputs(904);
    layer2_outputs(1051) <= layer1_outputs(1096);
    layer2_outputs(1052) <= layer1_outputs(2416);
    layer2_outputs(1053) <= not((layer1_outputs(1705)) and (layer1_outputs(1936)));
    layer2_outputs(1054) <= '1';
    layer2_outputs(1055) <= not(layer1_outputs(1324)) or (layer1_outputs(889));
    layer2_outputs(1056) <= not(layer1_outputs(78));
    layer2_outputs(1057) <= layer1_outputs(1190);
    layer2_outputs(1058) <= layer1_outputs(2208);
    layer2_outputs(1059) <= '1';
    layer2_outputs(1060) <= not(layer1_outputs(862));
    layer2_outputs(1061) <= layer1_outputs(2263);
    layer2_outputs(1062) <= not(layer1_outputs(2369));
    layer2_outputs(1063) <= not(layer1_outputs(1999));
    layer2_outputs(1064) <= '1';
    layer2_outputs(1065) <= (layer1_outputs(294)) and not (layer1_outputs(599));
    layer2_outputs(1066) <= not(layer1_outputs(1446));
    layer2_outputs(1067) <= layer1_outputs(2252);
    layer2_outputs(1068) <= '0';
    layer2_outputs(1069) <= (layer1_outputs(946)) and not (layer1_outputs(115));
    layer2_outputs(1070) <= layer1_outputs(1733);
    layer2_outputs(1071) <= '1';
    layer2_outputs(1072) <= not(layer1_outputs(1317));
    layer2_outputs(1073) <= not((layer1_outputs(1425)) or (layer1_outputs(2542)));
    layer2_outputs(1074) <= layer1_outputs(2384);
    layer2_outputs(1075) <= (layer1_outputs(1192)) or (layer1_outputs(1960));
    layer2_outputs(1076) <= not(layer1_outputs(1788));
    layer2_outputs(1077) <= layer1_outputs(2117);
    layer2_outputs(1078) <= (layer1_outputs(1165)) or (layer1_outputs(1271));
    layer2_outputs(1079) <= not((layer1_outputs(1473)) or (layer1_outputs(2385)));
    layer2_outputs(1080) <= (layer1_outputs(221)) and not (layer1_outputs(1234));
    layer2_outputs(1081) <= not((layer1_outputs(1971)) and (layer1_outputs(1159)));
    layer2_outputs(1082) <= '1';
    layer2_outputs(1083) <= layer1_outputs(1251);
    layer2_outputs(1084) <= layer1_outputs(2405);
    layer2_outputs(1085) <= not(layer1_outputs(776)) or (layer1_outputs(334));
    layer2_outputs(1086) <= not((layer1_outputs(212)) or (layer1_outputs(257)));
    layer2_outputs(1087) <= not((layer1_outputs(888)) and (layer1_outputs(1330)));
    layer2_outputs(1088) <= '0';
    layer2_outputs(1089) <= not(layer1_outputs(513));
    layer2_outputs(1090) <= not((layer1_outputs(738)) xor (layer1_outputs(1862)));
    layer2_outputs(1091) <= layer1_outputs(1416);
    layer2_outputs(1092) <= (layer1_outputs(2007)) and (layer1_outputs(477));
    layer2_outputs(1093) <= not(layer1_outputs(2280));
    layer2_outputs(1094) <= not((layer1_outputs(2407)) or (layer1_outputs(846)));
    layer2_outputs(1095) <= layer1_outputs(1308);
    layer2_outputs(1096) <= (layer1_outputs(2405)) and not (layer1_outputs(1840));
    layer2_outputs(1097) <= not(layer1_outputs(1613));
    layer2_outputs(1098) <= not(layer1_outputs(1496));
    layer2_outputs(1099) <= not((layer1_outputs(1727)) or (layer1_outputs(348)));
    layer2_outputs(1100) <= not(layer1_outputs(2281));
    layer2_outputs(1101) <= not(layer1_outputs(2294));
    layer2_outputs(1102) <= (layer1_outputs(1542)) or (layer1_outputs(1931));
    layer2_outputs(1103) <= layer1_outputs(2378);
    layer2_outputs(1104) <= (layer1_outputs(174)) xor (layer1_outputs(613));
    layer2_outputs(1105) <= not(layer1_outputs(264));
    layer2_outputs(1106) <= not(layer1_outputs(51)) or (layer1_outputs(1782));
    layer2_outputs(1107) <= (layer1_outputs(47)) xor (layer1_outputs(2188));
    layer2_outputs(1108) <= not(layer1_outputs(276));
    layer2_outputs(1109) <= layer1_outputs(229);
    layer2_outputs(1110) <= '1';
    layer2_outputs(1111) <= layer1_outputs(1154);
    layer2_outputs(1112) <= not(layer1_outputs(871));
    layer2_outputs(1113) <= not((layer1_outputs(1037)) xor (layer1_outputs(407)));
    layer2_outputs(1114) <= not(layer1_outputs(687)) or (layer1_outputs(1607));
    layer2_outputs(1115) <= layer1_outputs(1528);
    layer2_outputs(1116) <= (layer1_outputs(2450)) xor (layer1_outputs(431));
    layer2_outputs(1117) <= not(layer1_outputs(30)) or (layer1_outputs(773));
    layer2_outputs(1118) <= not(layer1_outputs(1205));
    layer2_outputs(1119) <= not(layer1_outputs(1850)) or (layer1_outputs(1161));
    layer2_outputs(1120) <= not(layer1_outputs(2154));
    layer2_outputs(1121) <= (layer1_outputs(138)) and (layer1_outputs(950));
    layer2_outputs(1122) <= not(layer1_outputs(417));
    layer2_outputs(1123) <= not((layer1_outputs(2082)) and (layer1_outputs(2355)));
    layer2_outputs(1124) <= (layer1_outputs(651)) or (layer1_outputs(2420));
    layer2_outputs(1125) <= (layer1_outputs(2530)) and not (layer1_outputs(776));
    layer2_outputs(1126) <= layer1_outputs(2524);
    layer2_outputs(1127) <= not(layer1_outputs(700));
    layer2_outputs(1128) <= (layer1_outputs(1929)) and not (layer1_outputs(206));
    layer2_outputs(1129) <= not(layer1_outputs(1499)) or (layer1_outputs(1209));
    layer2_outputs(1130) <= not((layer1_outputs(2110)) or (layer1_outputs(2328)));
    layer2_outputs(1131) <= not(layer1_outputs(818));
    layer2_outputs(1132) <= not(layer1_outputs(434));
    layer2_outputs(1133) <= not(layer1_outputs(1648));
    layer2_outputs(1134) <= (layer1_outputs(1146)) and (layer1_outputs(1423));
    layer2_outputs(1135) <= not(layer1_outputs(2545));
    layer2_outputs(1136) <= not(layer1_outputs(372));
    layer2_outputs(1137) <= layer1_outputs(707);
    layer2_outputs(1138) <= not(layer1_outputs(1643));
    layer2_outputs(1139) <= layer1_outputs(547);
    layer2_outputs(1140) <= not((layer1_outputs(1349)) or (layer1_outputs(82)));
    layer2_outputs(1141) <= not(layer1_outputs(2329));
    layer2_outputs(1142) <= not((layer1_outputs(2430)) xor (layer1_outputs(1486)));
    layer2_outputs(1143) <= (layer1_outputs(86)) and (layer1_outputs(2216));
    layer2_outputs(1144) <= not(layer1_outputs(2478));
    layer2_outputs(1145) <= (layer1_outputs(2050)) and not (layer1_outputs(2006));
    layer2_outputs(1146) <= layer1_outputs(1126);
    layer2_outputs(1147) <= not(layer1_outputs(467));
    layer2_outputs(1148) <= (layer1_outputs(1263)) and not (layer1_outputs(2493));
    layer2_outputs(1149) <= (layer1_outputs(1430)) and not (layer1_outputs(2348));
    layer2_outputs(1150) <= layer1_outputs(2537);
    layer2_outputs(1151) <= (layer1_outputs(1350)) and not (layer1_outputs(228));
    layer2_outputs(1152) <= not(layer1_outputs(868));
    layer2_outputs(1153) <= (layer1_outputs(401)) and not (layer1_outputs(902));
    layer2_outputs(1154) <= (layer1_outputs(2301)) and not (layer1_outputs(898));
    layer2_outputs(1155) <= not((layer1_outputs(1948)) xor (layer1_outputs(930)));
    layer2_outputs(1156) <= layer1_outputs(57);
    layer2_outputs(1157) <= not(layer1_outputs(1926));
    layer2_outputs(1158) <= not((layer1_outputs(277)) and (layer1_outputs(2478)));
    layer2_outputs(1159) <= not(layer1_outputs(1095));
    layer2_outputs(1160) <= layer1_outputs(855);
    layer2_outputs(1161) <= not(layer1_outputs(206));
    layer2_outputs(1162) <= '1';
    layer2_outputs(1163) <= not((layer1_outputs(1895)) and (layer1_outputs(781)));
    layer2_outputs(1164) <= not(layer1_outputs(1527)) or (layer1_outputs(243));
    layer2_outputs(1165) <= not(layer1_outputs(1599));
    layer2_outputs(1166) <= '1';
    layer2_outputs(1167) <= not((layer1_outputs(464)) and (layer1_outputs(820)));
    layer2_outputs(1168) <= layer1_outputs(381);
    layer2_outputs(1169) <= (layer1_outputs(322)) and (layer1_outputs(1223));
    layer2_outputs(1170) <= not(layer1_outputs(866));
    layer2_outputs(1171) <= not((layer1_outputs(1175)) or (layer1_outputs(721)));
    layer2_outputs(1172) <= layer1_outputs(511);
    layer2_outputs(1173) <= (layer1_outputs(752)) and not (layer1_outputs(1372));
    layer2_outputs(1174) <= layer1_outputs(1756);
    layer2_outputs(1175) <= '0';
    layer2_outputs(1176) <= not(layer1_outputs(600));
    layer2_outputs(1177) <= not(layer1_outputs(2066));
    layer2_outputs(1178) <= (layer1_outputs(2228)) or (layer1_outputs(1486));
    layer2_outputs(1179) <= '1';
    layer2_outputs(1180) <= '1';
    layer2_outputs(1181) <= layer1_outputs(131);
    layer2_outputs(1182) <= (layer1_outputs(2446)) xor (layer1_outputs(2061));
    layer2_outputs(1183) <= (layer1_outputs(420)) and not (layer1_outputs(680));
    layer2_outputs(1184) <= not(layer1_outputs(886)) or (layer1_outputs(210));
    layer2_outputs(1185) <= not(layer1_outputs(1721));
    layer2_outputs(1186) <= not(layer1_outputs(111)) or (layer1_outputs(266));
    layer2_outputs(1187) <= (layer1_outputs(607)) and not (layer1_outputs(1407));
    layer2_outputs(1188) <= (layer1_outputs(1169)) and (layer1_outputs(1217));
    layer2_outputs(1189) <= (layer1_outputs(1678)) and not (layer1_outputs(1716));
    layer2_outputs(1190) <= not((layer1_outputs(10)) and (layer1_outputs(352)));
    layer2_outputs(1191) <= '1';
    layer2_outputs(1192) <= not(layer1_outputs(2357));
    layer2_outputs(1193) <= layer1_outputs(533);
    layer2_outputs(1194) <= not(layer1_outputs(523)) or (layer1_outputs(866));
    layer2_outputs(1195) <= not((layer1_outputs(730)) and (layer1_outputs(962)));
    layer2_outputs(1196) <= layer1_outputs(2442);
    layer2_outputs(1197) <= (layer1_outputs(1170)) and not (layer1_outputs(2054));
    layer2_outputs(1198) <= not(layer1_outputs(1473));
    layer2_outputs(1199) <= (layer1_outputs(225)) or (layer1_outputs(2540));
    layer2_outputs(1200) <= layer1_outputs(2419);
    layer2_outputs(1201) <= layer1_outputs(1427);
    layer2_outputs(1202) <= not(layer1_outputs(199)) or (layer1_outputs(382));
    layer2_outputs(1203) <= '0';
    layer2_outputs(1204) <= not(layer1_outputs(107)) or (layer1_outputs(848));
    layer2_outputs(1205) <= '1';
    layer2_outputs(1206) <= not(layer1_outputs(1966));
    layer2_outputs(1207) <= '0';
    layer2_outputs(1208) <= not(layer1_outputs(1157)) or (layer1_outputs(2368));
    layer2_outputs(1209) <= not(layer1_outputs(944));
    layer2_outputs(1210) <= (layer1_outputs(2185)) and not (layer1_outputs(1654));
    layer2_outputs(1211) <= not(layer1_outputs(601));
    layer2_outputs(1212) <= layer1_outputs(1968);
    layer2_outputs(1213) <= (layer1_outputs(1513)) or (layer1_outputs(2512));
    layer2_outputs(1214) <= not(layer1_outputs(692));
    layer2_outputs(1215) <= (layer1_outputs(798)) and not (layer1_outputs(102));
    layer2_outputs(1216) <= (layer1_outputs(1276)) or (layer1_outputs(720));
    layer2_outputs(1217) <= (layer1_outputs(909)) and (layer1_outputs(1943));
    layer2_outputs(1218) <= not(layer1_outputs(484));
    layer2_outputs(1219) <= (layer1_outputs(468)) or (layer1_outputs(577));
    layer2_outputs(1220) <= '0';
    layer2_outputs(1221) <= (layer1_outputs(1130)) or (layer1_outputs(239));
    layer2_outputs(1222) <= not((layer1_outputs(2314)) and (layer1_outputs(1585)));
    layer2_outputs(1223) <= '0';
    layer2_outputs(1224) <= not(layer1_outputs(149)) or (layer1_outputs(992));
    layer2_outputs(1225) <= not(layer1_outputs(2195));
    layer2_outputs(1226) <= '1';
    layer2_outputs(1227) <= not(layer1_outputs(1420));
    layer2_outputs(1228) <= (layer1_outputs(1286)) and (layer1_outputs(380));
    layer2_outputs(1229) <= not(layer1_outputs(575));
    layer2_outputs(1230) <= not(layer1_outputs(1953));
    layer2_outputs(1231) <= not(layer1_outputs(1063));
    layer2_outputs(1232) <= not((layer1_outputs(1976)) or (layer1_outputs(1641)));
    layer2_outputs(1233) <= '1';
    layer2_outputs(1234) <= not(layer1_outputs(1858));
    layer2_outputs(1235) <= layer1_outputs(913);
    layer2_outputs(1236) <= not(layer1_outputs(2484));
    layer2_outputs(1237) <= not(layer1_outputs(701)) or (layer1_outputs(1077));
    layer2_outputs(1238) <= (layer1_outputs(1410)) and (layer1_outputs(2192));
    layer2_outputs(1239) <= layer1_outputs(2428);
    layer2_outputs(1240) <= not(layer1_outputs(1633));
    layer2_outputs(1241) <= not(layer1_outputs(1684));
    layer2_outputs(1242) <= (layer1_outputs(118)) and not (layer1_outputs(1748));
    layer2_outputs(1243) <= layer1_outputs(21);
    layer2_outputs(1244) <= not((layer1_outputs(509)) and (layer1_outputs(1304)));
    layer2_outputs(1245) <= not(layer1_outputs(2112));
    layer2_outputs(1246) <= '1';
    layer2_outputs(1247) <= layer1_outputs(265);
    layer2_outputs(1248) <= not((layer1_outputs(2028)) xor (layer1_outputs(2434)));
    layer2_outputs(1249) <= '0';
    layer2_outputs(1250) <= not(layer1_outputs(475));
    layer2_outputs(1251) <= not((layer1_outputs(2072)) or (layer1_outputs(1672)));
    layer2_outputs(1252) <= not(layer1_outputs(2407));
    layer2_outputs(1253) <= (layer1_outputs(1768)) and not (layer1_outputs(92));
    layer2_outputs(1254) <= not((layer1_outputs(1456)) or (layer1_outputs(2400)));
    layer2_outputs(1255) <= layer1_outputs(1164);
    layer2_outputs(1256) <= layer1_outputs(503);
    layer2_outputs(1257) <= not(layer1_outputs(1027));
    layer2_outputs(1258) <= layer1_outputs(1083);
    layer2_outputs(1259) <= not(layer1_outputs(2330)) or (layer1_outputs(635));
    layer2_outputs(1260) <= (layer1_outputs(830)) and not (layer1_outputs(490));
    layer2_outputs(1261) <= layer1_outputs(378);
    layer2_outputs(1262) <= '0';
    layer2_outputs(1263) <= (layer1_outputs(2077)) or (layer1_outputs(616));
    layer2_outputs(1264) <= not(layer1_outputs(1134));
    layer2_outputs(1265) <= (layer1_outputs(227)) and not (layer1_outputs(1724));
    layer2_outputs(1266) <= '1';
    layer2_outputs(1267) <= layer1_outputs(1076);
    layer2_outputs(1268) <= not(layer1_outputs(659));
    layer2_outputs(1269) <= (layer1_outputs(95)) or (layer1_outputs(2244));
    layer2_outputs(1270) <= not(layer1_outputs(2177)) or (layer1_outputs(445));
    layer2_outputs(1271) <= layer1_outputs(899);
    layer2_outputs(1272) <= layer1_outputs(785);
    layer2_outputs(1273) <= layer1_outputs(98);
    layer2_outputs(1274) <= (layer1_outputs(606)) and not (layer1_outputs(531));
    layer2_outputs(1275) <= layer1_outputs(660);
    layer2_outputs(1276) <= (layer1_outputs(700)) and not (layer1_outputs(991));
    layer2_outputs(1277) <= (layer1_outputs(1839)) and not (layer1_outputs(2113));
    layer2_outputs(1278) <= layer1_outputs(1786);
    layer2_outputs(1279) <= not((layer1_outputs(2055)) or (layer1_outputs(2543)));
    layer2_outputs(1280) <= (layer1_outputs(550)) and not (layer1_outputs(104));
    layer2_outputs(1281) <= not(layer1_outputs(2118)) or (layer1_outputs(1584));
    layer2_outputs(1282) <= layer1_outputs(2180);
    layer2_outputs(1283) <= not(layer1_outputs(1490));
    layer2_outputs(1284) <= (layer1_outputs(703)) or (layer1_outputs(213));
    layer2_outputs(1285) <= (layer1_outputs(2154)) and not (layer1_outputs(572));
    layer2_outputs(1286) <= not(layer1_outputs(954)) or (layer1_outputs(749));
    layer2_outputs(1287) <= not((layer1_outputs(28)) or (layer1_outputs(2246)));
    layer2_outputs(1288) <= layer1_outputs(2052);
    layer2_outputs(1289) <= not(layer1_outputs(1519));
    layer2_outputs(1290) <= not(layer1_outputs(685));
    layer2_outputs(1291) <= layer1_outputs(1206);
    layer2_outputs(1292) <= not(layer1_outputs(862));
    layer2_outputs(1293) <= '0';
    layer2_outputs(1294) <= (layer1_outputs(63)) and (layer1_outputs(2322));
    layer2_outputs(1295) <= layer1_outputs(1613);
    layer2_outputs(1296) <= (layer1_outputs(1203)) and not (layer1_outputs(377));
    layer2_outputs(1297) <= (layer1_outputs(832)) or (layer1_outputs(2123));
    layer2_outputs(1298) <= not(layer1_outputs(942)) or (layer1_outputs(2418));
    layer2_outputs(1299) <= not(layer1_outputs(1138)) or (layer1_outputs(535));
    layer2_outputs(1300) <= '1';
    layer2_outputs(1301) <= (layer1_outputs(1657)) or (layer1_outputs(2316));
    layer2_outputs(1302) <= (layer1_outputs(1546)) or (layer1_outputs(75));
    layer2_outputs(1303) <= not(layer1_outputs(1290));
    layer2_outputs(1304) <= layer1_outputs(1722);
    layer2_outputs(1305) <= not((layer1_outputs(2455)) and (layer1_outputs(297)));
    layer2_outputs(1306) <= (layer1_outputs(2464)) and not (layer1_outputs(579));
    layer2_outputs(1307) <= (layer1_outputs(1728)) and (layer1_outputs(1266));
    layer2_outputs(1308) <= '0';
    layer2_outputs(1309) <= not(layer1_outputs(1060));
    layer2_outputs(1310) <= not(layer1_outputs(1210));
    layer2_outputs(1311) <= not((layer1_outputs(2014)) and (layer1_outputs(246)));
    layer2_outputs(1312) <= '0';
    layer2_outputs(1313) <= layer1_outputs(787);
    layer2_outputs(1314) <= not((layer1_outputs(688)) or (layer1_outputs(2283)));
    layer2_outputs(1315) <= not(layer1_outputs(602)) or (layer1_outputs(1207));
    layer2_outputs(1316) <= (layer1_outputs(580)) and not (layer1_outputs(1644));
    layer2_outputs(1317) <= (layer1_outputs(112)) and not (layer1_outputs(367));
    layer2_outputs(1318) <= not(layer1_outputs(1471)) or (layer1_outputs(1281));
    layer2_outputs(1319) <= (layer1_outputs(1988)) and not (layer1_outputs(2076));
    layer2_outputs(1320) <= not(layer1_outputs(1450)) or (layer1_outputs(1910));
    layer2_outputs(1321) <= not(layer1_outputs(841));
    layer2_outputs(1322) <= not(layer1_outputs(347));
    layer2_outputs(1323) <= '1';
    layer2_outputs(1324) <= (layer1_outputs(871)) and (layer1_outputs(1352));
    layer2_outputs(1325) <= (layer1_outputs(1413)) and not (layer1_outputs(2059));
    layer2_outputs(1326) <= layer1_outputs(1008);
    layer2_outputs(1327) <= not(layer1_outputs(2494)) or (layer1_outputs(1335));
    layer2_outputs(1328) <= not(layer1_outputs(811)) or (layer1_outputs(1699));
    layer2_outputs(1329) <= not(layer1_outputs(2026));
    layer2_outputs(1330) <= layer1_outputs(845);
    layer2_outputs(1331) <= not(layer1_outputs(340));
    layer2_outputs(1332) <= not(layer1_outputs(249)) or (layer1_outputs(704));
    layer2_outputs(1333) <= not(layer1_outputs(330)) or (layer1_outputs(244));
    layer2_outputs(1334) <= not(layer1_outputs(1252)) or (layer1_outputs(870));
    layer2_outputs(1335) <= not(layer1_outputs(2165));
    layer2_outputs(1336) <= not(layer1_outputs(790));
    layer2_outputs(1337) <= not((layer1_outputs(2400)) xor (layer1_outputs(1541)));
    layer2_outputs(1338) <= layer1_outputs(2110);
    layer2_outputs(1339) <= not(layer1_outputs(1294)) or (layer1_outputs(430));
    layer2_outputs(1340) <= '0';
    layer2_outputs(1341) <= '0';
    layer2_outputs(1342) <= not(layer1_outputs(1198));
    layer2_outputs(1343) <= layer1_outputs(1135);
    layer2_outputs(1344) <= '1';
    layer2_outputs(1345) <= layer1_outputs(1714);
    layer2_outputs(1346) <= not((layer1_outputs(1766)) and (layer1_outputs(694)));
    layer2_outputs(1347) <= (layer1_outputs(2086)) and not (layer1_outputs(263));
    layer2_outputs(1348) <= layer1_outputs(1648);
    layer2_outputs(1349) <= layer1_outputs(1382);
    layer2_outputs(1350) <= layer1_outputs(2480);
    layer2_outputs(1351) <= (layer1_outputs(764)) and not (layer1_outputs(105));
    layer2_outputs(1352) <= not(layer1_outputs(874));
    layer2_outputs(1353) <= not(layer1_outputs(23)) or (layer1_outputs(2099));
    layer2_outputs(1354) <= (layer1_outputs(103)) and not (layer1_outputs(87));
    layer2_outputs(1355) <= not(layer1_outputs(426)) or (layer1_outputs(1437));
    layer2_outputs(1356) <= layer1_outputs(2018);
    layer2_outputs(1357) <= (layer1_outputs(1854)) and not (layer1_outputs(1116));
    layer2_outputs(1358) <= (layer1_outputs(510)) and not (layer1_outputs(2055));
    layer2_outputs(1359) <= not(layer1_outputs(1764)) or (layer1_outputs(635));
    layer2_outputs(1360) <= '1';
    layer2_outputs(1361) <= (layer1_outputs(2429)) and (layer1_outputs(2414));
    layer2_outputs(1362) <= not(layer1_outputs(1631));
    layer2_outputs(1363) <= '0';
    layer2_outputs(1364) <= (layer1_outputs(172)) and not (layer1_outputs(1075));
    layer2_outputs(1365) <= not((layer1_outputs(719)) or (layer1_outputs(311)));
    layer2_outputs(1366) <= not((layer1_outputs(275)) and (layer1_outputs(819)));
    layer2_outputs(1367) <= not(layer1_outputs(139));
    layer2_outputs(1368) <= layer1_outputs(1796);
    layer2_outputs(1369) <= (layer1_outputs(1454)) and not (layer1_outputs(80));
    layer2_outputs(1370) <= (layer1_outputs(376)) and (layer1_outputs(1332));
    layer2_outputs(1371) <= layer1_outputs(783);
    layer2_outputs(1372) <= not((layer1_outputs(1225)) or (layer1_outputs(552)));
    layer2_outputs(1373) <= not(layer1_outputs(229));
    layer2_outputs(1374) <= layer1_outputs(174);
    layer2_outputs(1375) <= not((layer1_outputs(45)) or (layer1_outputs(718)));
    layer2_outputs(1376) <= not(layer1_outputs(505)) or (layer1_outputs(1162));
    layer2_outputs(1377) <= (layer1_outputs(441)) and not (layer1_outputs(581));
    layer2_outputs(1378) <= layer1_outputs(259);
    layer2_outputs(1379) <= not(layer1_outputs(739)) or (layer1_outputs(2101));
    layer2_outputs(1380) <= (layer1_outputs(1075)) or (layer1_outputs(1301));
    layer2_outputs(1381) <= layer1_outputs(382);
    layer2_outputs(1382) <= not((layer1_outputs(1315)) and (layer1_outputs(689)));
    layer2_outputs(1383) <= '0';
    layer2_outputs(1384) <= not(layer1_outputs(2062));
    layer2_outputs(1385) <= (layer1_outputs(492)) and (layer1_outputs(264));
    layer2_outputs(1386) <= '1';
    layer2_outputs(1387) <= (layer1_outputs(238)) xor (layer1_outputs(1904));
    layer2_outputs(1388) <= not(layer1_outputs(2441));
    layer2_outputs(1389) <= (layer1_outputs(1914)) and not (layer1_outputs(1833));
    layer2_outputs(1390) <= not(layer1_outputs(1753));
    layer2_outputs(1391) <= not(layer1_outputs(704)) or (layer1_outputs(2334));
    layer2_outputs(1392) <= not(layer1_outputs(1503));
    layer2_outputs(1393) <= layer1_outputs(2184);
    layer2_outputs(1394) <= not((layer1_outputs(455)) or (layer1_outputs(2297)));
    layer2_outputs(1395) <= not(layer1_outputs(2498)) or (layer1_outputs(740));
    layer2_outputs(1396) <= '1';
    layer2_outputs(1397) <= not(layer1_outputs(2188)) or (layer1_outputs(312));
    layer2_outputs(1398) <= (layer1_outputs(1890)) and not (layer1_outputs(2079));
    layer2_outputs(1399) <= (layer1_outputs(1201)) and not (layer1_outputs(1942));
    layer2_outputs(1400) <= not(layer1_outputs(186)) or (layer1_outputs(45));
    layer2_outputs(1401) <= (layer1_outputs(37)) and not (layer1_outputs(1723));
    layer2_outputs(1402) <= not((layer1_outputs(604)) or (layer1_outputs(1653)));
    layer2_outputs(1403) <= not(layer1_outputs(118)) or (layer1_outputs(713));
    layer2_outputs(1404) <= not(layer1_outputs(1099));
    layer2_outputs(1405) <= layer1_outputs(2211);
    layer2_outputs(1406) <= not((layer1_outputs(2469)) or (layer1_outputs(62)));
    layer2_outputs(1407) <= '0';
    layer2_outputs(1408) <= '0';
    layer2_outputs(1409) <= not((layer1_outputs(100)) or (layer1_outputs(1562)));
    layer2_outputs(1410) <= '0';
    layer2_outputs(1411) <= not((layer1_outputs(1257)) or (layer1_outputs(1839)));
    layer2_outputs(1412) <= not((layer1_outputs(595)) xor (layer1_outputs(1183)));
    layer2_outputs(1413) <= not(layer1_outputs(181));
    layer2_outputs(1414) <= not(layer1_outputs(716));
    layer2_outputs(1415) <= not(layer1_outputs(365)) or (layer1_outputs(232));
    layer2_outputs(1416) <= (layer1_outputs(1467)) and not (layer1_outputs(221));
    layer2_outputs(1417) <= not((layer1_outputs(2166)) and (layer1_outputs(2288)));
    layer2_outputs(1418) <= layer1_outputs(646);
    layer2_outputs(1419) <= layer1_outputs(1843);
    layer2_outputs(1420) <= not((layer1_outputs(1048)) and (layer1_outputs(616)));
    layer2_outputs(1421) <= not(layer1_outputs(1056));
    layer2_outputs(1422) <= layer1_outputs(2201);
    layer2_outputs(1423) <= layer1_outputs(2515);
    layer2_outputs(1424) <= (layer1_outputs(1177)) or (layer1_outputs(1087));
    layer2_outputs(1425) <= not(layer1_outputs(2002));
    layer2_outputs(1426) <= layer1_outputs(1475);
    layer2_outputs(1427) <= not(layer1_outputs(334)) or (layer1_outputs(2273));
    layer2_outputs(1428) <= not((layer1_outputs(708)) and (layer1_outputs(344)));
    layer2_outputs(1429) <= (layer1_outputs(2103)) and not (layer1_outputs(539));
    layer2_outputs(1430) <= '0';
    layer2_outputs(1431) <= not(layer1_outputs(1967)) or (layer1_outputs(2490));
    layer2_outputs(1432) <= '1';
    layer2_outputs(1433) <= not(layer1_outputs(2275));
    layer2_outputs(1434) <= not(layer1_outputs(261)) or (layer1_outputs(1609));
    layer2_outputs(1435) <= not((layer1_outputs(2276)) xor (layer1_outputs(1754)));
    layer2_outputs(1436) <= not(layer1_outputs(728));
    layer2_outputs(1437) <= not((layer1_outputs(369)) and (layer1_outputs(1535)));
    layer2_outputs(1438) <= not(layer1_outputs(53));
    layer2_outputs(1439) <= not((layer1_outputs(1822)) and (layer1_outputs(2271)));
    layer2_outputs(1440) <= not(layer1_outputs(565)) or (layer1_outputs(1466));
    layer2_outputs(1441) <= '1';
    layer2_outputs(1442) <= not((layer1_outputs(571)) and (layer1_outputs(2385)));
    layer2_outputs(1443) <= layer1_outputs(1775);
    layer2_outputs(1444) <= not((layer1_outputs(163)) or (layer1_outputs(1214)));
    layer2_outputs(1445) <= '0';
    layer2_outputs(1446) <= not(layer1_outputs(384));
    layer2_outputs(1447) <= '0';
    layer2_outputs(1448) <= not((layer1_outputs(1543)) and (layer1_outputs(2197)));
    layer2_outputs(1449) <= not(layer1_outputs(943));
    layer2_outputs(1450) <= (layer1_outputs(913)) or (layer1_outputs(1394));
    layer2_outputs(1451) <= not(layer1_outputs(437));
    layer2_outputs(1452) <= layer1_outputs(1711);
    layer2_outputs(1453) <= not(layer1_outputs(1211));
    layer2_outputs(1454) <= layer1_outputs(701);
    layer2_outputs(1455) <= '0';
    layer2_outputs(1456) <= layer1_outputs(2125);
    layer2_outputs(1457) <= not(layer1_outputs(881));
    layer2_outputs(1458) <= not(layer1_outputs(1909)) or (layer1_outputs(1313));
    layer2_outputs(1459) <= layer1_outputs(1132);
    layer2_outputs(1460) <= (layer1_outputs(1003)) and (layer1_outputs(1093));
    layer2_outputs(1461) <= layer1_outputs(2483);
    layer2_outputs(1462) <= '1';
    layer2_outputs(1463) <= '0';
    layer2_outputs(1464) <= (layer1_outputs(1697)) and (layer1_outputs(1583));
    layer2_outputs(1465) <= (layer1_outputs(1734)) and not (layer1_outputs(488));
    layer2_outputs(1466) <= (layer1_outputs(925)) and not (layer1_outputs(566));
    layer2_outputs(1467) <= '1';
    layer2_outputs(1468) <= not(layer1_outputs(2332));
    layer2_outputs(1469) <= not((layer1_outputs(383)) and (layer1_outputs(1905)));
    layer2_outputs(1470) <= not(layer1_outputs(778)) or (layer1_outputs(1538));
    layer2_outputs(1471) <= not(layer1_outputs(1618));
    layer2_outputs(1472) <= (layer1_outputs(2182)) and not (layer1_outputs(1550));
    layer2_outputs(1473) <= not(layer1_outputs(1212));
    layer2_outputs(1474) <= not(layer1_outputs(1176));
    layer2_outputs(1475) <= layer1_outputs(2217);
    layer2_outputs(1476) <= not(layer1_outputs(551)) or (layer1_outputs(218));
    layer2_outputs(1477) <= not(layer1_outputs(723)) or (layer1_outputs(1559));
    layer2_outputs(1478) <= (layer1_outputs(241)) and not (layer1_outputs(622));
    layer2_outputs(1479) <= '1';
    layer2_outputs(1480) <= (layer1_outputs(195)) and (layer1_outputs(537));
    layer2_outputs(1481) <= not(layer1_outputs(2474));
    layer2_outputs(1482) <= layer1_outputs(2506);
    layer2_outputs(1483) <= (layer1_outputs(534)) and not (layer1_outputs(757));
    layer2_outputs(1484) <= '1';
    layer2_outputs(1485) <= not(layer1_outputs(1750));
    layer2_outputs(1486) <= '0';
    layer2_outputs(1487) <= not((layer1_outputs(956)) xor (layer1_outputs(499)));
    layer2_outputs(1488) <= (layer1_outputs(277)) and (layer1_outputs(275));
    layer2_outputs(1489) <= (layer1_outputs(2309)) and not (layer1_outputs(1684));
    layer2_outputs(1490) <= layer1_outputs(2026);
    layer2_outputs(1491) <= layer1_outputs(116);
    layer2_outputs(1492) <= not(layer1_outputs(715)) or (layer1_outputs(1243));
    layer2_outputs(1493) <= not(layer1_outputs(1757));
    layer2_outputs(1494) <= layer1_outputs(1177);
    layer2_outputs(1495) <= (layer1_outputs(2341)) and (layer1_outputs(1301));
    layer2_outputs(1496) <= '0';
    layer2_outputs(1497) <= not(layer1_outputs(1563));
    layer2_outputs(1498) <= not((layer1_outputs(1461)) and (layer1_outputs(1453)));
    layer2_outputs(1499) <= (layer1_outputs(2473)) and not (layer1_outputs(1927));
    layer2_outputs(1500) <= not((layer1_outputs(1883)) and (layer1_outputs(914)));
    layer2_outputs(1501) <= layer1_outputs(960);
    layer2_outputs(1502) <= not(layer1_outputs(497));
    layer2_outputs(1503) <= not(layer1_outputs(2243));
    layer2_outputs(1504) <= (layer1_outputs(758)) and not (layer1_outputs(129));
    layer2_outputs(1505) <= layer1_outputs(613);
    layer2_outputs(1506) <= not(layer1_outputs(1973));
    layer2_outputs(1507) <= layer1_outputs(2038);
    layer2_outputs(1508) <= (layer1_outputs(919)) and (layer1_outputs(1532));
    layer2_outputs(1509) <= layer1_outputs(1917);
    layer2_outputs(1510) <= not(layer1_outputs(2518));
    layer2_outputs(1511) <= layer1_outputs(2263);
    layer2_outputs(1512) <= not(layer1_outputs(698));
    layer2_outputs(1513) <= (layer1_outputs(200)) and not (layer1_outputs(2214));
    layer2_outputs(1514) <= (layer1_outputs(2470)) and not (layer1_outputs(14));
    layer2_outputs(1515) <= layer1_outputs(42);
    layer2_outputs(1516) <= not(layer1_outputs(357)) or (layer1_outputs(2000));
    layer2_outputs(1517) <= not(layer1_outputs(1866));
    layer2_outputs(1518) <= not((layer1_outputs(1601)) and (layer1_outputs(702)));
    layer2_outputs(1519) <= layer1_outputs(2491);
    layer2_outputs(1520) <= (layer1_outputs(2552)) or (layer1_outputs(43));
    layer2_outputs(1521) <= not((layer1_outputs(824)) xor (layer1_outputs(365)));
    layer2_outputs(1522) <= (layer1_outputs(1696)) or (layer1_outputs(515));
    layer2_outputs(1523) <= '0';
    layer2_outputs(1524) <= '0';
    layer2_outputs(1525) <= '0';
    layer2_outputs(1526) <= not((layer1_outputs(1593)) and (layer1_outputs(828)));
    layer2_outputs(1527) <= not(layer1_outputs(1289));
    layer2_outputs(1528) <= layer1_outputs(14);
    layer2_outputs(1529) <= (layer1_outputs(1202)) and not (layer1_outputs(1784));
    layer2_outputs(1530) <= layer1_outputs(1364);
    layer2_outputs(1531) <= not((layer1_outputs(1338)) and (layer1_outputs(1738)));
    layer2_outputs(1532) <= (layer1_outputs(1086)) and not (layer1_outputs(1918));
    layer2_outputs(1533) <= (layer1_outputs(2372)) and not (layer1_outputs(1202));
    layer2_outputs(1534) <= not(layer1_outputs(1655));
    layer2_outputs(1535) <= (layer1_outputs(542)) and (layer1_outputs(1417));
    layer2_outputs(1536) <= not((layer1_outputs(1595)) or (layer1_outputs(1479)));
    layer2_outputs(1537) <= (layer1_outputs(72)) and (layer1_outputs(88));
    layer2_outputs(1538) <= layer1_outputs(988);
    layer2_outputs(1539) <= not(layer1_outputs(1343));
    layer2_outputs(1540) <= not((layer1_outputs(1002)) or (layer1_outputs(2350)));
    layer2_outputs(1541) <= not(layer1_outputs(587)) or (layer1_outputs(2210));
    layer2_outputs(1542) <= layer1_outputs(783);
    layer2_outputs(1543) <= '1';
    layer2_outputs(1544) <= layer1_outputs(1798);
    layer2_outputs(1545) <= not(layer1_outputs(2344)) or (layer1_outputs(1833));
    layer2_outputs(1546) <= (layer1_outputs(1119)) and not (layer1_outputs(773));
    layer2_outputs(1547) <= (layer1_outputs(845)) or (layer1_outputs(175));
    layer2_outputs(1548) <= layer1_outputs(1250);
    layer2_outputs(1549) <= layer1_outputs(695);
    layer2_outputs(1550) <= layer1_outputs(645);
    layer2_outputs(1551) <= '1';
    layer2_outputs(1552) <= not((layer1_outputs(363)) and (layer1_outputs(1184)));
    layer2_outputs(1553) <= '0';
    layer2_outputs(1554) <= not(layer1_outputs(978));
    layer2_outputs(1555) <= '0';
    layer2_outputs(1556) <= layer1_outputs(42);
    layer2_outputs(1557) <= not((layer1_outputs(658)) and (layer1_outputs(1515)));
    layer2_outputs(1558) <= (layer1_outputs(1533)) or (layer1_outputs(164));
    layer2_outputs(1559) <= layer1_outputs(2485);
    layer2_outputs(1560) <= not(layer1_outputs(730));
    layer2_outputs(1561) <= (layer1_outputs(1373)) and not (layer1_outputs(1372));
    layer2_outputs(1562) <= '1';
    layer2_outputs(1563) <= (layer1_outputs(255)) and (layer1_outputs(1664));
    layer2_outputs(1564) <= not((layer1_outputs(1906)) or (layer1_outputs(240)));
    layer2_outputs(1565) <= (layer1_outputs(2063)) and not (layer1_outputs(2550));
    layer2_outputs(1566) <= not((layer1_outputs(1853)) and (layer1_outputs(466)));
    layer2_outputs(1567) <= (layer1_outputs(1626)) and (layer1_outputs(989));
    layer2_outputs(1568) <= '0';
    layer2_outputs(1569) <= not(layer1_outputs(864)) or (layer1_outputs(1690));
    layer2_outputs(1570) <= layer1_outputs(2425);
    layer2_outputs(1571) <= layer1_outputs(2246);
    layer2_outputs(1572) <= not((layer1_outputs(632)) or (layer1_outputs(1170)));
    layer2_outputs(1573) <= not((layer1_outputs(742)) and (layer1_outputs(1484)));
    layer2_outputs(1574) <= not(layer1_outputs(1908));
    layer2_outputs(1575) <= (layer1_outputs(1195)) or (layer1_outputs(1812));
    layer2_outputs(1576) <= not(layer1_outputs(768));
    layer2_outputs(1577) <= (layer1_outputs(1295)) or (layer1_outputs(2411));
    layer2_outputs(1578) <= layer1_outputs(1405);
    layer2_outputs(1579) <= (layer1_outputs(2469)) or (layer1_outputs(1352));
    layer2_outputs(1580) <= not((layer1_outputs(1007)) and (layer1_outputs(1831)));
    layer2_outputs(1581) <= not(layer1_outputs(2249)) or (layer1_outputs(1641));
    layer2_outputs(1582) <= not(layer1_outputs(1647)) or (layer1_outputs(1194));
    layer2_outputs(1583) <= layer1_outputs(427);
    layer2_outputs(1584) <= layer1_outputs(308);
    layer2_outputs(1585) <= not(layer1_outputs(1196)) or (layer1_outputs(2076));
    layer2_outputs(1586) <= '0';
    layer2_outputs(1587) <= not((layer1_outputs(950)) and (layer1_outputs(1744)));
    layer2_outputs(1588) <= (layer1_outputs(2408)) and (layer1_outputs(2373));
    layer2_outputs(1589) <= (layer1_outputs(209)) or (layer1_outputs(2093));
    layer2_outputs(1590) <= not(layer1_outputs(2356));
    layer2_outputs(1591) <= '0';
    layer2_outputs(1592) <= not((layer1_outputs(398)) or (layer1_outputs(63)));
    layer2_outputs(1593) <= (layer1_outputs(986)) or (layer1_outputs(1577));
    layer2_outputs(1594) <= not((layer1_outputs(1847)) or (layer1_outputs(1636)));
    layer2_outputs(1595) <= (layer1_outputs(990)) and not (layer1_outputs(2237));
    layer2_outputs(1596) <= not(layer1_outputs(1226)) or (layer1_outputs(1221));
    layer2_outputs(1597) <= not(layer1_outputs(2554));
    layer2_outputs(1598) <= not(layer1_outputs(2138));
    layer2_outputs(1599) <= '0';
    layer2_outputs(1600) <= '1';
    layer2_outputs(1601) <= not((layer1_outputs(8)) and (layer1_outputs(1548)));
    layer2_outputs(1602) <= (layer1_outputs(1823)) and not (layer1_outputs(1052));
    layer2_outputs(1603) <= (layer1_outputs(121)) and not (layer1_outputs(70));
    layer2_outputs(1604) <= not((layer1_outputs(1287)) or (layer1_outputs(2074)));
    layer2_outputs(1605) <= not((layer1_outputs(1908)) or (layer1_outputs(2057)));
    layer2_outputs(1606) <= layer1_outputs(596);
    layer2_outputs(1607) <= not(layer1_outputs(1229));
    layer2_outputs(1608) <= layer1_outputs(1195);
    layer2_outputs(1609) <= not(layer1_outputs(855)) or (layer1_outputs(321));
    layer2_outputs(1610) <= layer1_outputs(1907);
    layer2_outputs(1611) <= (layer1_outputs(2390)) and not (layer1_outputs(1585));
    layer2_outputs(1612) <= layer1_outputs(451);
    layer2_outputs(1613) <= layer1_outputs(573);
    layer2_outputs(1614) <= (layer1_outputs(452)) and (layer1_outputs(1972));
    layer2_outputs(1615) <= '1';
    layer2_outputs(1616) <= (layer1_outputs(1447)) or (layer1_outputs(1587));
    layer2_outputs(1617) <= (layer1_outputs(1898)) or (layer1_outputs(1610));
    layer2_outputs(1618) <= layer1_outputs(2368);
    layer2_outputs(1619) <= layer1_outputs(438);
    layer2_outputs(1620) <= not(layer1_outputs(686)) or (layer1_outputs(2138));
    layer2_outputs(1621) <= (layer1_outputs(2165)) or (layer1_outputs(1828));
    layer2_outputs(1622) <= layer1_outputs(2205);
    layer2_outputs(1623) <= layer1_outputs(543);
    layer2_outputs(1624) <= layer1_outputs(1061);
    layer2_outputs(1625) <= not(layer1_outputs(309));
    layer2_outputs(1626) <= not(layer1_outputs(1959));
    layer2_outputs(1627) <= '1';
    layer2_outputs(1628) <= not(layer1_outputs(1235));
    layer2_outputs(1629) <= '1';
    layer2_outputs(1630) <= layer1_outputs(983);
    layer2_outputs(1631) <= '0';
    layer2_outputs(1632) <= layer1_outputs(1438);
    layer2_outputs(1633) <= not(layer1_outputs(1015));
    layer2_outputs(1634) <= not(layer1_outputs(1027)) or (layer1_outputs(1789));
    layer2_outputs(1635) <= (layer1_outputs(2139)) and (layer1_outputs(1731));
    layer2_outputs(1636) <= not((layer1_outputs(226)) or (layer1_outputs(557)));
    layer2_outputs(1637) <= layer1_outputs(1730);
    layer2_outputs(1638) <= layer1_outputs(2042);
    layer2_outputs(1639) <= (layer1_outputs(135)) and not (layer1_outputs(869));
    layer2_outputs(1640) <= not(layer1_outputs(2520));
    layer2_outputs(1641) <= (layer1_outputs(1686)) and (layer1_outputs(405));
    layer2_outputs(1642) <= layer1_outputs(1189);
    layer2_outputs(1643) <= not((layer1_outputs(1480)) and (layer1_outputs(2183)));
    layer2_outputs(1644) <= (layer1_outputs(556)) and not (layer1_outputs(1781));
    layer2_outputs(1645) <= (layer1_outputs(1887)) and not (layer1_outputs(1461));
    layer2_outputs(1646) <= '1';
    layer2_outputs(1647) <= (layer1_outputs(181)) and (layer1_outputs(187));
    layer2_outputs(1648) <= not((layer1_outputs(524)) or (layer1_outputs(1235)));
    layer2_outputs(1649) <= not(layer1_outputs(2253)) or (layer1_outputs(2430));
    layer2_outputs(1650) <= not((layer1_outputs(1533)) or (layer1_outputs(1912)));
    layer2_outputs(1651) <= (layer1_outputs(2463)) and not (layer1_outputs(2048));
    layer2_outputs(1652) <= not(layer1_outputs(202));
    layer2_outputs(1653) <= not((layer1_outputs(1398)) and (layer1_outputs(489)));
    layer2_outputs(1654) <= '0';
    layer2_outputs(1655) <= layer1_outputs(113);
    layer2_outputs(1656) <= '0';
    layer2_outputs(1657) <= not(layer1_outputs(1510));
    layer2_outputs(1658) <= layer1_outputs(788);
    layer2_outputs(1659) <= not(layer1_outputs(1972));
    layer2_outputs(1660) <= '1';
    layer2_outputs(1661) <= (layer1_outputs(48)) and not (layer1_outputs(614));
    layer2_outputs(1662) <= (layer1_outputs(1857)) and (layer1_outputs(589));
    layer2_outputs(1663) <= (layer1_outputs(900)) and not (layer1_outputs(2073));
    layer2_outputs(1664) <= layer1_outputs(2452);
    layer2_outputs(1665) <= not(layer1_outputs(2454));
    layer2_outputs(1666) <= not(layer1_outputs(450)) or (layer1_outputs(41));
    layer2_outputs(1667) <= not(layer1_outputs(1376));
    layer2_outputs(1668) <= '0';
    layer2_outputs(1669) <= (layer1_outputs(54)) and not (layer1_outputs(1392));
    layer2_outputs(1670) <= (layer1_outputs(1127)) and not (layer1_outputs(2342));
    layer2_outputs(1671) <= not(layer1_outputs(2255));
    layer2_outputs(1672) <= (layer1_outputs(59)) or (layer1_outputs(1709));
    layer2_outputs(1673) <= not(layer1_outputs(2005)) or (layer1_outputs(1995));
    layer2_outputs(1674) <= layer1_outputs(1920);
    layer2_outputs(1675) <= layer1_outputs(2316);
    layer2_outputs(1676) <= layer1_outputs(2174);
    layer2_outputs(1677) <= not(layer1_outputs(1619)) or (layer1_outputs(1655));
    layer2_outputs(1678) <= not(layer1_outputs(833));
    layer2_outputs(1679) <= not(layer1_outputs(2095));
    layer2_outputs(1680) <= (layer1_outputs(1671)) or (layer1_outputs(1047));
    layer2_outputs(1681) <= '0';
    layer2_outputs(1682) <= not(layer1_outputs(1779));
    layer2_outputs(1683) <= not(layer1_outputs(2438)) or (layer1_outputs(1815));
    layer2_outputs(1684) <= (layer1_outputs(930)) and not (layer1_outputs(2287));
    layer2_outputs(1685) <= not(layer1_outputs(2179)) or (layer1_outputs(563));
    layer2_outputs(1686) <= not(layer1_outputs(1148));
    layer2_outputs(1687) <= (layer1_outputs(1188)) and (layer1_outputs(2456));
    layer2_outputs(1688) <= layer1_outputs(1761);
    layer2_outputs(1689) <= layer1_outputs(295);
    layer2_outputs(1690) <= not(layer1_outputs(1634)) or (layer1_outputs(2477));
    layer2_outputs(1691) <= layer1_outputs(878);
    layer2_outputs(1692) <= (layer1_outputs(1180)) and not (layer1_outputs(1670));
    layer2_outputs(1693) <= not(layer1_outputs(1898));
    layer2_outputs(1694) <= not((layer1_outputs(2114)) and (layer1_outputs(2312)));
    layer2_outputs(1695) <= not(layer1_outputs(709));
    layer2_outputs(1696) <= '0';
    layer2_outputs(1697) <= (layer1_outputs(561)) and (layer1_outputs(2529));
    layer2_outputs(1698) <= not(layer1_outputs(38)) or (layer1_outputs(73));
    layer2_outputs(1699) <= not(layer1_outputs(754));
    layer2_outputs(1700) <= layer1_outputs(826);
    layer2_outputs(1701) <= not((layer1_outputs(2493)) or (layer1_outputs(1292)));
    layer2_outputs(1702) <= not((layer1_outputs(2009)) or (layer1_outputs(1920)));
    layer2_outputs(1703) <= not((layer1_outputs(1886)) and (layer1_outputs(1354)));
    layer2_outputs(1704) <= not(layer1_outputs(1397)) or (layer1_outputs(2433));
    layer2_outputs(1705) <= (layer1_outputs(301)) and not (layer1_outputs(1555));
    layer2_outputs(1706) <= layer1_outputs(412);
    layer2_outputs(1707) <= not(layer1_outputs(1959));
    layer2_outputs(1708) <= not(layer1_outputs(396));
    layer2_outputs(1709) <= (layer1_outputs(1101)) and not (layer1_outputs(1492));
    layer2_outputs(1710) <= not(layer1_outputs(1541)) or (layer1_outputs(211));
    layer2_outputs(1711) <= (layer1_outputs(153)) and not (layer1_outputs(2339));
    layer2_outputs(1712) <= '0';
    layer2_outputs(1713) <= '1';
    layer2_outputs(1714) <= (layer1_outputs(415)) xor (layer1_outputs(672));
    layer2_outputs(1715) <= (layer1_outputs(2205)) and (layer1_outputs(746));
    layer2_outputs(1716) <= not(layer1_outputs(1246));
    layer2_outputs(1717) <= layer1_outputs(683);
    layer2_outputs(1718) <= layer1_outputs(284);
    layer2_outputs(1719) <= not(layer1_outputs(2517));
    layer2_outputs(1720) <= not((layer1_outputs(2208)) and (layer1_outputs(99)));
    layer2_outputs(1721) <= not(layer1_outputs(2081));
    layer2_outputs(1722) <= not(layer1_outputs(1006)) or (layer1_outputs(1016));
    layer2_outputs(1723) <= layer1_outputs(153);
    layer2_outputs(1724) <= layer1_outputs(1863);
    layer2_outputs(1725) <= not(layer1_outputs(1881));
    layer2_outputs(1726) <= not(layer1_outputs(1875)) or (layer1_outputs(1118));
    layer2_outputs(1727) <= layer1_outputs(1156);
    layer2_outputs(1728) <= not(layer1_outputs(157)) or (layer1_outputs(605));
    layer2_outputs(1729) <= layer1_outputs(1337);
    layer2_outputs(1730) <= not(layer1_outputs(2462)) or (layer1_outputs(1404));
    layer2_outputs(1731) <= layer1_outputs(290);
    layer2_outputs(1732) <= layer1_outputs(1913);
    layer2_outputs(1733) <= layer1_outputs(1409);
    layer2_outputs(1734) <= not(layer1_outputs(1623));
    layer2_outputs(1735) <= (layer1_outputs(1477)) xor (layer1_outputs(2259));
    layer2_outputs(1736) <= '0';
    layer2_outputs(1737) <= not(layer1_outputs(2313)) or (layer1_outputs(123));
    layer2_outputs(1738) <= not(layer1_outputs(196));
    layer2_outputs(1739) <= not(layer1_outputs(805));
    layer2_outputs(1740) <= layer1_outputs(2377);
    layer2_outputs(1741) <= '1';
    layer2_outputs(1742) <= (layer1_outputs(1569)) and not (layer1_outputs(1873));
    layer2_outputs(1743) <= not(layer1_outputs(1700)) or (layer1_outputs(1038));
    layer2_outputs(1744) <= (layer1_outputs(626)) and (layer1_outputs(2466));
    layer2_outputs(1745) <= layer1_outputs(85);
    layer2_outputs(1746) <= (layer1_outputs(1780)) or (layer1_outputs(108));
    layer2_outputs(1747) <= layer1_outputs(708);
    layer2_outputs(1748) <= not(layer1_outputs(1144)) or (layer1_outputs(67));
    layer2_outputs(1749) <= not(layer1_outputs(2427)) or (layer1_outputs(1540));
    layer2_outputs(1750) <= not((layer1_outputs(2253)) and (layer1_outputs(657)));
    layer2_outputs(1751) <= not(layer1_outputs(1091)) or (layer1_outputs(145));
    layer2_outputs(1752) <= not((layer1_outputs(527)) xor (layer1_outputs(1531)));
    layer2_outputs(1753) <= not(layer1_outputs(135)) or (layer1_outputs(60));
    layer2_outputs(1754) <= '0';
    layer2_outputs(1755) <= (layer1_outputs(793)) or (layer1_outputs(2149));
    layer2_outputs(1756) <= (layer1_outputs(2310)) and (layer1_outputs(1142));
    layer2_outputs(1757) <= not((layer1_outputs(1867)) and (layer1_outputs(540)));
    layer2_outputs(1758) <= not(layer1_outputs(1325)) or (layer1_outputs(1923));
    layer2_outputs(1759) <= layer1_outputs(355);
    layer2_outputs(1760) <= not(layer1_outputs(2102));
    layer2_outputs(1761) <= not(layer1_outputs(1296));
    layer2_outputs(1762) <= not((layer1_outputs(453)) and (layer1_outputs(720)));
    layer2_outputs(1763) <= (layer1_outputs(286)) and (layer1_outputs(404));
    layer2_outputs(1764) <= (layer1_outputs(1006)) and not (layer1_outputs(156));
    layer2_outputs(1765) <= layer1_outputs(2304);
    layer2_outputs(1766) <= not(layer1_outputs(2139)) or (layer1_outputs(1511));
    layer2_outputs(1767) <= (layer1_outputs(1139)) and (layer1_outputs(1878));
    layer2_outputs(1768) <= not(layer1_outputs(727));
    layer2_outputs(1769) <= (layer1_outputs(6)) or (layer1_outputs(1490));
    layer2_outputs(1770) <= not(layer1_outputs(46));
    layer2_outputs(1771) <= (layer1_outputs(1841)) and not (layer1_outputs(1725));
    layer2_outputs(1772) <= (layer1_outputs(2487)) and not (layer1_outputs(1046));
    layer2_outputs(1773) <= not(layer1_outputs(889));
    layer2_outputs(1774) <= not(layer1_outputs(865));
    layer2_outputs(1775) <= not(layer1_outputs(147));
    layer2_outputs(1776) <= (layer1_outputs(627)) xor (layer1_outputs(384));
    layer2_outputs(1777) <= (layer1_outputs(673)) or (layer1_outputs(757));
    layer2_outputs(1778) <= '1';
    layer2_outputs(1779) <= (layer1_outputs(2297)) and not (layer1_outputs(252));
    layer2_outputs(1780) <= not(layer1_outputs(1283));
    layer2_outputs(1781) <= not(layer1_outputs(1800)) or (layer1_outputs(1079));
    layer2_outputs(1782) <= '1';
    layer2_outputs(1783) <= (layer1_outputs(905)) xor (layer1_outputs(980));
    layer2_outputs(1784) <= '1';
    layer2_outputs(1785) <= '1';
    layer2_outputs(1786) <= not(layer1_outputs(528));
    layer2_outputs(1787) <= not((layer1_outputs(2164)) or (layer1_outputs(803)));
    layer2_outputs(1788) <= layer1_outputs(1225);
    layer2_outputs(1789) <= layer1_outputs(911);
    layer2_outputs(1790) <= not(layer1_outputs(2376));
    layer2_outputs(1791) <= (layer1_outputs(210)) and not (layer1_outputs(479));
    layer2_outputs(1792) <= (layer1_outputs(692)) and not (layer1_outputs(610));
    layer2_outputs(1793) <= not(layer1_outputs(2303)) or (layer1_outputs(120));
    layer2_outputs(1794) <= '1';
    layer2_outputs(1795) <= (layer1_outputs(1240)) or (layer1_outputs(1848));
    layer2_outputs(1796) <= layer1_outputs(1676);
    layer2_outputs(1797) <= not(layer1_outputs(2124)) or (layer1_outputs(362));
    layer2_outputs(1798) <= not((layer1_outputs(996)) and (layer1_outputs(1136)));
    layer2_outputs(1799) <= (layer1_outputs(1217)) and (layer1_outputs(2406));
    layer2_outputs(1800) <= not(layer1_outputs(2307));
    layer2_outputs(1801) <= not(layer1_outputs(909));
    layer2_outputs(1802) <= not(layer1_outputs(2505));
    layer2_outputs(1803) <= not(layer1_outputs(867));
    layer2_outputs(1804) <= layer1_outputs(1427);
    layer2_outputs(1805) <= (layer1_outputs(942)) and (layer1_outputs(2142));
    layer2_outputs(1806) <= not(layer1_outputs(2502)) or (layer1_outputs(1436));
    layer2_outputs(1807) <= '0';
    layer2_outputs(1808) <= not(layer1_outputs(1429));
    layer2_outputs(1809) <= (layer1_outputs(1449)) and not (layer1_outputs(1342));
    layer2_outputs(1810) <= (layer1_outputs(1889)) and (layer1_outputs(241));
    layer2_outputs(1811) <= not(layer1_outputs(1117));
    layer2_outputs(1812) <= not(layer1_outputs(947));
    layer2_outputs(1813) <= not(layer1_outputs(853));
    layer2_outputs(1814) <= (layer1_outputs(679)) and (layer1_outputs(2032));
    layer2_outputs(1815) <= not(layer1_outputs(345));
    layer2_outputs(1816) <= layer1_outputs(2461);
    layer2_outputs(1817) <= not(layer1_outputs(1687));
    layer2_outputs(1818) <= '1';
    layer2_outputs(1819) <= not(layer1_outputs(281));
    layer2_outputs(1820) <= not((layer1_outputs(1504)) or (layer1_outputs(1885)));
    layer2_outputs(1821) <= layer1_outputs(1439);
    layer2_outputs(1822) <= layer1_outputs(1787);
    layer2_outputs(1823) <= not(layer1_outputs(76)) or (layer1_outputs(1590));
    layer2_outputs(1824) <= not((layer1_outputs(2168)) or (layer1_outputs(1952)));
    layer2_outputs(1825) <= layer1_outputs(2377);
    layer2_outputs(1826) <= not(layer1_outputs(1606));
    layer2_outputs(1827) <= not(layer1_outputs(291));
    layer2_outputs(1828) <= (layer1_outputs(811)) or (layer1_outputs(1390));
    layer2_outputs(1829) <= (layer1_outputs(931)) and (layer1_outputs(1563));
    layer2_outputs(1830) <= not(layer1_outputs(1381));
    layer2_outputs(1831) <= (layer1_outputs(640)) or (layer1_outputs(1051));
    layer2_outputs(1832) <= not((layer1_outputs(542)) and (layer1_outputs(759)));
    layer2_outputs(1833) <= not(layer1_outputs(2080));
    layer2_outputs(1834) <= not(layer1_outputs(236));
    layer2_outputs(1835) <= not((layer1_outputs(2292)) or (layer1_outputs(1624)));
    layer2_outputs(1836) <= (layer1_outputs(96)) and not (layer1_outputs(2508));
    layer2_outputs(1837) <= (layer1_outputs(2444)) and (layer1_outputs(661));
    layer2_outputs(1838) <= layer1_outputs(1584);
    layer2_outputs(1839) <= '1';
    layer2_outputs(1840) <= not(layer1_outputs(690));
    layer2_outputs(1841) <= layer1_outputs(1243);
    layer2_outputs(1842) <= not((layer1_outputs(82)) or (layer1_outputs(1544)));
    layer2_outputs(1843) <= (layer1_outputs(2484)) and not (layer1_outputs(806));
    layer2_outputs(1844) <= '1';
    layer2_outputs(1845) <= (layer1_outputs(2085)) or (layer1_outputs(470));
    layer2_outputs(1846) <= not((layer1_outputs(519)) and (layer1_outputs(386)));
    layer2_outputs(1847) <= '0';
    layer2_outputs(1848) <= not(layer1_outputs(1512)) or (layer1_outputs(998));
    layer2_outputs(1849) <= not(layer1_outputs(1666));
    layer2_outputs(1850) <= '1';
    layer2_outputs(1851) <= not(layer1_outputs(1255));
    layer2_outputs(1852) <= not((layer1_outputs(1109)) and (layer1_outputs(1268)));
    layer2_outputs(1853) <= layer1_outputs(884);
    layer2_outputs(1854) <= (layer1_outputs(1747)) and not (layer1_outputs(1530));
    layer2_outputs(1855) <= (layer1_outputs(2229)) and not (layer1_outputs(148));
    layer2_outputs(1856) <= not(layer1_outputs(105)) or (layer1_outputs(504));
    layer2_outputs(1857) <= not((layer1_outputs(1212)) or (layer1_outputs(1785)));
    layer2_outputs(1858) <= '1';
    layer2_outputs(1859) <= (layer1_outputs(1494)) and not (layer1_outputs(395));
    layer2_outputs(1860) <= '1';
    layer2_outputs(1861) <= not(layer1_outputs(1351)) or (layer1_outputs(64));
    layer2_outputs(1862) <= not(layer1_outputs(725)) or (layer1_outputs(552));
    layer2_outputs(1863) <= (layer1_outputs(564)) and (layer1_outputs(428));
    layer2_outputs(1864) <= layer1_outputs(2175);
    layer2_outputs(1865) <= (layer1_outputs(1743)) and not (layer1_outputs(2092));
    layer2_outputs(1866) <= (layer1_outputs(1679)) and not (layer1_outputs(1594));
    layer2_outputs(1867) <= not(layer1_outputs(2448));
    layer2_outputs(1868) <= (layer1_outputs(2290)) or (layer1_outputs(1384));
    layer2_outputs(1869) <= (layer1_outputs(2558)) and not (layer1_outputs(2248));
    layer2_outputs(1870) <= layer1_outputs(301);
    layer2_outputs(1871) <= not(layer1_outputs(442)) or (layer1_outputs(2543));
    layer2_outputs(1872) <= not(layer1_outputs(967)) or (layer1_outputs(956));
    layer2_outputs(1873) <= (layer1_outputs(1067)) and not (layer1_outputs(620));
    layer2_outputs(1874) <= layer1_outputs(2534);
    layer2_outputs(1875) <= not(layer1_outputs(1321));
    layer2_outputs(1876) <= not(layer1_outputs(364)) or (layer1_outputs(179));
    layer2_outputs(1877) <= (layer1_outputs(1800)) or (layer1_outputs(1602));
    layer2_outputs(1878) <= (layer1_outputs(1367)) and (layer1_outputs(1505));
    layer2_outputs(1879) <= layer1_outputs(847);
    layer2_outputs(1880) <= (layer1_outputs(529)) xor (layer1_outputs(2287));
    layer2_outputs(1881) <= layer1_outputs(2090);
    layer2_outputs(1882) <= not((layer1_outputs(562)) or (layer1_outputs(1030)));
    layer2_outputs(1883) <= not(layer1_outputs(1732));
    layer2_outputs(1884) <= layer1_outputs(536);
    layer2_outputs(1885) <= layer1_outputs(860);
    layer2_outputs(1886) <= (layer1_outputs(1691)) and not (layer1_outputs(1984));
    layer2_outputs(1887) <= not((layer1_outputs(1434)) or (layer1_outputs(2505)));
    layer2_outputs(1888) <= not(layer1_outputs(492)) or (layer1_outputs(877));
    layer2_outputs(1889) <= '0';
    layer2_outputs(1890) <= (layer1_outputs(122)) and not (layer1_outputs(702));
    layer2_outputs(1891) <= (layer1_outputs(990)) and not (layer1_outputs(1144));
    layer2_outputs(1892) <= layer1_outputs(134);
    layer2_outputs(1893) <= not(layer1_outputs(39));
    layer2_outputs(1894) <= (layer1_outputs(2221)) and (layer1_outputs(2266));
    layer2_outputs(1895) <= '1';
    layer2_outputs(1896) <= (layer1_outputs(1069)) and not (layer1_outputs(1290));
    layer2_outputs(1897) <= (layer1_outputs(852)) and not (layer1_outputs(437));
    layer2_outputs(1898) <= (layer1_outputs(235)) xor (layer1_outputs(1422));
    layer2_outputs(1899) <= (layer1_outputs(1745)) and not (layer1_outputs(1692));
    layer2_outputs(1900) <= '0';
    layer2_outputs(1901) <= (layer1_outputs(1296)) and not (layer1_outputs(1916));
    layer2_outputs(1902) <= not(layer1_outputs(2446));
    layer2_outputs(1903) <= not(layer1_outputs(403)) or (layer1_outputs(2223));
    layer2_outputs(1904) <= layer1_outputs(891);
    layer2_outputs(1905) <= layer1_outputs(1593);
    layer2_outputs(1906) <= not(layer1_outputs(65)) or (layer1_outputs(1349));
    layer2_outputs(1907) <= not(layer1_outputs(339)) or (layer1_outputs(726));
    layer2_outputs(1908) <= layer1_outputs(331);
    layer2_outputs(1909) <= not((layer1_outputs(1748)) and (layer1_outputs(958)));
    layer2_outputs(1910) <= (layer1_outputs(594)) and not (layer1_outputs(402));
    layer2_outputs(1911) <= not(layer1_outputs(1675));
    layer2_outputs(1912) <= layer1_outputs(999);
    layer2_outputs(1913) <= not(layer1_outputs(548));
    layer2_outputs(1914) <= '1';
    layer2_outputs(1915) <= (layer1_outputs(218)) or (layer1_outputs(2394));
    layer2_outputs(1916) <= not((layer1_outputs(373)) and (layer1_outputs(86)));
    layer2_outputs(1917) <= layer1_outputs(1115);
    layer2_outputs(1918) <= not(layer1_outputs(38));
    layer2_outputs(1919) <= '1';
    layer2_outputs(1920) <= '0';
    layer2_outputs(1921) <= (layer1_outputs(230)) and (layer1_outputs(230));
    layer2_outputs(1922) <= layer1_outputs(2240);
    layer2_outputs(1923) <= layer1_outputs(2043);
    layer2_outputs(1924) <= not(layer1_outputs(56)) or (layer1_outputs(1939));
    layer2_outputs(1925) <= layer1_outputs(2216);
    layer2_outputs(1926) <= layer1_outputs(1572);
    layer2_outputs(1927) <= layer1_outputs(224);
    layer2_outputs(1928) <= (layer1_outputs(1572)) and not (layer1_outputs(760));
    layer2_outputs(1929) <= '1';
    layer2_outputs(1930) <= not(layer1_outputs(521)) or (layer1_outputs(1579));
    layer2_outputs(1931) <= not(layer1_outputs(141));
    layer2_outputs(1932) <= '1';
    layer2_outputs(1933) <= layer1_outputs(493);
    layer2_outputs(1934) <= layer1_outputs(1639);
    layer2_outputs(1935) <= (layer1_outputs(371)) or (layer1_outputs(2198));
    layer2_outputs(1936) <= layer1_outputs(2264);
    layer2_outputs(1937) <= layer1_outputs(780);
    layer2_outputs(1938) <= (layer1_outputs(1319)) and (layer1_outputs(981));
    layer2_outputs(1939) <= layer1_outputs(1026);
    layer2_outputs(1940) <= (layer1_outputs(1539)) and not (layer1_outputs(348));
    layer2_outputs(1941) <= (layer1_outputs(1930)) and not (layer1_outputs(134));
    layer2_outputs(1942) <= (layer1_outputs(1892)) and (layer1_outputs(83));
    layer2_outputs(1943) <= (layer1_outputs(939)) and not (layer1_outputs(93));
    layer2_outputs(1944) <= (layer1_outputs(1238)) and not (layer1_outputs(2318));
    layer2_outputs(1945) <= layer1_outputs(1852);
    layer2_outputs(1946) <= not((layer1_outputs(1000)) and (layer1_outputs(2288)));
    layer2_outputs(1947) <= (layer1_outputs(1805)) or (layer1_outputs(893));
    layer2_outputs(1948) <= (layer1_outputs(1637)) and not (layer1_outputs(938));
    layer2_outputs(1949) <= layer1_outputs(432);
    layer2_outputs(1950) <= not(layer1_outputs(233));
    layer2_outputs(1951) <= (layer1_outputs(1917)) and not (layer1_outputs(706));
    layer2_outputs(1952) <= not((layer1_outputs(1520)) or (layer1_outputs(822)));
    layer2_outputs(1953) <= not((layer1_outputs(1566)) and (layer1_outputs(268)));
    layer2_outputs(1954) <= not(layer1_outputs(1412));
    layer2_outputs(1955) <= (layer1_outputs(2140)) xor (layer1_outputs(1617));
    layer2_outputs(1956) <= layer1_outputs(1088);
    layer2_outputs(1957) <= (layer1_outputs(558)) and (layer1_outputs(35));
    layer2_outputs(1958) <= not((layer1_outputs(2509)) or (layer1_outputs(1480)));
    layer2_outputs(1959) <= '1';
    layer2_outputs(1960) <= not((layer1_outputs(346)) xor (layer1_outputs(2516)));
    layer2_outputs(1961) <= (layer1_outputs(2226)) or (layer1_outputs(2379));
    layer2_outputs(1962) <= not(layer1_outputs(1561));
    layer2_outputs(1963) <= not(layer1_outputs(1185)) or (layer1_outputs(411));
    layer2_outputs(1964) <= not(layer1_outputs(2075));
    layer2_outputs(1965) <= '1';
    layer2_outputs(1966) <= (layer1_outputs(2375)) and not (layer1_outputs(1871));
    layer2_outputs(1967) <= not(layer1_outputs(376));
    layer2_outputs(1968) <= not((layer1_outputs(1141)) or (layer1_outputs(972)));
    layer2_outputs(1969) <= layer1_outputs(622);
    layer2_outputs(1970) <= '1';
    layer2_outputs(1971) <= not((layer1_outputs(288)) or (layer1_outputs(655)));
    layer2_outputs(1972) <= layer1_outputs(398);
    layer2_outputs(1973) <= (layer1_outputs(928)) or (layer1_outputs(191));
    layer2_outputs(1974) <= layer1_outputs(685);
    layer2_outputs(1975) <= layer1_outputs(2374);
    layer2_outputs(1976) <= layer1_outputs(482);
    layer2_outputs(1977) <= (layer1_outputs(2012)) and (layer1_outputs(2059));
    layer2_outputs(1978) <= layer1_outputs(1855);
    layer2_outputs(1979) <= not(layer1_outputs(331));
    layer2_outputs(1980) <= not(layer1_outputs(1076));
    layer2_outputs(1981) <= not(layer1_outputs(2513)) or (layer1_outputs(138));
    layer2_outputs(1982) <= (layer1_outputs(1915)) and (layer1_outputs(1882));
    layer2_outputs(1983) <= (layer1_outputs(1867)) and not (layer1_outputs(682));
    layer2_outputs(1984) <= not(layer1_outputs(1057));
    layer2_outputs(1985) <= (layer1_outputs(854)) and not (layer1_outputs(1955));
    layer2_outputs(1986) <= not((layer1_outputs(1755)) and (layer1_outputs(481)));
    layer2_outputs(1987) <= layer1_outputs(1280);
    layer2_outputs(1988) <= layer1_outputs(172);
    layer2_outputs(1989) <= layer1_outputs(84);
    layer2_outputs(1990) <= not(layer1_outputs(924));
    layer2_outputs(1991) <= (layer1_outputs(1557)) and not (layer1_outputs(851));
    layer2_outputs(1992) <= not((layer1_outputs(882)) and (layer1_outputs(164)));
    layer2_outputs(1993) <= (layer1_outputs(837)) and not (layer1_outputs(1822));
    layer2_outputs(1994) <= not(layer1_outputs(826));
    layer2_outputs(1995) <= layer1_outputs(2282);
    layer2_outputs(1996) <= not((layer1_outputs(1094)) or (layer1_outputs(93)));
    layer2_outputs(1997) <= layer1_outputs(2046);
    layer2_outputs(1998) <= '1';
    layer2_outputs(1999) <= layer1_outputs(155);
    layer2_outputs(2000) <= layer1_outputs(1588);
    layer2_outputs(2001) <= '0';
    layer2_outputs(2002) <= not(layer1_outputs(1726));
    layer2_outputs(2003) <= not((layer1_outputs(1293)) or (layer1_outputs(163)));
    layer2_outputs(2004) <= not((layer1_outputs(1259)) xor (layer1_outputs(1267)));
    layer2_outputs(2005) <= not(layer1_outputs(1444));
    layer2_outputs(2006) <= not(layer1_outputs(91));
    layer2_outputs(2007) <= layer1_outputs(119);
    layer2_outputs(2008) <= (layer1_outputs(2465)) and (layer1_outputs(159));
    layer2_outputs(2009) <= not((layer1_outputs(2531)) xor (layer1_outputs(751)));
    layer2_outputs(2010) <= layer1_outputs(2058);
    layer2_outputs(2011) <= not((layer1_outputs(2465)) or (layer1_outputs(2193)));
    layer2_outputs(2012) <= not(layer1_outputs(289));
    layer2_outputs(2013) <= (layer1_outputs(985)) or (layer1_outputs(789));
    layer2_outputs(2014) <= not(layer1_outputs(2272));
    layer2_outputs(2015) <= (layer1_outputs(1491)) or (layer1_outputs(1672));
    layer2_outputs(2016) <= layer1_outputs(1869);
    layer2_outputs(2017) <= not(layer1_outputs(2383));
    layer2_outputs(2018) <= '0';
    layer2_outputs(2019) <= not(layer1_outputs(1692));
    layer2_outputs(2020) <= not((layer1_outputs(1900)) and (layer1_outputs(74)));
    layer2_outputs(2021) <= layer1_outputs(2207);
    layer2_outputs(2022) <= not((layer1_outputs(1674)) or (layer1_outputs(1834)));
    layer2_outputs(2023) <= (layer1_outputs(745)) and not (layer1_outputs(1140));
    layer2_outputs(2024) <= (layer1_outputs(670)) and not (layer1_outputs(2135));
    layer2_outputs(2025) <= (layer1_outputs(2517)) and not (layer1_outputs(836));
    layer2_outputs(2026) <= layer1_outputs(1561);
    layer2_outputs(2027) <= (layer1_outputs(441)) and (layer1_outputs(2510));
    layer2_outputs(2028) <= layer1_outputs(1518);
    layer2_outputs(2029) <= not((layer1_outputs(262)) or (layer1_outputs(386)));
    layer2_outputs(2030) <= (layer1_outputs(914)) and not (layer1_outputs(681));
    layer2_outputs(2031) <= layer1_outputs(901);
    layer2_outputs(2032) <= (layer1_outputs(101)) or (layer1_outputs(1360));
    layer2_outputs(2033) <= '0';
    layer2_outputs(2034) <= (layer1_outputs(2209)) and (layer1_outputs(2040));
    layer2_outputs(2035) <= not(layer1_outputs(1271)) or (layer1_outputs(1530));
    layer2_outputs(2036) <= (layer1_outputs(1935)) or (layer1_outputs(429));
    layer2_outputs(2037) <= '1';
    layer2_outputs(2038) <= not(layer1_outputs(2425));
    layer2_outputs(2039) <= not(layer1_outputs(959));
    layer2_outputs(2040) <= (layer1_outputs(994)) and not (layer1_outputs(2537));
    layer2_outputs(2041) <= '0';
    layer2_outputs(2042) <= not(layer1_outputs(392));
    layer2_outputs(2043) <= layer1_outputs(1913);
    layer2_outputs(2044) <= (layer1_outputs(1060)) or (layer1_outputs(1549));
    layer2_outputs(2045) <= not(layer1_outputs(1371)) or (layer1_outputs(1534));
    layer2_outputs(2046) <= layer1_outputs(2147);
    layer2_outputs(2047) <= not(layer1_outputs(610));
    layer2_outputs(2048) <= not(layer1_outputs(2142));
    layer2_outputs(2049) <= (layer1_outputs(771)) and not (layer1_outputs(1197));
    layer2_outputs(2050) <= not(layer1_outputs(1013));
    layer2_outputs(2051) <= not(layer1_outputs(2219));
    layer2_outputs(2052) <= not(layer1_outputs(1896));
    layer2_outputs(2053) <= not((layer1_outputs(2401)) or (layer1_outputs(546)));
    layer2_outputs(2054) <= layer1_outputs(753);
    layer2_outputs(2055) <= (layer1_outputs(588)) or (layer1_outputs(1668));
    layer2_outputs(2056) <= not(layer1_outputs(260));
    layer2_outputs(2057) <= (layer1_outputs(1847)) or (layer1_outputs(1914));
    layer2_outputs(2058) <= layer1_outputs(1405);
    layer2_outputs(2059) <= (layer1_outputs(611)) and not (layer1_outputs(271));
    layer2_outputs(2060) <= '0';
    layer2_outputs(2061) <= not(layer1_outputs(1497));
    layer2_outputs(2062) <= (layer1_outputs(1163)) and not (layer1_outputs(1063));
    layer2_outputs(2063) <= (layer1_outputs(619)) and not (layer1_outputs(1285));
    layer2_outputs(2064) <= (layer1_outputs(2278)) and (layer1_outputs(916));
    layer2_outputs(2065) <= layer1_outputs(77);
    layer2_outputs(2066) <= (layer1_outputs(1256)) and not (layer1_outputs(2225));
    layer2_outputs(2067) <= not(layer1_outputs(576));
    layer2_outputs(2068) <= not((layer1_outputs(547)) xor (layer1_outputs(2013)));
    layer2_outputs(2069) <= not((layer1_outputs(282)) or (layer1_outputs(344)));
    layer2_outputs(2070) <= (layer1_outputs(2070)) or (layer1_outputs(1603));
    layer2_outputs(2071) <= not(layer1_outputs(1051));
    layer2_outputs(2072) <= not(layer1_outputs(2104));
    layer2_outputs(2073) <= not(layer1_outputs(125)) or (layer1_outputs(1414));
    layer2_outputs(2074) <= layer1_outputs(493);
    layer2_outputs(2075) <= not((layer1_outputs(1196)) or (layer1_outputs(2131)));
    layer2_outputs(2076) <= not(layer1_outputs(903)) or (layer1_outputs(1258));
    layer2_outputs(2077) <= (layer1_outputs(849)) and not (layer1_outputs(589));
    layer2_outputs(2078) <= layer1_outputs(936);
    layer2_outputs(2079) <= not(layer1_outputs(2393));
    layer2_outputs(2080) <= not(layer1_outputs(1773));
    layer2_outputs(2081) <= not((layer1_outputs(2129)) xor (layer1_outputs(892)));
    layer2_outputs(2082) <= not((layer1_outputs(1261)) and (layer1_outputs(322)));
    layer2_outputs(2083) <= (layer1_outputs(1796)) and not (layer1_outputs(796));
    layer2_outputs(2084) <= '1';
    layer2_outputs(2085) <= '0';
    layer2_outputs(2086) <= not((layer1_outputs(2496)) or (layer1_outputs(2418)));
    layer2_outputs(2087) <= not(layer1_outputs(274)) or (layer1_outputs(971));
    layer2_outputs(2088) <= (layer1_outputs(951)) and (layer1_outputs(1662));
    layer2_outputs(2089) <= not((layer1_outputs(799)) and (layer1_outputs(1143)));
    layer2_outputs(2090) <= (layer1_outputs(813)) and not (layer1_outputs(2250));
    layer2_outputs(2091) <= not(layer1_outputs(1644));
    layer2_outputs(2092) <= '0';
    layer2_outputs(2093) <= layer1_outputs(2124);
    layer2_outputs(2094) <= (layer1_outputs(1514)) and not (layer1_outputs(236));
    layer2_outputs(2095) <= not((layer1_outputs(1528)) or (layer1_outputs(513)));
    layer2_outputs(2096) <= (layer1_outputs(2506)) and not (layer1_outputs(1612));
    layer2_outputs(2097) <= not(layer1_outputs(724));
    layer2_outputs(2098) <= not(layer1_outputs(1587)) or (layer1_outputs(908));
    layer2_outputs(2099) <= (layer1_outputs(2345)) and not (layer1_outputs(1554));
    layer2_outputs(2100) <= not(layer1_outputs(274)) or (layer1_outputs(779));
    layer2_outputs(2101) <= layer1_outputs(310);
    layer2_outputs(2102) <= not((layer1_outputs(2160)) or (layer1_outputs(2411)));
    layer2_outputs(2103) <= (layer1_outputs(1890)) and not (layer1_outputs(1934));
    layer2_outputs(2104) <= not((layer1_outputs(887)) or (layer1_outputs(2422)));
    layer2_outputs(2105) <= layer1_outputs(1579);
    layer2_outputs(2106) <= (layer1_outputs(569)) and not (layer1_outputs(186));
    layer2_outputs(2107) <= (layer1_outputs(1309)) and not (layer1_outputs(897));
    layer2_outputs(2108) <= (layer1_outputs(2163)) or (layer1_outputs(1879));
    layer2_outputs(2109) <= not(layer1_outputs(1451)) or (layer1_outputs(1992));
    layer2_outputs(2110) <= '1';
    layer2_outputs(2111) <= layer1_outputs(815);
    layer2_outputs(2112) <= not(layer1_outputs(248));
    layer2_outputs(2113) <= not(layer1_outputs(1592)) or (layer1_outputs(507));
    layer2_outputs(2114) <= layer1_outputs(303);
    layer2_outputs(2115) <= '0';
    layer2_outputs(2116) <= not(layer1_outputs(1508));
    layer2_outputs(2117) <= not(layer1_outputs(2509));
    layer2_outputs(2118) <= layer1_outputs(2215);
    layer2_outputs(2119) <= not(layer1_outputs(687)) or (layer1_outputs(2438));
    layer2_outputs(2120) <= layer1_outputs(1970);
    layer2_outputs(2121) <= not(layer1_outputs(519));
    layer2_outputs(2122) <= (layer1_outputs(1292)) or (layer1_outputs(2264));
    layer2_outputs(2123) <= not(layer1_outputs(1507)) or (layer1_outputs(2187));
    layer2_outputs(2124) <= layer1_outputs(1269);
    layer2_outputs(2125) <= (layer1_outputs(733)) and (layer1_outputs(423));
    layer2_outputs(2126) <= '1';
    layer2_outputs(2127) <= layer1_outputs(1065);
    layer2_outputs(2128) <= layer1_outputs(1911);
    layer2_outputs(2129) <= '0';
    layer2_outputs(2130) <= not(layer1_outputs(1270));
    layer2_outputs(2131) <= '1';
    layer2_outputs(2132) <= not((layer1_outputs(1067)) and (layer1_outputs(541)));
    layer2_outputs(2133) <= layer1_outputs(684);
    layer2_outputs(2134) <= not(layer1_outputs(1114));
    layer2_outputs(2135) <= layer1_outputs(782);
    layer2_outputs(2136) <= '0';
    layer2_outputs(2137) <= layer1_outputs(306);
    layer2_outputs(2138) <= (layer1_outputs(2014)) and (layer1_outputs(852));
    layer2_outputs(2139) <= not((layer1_outputs(1499)) and (layer1_outputs(1445)));
    layer2_outputs(2140) <= not(layer1_outputs(678));
    layer2_outputs(2141) <= not(layer1_outputs(1607));
    layer2_outputs(2142) <= '0';
    layer2_outputs(2143) <= (layer1_outputs(390)) and (layer1_outputs(200));
    layer2_outputs(2144) <= not(layer1_outputs(1701)) or (layer1_outputs(1485));
    layer2_outputs(2145) <= (layer1_outputs(2029)) and not (layer1_outputs(898));
    layer2_outputs(2146) <= not((layer1_outputs(804)) and (layer1_outputs(863)));
    layer2_outputs(2147) <= (layer1_outputs(2196)) and (layer1_outputs(920));
    layer2_outputs(2148) <= not(layer1_outputs(2526)) or (layer1_outputs(647));
    layer2_outputs(2149) <= (layer1_outputs(2268)) or (layer1_outputs(317));
    layer2_outputs(2150) <= layer1_outputs(2172);
    layer2_outputs(2151) <= (layer1_outputs(99)) and not (layer1_outputs(1285));
    layer2_outputs(2152) <= '0';
    layer2_outputs(2153) <= not(layer1_outputs(1754));
    layer2_outputs(2154) <= not(layer1_outputs(1717)) or (layer1_outputs(162));
    layer2_outputs(2155) <= not(layer1_outputs(2232));
    layer2_outputs(2156) <= layer1_outputs(634);
    layer2_outputs(2157) <= (layer1_outputs(2559)) and (layer1_outputs(1883));
    layer2_outputs(2158) <= layer1_outputs(817);
    layer2_outputs(2159) <= layer1_outputs(1663);
    layer2_outputs(2160) <= not((layer1_outputs(974)) and (layer1_outputs(2031)));
    layer2_outputs(2161) <= not((layer1_outputs(2148)) and (layer1_outputs(1525)));
    layer2_outputs(2162) <= layer1_outputs(2551);
    layer2_outputs(2163) <= layer1_outputs(37);
    layer2_outputs(2164) <= (layer1_outputs(51)) or (layer1_outputs(2109));
    layer2_outputs(2165) <= '1';
    layer2_outputs(2166) <= (layer1_outputs(735)) and not (layer1_outputs(2559));
    layer2_outputs(2167) <= not((layer1_outputs(641)) xor (layer1_outputs(1896)));
    layer2_outputs(2168) <= not((layer1_outputs(1322)) and (layer1_outputs(2136)));
    layer2_outputs(2169) <= not(layer1_outputs(766)) or (layer1_outputs(717));
    layer2_outputs(2170) <= not(layer1_outputs(626)) or (layer1_outputs(850));
    layer2_outputs(2171) <= not((layer1_outputs(1524)) and (layer1_outputs(132)));
    layer2_outputs(2172) <= layer1_outputs(247);
    layer2_outputs(2173) <= '1';
    layer2_outputs(2174) <= not(layer1_outputs(1402)) or (layer1_outputs(1436));
    layer2_outputs(2175) <= not(layer1_outputs(1443));
    layer2_outputs(2176) <= layer1_outputs(2019);
    layer2_outputs(2177) <= not((layer1_outputs(710)) and (layer1_outputs(2415)));
    layer2_outputs(2178) <= (layer1_outputs(748)) or (layer1_outputs(675));
    layer2_outputs(2179) <= layer1_outputs(1447);
    layer2_outputs(2180) <= not(layer1_outputs(50)) or (layer1_outputs(460));
    layer2_outputs(2181) <= (layer1_outputs(2399)) and not (layer1_outputs(2365));
    layer2_outputs(2182) <= not((layer1_outputs(471)) and (layer1_outputs(543)));
    layer2_outputs(2183) <= layer1_outputs(918);
    layer2_outputs(2184) <= not((layer1_outputs(1936)) or (layer1_outputs(187)));
    layer2_outputs(2185) <= layer1_outputs(1442);
    layer2_outputs(2186) <= layer1_outputs(85);
    layer2_outputs(2187) <= not(layer1_outputs(0));
    layer2_outputs(2188) <= (layer1_outputs(498)) xor (layer1_outputs(1856));
    layer2_outputs(2189) <= layer1_outputs(1458);
    layer2_outputs(2190) <= layer1_outputs(406);
    layer2_outputs(2191) <= '1';
    layer2_outputs(2192) <= layer1_outputs(2126);
    layer2_outputs(2193) <= layer1_outputs(1363);
    layer2_outputs(2194) <= (layer1_outputs(1404)) and not (layer1_outputs(2064));
    layer2_outputs(2195) <= (layer1_outputs(487)) and not (layer1_outputs(2050));
    layer2_outputs(2196) <= not(layer1_outputs(915));
    layer2_outputs(2197) <= not(layer1_outputs(569)) or (layer1_outputs(446));
    layer2_outputs(2198) <= (layer1_outputs(1907)) and (layer1_outputs(1305));
    layer2_outputs(2199) <= not(layer1_outputs(20));
    layer2_outputs(2200) <= (layer1_outputs(1841)) or (layer1_outputs(1651));
    layer2_outputs(2201) <= not(layer1_outputs(1866));
    layer2_outputs(2202) <= (layer1_outputs(110)) and (layer1_outputs(337));
    layer2_outputs(2203) <= layer1_outputs(25);
    layer2_outputs(2204) <= (layer1_outputs(460)) and (layer1_outputs(2523));
    layer2_outputs(2205) <= '1';
    layer2_outputs(2206) <= not(layer1_outputs(992));
    layer2_outputs(2207) <= (layer1_outputs(278)) or (layer1_outputs(2170));
    layer2_outputs(2208) <= not(layer1_outputs(1947)) or (layer1_outputs(977));
    layer2_outputs(2209) <= not(layer1_outputs(1962));
    layer2_outputs(2210) <= (layer1_outputs(1268)) and not (layer1_outputs(18));
    layer2_outputs(2211) <= layer1_outputs(1812);
    layer2_outputs(2212) <= layer1_outputs(2326);
    layer2_outputs(2213) <= not(layer1_outputs(1524)) or (layer1_outputs(1246));
    layer2_outputs(2214) <= not((layer1_outputs(1826)) xor (layer1_outputs(39)));
    layer2_outputs(2215) <= layer1_outputs(1476);
    layer2_outputs(2216) <= not(layer1_outputs(586)) or (layer1_outputs(1600));
    layer2_outputs(2217) <= not((layer1_outputs(2213)) or (layer1_outputs(433)));
    layer2_outputs(2218) <= '1';
    layer2_outputs(2219) <= not(layer1_outputs(2332));
    layer2_outputs(2220) <= not(layer1_outputs(535));
    layer2_outputs(2221) <= not(layer1_outputs(923));
    layer2_outputs(2222) <= not(layer1_outputs(471));
    layer2_outputs(2223) <= (layer1_outputs(1318)) and not (layer1_outputs(1358));
    layer2_outputs(2224) <= (layer1_outputs(354)) and not (layer1_outputs(1591));
    layer2_outputs(2225) <= layer1_outputs(326);
    layer2_outputs(2226) <= not(layer1_outputs(154));
    layer2_outputs(2227) <= not((layer1_outputs(1440)) or (layer1_outputs(2001)));
    layer2_outputs(2228) <= (layer1_outputs(2122)) or (layer1_outputs(2356));
    layer2_outputs(2229) <= (layer1_outputs(2063)) xor (layer1_outputs(555));
    layer2_outputs(2230) <= not((layer1_outputs(1039)) or (layer1_outputs(490)));
    layer2_outputs(2231) <= '1';
    layer2_outputs(2232) <= '1';
    layer2_outputs(2233) <= (layer1_outputs(2535)) and not (layer1_outputs(1182));
    layer2_outputs(2234) <= not(layer1_outputs(2015)) or (layer1_outputs(26));
    layer2_outputs(2235) <= (layer1_outputs(1996)) and not (layer1_outputs(1407));
    layer2_outputs(2236) <= (layer1_outputs(1380)) and (layer1_outputs(910));
    layer2_outputs(2237) <= '1';
    layer2_outputs(2238) <= '0';
    layer2_outputs(2239) <= layer1_outputs(1187);
    layer2_outputs(2240) <= not((layer1_outputs(838)) and (layer1_outputs(1180)));
    layer2_outputs(2241) <= layer1_outputs(2);
    layer2_outputs(2242) <= not(layer1_outputs(743)) or (layer1_outputs(184));
    layer2_outputs(2243) <= not(layer1_outputs(2096)) or (layer1_outputs(1544));
    layer2_outputs(2244) <= (layer1_outputs(721)) and not (layer1_outputs(1043));
    layer2_outputs(2245) <= '0';
    layer2_outputs(2246) <= not((layer1_outputs(1994)) and (layer1_outputs(612)));
    layer2_outputs(2247) <= layer1_outputs(847);
    layer2_outputs(2248) <= not(layer1_outputs(921));
    layer2_outputs(2249) <= not(layer1_outputs(2477)) or (layer1_outputs(1092));
    layer2_outputs(2250) <= layer1_outputs(436);
    layer2_outputs(2251) <= layer1_outputs(1766);
    layer2_outputs(2252) <= '1';
    layer2_outputs(2253) <= not(layer1_outputs(1865));
    layer2_outputs(2254) <= not(layer1_outputs(1055));
    layer2_outputs(2255) <= layer1_outputs(1163);
    layer2_outputs(2256) <= '0';
    layer2_outputs(2257) <= not(layer1_outputs(1940)) or (layer1_outputs(2354));
    layer2_outputs(2258) <= (layer1_outputs(1064)) or (layer1_outputs(2333));
    layer2_outputs(2259) <= not((layer1_outputs(508)) or (layer1_outputs(2071)));
    layer2_outputs(2260) <= layer1_outputs(1998);
    layer2_outputs(2261) <= (layer1_outputs(108)) and not (layer1_outputs(2151));
    layer2_outputs(2262) <= '1';
    layer2_outputs(2263) <= not(layer1_outputs(2035));
    layer2_outputs(2264) <= not((layer1_outputs(2503)) and (layer1_outputs(2144)));
    layer2_outputs(2265) <= not(layer1_outputs(270));
    layer2_outputs(2266) <= (layer1_outputs(49)) and not (layer1_outputs(1736));
    layer2_outputs(2267) <= not((layer1_outputs(1462)) and (layer1_outputs(2056)));
    layer2_outputs(2268) <= (layer1_outputs(1696)) and not (layer1_outputs(150));
    layer2_outputs(2269) <= (layer1_outputs(482)) and not (layer1_outputs(1542));
    layer2_outputs(2270) <= not((layer1_outputs(1098)) or (layer1_outputs(1630)));
    layer2_outputs(2271) <= layer1_outputs(2334);
    layer2_outputs(2272) <= '0';
    layer2_outputs(2273) <= (layer1_outputs(388)) and (layer1_outputs(175));
    layer2_outputs(2274) <= layer1_outputs(353);
    layer2_outputs(2275) <= not(layer1_outputs(2250));
    layer2_outputs(2276) <= not(layer1_outputs(2030)) or (layer1_outputs(252));
    layer2_outputs(2277) <= layer1_outputs(1131);
    layer2_outputs(2278) <= '1';
    layer2_outputs(2279) <= not(layer1_outputs(525));
    layer2_outputs(2280) <= not(layer1_outputs(1570)) or (layer1_outputs(2156));
    layer2_outputs(2281) <= layer1_outputs(1718);
    layer2_outputs(2282) <= '0';
    layer2_outputs(2283) <= (layer1_outputs(157)) and (layer1_outputs(986));
    layer2_outputs(2284) <= not(layer1_outputs(917));
    layer2_outputs(2285) <= layer1_outputs(2298);
    layer2_outputs(2286) <= layer1_outputs(1187);
    layer2_outputs(2287) <= (layer1_outputs(595)) and not (layer1_outputs(1886));
    layer2_outputs(2288) <= (layer1_outputs(2514)) and (layer1_outputs(2353));
    layer2_outputs(2289) <= not(layer1_outputs(674));
    layer2_outputs(2290) <= layer1_outputs(2227);
    layer2_outputs(2291) <= layer1_outputs(2546);
    layer2_outputs(2292) <= '1';
    layer2_outputs(2293) <= layer1_outputs(1042);
    layer2_outputs(2294) <= not(layer1_outputs(1988));
    layer2_outputs(2295) <= not((layer1_outputs(597)) and (layer1_outputs(2406)));
    layer2_outputs(2296) <= not(layer1_outputs(1901)) or (layer1_outputs(78));
    layer2_outputs(2297) <= layer1_outputs(755);
    layer2_outputs(2298) <= not((layer1_outputs(1130)) or (layer1_outputs(126)));
    layer2_outputs(2299) <= (layer1_outputs(924)) and not (layer1_outputs(185));
    layer2_outputs(2300) <= not(layer1_outputs(1411));
    layer2_outputs(2301) <= not((layer1_outputs(2202)) or (layer1_outputs(1)));
    layer2_outputs(2302) <= (layer1_outputs(1982)) and (layer1_outputs(968));
    layer2_outputs(2303) <= '1';
    layer2_outputs(2304) <= '1';
    layer2_outputs(2305) <= not(layer1_outputs(1735));
    layer2_outputs(2306) <= '1';
    layer2_outputs(2307) <= (layer1_outputs(1963)) and not (layer1_outputs(1511));
    layer2_outputs(2308) <= '0';
    layer2_outputs(2309) <= layer1_outputs(1326);
    layer2_outputs(2310) <= not((layer1_outputs(1808)) and (layer1_outputs(837)));
    layer2_outputs(2311) <= not(layer1_outputs(1580));
    layer2_outputs(2312) <= layer1_outputs(1604);
    layer2_outputs(2313) <= layer1_outputs(1347);
    layer2_outputs(2314) <= layer1_outputs(729);
    layer2_outputs(2315) <= (layer1_outputs(502)) and (layer1_outputs(2557));
    layer2_outputs(2316) <= (layer1_outputs(180)) or (layer1_outputs(1598));
    layer2_outputs(2317) <= not((layer1_outputs(1390)) and (layer1_outputs(949)));
    layer2_outputs(2318) <= not((layer1_outputs(496)) or (layer1_outputs(1171)));
    layer2_outputs(2319) <= '1';
    layer2_outputs(2320) <= not(layer1_outputs(1532)) or (layer1_outputs(671));
    layer2_outputs(2321) <= not(layer1_outputs(2256));
    layer2_outputs(2322) <= not(layer1_outputs(2533));
    layer2_outputs(2323) <= (layer1_outputs(937)) and not (layer1_outputs(978));
    layer2_outputs(2324) <= not(layer1_outputs(205)) or (layer1_outputs(456));
    layer2_outputs(2325) <= not((layer1_outputs(1437)) xor (layer1_outputs(2347)));
    layer2_outputs(2326) <= '1';
    layer2_outputs(2327) <= (layer1_outputs(1179)) and (layer1_outputs(1594));
    layer2_outputs(2328) <= layer1_outputs(177);
    layer2_outputs(2329) <= not((layer1_outputs(1359)) or (layer1_outputs(553)));
    layer2_outputs(2330) <= (layer1_outputs(935)) and not (layer1_outputs(150));
    layer2_outputs(2331) <= layer1_outputs(2325);
    layer2_outputs(2332) <= (layer1_outputs(265)) and not (layer1_outputs(2178));
    layer2_outputs(2333) <= not(layer1_outputs(1573));
    layer2_outputs(2334) <= '0';
    layer2_outputs(2335) <= layer1_outputs(714);
    layer2_outputs(2336) <= not(layer1_outputs(171));
    layer2_outputs(2337) <= not(layer1_outputs(1821));
    layer2_outputs(2338) <= '0';
    layer2_outputs(2339) <= '0';
    layer2_outputs(2340) <= layer1_outputs(1615);
    layer2_outputs(2341) <= not(layer1_outputs(409));
    layer2_outputs(2342) <= layer1_outputs(637);
    layer2_outputs(2343) <= '0';
    layer2_outputs(2344) <= layer1_outputs(526);
    layer2_outputs(2345) <= not((layer1_outputs(404)) and (layer1_outputs(1676)));
    layer2_outputs(2346) <= not((layer1_outputs(2324)) or (layer1_outputs(1119)));
    layer2_outputs(2347) <= (layer1_outputs(1475)) and not (layer1_outputs(1391));
    layer2_outputs(2348) <= not(layer1_outputs(2384)) or (layer1_outputs(1687));
    layer2_outputs(2349) <= (layer1_outputs(1399)) and not (layer1_outputs(319));
    layer2_outputs(2350) <= layer1_outputs(1172);
    layer2_outputs(2351) <= not(layer1_outputs(1853)) or (layer1_outputs(160));
    layer2_outputs(2352) <= not((layer1_outputs(2408)) and (layer1_outputs(2299)));
    layer2_outputs(2353) <= not(layer1_outputs(2033)) or (layer1_outputs(670));
    layer2_outputs(2354) <= (layer1_outputs(2087)) and not (layer1_outputs(1419));
    layer2_outputs(2355) <= (layer1_outputs(168)) and not (layer1_outputs(1602));
    layer2_outputs(2356) <= layer1_outputs(65);
    layer2_outputs(2357) <= not(layer1_outputs(2353));
    layer2_outputs(2358) <= not(layer1_outputs(1665));
    layer2_outputs(2359) <= (layer1_outputs(1899)) and not (layer1_outputs(1284));
    layer2_outputs(2360) <= '1';
    layer2_outputs(2361) <= '1';
    layer2_outputs(2362) <= '1';
    layer2_outputs(2363) <= layer1_outputs(965);
    layer2_outputs(2364) <= (layer1_outputs(287)) and not (layer1_outputs(2314));
    layer2_outputs(2365) <= not(layer1_outputs(1864)) or (layer1_outputs(1956));
    layer2_outputs(2366) <= (layer1_outputs(1219)) and not (layer1_outputs(666));
    layer2_outputs(2367) <= '0';
    layer2_outputs(2368) <= not((layer1_outputs(2391)) and (layer1_outputs(1838)));
    layer2_outputs(2369) <= not(layer1_outputs(975)) or (layer1_outputs(1469));
    layer2_outputs(2370) <= (layer1_outputs(1487)) xor (layer1_outputs(1229));
    layer2_outputs(2371) <= '0';
    layer2_outputs(2372) <= '0';
    layer2_outputs(2373) <= (layer1_outputs(207)) and not (layer1_outputs(1742));
    layer2_outputs(2374) <= '1';
    layer2_outputs(2375) <= not(layer1_outputs(68)) or (layer1_outputs(1186));
    layer2_outputs(2376) <= (layer1_outputs(2426)) and (layer1_outputs(133));
    layer2_outputs(2377) <= not(layer1_outputs(1932));
    layer2_outputs(2378) <= not(layer1_outputs(729)) or (layer1_outputs(1173));
    layer2_outputs(2379) <= layer1_outputs(1734);
    layer2_outputs(2380) <= layer1_outputs(340);
    layer2_outputs(2381) <= layer1_outputs(639);
    layer2_outputs(2382) <= '1';
    layer2_outputs(2383) <= (layer1_outputs(171)) and not (layer1_outputs(25));
    layer2_outputs(2384) <= not((layer1_outputs(2249)) and (layer1_outputs(286)));
    layer2_outputs(2385) <= '0';
    layer2_outputs(2386) <= (layer1_outputs(2521)) and not (layer1_outputs(1876));
    layer2_outputs(2387) <= layer1_outputs(2303);
    layer2_outputs(2388) <= not(layer1_outputs(929)) or (layer1_outputs(1255));
    layer2_outputs(2389) <= layer1_outputs(644);
    layer2_outputs(2390) <= not(layer1_outputs(2318));
    layer2_outputs(2391) <= layer1_outputs(1525);
    layer2_outputs(2392) <= (layer1_outputs(1478)) or (layer1_outputs(1348));
    layer2_outputs(2393) <= layer1_outputs(693);
    layer2_outputs(2394) <= not(layer1_outputs(1154));
    layer2_outputs(2395) <= (layer1_outputs(1806)) and not (layer1_outputs(966));
    layer2_outputs(2396) <= (layer1_outputs(2134)) and not (layer1_outputs(1099));
    layer2_outputs(2397) <= not(layer1_outputs(2206));
    layer2_outputs(2398) <= layer1_outputs(2052);
    layer2_outputs(2399) <= not(layer1_outputs(1537));
    layer2_outputs(2400) <= not((layer1_outputs(925)) or (layer1_outputs(888)));
    layer2_outputs(2401) <= layer1_outputs(419);
    layer2_outputs(2402) <= not((layer1_outputs(573)) and (layer1_outputs(2323)));
    layer2_outputs(2403) <= layer1_outputs(722);
    layer2_outputs(2404) <= not(layer1_outputs(1565));
    layer2_outputs(2405) <= not(layer1_outputs(918));
    layer2_outputs(2406) <= not(layer1_outputs(1582));
    layer2_outputs(2407) <= '0';
    layer2_outputs(2408) <= layer1_outputs(253);
    layer2_outputs(2409) <= not(layer1_outputs(49));
    layer2_outputs(2410) <= '0';
    layer2_outputs(2411) <= layer1_outputs(79);
    layer2_outputs(2412) <= not(layer1_outputs(448));
    layer2_outputs(2413) <= (layer1_outputs(784)) and not (layer1_outputs(1565));
    layer2_outputs(2414) <= (layer1_outputs(1520)) or (layer1_outputs(305));
    layer2_outputs(2415) <= layer1_outputs(1905);
    layer2_outputs(2416) <= '1';
    layer2_outputs(2417) <= layer1_outputs(1474);
    layer2_outputs(2418) <= (layer1_outputs(2271)) and (layer1_outputs(148));
    layer2_outputs(2419) <= '0';
    layer2_outputs(2420) <= (layer1_outputs(2306)) and not (layer1_outputs(497));
    layer2_outputs(2421) <= not((layer1_outputs(1275)) and (layer1_outputs(35)));
    layer2_outputs(2422) <= (layer1_outputs(1937)) and not (layer1_outputs(907));
    layer2_outputs(2423) <= layer1_outputs(190);
    layer2_outputs(2424) <= (layer1_outputs(416)) and not (layer1_outputs(1715));
    layer2_outputs(2425) <= not(layer1_outputs(1364));
    layer2_outputs(2426) <= (layer1_outputs(1677)) and not (layer1_outputs(1900));
    layer2_outputs(2427) <= (layer1_outputs(662)) and (layer1_outputs(2001));
    layer2_outputs(2428) <= '0';
    layer2_outputs(2429) <= not(layer1_outputs(735)) or (layer1_outputs(1943));
    layer2_outputs(2430) <= not(layer1_outputs(1055));
    layer2_outputs(2431) <= not(layer1_outputs(574));
    layer2_outputs(2432) <= not(layer1_outputs(711));
    layer2_outputs(2433) <= '1';
    layer2_outputs(2434) <= not(layer1_outputs(2037)) or (layer1_outputs(48));
    layer2_outputs(2435) <= '0';
    layer2_outputs(2436) <= (layer1_outputs(883)) and (layer1_outputs(214));
    layer2_outputs(2437) <= not((layer1_outputs(630)) and (layer1_outputs(1340)));
    layer2_outputs(2438) <= (layer1_outputs(1004)) xor (layer1_outputs(452));
    layer2_outputs(2439) <= not(layer1_outputs(69));
    layer2_outputs(2440) <= (layer1_outputs(1222)) and not (layer1_outputs(2482));
    layer2_outputs(2441) <= not(layer1_outputs(79));
    layer2_outputs(2442) <= not((layer1_outputs(2439)) or (layer1_outputs(786)));
    layer2_outputs(2443) <= not(layer1_outputs(877));
    layer2_outputs(2444) <= (layer1_outputs(146)) and (layer1_outputs(173));
    layer2_outputs(2445) <= not(layer1_outputs(661)) or (layer1_outputs(2420));
    layer2_outputs(2446) <= not(layer1_outputs(2212));
    layer2_outputs(2447) <= not(layer1_outputs(1481));
    layer2_outputs(2448) <= not((layer1_outputs(1474)) or (layer1_outputs(1992)));
    layer2_outputs(2449) <= (layer1_outputs(1777)) and not (layer1_outputs(810));
    layer2_outputs(2450) <= '0';
    layer2_outputs(2451) <= layer1_outputs(248);
    layer2_outputs(2452) <= not(layer1_outputs(1093));
    layer2_outputs(2453) <= '0';
    layer2_outputs(2454) <= layer1_outputs(1809);
    layer2_outputs(2455) <= layer1_outputs(1205);
    layer2_outputs(2456) <= layer1_outputs(1089);
    layer2_outputs(2457) <= layer1_outputs(2158);
    layer2_outputs(2458) <= layer1_outputs(270);
    layer2_outputs(2459) <= (layer1_outputs(945)) or (layer1_outputs(537));
    layer2_outputs(2460) <= (layer1_outputs(57)) and not (layer1_outputs(1141));
    layer2_outputs(2461) <= layer1_outputs(5);
    layer2_outputs(2462) <= (layer1_outputs(1576)) and (layer1_outputs(1650));
    layer2_outputs(2463) <= not(layer1_outputs(107)) or (layer1_outputs(784));
    layer2_outputs(2464) <= not(layer1_outputs(394)) or (layer1_outputs(2104));
    layer2_outputs(2465) <= layer1_outputs(1232);
    layer2_outputs(2466) <= not(layer1_outputs(973));
    layer2_outputs(2467) <= (layer1_outputs(2234)) and not (layer1_outputs(1661));
    layer2_outputs(2468) <= not(layer1_outputs(1762)) or (layer1_outputs(1013));
    layer2_outputs(2469) <= not(layer1_outputs(2231));
    layer2_outputs(2470) <= '0';
    layer2_outputs(2471) <= layer1_outputs(1382);
    layer2_outputs(2472) <= layer1_outputs(2146);
    layer2_outputs(2473) <= (layer1_outputs(2409)) and not (layer1_outputs(1232));
    layer2_outputs(2474) <= layer1_outputs(788);
    layer2_outputs(2475) <= not(layer1_outputs(2391));
    layer2_outputs(2476) <= (layer1_outputs(1167)) and not (layer1_outputs(2108));
    layer2_outputs(2477) <= not(layer1_outputs(1249)) or (layer1_outputs(1794));
    layer2_outputs(2478) <= layer1_outputs(1083);
    layer2_outputs(2479) <= '0';
    layer2_outputs(2480) <= not(layer1_outputs(1150)) or (layer1_outputs(1693));
    layer2_outputs(2481) <= '0';
    layer2_outputs(2482) <= (layer1_outputs(1311)) and not (layer1_outputs(2119));
    layer2_outputs(2483) <= layer1_outputs(1662);
    layer2_outputs(2484) <= layer1_outputs(213);
    layer2_outputs(2485) <= not(layer1_outputs(1001)) or (layer1_outputs(1464));
    layer2_outputs(2486) <= not((layer1_outputs(1471)) and (layer1_outputs(170)));
    layer2_outputs(2487) <= layer1_outputs(314);
    layer2_outputs(2488) <= layer1_outputs(54);
    layer2_outputs(2489) <= not(layer1_outputs(1811));
    layer2_outputs(2490) <= layer1_outputs(1955);
    layer2_outputs(2491) <= (layer1_outputs(399)) and not (layer1_outputs(1377));
    layer2_outputs(2492) <= layer1_outputs(375);
    layer2_outputs(2493) <= (layer1_outputs(841)) or (layer1_outputs(578));
    layer2_outputs(2494) <= not(layer1_outputs(1293)) or (layer1_outputs(345));
    layer2_outputs(2495) <= not(layer1_outputs(775));
    layer2_outputs(2496) <= not((layer1_outputs(2392)) or (layer1_outputs(669)));
    layer2_outputs(2497) <= (layer1_outputs(478)) and not (layer1_outputs(1848));
    layer2_outputs(2498) <= not(layer1_outputs(2232)) or (layer1_outputs(1200));
    layer2_outputs(2499) <= not(layer1_outputs(1155));
    layer2_outputs(2500) <= layer1_outputs(2000);
    layer2_outputs(2501) <= not(layer1_outputs(1793)) or (layer1_outputs(2251));
    layer2_outputs(2502) <= not((layer1_outputs(894)) or (layer1_outputs(2354)));
    layer2_outputs(2503) <= (layer1_outputs(1439)) and (layer1_outputs(981));
    layer2_outputs(2504) <= not((layer1_outputs(755)) or (layer1_outputs(2025)));
    layer2_outputs(2505) <= layer1_outputs(1276);
    layer2_outputs(2506) <= (layer1_outputs(332)) and (layer1_outputs(197));
    layer2_outputs(2507) <= layer1_outputs(117);
    layer2_outputs(2508) <= layer1_outputs(2443);
    layer2_outputs(2509) <= (layer1_outputs(1806)) and not (layer1_outputs(182));
    layer2_outputs(2510) <= not((layer1_outputs(1265)) or (layer1_outputs(204)));
    layer2_outputs(2511) <= not(layer1_outputs(2145));
    layer2_outputs(2512) <= (layer1_outputs(1535)) and not (layer1_outputs(1426));
    layer2_outputs(2513) <= '1';
    layer2_outputs(2514) <= layer1_outputs(544);
    layer2_outputs(2515) <= layer1_outputs(1816);
    layer2_outputs(2516) <= not((layer1_outputs(2538)) and (layer1_outputs(1540)));
    layer2_outputs(2517) <= not(layer1_outputs(2333)) or (layer1_outputs(2274));
    layer2_outputs(2518) <= not(layer1_outputs(1924));
    layer2_outputs(2519) <= not(layer1_outputs(665));
    layer2_outputs(2520) <= (layer1_outputs(1406)) and not (layer1_outputs(896));
    layer2_outputs(2521) <= not(layer1_outputs(325));
    layer2_outputs(2522) <= not(layer1_outputs(2504));
    layer2_outputs(2523) <= '0';
    layer2_outputs(2524) <= not((layer1_outputs(1635)) or (layer1_outputs(819)));
    layer2_outputs(2525) <= not(layer1_outputs(1537));
    layer2_outputs(2526) <= not(layer1_outputs(2312));
    layer2_outputs(2527) <= not(layer1_outputs(892));
    layer2_outputs(2528) <= not(layer1_outputs(829));
    layer2_outputs(2529) <= (layer1_outputs(2320)) xor (layer1_outputs(2404));
    layer2_outputs(2530) <= not((layer1_outputs(1502)) and (layer1_outputs(320)));
    layer2_outputs(2531) <= not(layer1_outputs(1483));
    layer2_outputs(2532) <= '1';
    layer2_outputs(2533) <= not((layer1_outputs(2305)) and (layer1_outputs(827)));
    layer2_outputs(2534) <= layer1_outputs(1736);
    layer2_outputs(2535) <= '0';
    layer2_outputs(2536) <= layer1_outputs(1832);
    layer2_outputs(2537) <= not((layer1_outputs(1045)) and (layer1_outputs(464)));
    layer2_outputs(2538) <= layer1_outputs(1078);
    layer2_outputs(2539) <= not(layer1_outputs(1649));
    layer2_outputs(2540) <= not((layer1_outputs(113)) and (layer1_outputs(2141)));
    layer2_outputs(2541) <= (layer1_outputs(1577)) xor (layer1_outputs(2399));
    layer2_outputs(2542) <= not((layer1_outputs(1815)) or (layer1_outputs(136)));
    layer2_outputs(2543) <= not(layer1_outputs(1328));
    layer2_outputs(2544) <= not(layer1_outputs(1234)) or (layer1_outputs(870));
    layer2_outputs(2545) <= not(layer1_outputs(1501));
    layer2_outputs(2546) <= not((layer1_outputs(1902)) xor (layer1_outputs(2444)));
    layer2_outputs(2547) <= (layer1_outputs(679)) and (layer1_outputs(1368));
    layer2_outputs(2548) <= (layer1_outputs(1454)) and not (layer1_outputs(1505));
    layer2_outputs(2549) <= not(layer1_outputs(1884));
    layer2_outputs(2550) <= layer1_outputs(1835);
    layer2_outputs(2551) <= (layer1_outputs(2295)) and (layer1_outputs(1360));
    layer2_outputs(2552) <= not(layer1_outputs(263));
    layer2_outputs(2553) <= not(layer1_outputs(1421));
    layer2_outputs(2554) <= (layer1_outputs(413)) or (layer1_outputs(2481));
    layer2_outputs(2555) <= '1';
    layer2_outputs(2556) <= not(layer1_outputs(911)) or (layer1_outputs(1110));
    layer2_outputs(2557) <= not(layer1_outputs(1893)) or (layer1_outputs(410));
    layer2_outputs(2558) <= not(layer1_outputs(927));
    layer2_outputs(2559) <= layer1_outputs(633);
    layer3_outputs(0) <= not((layer2_outputs(379)) and (layer2_outputs(1833)));
    layer3_outputs(1) <= (layer2_outputs(2305)) and not (layer2_outputs(1477));
    layer3_outputs(2) <= (layer2_outputs(1351)) or (layer2_outputs(1461));
    layer3_outputs(3) <= layer2_outputs(52);
    layer3_outputs(4) <= not((layer2_outputs(2410)) xor (layer2_outputs(529)));
    layer3_outputs(5) <= not(layer2_outputs(256));
    layer3_outputs(6) <= not(layer2_outputs(1723));
    layer3_outputs(7) <= (layer2_outputs(1779)) or (layer2_outputs(731));
    layer3_outputs(8) <= not(layer2_outputs(2266));
    layer3_outputs(9) <= not(layer2_outputs(125));
    layer3_outputs(10) <= not(layer2_outputs(636));
    layer3_outputs(11) <= layer2_outputs(1584);
    layer3_outputs(12) <= (layer2_outputs(2028)) and not (layer2_outputs(201));
    layer3_outputs(13) <= not(layer2_outputs(2015));
    layer3_outputs(14) <= not(layer2_outputs(158));
    layer3_outputs(15) <= not(layer2_outputs(1280));
    layer3_outputs(16) <= (layer2_outputs(364)) and not (layer2_outputs(1695));
    layer3_outputs(17) <= (layer2_outputs(520)) and not (layer2_outputs(31));
    layer3_outputs(18) <= not(layer2_outputs(1075)) or (layer2_outputs(1214));
    layer3_outputs(19) <= not(layer2_outputs(1503));
    layer3_outputs(20) <= layer2_outputs(494);
    layer3_outputs(21) <= (layer2_outputs(1333)) and not (layer2_outputs(2318));
    layer3_outputs(22) <= (layer2_outputs(2556)) or (layer2_outputs(815));
    layer3_outputs(23) <= layer2_outputs(235);
    layer3_outputs(24) <= layer2_outputs(206);
    layer3_outputs(25) <= not((layer2_outputs(493)) or (layer2_outputs(1869)));
    layer3_outputs(26) <= (layer2_outputs(2160)) and (layer2_outputs(1289));
    layer3_outputs(27) <= not((layer2_outputs(1647)) or (layer2_outputs(198)));
    layer3_outputs(28) <= layer2_outputs(2486);
    layer3_outputs(29) <= not(layer2_outputs(1070)) or (layer2_outputs(597));
    layer3_outputs(30) <= not((layer2_outputs(816)) xor (layer2_outputs(656)));
    layer3_outputs(31) <= not((layer2_outputs(97)) and (layer2_outputs(2146)));
    layer3_outputs(32) <= layer2_outputs(841);
    layer3_outputs(33) <= not((layer2_outputs(2004)) and (layer2_outputs(2079)));
    layer3_outputs(34) <= not(layer2_outputs(2399)) or (layer2_outputs(1907));
    layer3_outputs(35) <= not(layer2_outputs(732));
    layer3_outputs(36) <= not(layer2_outputs(857));
    layer3_outputs(37) <= not(layer2_outputs(2082)) or (layer2_outputs(1084));
    layer3_outputs(38) <= not(layer2_outputs(2493));
    layer3_outputs(39) <= (layer2_outputs(1100)) or (layer2_outputs(2143));
    layer3_outputs(40) <= not(layer2_outputs(2));
    layer3_outputs(41) <= not(layer2_outputs(1550));
    layer3_outputs(42) <= not(layer2_outputs(2056));
    layer3_outputs(43) <= not(layer2_outputs(1209)) or (layer2_outputs(1540));
    layer3_outputs(44) <= not(layer2_outputs(1565)) or (layer2_outputs(222));
    layer3_outputs(45) <= not((layer2_outputs(1008)) and (layer2_outputs(1426)));
    layer3_outputs(46) <= layer2_outputs(559);
    layer3_outputs(47) <= not(layer2_outputs(2490));
    layer3_outputs(48) <= not(layer2_outputs(279)) or (layer2_outputs(1132));
    layer3_outputs(49) <= not(layer2_outputs(578));
    layer3_outputs(50) <= (layer2_outputs(981)) xor (layer2_outputs(2378));
    layer3_outputs(51) <= not((layer2_outputs(626)) and (layer2_outputs(460)));
    layer3_outputs(52) <= not(layer2_outputs(1624)) or (layer2_outputs(447));
    layer3_outputs(53) <= (layer2_outputs(1465)) and not (layer2_outputs(1732));
    layer3_outputs(54) <= layer2_outputs(1156);
    layer3_outputs(55) <= (layer2_outputs(2415)) or (layer2_outputs(1835));
    layer3_outputs(56) <= layer2_outputs(2365);
    layer3_outputs(57) <= not(layer2_outputs(620));
    layer3_outputs(58) <= not(layer2_outputs(1101));
    layer3_outputs(59) <= layer2_outputs(1804);
    layer3_outputs(60) <= not(layer2_outputs(192)) or (layer2_outputs(1518));
    layer3_outputs(61) <= not(layer2_outputs(2331)) or (layer2_outputs(1406));
    layer3_outputs(62) <= not((layer2_outputs(305)) or (layer2_outputs(1662)));
    layer3_outputs(63) <= (layer2_outputs(196)) or (layer2_outputs(794));
    layer3_outputs(64) <= not(layer2_outputs(1319)) or (layer2_outputs(1463));
    layer3_outputs(65) <= '1';
    layer3_outputs(66) <= not(layer2_outputs(1259));
    layer3_outputs(67) <= layer2_outputs(1261);
    layer3_outputs(68) <= (layer2_outputs(2093)) and not (layer2_outputs(146));
    layer3_outputs(69) <= not(layer2_outputs(427));
    layer3_outputs(70) <= layer2_outputs(562);
    layer3_outputs(71) <= not(layer2_outputs(1906));
    layer3_outputs(72) <= not((layer2_outputs(1397)) or (layer2_outputs(2282)));
    layer3_outputs(73) <= layer2_outputs(612);
    layer3_outputs(74) <= layer2_outputs(1701);
    layer3_outputs(75) <= not((layer2_outputs(1808)) or (layer2_outputs(2303)));
    layer3_outputs(76) <= not(layer2_outputs(1353));
    layer3_outputs(77) <= (layer2_outputs(490)) and not (layer2_outputs(1258));
    layer3_outputs(78) <= not(layer2_outputs(1089));
    layer3_outputs(79) <= not(layer2_outputs(569));
    layer3_outputs(80) <= layer2_outputs(327);
    layer3_outputs(81) <= not(layer2_outputs(1310));
    layer3_outputs(82) <= (layer2_outputs(1765)) and not (layer2_outputs(1802));
    layer3_outputs(83) <= not(layer2_outputs(2277)) or (layer2_outputs(559));
    layer3_outputs(84) <= (layer2_outputs(2208)) or (layer2_outputs(2530));
    layer3_outputs(85) <= (layer2_outputs(926)) and not (layer2_outputs(306));
    layer3_outputs(86) <= not((layer2_outputs(877)) xor (layer2_outputs(1537)));
    layer3_outputs(87) <= layer2_outputs(2034);
    layer3_outputs(88) <= (layer2_outputs(2189)) and not (layer2_outputs(1692));
    layer3_outputs(89) <= not((layer2_outputs(370)) and (layer2_outputs(740)));
    layer3_outputs(90) <= '1';
    layer3_outputs(91) <= '1';
    layer3_outputs(92) <= layer2_outputs(525);
    layer3_outputs(93) <= layer2_outputs(771);
    layer3_outputs(94) <= not(layer2_outputs(32));
    layer3_outputs(95) <= '0';
    layer3_outputs(96) <= not((layer2_outputs(1787)) or (layer2_outputs(252)));
    layer3_outputs(97) <= layer2_outputs(535);
    layer3_outputs(98) <= not(layer2_outputs(2480));
    layer3_outputs(99) <= not(layer2_outputs(2052));
    layer3_outputs(100) <= layer2_outputs(1097);
    layer3_outputs(101) <= not(layer2_outputs(1553));
    layer3_outputs(102) <= '1';
    layer3_outputs(103) <= layer2_outputs(614);
    layer3_outputs(104) <= not((layer2_outputs(898)) and (layer2_outputs(2376)));
    layer3_outputs(105) <= layer2_outputs(1872);
    layer3_outputs(106) <= layer2_outputs(153);
    layer3_outputs(107) <= layer2_outputs(837);
    layer3_outputs(108) <= not(layer2_outputs(582));
    layer3_outputs(109) <= not(layer2_outputs(1659));
    layer3_outputs(110) <= not(layer2_outputs(1287));
    layer3_outputs(111) <= (layer2_outputs(888)) and not (layer2_outputs(576));
    layer3_outputs(112) <= not(layer2_outputs(152)) or (layer2_outputs(228));
    layer3_outputs(113) <= '1';
    layer3_outputs(114) <= '1';
    layer3_outputs(115) <= layer2_outputs(1533);
    layer3_outputs(116) <= (layer2_outputs(526)) and not (layer2_outputs(677));
    layer3_outputs(117) <= layer2_outputs(1245);
    layer3_outputs(118) <= (layer2_outputs(1776)) and not (layer2_outputs(433));
    layer3_outputs(119) <= not(layer2_outputs(1023));
    layer3_outputs(120) <= (layer2_outputs(2274)) and not (layer2_outputs(19));
    layer3_outputs(121) <= not(layer2_outputs(1597));
    layer3_outputs(122) <= not((layer2_outputs(1675)) and (layer2_outputs(659)));
    layer3_outputs(123) <= not(layer2_outputs(2234)) or (layer2_outputs(235));
    layer3_outputs(124) <= not(layer2_outputs(1512));
    layer3_outputs(125) <= layer2_outputs(2149);
    layer3_outputs(126) <= (layer2_outputs(541)) and not (layer2_outputs(1215));
    layer3_outputs(127) <= (layer2_outputs(1983)) and (layer2_outputs(1618));
    layer3_outputs(128) <= not(layer2_outputs(2511));
    layer3_outputs(129) <= not(layer2_outputs(1720));
    layer3_outputs(130) <= not(layer2_outputs(659));
    layer3_outputs(131) <= layer2_outputs(641);
    layer3_outputs(132) <= layer2_outputs(537);
    layer3_outputs(133) <= (layer2_outputs(749)) and not (layer2_outputs(499));
    layer3_outputs(134) <= (layer2_outputs(1069)) and not (layer2_outputs(2388));
    layer3_outputs(135) <= not(layer2_outputs(530)) or (layer2_outputs(1310));
    layer3_outputs(136) <= not((layer2_outputs(631)) and (layer2_outputs(267)));
    layer3_outputs(137) <= (layer2_outputs(2300)) or (layer2_outputs(1130));
    layer3_outputs(138) <= not((layer2_outputs(2188)) or (layer2_outputs(1975)));
    layer3_outputs(139) <= layer2_outputs(1728);
    layer3_outputs(140) <= layer2_outputs(357);
    layer3_outputs(141) <= not(layer2_outputs(1697));
    layer3_outputs(142) <= not((layer2_outputs(1400)) or (layer2_outputs(268)));
    layer3_outputs(143) <= (layer2_outputs(1902)) or (layer2_outputs(2013));
    layer3_outputs(144) <= (layer2_outputs(1843)) and not (layer2_outputs(954));
    layer3_outputs(145) <= layer2_outputs(1689);
    layer3_outputs(146) <= not((layer2_outputs(307)) and (layer2_outputs(774)));
    layer3_outputs(147) <= (layer2_outputs(1266)) and (layer2_outputs(1958));
    layer3_outputs(148) <= (layer2_outputs(775)) and not (layer2_outputs(261));
    layer3_outputs(149) <= not(layer2_outputs(1075));
    layer3_outputs(150) <= not((layer2_outputs(1296)) and (layer2_outputs(1534)));
    layer3_outputs(151) <= not(layer2_outputs(348));
    layer3_outputs(152) <= not(layer2_outputs(2240)) or (layer2_outputs(1563));
    layer3_outputs(153) <= not((layer2_outputs(2497)) or (layer2_outputs(556)));
    layer3_outputs(154) <= layer2_outputs(1962);
    layer3_outputs(155) <= layer2_outputs(1052);
    layer3_outputs(156) <= layer2_outputs(573);
    layer3_outputs(157) <= not(layer2_outputs(310));
    layer3_outputs(158) <= not(layer2_outputs(2386)) or (layer2_outputs(1479));
    layer3_outputs(159) <= not((layer2_outputs(2055)) and (layer2_outputs(2375)));
    layer3_outputs(160) <= layer2_outputs(1425);
    layer3_outputs(161) <= not(layer2_outputs(2270));
    layer3_outputs(162) <= not(layer2_outputs(1080));
    layer3_outputs(163) <= not((layer2_outputs(398)) and (layer2_outputs(1419)));
    layer3_outputs(164) <= not(layer2_outputs(1858));
    layer3_outputs(165) <= not(layer2_outputs(1898)) or (layer2_outputs(508));
    layer3_outputs(166) <= not((layer2_outputs(991)) xor (layer2_outputs(1181)));
    layer3_outputs(167) <= (layer2_outputs(1686)) or (layer2_outputs(435));
    layer3_outputs(168) <= layer2_outputs(233);
    layer3_outputs(169) <= not(layer2_outputs(1193));
    layer3_outputs(170) <= not((layer2_outputs(2467)) and (layer2_outputs(356)));
    layer3_outputs(171) <= not(layer2_outputs(392));
    layer3_outputs(172) <= layer2_outputs(365);
    layer3_outputs(173) <= layer2_outputs(289);
    layer3_outputs(174) <= not(layer2_outputs(955)) or (layer2_outputs(2010));
    layer3_outputs(175) <= (layer2_outputs(1356)) and not (layer2_outputs(2304));
    layer3_outputs(176) <= (layer2_outputs(1155)) and (layer2_outputs(1082));
    layer3_outputs(177) <= layer2_outputs(226);
    layer3_outputs(178) <= (layer2_outputs(766)) and not (layer2_outputs(1560));
    layer3_outputs(179) <= layer2_outputs(552);
    layer3_outputs(180) <= not(layer2_outputs(1875));
    layer3_outputs(181) <= layer2_outputs(1090);
    layer3_outputs(182) <= not(layer2_outputs(294));
    layer3_outputs(183) <= not(layer2_outputs(403)) or (layer2_outputs(1240));
    layer3_outputs(184) <= layer2_outputs(722);
    layer3_outputs(185) <= not((layer2_outputs(1593)) and (layer2_outputs(2093)));
    layer3_outputs(186) <= not(layer2_outputs(855));
    layer3_outputs(187) <= not(layer2_outputs(1227)) or (layer2_outputs(589));
    layer3_outputs(188) <= layer2_outputs(2073);
    layer3_outputs(189) <= layer2_outputs(1891);
    layer3_outputs(190) <= not((layer2_outputs(153)) or (layer2_outputs(113)));
    layer3_outputs(191) <= layer2_outputs(1960);
    layer3_outputs(192) <= layer2_outputs(1885);
    layer3_outputs(193) <= layer2_outputs(1028);
    layer3_outputs(194) <= '0';
    layer3_outputs(195) <= not(layer2_outputs(204));
    layer3_outputs(196) <= layer2_outputs(1022);
    layer3_outputs(197) <= not(layer2_outputs(1607)) or (layer2_outputs(338));
    layer3_outputs(198) <= layer2_outputs(1789);
    layer3_outputs(199) <= layer2_outputs(2390);
    layer3_outputs(200) <= not(layer2_outputs(1947));
    layer3_outputs(201) <= not(layer2_outputs(229)) or (layer2_outputs(768));
    layer3_outputs(202) <= layer2_outputs(2555);
    layer3_outputs(203) <= not((layer2_outputs(1735)) and (layer2_outputs(1488)));
    layer3_outputs(204) <= not(layer2_outputs(2302));
    layer3_outputs(205) <= layer2_outputs(2072);
    layer3_outputs(206) <= not(layer2_outputs(2351));
    layer3_outputs(207) <= layer2_outputs(260);
    layer3_outputs(208) <= (layer2_outputs(1120)) or (layer2_outputs(644));
    layer3_outputs(209) <= not(layer2_outputs(2363));
    layer3_outputs(210) <= not(layer2_outputs(1048));
    layer3_outputs(211) <= not(layer2_outputs(804));
    layer3_outputs(212) <= not(layer2_outputs(1632));
    layer3_outputs(213) <= not(layer2_outputs(1707));
    layer3_outputs(214) <= not(layer2_outputs(386));
    layer3_outputs(215) <= '1';
    layer3_outputs(216) <= not(layer2_outputs(1752));
    layer3_outputs(217) <= (layer2_outputs(2137)) and not (layer2_outputs(2021));
    layer3_outputs(218) <= layer2_outputs(469);
    layer3_outputs(219) <= not(layer2_outputs(1983));
    layer3_outputs(220) <= not(layer2_outputs(452));
    layer3_outputs(221) <= not(layer2_outputs(1948));
    layer3_outputs(222) <= layer2_outputs(305);
    layer3_outputs(223) <= not(layer2_outputs(2127));
    layer3_outputs(224) <= layer2_outputs(1452);
    layer3_outputs(225) <= '0';
    layer3_outputs(226) <= not(layer2_outputs(622)) or (layer2_outputs(1634));
    layer3_outputs(227) <= layer2_outputs(2432);
    layer3_outputs(228) <= (layer2_outputs(2121)) and not (layer2_outputs(2057));
    layer3_outputs(229) <= '0';
    layer3_outputs(230) <= layer2_outputs(2464);
    layer3_outputs(231) <= (layer2_outputs(462)) and not (layer2_outputs(1107));
    layer3_outputs(232) <= (layer2_outputs(1938)) and not (layer2_outputs(1292));
    layer3_outputs(233) <= not(layer2_outputs(367)) or (layer2_outputs(22));
    layer3_outputs(234) <= not(layer2_outputs(1099));
    layer3_outputs(235) <= layer2_outputs(2553);
    layer3_outputs(236) <= layer2_outputs(1862);
    layer3_outputs(237) <= layer2_outputs(1621);
    layer3_outputs(238) <= (layer2_outputs(726)) and not (layer2_outputs(187));
    layer3_outputs(239) <= not((layer2_outputs(1675)) or (layer2_outputs(834)));
    layer3_outputs(240) <= layer2_outputs(1102);
    layer3_outputs(241) <= not(layer2_outputs(36));
    layer3_outputs(242) <= (layer2_outputs(1357)) and not (layer2_outputs(2046));
    layer3_outputs(243) <= layer2_outputs(2109);
    layer3_outputs(244) <= not(layer2_outputs(1570));
    layer3_outputs(245) <= '0';
    layer3_outputs(246) <= layer2_outputs(1756);
    layer3_outputs(247) <= layer2_outputs(45);
    layer3_outputs(248) <= not(layer2_outputs(417));
    layer3_outputs(249) <= layer2_outputs(399);
    layer3_outputs(250) <= not(layer2_outputs(295)) or (layer2_outputs(2183));
    layer3_outputs(251) <= layer2_outputs(1424);
    layer3_outputs(252) <= not(layer2_outputs(278)) or (layer2_outputs(2551));
    layer3_outputs(253) <= '1';
    layer3_outputs(254) <= layer2_outputs(2296);
    layer3_outputs(255) <= not(layer2_outputs(625));
    layer3_outputs(256) <= layer2_outputs(2434);
    layer3_outputs(257) <= not(layer2_outputs(1190));
    layer3_outputs(258) <= not(layer2_outputs(1717));
    layer3_outputs(259) <= not((layer2_outputs(1306)) or (layer2_outputs(1911)));
    layer3_outputs(260) <= not(layer2_outputs(177));
    layer3_outputs(261) <= (layer2_outputs(952)) or (layer2_outputs(2552));
    layer3_outputs(262) <= layer2_outputs(1884);
    layer3_outputs(263) <= layer2_outputs(1223);
    layer3_outputs(264) <= not((layer2_outputs(1850)) and (layer2_outputs(2501)));
    layer3_outputs(265) <= not(layer2_outputs(2342)) or (layer2_outputs(441));
    layer3_outputs(266) <= (layer2_outputs(2548)) and not (layer2_outputs(1800));
    layer3_outputs(267) <= layer2_outputs(2333);
    layer3_outputs(268) <= not((layer2_outputs(768)) and (layer2_outputs(1523)));
    layer3_outputs(269) <= not(layer2_outputs(197));
    layer3_outputs(270) <= (layer2_outputs(912)) and (layer2_outputs(911));
    layer3_outputs(271) <= not(layer2_outputs(946)) or (layer2_outputs(1729));
    layer3_outputs(272) <= not(layer2_outputs(257)) or (layer2_outputs(180));
    layer3_outputs(273) <= layer2_outputs(1385);
    layer3_outputs(274) <= not(layer2_outputs(1010)) or (layer2_outputs(701));
    layer3_outputs(275) <= (layer2_outputs(1216)) or (layer2_outputs(527));
    layer3_outputs(276) <= '1';
    layer3_outputs(277) <= not(layer2_outputs(468));
    layer3_outputs(278) <= not((layer2_outputs(1066)) and (layer2_outputs(2559)));
    layer3_outputs(279) <= '1';
    layer3_outputs(280) <= layer2_outputs(1427);
    layer3_outputs(281) <= not(layer2_outputs(727));
    layer3_outputs(282) <= (layer2_outputs(1951)) and (layer2_outputs(1316));
    layer3_outputs(283) <= (layer2_outputs(1317)) and not (layer2_outputs(1966));
    layer3_outputs(284) <= not(layer2_outputs(946));
    layer3_outputs(285) <= not((layer2_outputs(456)) or (layer2_outputs(2360)));
    layer3_outputs(286) <= not(layer2_outputs(601));
    layer3_outputs(287) <= not((layer2_outputs(449)) xor (layer2_outputs(1014)));
    layer3_outputs(288) <= layer2_outputs(919);
    layer3_outputs(289) <= not(layer2_outputs(1756));
    layer3_outputs(290) <= not(layer2_outputs(1014)) or (layer2_outputs(1475));
    layer3_outputs(291) <= (layer2_outputs(2163)) and (layer2_outputs(2077));
    layer3_outputs(292) <= not(layer2_outputs(303)) or (layer2_outputs(1682));
    layer3_outputs(293) <= not(layer2_outputs(2406)) or (layer2_outputs(1450));
    layer3_outputs(294) <= not(layer2_outputs(1247));
    layer3_outputs(295) <= (layer2_outputs(227)) or (layer2_outputs(1242));
    layer3_outputs(296) <= not((layer2_outputs(2213)) xor (layer2_outputs(242)));
    layer3_outputs(297) <= not(layer2_outputs(2319));
    layer3_outputs(298) <= '0';
    layer3_outputs(299) <= not(layer2_outputs(1516)) or (layer2_outputs(1722));
    layer3_outputs(300) <= not((layer2_outputs(2168)) or (layer2_outputs(1439)));
    layer3_outputs(301) <= (layer2_outputs(2392)) and not (layer2_outputs(297));
    layer3_outputs(302) <= layer2_outputs(1643);
    layer3_outputs(303) <= (layer2_outputs(1745)) xor (layer2_outputs(345));
    layer3_outputs(304) <= layer2_outputs(1896);
    layer3_outputs(305) <= not(layer2_outputs(1231));
    layer3_outputs(306) <= not(layer2_outputs(63)) or (layer2_outputs(797));
    layer3_outputs(307) <= layer2_outputs(1282);
    layer3_outputs(308) <= layer2_outputs(1960);
    layer3_outputs(309) <= not(layer2_outputs(603)) or (layer2_outputs(1763));
    layer3_outputs(310) <= not(layer2_outputs(270));
    layer3_outputs(311) <= (layer2_outputs(778)) or (layer2_outputs(1152));
    layer3_outputs(312) <= not(layer2_outputs(709));
    layer3_outputs(313) <= not(layer2_outputs(2415));
    layer3_outputs(314) <= layer2_outputs(1752);
    layer3_outputs(315) <= layer2_outputs(535);
    layer3_outputs(316) <= not(layer2_outputs(288)) or (layer2_outputs(1652));
    layer3_outputs(317) <= not((layer2_outputs(1547)) or (layer2_outputs(1085)));
    layer3_outputs(318) <= not(layer2_outputs(937));
    layer3_outputs(319) <= not(layer2_outputs(2120));
    layer3_outputs(320) <= not(layer2_outputs(717)) or (layer2_outputs(2413));
    layer3_outputs(321) <= layer2_outputs(2396);
    layer3_outputs(322) <= (layer2_outputs(2175)) and (layer2_outputs(2478));
    layer3_outputs(323) <= layer2_outputs(1524);
    layer3_outputs(324) <= not(layer2_outputs(2533));
    layer3_outputs(325) <= not(layer2_outputs(505));
    layer3_outputs(326) <= not(layer2_outputs(1362));
    layer3_outputs(327) <= not(layer2_outputs(1932)) or (layer2_outputs(220));
    layer3_outputs(328) <= layer2_outputs(2281);
    layer3_outputs(329) <= layer2_outputs(384);
    layer3_outputs(330) <= layer2_outputs(1996);
    layer3_outputs(331) <= (layer2_outputs(2100)) and not (layer2_outputs(2273));
    layer3_outputs(332) <= (layer2_outputs(2202)) and (layer2_outputs(140));
    layer3_outputs(333) <= not(layer2_outputs(1382));
    layer3_outputs(334) <= layer2_outputs(872);
    layer3_outputs(335) <= layer2_outputs(766);
    layer3_outputs(336) <= layer2_outputs(2290);
    layer3_outputs(337) <= (layer2_outputs(2485)) and (layer2_outputs(2334));
    layer3_outputs(338) <= not(layer2_outputs(2005)) or (layer2_outputs(2361));
    layer3_outputs(339) <= layer2_outputs(2230);
    layer3_outputs(340) <= not(layer2_outputs(1168)) or (layer2_outputs(2115));
    layer3_outputs(341) <= not(layer2_outputs(1604)) or (layer2_outputs(2470));
    layer3_outputs(342) <= not((layer2_outputs(1272)) and (layer2_outputs(1694)));
    layer3_outputs(343) <= (layer2_outputs(1668)) or (layer2_outputs(827));
    layer3_outputs(344) <= not((layer2_outputs(1145)) and (layer2_outputs(1943)));
    layer3_outputs(345) <= layer2_outputs(66);
    layer3_outputs(346) <= layer2_outputs(1366);
    layer3_outputs(347) <= (layer2_outputs(1954)) and not (layer2_outputs(1544));
    layer3_outputs(348) <= not((layer2_outputs(320)) or (layer2_outputs(763)));
    layer3_outputs(349) <= not(layer2_outputs(1480)) or (layer2_outputs(1467));
    layer3_outputs(350) <= not((layer2_outputs(2221)) and (layer2_outputs(1636)));
    layer3_outputs(351) <= not(layer2_outputs(599));
    layer3_outputs(352) <= layer2_outputs(418);
    layer3_outputs(353) <= layer2_outputs(1761);
    layer3_outputs(354) <= (layer2_outputs(1192)) or (layer2_outputs(1957));
    layer3_outputs(355) <= not(layer2_outputs(2020)) or (layer2_outputs(2459));
    layer3_outputs(356) <= not(layer2_outputs(2228)) or (layer2_outputs(996));
    layer3_outputs(357) <= not(layer2_outputs(776)) or (layer2_outputs(123));
    layer3_outputs(358) <= (layer2_outputs(1661)) and not (layer2_outputs(896));
    layer3_outputs(359) <= '1';
    layer3_outputs(360) <= layer2_outputs(119);
    layer3_outputs(361) <= (layer2_outputs(1065)) and not (layer2_outputs(1342));
    layer3_outputs(362) <= layer2_outputs(311);
    layer3_outputs(363) <= not(layer2_outputs(1793));
    layer3_outputs(364) <= not(layer2_outputs(1178));
    layer3_outputs(365) <= (layer2_outputs(710)) and not (layer2_outputs(163));
    layer3_outputs(366) <= layer2_outputs(891);
    layer3_outputs(367) <= layer2_outputs(6);
    layer3_outputs(368) <= not((layer2_outputs(387)) and (layer2_outputs(1011)));
    layer3_outputs(369) <= not(layer2_outputs(729)) or (layer2_outputs(1294));
    layer3_outputs(370) <= not(layer2_outputs(2025));
    layer3_outputs(371) <= not(layer2_outputs(1336));
    layer3_outputs(372) <= (layer2_outputs(963)) and not (layer2_outputs(1820));
    layer3_outputs(373) <= '1';
    layer3_outputs(374) <= not(layer2_outputs(2244));
    layer3_outputs(375) <= (layer2_outputs(1060)) or (layer2_outputs(2063));
    layer3_outputs(376) <= not(layer2_outputs(381)) or (layer2_outputs(603));
    layer3_outputs(377) <= layer2_outputs(1765);
    layer3_outputs(378) <= not(layer2_outputs(2047));
    layer3_outputs(379) <= '0';
    layer3_outputs(380) <= layer2_outputs(1608);
    layer3_outputs(381) <= layer2_outputs(2392);
    layer3_outputs(382) <= layer2_outputs(203);
    layer3_outputs(383) <= layer2_outputs(1003);
    layer3_outputs(384) <= (layer2_outputs(1339)) and not (layer2_outputs(1963));
    layer3_outputs(385) <= not(layer2_outputs(467));
    layer3_outputs(386) <= layer2_outputs(1051);
    layer3_outputs(387) <= not((layer2_outputs(606)) xor (layer2_outputs(931)));
    layer3_outputs(388) <= layer2_outputs(1045);
    layer3_outputs(389) <= not(layer2_outputs(43));
    layer3_outputs(390) <= not((layer2_outputs(1829)) and (layer2_outputs(588)));
    layer3_outputs(391) <= (layer2_outputs(1891)) or (layer2_outputs(1955));
    layer3_outputs(392) <= not(layer2_outputs(1650)) or (layer2_outputs(1212));
    layer3_outputs(393) <= not(layer2_outputs(1167));
    layer3_outputs(394) <= (layer2_outputs(1614)) and not (layer2_outputs(84));
    layer3_outputs(395) <= not(layer2_outputs(215)) or (layer2_outputs(780));
    layer3_outputs(396) <= not(layer2_outputs(1361)) or (layer2_outputs(1013));
    layer3_outputs(397) <= not((layer2_outputs(2468)) or (layer2_outputs(2110)));
    layer3_outputs(398) <= layer2_outputs(347);
    layer3_outputs(399) <= (layer2_outputs(765)) and (layer2_outputs(2460));
    layer3_outputs(400) <= layer2_outputs(758);
    layer3_outputs(401) <= layer2_outputs(1532);
    layer3_outputs(402) <= not(layer2_outputs(337));
    layer3_outputs(403) <= not(layer2_outputs(192)) or (layer2_outputs(1054));
    layer3_outputs(404) <= not(layer2_outputs(1644));
    layer3_outputs(405) <= not(layer2_outputs(772));
    layer3_outputs(406) <= not(layer2_outputs(546));
    layer3_outputs(407) <= layer2_outputs(2201);
    layer3_outputs(408) <= (layer2_outputs(2151)) and (layer2_outputs(2424));
    layer3_outputs(409) <= '0';
    layer3_outputs(410) <= not((layer2_outputs(1791)) and (layer2_outputs(2344)));
    layer3_outputs(411) <= (layer2_outputs(350)) and not (layer2_outputs(1405));
    layer3_outputs(412) <= (layer2_outputs(1163)) and not (layer2_outputs(2080));
    layer3_outputs(413) <= (layer2_outputs(724)) and (layer2_outputs(9));
    layer3_outputs(414) <= (layer2_outputs(2399)) and not (layer2_outputs(343));
    layer3_outputs(415) <= (layer2_outputs(1451)) and not (layer2_outputs(2444));
    layer3_outputs(416) <= layer2_outputs(651);
    layer3_outputs(417) <= not(layer2_outputs(1450)) or (layer2_outputs(864));
    layer3_outputs(418) <= (layer2_outputs(1297)) and (layer2_outputs(2384));
    layer3_outputs(419) <= not(layer2_outputs(412));
    layer3_outputs(420) <= layer2_outputs(1487);
    layer3_outputs(421) <= (layer2_outputs(1681)) and not (layer2_outputs(1183));
    layer3_outputs(422) <= not(layer2_outputs(2273));
    layer3_outputs(423) <= layer2_outputs(1916);
    layer3_outputs(424) <= not(layer2_outputs(1276));
    layer3_outputs(425) <= not(layer2_outputs(1530));
    layer3_outputs(426) <= not((layer2_outputs(2413)) or (layer2_outputs(745)));
    layer3_outputs(427) <= (layer2_outputs(705)) and not (layer2_outputs(1314));
    layer3_outputs(428) <= layer2_outputs(2107);
    layer3_outputs(429) <= layer2_outputs(2040);
    layer3_outputs(430) <= not(layer2_outputs(1165));
    layer3_outputs(431) <= not(layer2_outputs(1769));
    layer3_outputs(432) <= layer2_outputs(2497);
    layer3_outputs(433) <= not((layer2_outputs(911)) and (layer2_outputs(1377)));
    layer3_outputs(434) <= (layer2_outputs(580)) and not (layer2_outputs(2543));
    layer3_outputs(435) <= layer2_outputs(2214);
    layer3_outputs(436) <= (layer2_outputs(1307)) or (layer2_outputs(1361));
    layer3_outputs(437) <= not(layer2_outputs(981));
    layer3_outputs(438) <= not(layer2_outputs(992));
    layer3_outputs(439) <= layer2_outputs(450);
    layer3_outputs(440) <= (layer2_outputs(700)) or (layer2_outputs(2112));
    layer3_outputs(441) <= not(layer2_outputs(1472));
    layer3_outputs(442) <= '1';
    layer3_outputs(443) <= '0';
    layer3_outputs(444) <= (layer2_outputs(2209)) and not (layer2_outputs(245));
    layer3_outputs(445) <= not((layer2_outputs(553)) and (layer2_outputs(1397)));
    layer3_outputs(446) <= not((layer2_outputs(998)) or (layer2_outputs(1153)));
    layer3_outputs(447) <= layer2_outputs(1428);
    layer3_outputs(448) <= not(layer2_outputs(479));
    layer3_outputs(449) <= not(layer2_outputs(2423));
    layer3_outputs(450) <= (layer2_outputs(2437)) and not (layer2_outputs(68));
    layer3_outputs(451) <= not((layer2_outputs(683)) and (layer2_outputs(1228)));
    layer3_outputs(452) <= not(layer2_outputs(2065)) or (layer2_outputs(1143));
    layer3_outputs(453) <= not(layer2_outputs(124));
    layer3_outputs(454) <= (layer2_outputs(795)) and (layer2_outputs(2076));
    layer3_outputs(455) <= not((layer2_outputs(1731)) and (layer2_outputs(1442)));
    layer3_outputs(456) <= not(layer2_outputs(2043));
    layer3_outputs(457) <= layer2_outputs(1596);
    layer3_outputs(458) <= not(layer2_outputs(1605));
    layer3_outputs(459) <= not(layer2_outputs(1149)) or (layer2_outputs(844));
    layer3_outputs(460) <= layer2_outputs(2288);
    layer3_outputs(461) <= not((layer2_outputs(112)) and (layer2_outputs(1538)));
    layer3_outputs(462) <= not(layer2_outputs(1735)) or (layer2_outputs(2064));
    layer3_outputs(463) <= not(layer2_outputs(2555));
    layer3_outputs(464) <= not(layer2_outputs(2266));
    layer3_outputs(465) <= not(layer2_outputs(1685)) or (layer2_outputs(920));
    layer3_outputs(466) <= (layer2_outputs(223)) or (layer2_outputs(2315));
    layer3_outputs(467) <= (layer2_outputs(1069)) and not (layer2_outputs(675));
    layer3_outputs(468) <= not(layer2_outputs(1839)) or (layer2_outputs(1123));
    layer3_outputs(469) <= (layer2_outputs(262)) and not (layer2_outputs(2455));
    layer3_outputs(470) <= not(layer2_outputs(159));
    layer3_outputs(471) <= layer2_outputs(95);
    layer3_outputs(472) <= not(layer2_outputs(615)) or (layer2_outputs(118));
    layer3_outputs(473) <= layer2_outputs(906);
    layer3_outputs(474) <= not((layer2_outputs(1905)) and (layer2_outputs(371)));
    layer3_outputs(475) <= layer2_outputs(1688);
    layer3_outputs(476) <= layer2_outputs(1529);
    layer3_outputs(477) <= layer2_outputs(836);
    layer3_outputs(478) <= not(layer2_outputs(146));
    layer3_outputs(479) <= not(layer2_outputs(2009)) or (layer2_outputs(2074));
    layer3_outputs(480) <= (layer2_outputs(1947)) or (layer2_outputs(1146));
    layer3_outputs(481) <= (layer2_outputs(1102)) and not (layer2_outputs(1612));
    layer3_outputs(482) <= layer2_outputs(1109);
    layer3_outputs(483) <= not(layer2_outputs(1042));
    layer3_outputs(484) <= (layer2_outputs(807)) or (layer2_outputs(1711));
    layer3_outputs(485) <= layer2_outputs(587);
    layer3_outputs(486) <= not(layer2_outputs(915));
    layer3_outputs(487) <= layer2_outputs(2327);
    layer3_outputs(488) <= not((layer2_outputs(1577)) or (layer2_outputs(2126)));
    layer3_outputs(489) <= layer2_outputs(829);
    layer3_outputs(490) <= not(layer2_outputs(690)) or (layer2_outputs(1028));
    layer3_outputs(491) <= not(layer2_outputs(1972)) or (layer2_outputs(1636));
    layer3_outputs(492) <= not((layer2_outputs(2380)) or (layer2_outputs(689)));
    layer3_outputs(493) <= (layer2_outputs(1619)) or (layer2_outputs(416));
    layer3_outputs(494) <= not(layer2_outputs(2445));
    layer3_outputs(495) <= layer2_outputs(1796);
    layer3_outputs(496) <= layer2_outputs(1067);
    layer3_outputs(497) <= not(layer2_outputs(1363));
    layer3_outputs(498) <= not((layer2_outputs(195)) and (layer2_outputs(2423)));
    layer3_outputs(499) <= not(layer2_outputs(290)) or (layer2_outputs(501));
    layer3_outputs(500) <= (layer2_outputs(1824)) or (layer2_outputs(1272));
    layer3_outputs(501) <= not(layer2_outputs(1405)) or (layer2_outputs(2283));
    layer3_outputs(502) <= not(layer2_outputs(942)) or (layer2_outputs(859));
    layer3_outputs(503) <= not(layer2_outputs(2151));
    layer3_outputs(504) <= not((layer2_outputs(1888)) or (layer2_outputs(2200)));
    layer3_outputs(505) <= layer2_outputs(1582);
    layer3_outputs(506) <= layer2_outputs(1125);
    layer3_outputs(507) <= not((layer2_outputs(1747)) or (layer2_outputs(1256)));
    layer3_outputs(508) <= not(layer2_outputs(1781));
    layer3_outputs(509) <= layer2_outputs(292);
    layer3_outputs(510) <= not(layer2_outputs(2253));
    layer3_outputs(511) <= not(layer2_outputs(941));
    layer3_outputs(512) <= not(layer2_outputs(2247));
    layer3_outputs(513) <= layer2_outputs(686);
    layer3_outputs(514) <= (layer2_outputs(2132)) xor (layer2_outputs(2111));
    layer3_outputs(515) <= layer2_outputs(1471);
    layer3_outputs(516) <= not(layer2_outputs(858));
    layer3_outputs(517) <= not(layer2_outputs(728)) or (layer2_outputs(885));
    layer3_outputs(518) <= layer2_outputs(2006);
    layer3_outputs(519) <= not(layer2_outputs(1303)) or (layer2_outputs(1456));
    layer3_outputs(520) <= not(layer2_outputs(321));
    layer3_outputs(521) <= (layer2_outputs(1480)) or (layer2_outputs(497));
    layer3_outputs(522) <= layer2_outputs(653);
    layer3_outputs(523) <= layer2_outputs(865);
    layer3_outputs(524) <= layer2_outputs(2447);
    layer3_outputs(525) <= not(layer2_outputs(594)) or (layer2_outputs(1062));
    layer3_outputs(526) <= layer2_outputs(943);
    layer3_outputs(527) <= not(layer2_outputs(990));
    layer3_outputs(528) <= layer2_outputs(1510);
    layer3_outputs(529) <= layer2_outputs(2341);
    layer3_outputs(530) <= not((layer2_outputs(783)) or (layer2_outputs(2083)));
    layer3_outputs(531) <= not(layer2_outputs(1999));
    layer3_outputs(532) <= layer2_outputs(1403);
    layer3_outputs(533) <= (layer2_outputs(2084)) xor (layer2_outputs(1122));
    layer3_outputs(534) <= '0';
    layer3_outputs(535) <= not(layer2_outputs(1466));
    layer3_outputs(536) <= layer2_outputs(968);
    layer3_outputs(537) <= not(layer2_outputs(1835)) or (layer2_outputs(473));
    layer3_outputs(538) <= not(layer2_outputs(475));
    layer3_outputs(539) <= (layer2_outputs(1259)) and (layer2_outputs(1199));
    layer3_outputs(540) <= not(layer2_outputs(327)) or (layer2_outputs(43));
    layer3_outputs(541) <= '1';
    layer3_outputs(542) <= not((layer2_outputs(1002)) and (layer2_outputs(2461)));
    layer3_outputs(543) <= '0';
    layer3_outputs(544) <= not(layer2_outputs(1925));
    layer3_outputs(545) <= layer2_outputs(1205);
    layer3_outputs(546) <= not(layer2_outputs(1382)) or (layer2_outputs(29));
    layer3_outputs(547) <= not(layer2_outputs(916));
    layer3_outputs(548) <= '1';
    layer3_outputs(549) <= layer2_outputs(1403);
    layer3_outputs(550) <= not(layer2_outputs(1721));
    layer3_outputs(551) <= layer2_outputs(2235);
    layer3_outputs(552) <= not(layer2_outputs(737)) or (layer2_outputs(82));
    layer3_outputs(553) <= not(layer2_outputs(1256));
    layer3_outputs(554) <= layer2_outputs(1017);
    layer3_outputs(555) <= not(layer2_outputs(1032)) or (layer2_outputs(1407));
    layer3_outputs(556) <= (layer2_outputs(1281)) or (layer2_outputs(738));
    layer3_outputs(557) <= layer2_outputs(2534);
    layer3_outputs(558) <= not((layer2_outputs(492)) and (layer2_outputs(2332)));
    layer3_outputs(559) <= not(layer2_outputs(1036)) or (layer2_outputs(1593));
    layer3_outputs(560) <= layer2_outputs(392);
    layer3_outputs(561) <= layer2_outputs(1378);
    layer3_outputs(562) <= not(layer2_outputs(2506)) or (layer2_outputs(1249));
    layer3_outputs(563) <= not((layer2_outputs(757)) and (layer2_outputs(437)));
    layer3_outputs(564) <= not(layer2_outputs(2039)) or (layer2_outputs(224));
    layer3_outputs(565) <= '0';
    layer3_outputs(566) <= '1';
    layer3_outputs(567) <= layer2_outputs(1879);
    layer3_outputs(568) <= layer2_outputs(2412);
    layer3_outputs(569) <= not(layer2_outputs(549));
    layer3_outputs(570) <= not(layer2_outputs(624));
    layer3_outputs(571) <= not(layer2_outputs(843)) or (layer2_outputs(1644));
    layer3_outputs(572) <= not(layer2_outputs(314));
    layer3_outputs(573) <= layer2_outputs(1609);
    layer3_outputs(574) <= not(layer2_outputs(2)) or (layer2_outputs(120));
    layer3_outputs(575) <= not(layer2_outputs(1203));
    layer3_outputs(576) <= '0';
    layer3_outputs(577) <= not(layer2_outputs(1853));
    layer3_outputs(578) <= (layer2_outputs(106)) or (layer2_outputs(65));
    layer3_outputs(579) <= not(layer2_outputs(721));
    layer3_outputs(580) <= layer2_outputs(725);
    layer3_outputs(581) <= layer2_outputs(249);
    layer3_outputs(582) <= (layer2_outputs(1134)) or (layer2_outputs(359));
    layer3_outputs(583) <= layer2_outputs(1077);
    layer3_outputs(584) <= not(layer2_outputs(209)) or (layer2_outputs(260));
    layer3_outputs(585) <= not(layer2_outputs(1722));
    layer3_outputs(586) <= (layer2_outputs(2154)) and not (layer2_outputs(565));
    layer3_outputs(587) <= not(layer2_outputs(96));
    layer3_outputs(588) <= (layer2_outputs(116)) xor (layer2_outputs(1674));
    layer3_outputs(589) <= not((layer2_outputs(1022)) and (layer2_outputs(1771)));
    layer3_outputs(590) <= not(layer2_outputs(1548));
    layer3_outputs(591) <= not((layer2_outputs(2054)) or (layer2_outputs(1575)));
    layer3_outputs(592) <= not(layer2_outputs(1654)) or (layer2_outputs(1477));
    layer3_outputs(593) <= not((layer2_outputs(2349)) and (layer2_outputs(1363)));
    layer3_outputs(594) <= '0';
    layer3_outputs(595) <= (layer2_outputs(2344)) and not (layer2_outputs(1651));
    layer3_outputs(596) <= not(layer2_outputs(2494));
    layer3_outputs(597) <= (layer2_outputs(299)) or (layer2_outputs(1965));
    layer3_outputs(598) <= not((layer2_outputs(694)) and (layer2_outputs(66)));
    layer3_outputs(599) <= not(layer2_outputs(1874)) or (layer2_outputs(988));
    layer3_outputs(600) <= not(layer2_outputs(1591));
    layer3_outputs(601) <= layer2_outputs(524);
    layer3_outputs(602) <= not(layer2_outputs(2055));
    layer3_outputs(603) <= (layer2_outputs(68)) or (layer2_outputs(73));
    layer3_outputs(604) <= (layer2_outputs(2139)) and not (layer2_outputs(1695));
    layer3_outputs(605) <= (layer2_outputs(593)) or (layer2_outputs(394));
    layer3_outputs(606) <= not(layer2_outputs(2522));
    layer3_outputs(607) <= not(layer2_outputs(269));
    layer3_outputs(608) <= '0';
    layer3_outputs(609) <= (layer2_outputs(1250)) xor (layer2_outputs(147));
    layer3_outputs(610) <= layer2_outputs(647);
    layer3_outputs(611) <= (layer2_outputs(996)) and not (layer2_outputs(1670));
    layer3_outputs(612) <= not(layer2_outputs(627));
    layer3_outputs(613) <= layer2_outputs(1094);
    layer3_outputs(614) <= layer2_outputs(2337);
    layer3_outputs(615) <= not(layer2_outputs(1061));
    layer3_outputs(616) <= not(layer2_outputs(896)) or (layer2_outputs(892));
    layer3_outputs(617) <= not(layer2_outputs(1130));
    layer3_outputs(618) <= layer2_outputs(1857);
    layer3_outputs(619) <= not(layer2_outputs(1515));
    layer3_outputs(620) <= '0';
    layer3_outputs(621) <= layer2_outputs(463);
    layer3_outputs(622) <= not(layer2_outputs(770));
    layer3_outputs(623) <= not((layer2_outputs(1821)) and (layer2_outputs(1714)));
    layer3_outputs(624) <= layer2_outputs(2269);
    layer3_outputs(625) <= not((layer2_outputs(35)) xor (layer2_outputs(868)));
    layer3_outputs(626) <= '1';
    layer3_outputs(627) <= (layer2_outputs(1230)) and not (layer2_outputs(2109));
    layer3_outputs(628) <= layer2_outputs(2311);
    layer3_outputs(629) <= (layer2_outputs(1764)) and not (layer2_outputs(2312));
    layer3_outputs(630) <= not(layer2_outputs(1566));
    layer3_outputs(631) <= '1';
    layer3_outputs(632) <= layer2_outputs(2439);
    layer3_outputs(633) <= not(layer2_outputs(1105));
    layer3_outputs(634) <= (layer2_outputs(2056)) and not (layer2_outputs(2389));
    layer3_outputs(635) <= (layer2_outputs(2524)) and not (layer2_outputs(154));
    layer3_outputs(636) <= (layer2_outputs(1525)) and not (layer2_outputs(474));
    layer3_outputs(637) <= not(layer2_outputs(1159));
    layer3_outputs(638) <= (layer2_outputs(792)) and not (layer2_outputs(2146));
    layer3_outputs(639) <= not((layer2_outputs(789)) and (layer2_outputs(2030)));
    layer3_outputs(640) <= not(layer2_outputs(1665)) or (layer2_outputs(750));
    layer3_outputs(641) <= layer2_outputs(2166);
    layer3_outputs(642) <= layer2_outputs(991);
    layer3_outputs(643) <= layer2_outputs(1592);
    layer3_outputs(644) <= not(layer2_outputs(1669)) or (layer2_outputs(2346));
    layer3_outputs(645) <= not((layer2_outputs(698)) xor (layer2_outputs(1521)));
    layer3_outputs(646) <= (layer2_outputs(2345)) xor (layer2_outputs(587));
    layer3_outputs(647) <= layer2_outputs(205);
    layer3_outputs(648) <= (layer2_outputs(2113)) or (layer2_outputs(150));
    layer3_outputs(649) <= '0';
    layer3_outputs(650) <= not(layer2_outputs(1726));
    layer3_outputs(651) <= (layer2_outputs(429)) and not (layer2_outputs(715));
    layer3_outputs(652) <= not((layer2_outputs(1600)) or (layer2_outputs(45)));
    layer3_outputs(653) <= layer2_outputs(453);
    layer3_outputs(654) <= layer2_outputs(2019);
    layer3_outputs(655) <= (layer2_outputs(255)) and (layer2_outputs(371));
    layer3_outputs(656) <= not(layer2_outputs(430));
    layer3_outputs(657) <= not((layer2_outputs(632)) or (layer2_outputs(1430)));
    layer3_outputs(658) <= not(layer2_outputs(790)) or (layer2_outputs(653));
    layer3_outputs(659) <= (layer2_outputs(2208)) and not (layer2_outputs(2525));
    layer3_outputs(660) <= not((layer2_outputs(287)) xor (layer2_outputs(1995)));
    layer3_outputs(661) <= not(layer2_outputs(2520));
    layer3_outputs(662) <= (layer2_outputs(1046)) and not (layer2_outputs(2253));
    layer3_outputs(663) <= layer2_outputs(1892);
    layer3_outputs(664) <= layer2_outputs(2350);
    layer3_outputs(665) <= not(layer2_outputs(1666)) or (layer2_outputs(107));
    layer3_outputs(666) <= not(layer2_outputs(2235));
    layer3_outputs(667) <= (layer2_outputs(1216)) or (layer2_outputs(1704));
    layer3_outputs(668) <= not(layer2_outputs(1678));
    layer3_outputs(669) <= not(layer2_outputs(2216));
    layer3_outputs(670) <= layer2_outputs(1213);
    layer3_outputs(671) <= layer2_outputs(211);
    layer3_outputs(672) <= layer2_outputs(1055);
    layer3_outputs(673) <= not(layer2_outputs(283)) or (layer2_outputs(2546));
    layer3_outputs(674) <= not(layer2_outputs(2331));
    layer3_outputs(675) <= (layer2_outputs(1603)) or (layer2_outputs(753));
    layer3_outputs(676) <= not(layer2_outputs(2201));
    layer3_outputs(677) <= (layer2_outputs(1790)) and not (layer2_outputs(2219));
    layer3_outputs(678) <= (layer2_outputs(1387)) and (layer2_outputs(482));
    layer3_outputs(679) <= not(layer2_outputs(796)) or (layer2_outputs(1118));
    layer3_outputs(680) <= layer2_outputs(322);
    layer3_outputs(681) <= not(layer2_outputs(947));
    layer3_outputs(682) <= '1';
    layer3_outputs(683) <= not((layer2_outputs(2191)) or (layer2_outputs(1243)));
    layer3_outputs(684) <= not((layer2_outputs(1512)) and (layer2_outputs(1981)));
    layer3_outputs(685) <= not(layer2_outputs(410));
    layer3_outputs(686) <= (layer2_outputs(2124)) or (layer2_outputs(1492));
    layer3_outputs(687) <= not(layer2_outputs(2192));
    layer3_outputs(688) <= not(layer2_outputs(1691));
    layer3_outputs(689) <= (layer2_outputs(2365)) and (layer2_outputs(822));
    layer3_outputs(690) <= (layer2_outputs(279)) xor (layer2_outputs(2326));
    layer3_outputs(691) <= layer2_outputs(1701);
    layer3_outputs(692) <= (layer2_outputs(1208)) and not (layer2_outputs(1874));
    layer3_outputs(693) <= not(layer2_outputs(676));
    layer3_outputs(694) <= not(layer2_outputs(1556));
    layer3_outputs(695) <= layer2_outputs(1540);
    layer3_outputs(696) <= layer2_outputs(2010);
    layer3_outputs(697) <= not(layer2_outputs(1313));
    layer3_outputs(698) <= not(layer2_outputs(1944));
    layer3_outputs(699) <= not((layer2_outputs(1856)) or (layer2_outputs(965)));
    layer3_outputs(700) <= (layer2_outputs(1125)) and not (layer2_outputs(1346));
    layer3_outputs(701) <= not((layer2_outputs(1078)) xor (layer2_outputs(471)));
    layer3_outputs(702) <= not(layer2_outputs(602));
    layer3_outputs(703) <= '1';
    layer3_outputs(704) <= not((layer2_outputs(2317)) and (layer2_outputs(1030)));
    layer3_outputs(705) <= (layer2_outputs(2132)) and (layer2_outputs(383));
    layer3_outputs(706) <= layer2_outputs(1485);
    layer3_outputs(707) <= (layer2_outputs(1115)) and not (layer2_outputs(1831));
    layer3_outputs(708) <= not(layer2_outputs(1445));
    layer3_outputs(709) <= layer2_outputs(2426);
    layer3_outputs(710) <= not(layer2_outputs(1552));
    layer3_outputs(711) <= not(layer2_outputs(1727));
    layer3_outputs(712) <= (layer2_outputs(502)) or (layer2_outputs(1116));
    layer3_outputs(713) <= (layer2_outputs(2065)) and (layer2_outputs(2079));
    layer3_outputs(714) <= layer2_outputs(210);
    layer3_outputs(715) <= not(layer2_outputs(2528)) or (layer2_outputs(949));
    layer3_outputs(716) <= (layer2_outputs(48)) and (layer2_outputs(1472));
    layer3_outputs(717) <= layer2_outputs(303);
    layer3_outputs(718) <= not(layer2_outputs(2473));
    layer3_outputs(719) <= not(layer2_outputs(1385));
    layer3_outputs(720) <= not(layer2_outputs(1772)) or (layer2_outputs(1664));
    layer3_outputs(721) <= not(layer2_outputs(1091));
    layer3_outputs(722) <= (layer2_outputs(2430)) and not (layer2_outputs(220));
    layer3_outputs(723) <= '0';
    layer3_outputs(724) <= not((layer2_outputs(585)) and (layer2_outputs(1007)));
    layer3_outputs(725) <= layer2_outputs(2016);
    layer3_outputs(726) <= (layer2_outputs(1416)) or (layer2_outputs(1436));
    layer3_outputs(727) <= not((layer2_outputs(2364)) or (layer2_outputs(2136)));
    layer3_outputs(728) <= not((layer2_outputs(639)) xor (layer2_outputs(2521)));
    layer3_outputs(729) <= (layer2_outputs(707)) and (layer2_outputs(533));
    layer3_outputs(730) <= (layer2_outputs(813)) and not (layer2_outputs(1950));
    layer3_outputs(731) <= not(layer2_outputs(2357));
    layer3_outputs(732) <= not(layer2_outputs(247));
    layer3_outputs(733) <= (layer2_outputs(124)) and not (layer2_outputs(2531));
    layer3_outputs(734) <= not(layer2_outputs(1857));
    layer3_outputs(735) <= not((layer2_outputs(557)) or (layer2_outputs(1705)));
    layer3_outputs(736) <= layer2_outputs(365);
    layer3_outputs(737) <= layer2_outputs(1298);
    layer3_outputs(738) <= layer2_outputs(2161);
    layer3_outputs(739) <= not(layer2_outputs(1967)) or (layer2_outputs(59));
    layer3_outputs(740) <= not(layer2_outputs(1486)) or (layer2_outputs(1129));
    layer3_outputs(741) <= not(layer2_outputs(2217));
    layer3_outputs(742) <= layer2_outputs(1093);
    layer3_outputs(743) <= (layer2_outputs(2098)) and not (layer2_outputs(1127));
    layer3_outputs(744) <= (layer2_outputs(503)) xor (layer2_outputs(1544));
    layer3_outputs(745) <= not(layer2_outputs(2091));
    layer3_outputs(746) <= (layer2_outputs(253)) and not (layer2_outputs(1298));
    layer3_outputs(747) <= not(layer2_outputs(602));
    layer3_outputs(748) <= layer2_outputs(1268);
    layer3_outputs(749) <= not((layer2_outputs(434)) and (layer2_outputs(2282)));
    layer3_outputs(750) <= (layer2_outputs(1589)) and not (layer2_outputs(135));
    layer3_outputs(751) <= layer2_outputs(573);
    layer3_outputs(752) <= not((layer2_outputs(1738)) and (layer2_outputs(2153)));
    layer3_outputs(753) <= not((layer2_outputs(2061)) and (layer2_outputs(779)));
    layer3_outputs(754) <= layer2_outputs(542);
    layer3_outputs(755) <= not(layer2_outputs(1426)) or (layer2_outputs(1942));
    layer3_outputs(756) <= not(layer2_outputs(598)) or (layer2_outputs(2474));
    layer3_outputs(757) <= not((layer2_outputs(219)) and (layer2_outputs(1308)));
    layer3_outputs(758) <= not(layer2_outputs(2320));
    layer3_outputs(759) <= not(layer2_outputs(1498));
    layer3_outputs(760) <= not(layer2_outputs(1904));
    layer3_outputs(761) <= layer2_outputs(296);
    layer3_outputs(762) <= not(layer2_outputs(1217)) or (layer2_outputs(1859));
    layer3_outputs(763) <= not((layer2_outputs(139)) or (layer2_outputs(1224)));
    layer3_outputs(764) <= not(layer2_outputs(1994)) or (layer2_outputs(1950));
    layer3_outputs(765) <= not((layer2_outputs(2090)) or (layer2_outputs(1590)));
    layer3_outputs(766) <= layer2_outputs(736);
    layer3_outputs(767) <= layer2_outputs(2425);
    layer3_outputs(768) <= '0';
    layer3_outputs(769) <= not(layer2_outputs(2469));
    layer3_outputs(770) <= not(layer2_outputs(636));
    layer3_outputs(771) <= '1';
    layer3_outputs(772) <= (layer2_outputs(1181)) xor (layer2_outputs(1193));
    layer3_outputs(773) <= not(layer2_outputs(2114)) or (layer2_outputs(107));
    layer3_outputs(774) <= layer2_outputs(173);
    layer3_outputs(775) <= '0';
    layer3_outputs(776) <= not(layer2_outputs(265));
    layer3_outputs(777) <= not(layer2_outputs(2034));
    layer3_outputs(778) <= not((layer2_outputs(189)) xor (layer2_outputs(1599)));
    layer3_outputs(779) <= not(layer2_outputs(196)) or (layer2_outputs(1241));
    layer3_outputs(780) <= layer2_outputs(176);
    layer3_outputs(781) <= (layer2_outputs(1606)) and not (layer2_outputs(1415));
    layer3_outputs(782) <= layer2_outputs(2337);
    layer3_outputs(783) <= not(layer2_outputs(858));
    layer3_outputs(784) <= not(layer2_outputs(1806)) or (layer2_outputs(2120));
    layer3_outputs(785) <= not((layer2_outputs(1332)) or (layer2_outputs(1674)));
    layer3_outputs(786) <= (layer2_outputs(466)) xor (layer2_outputs(1218));
    layer3_outputs(787) <= not((layer2_outputs(1757)) and (layer2_outputs(2112)));
    layer3_outputs(788) <= (layer2_outputs(450)) and not (layer2_outputs(1804));
    layer3_outputs(789) <= layer2_outputs(67);
    layer3_outputs(790) <= layer2_outputs(241);
    layer3_outputs(791) <= (layer2_outputs(609)) and not (layer2_outputs(1334));
    layer3_outputs(792) <= not(layer2_outputs(835));
    layer3_outputs(793) <= layer2_outputs(616);
    layer3_outputs(794) <= not(layer2_outputs(1245)) or (layer2_outputs(253));
    layer3_outputs(795) <= layer2_outputs(642);
    layer3_outputs(796) <= layer2_outputs(2284);
    layer3_outputs(797) <= not((layer2_outputs(200)) or (layer2_outputs(1989)));
    layer3_outputs(798) <= layer2_outputs(1194);
    layer3_outputs(799) <= not(layer2_outputs(1056));
    layer3_outputs(800) <= not(layer2_outputs(985)) or (layer2_outputs(2066));
    layer3_outputs(801) <= not((layer2_outputs(916)) and (layer2_outputs(518)));
    layer3_outputs(802) <= not(layer2_outputs(812));
    layer3_outputs(803) <= layer2_outputs(243);
    layer3_outputs(804) <= layer2_outputs(713);
    layer3_outputs(805) <= not(layer2_outputs(292)) or (layer2_outputs(1646));
    layer3_outputs(806) <= not(layer2_outputs(2514)) or (layer2_outputs(1463));
    layer3_outputs(807) <= not(layer2_outputs(716));
    layer3_outputs(808) <= (layer2_outputs(1581)) and not (layer2_outputs(315));
    layer3_outputs(809) <= (layer2_outputs(1920)) and not (layer2_outputs(1961));
    layer3_outputs(810) <= layer2_outputs(1751);
    layer3_outputs(811) <= layer2_outputs(954);
    layer3_outputs(812) <= not(layer2_outputs(317));
    layer3_outputs(813) <= not((layer2_outputs(938)) or (layer2_outputs(2024)));
    layer3_outputs(814) <= (layer2_outputs(1576)) and (layer2_outputs(2086));
    layer3_outputs(815) <= not(layer2_outputs(614));
    layer3_outputs(816) <= not(layer2_outputs(994));
    layer3_outputs(817) <= not(layer2_outputs(2173)) or (layer2_outputs(1015));
    layer3_outputs(818) <= not(layer2_outputs(1759)) or (layer2_outputs(2042));
    layer3_outputs(819) <= layer2_outputs(2154);
    layer3_outputs(820) <= layer2_outputs(82);
    layer3_outputs(821) <= (layer2_outputs(421)) and not (layer2_outputs(28));
    layer3_outputs(822) <= not(layer2_outputs(422)) or (layer2_outputs(696));
    layer3_outputs(823) <= layer2_outputs(2404);
    layer3_outputs(824) <= (layer2_outputs(1931)) and not (layer2_outputs(622));
    layer3_outputs(825) <= not((layer2_outputs(1928)) or (layer2_outputs(2329)));
    layer3_outputs(826) <= layer2_outputs(781);
    layer3_outputs(827) <= layer2_outputs(1304);
    layer3_outputs(828) <= (layer2_outputs(530)) and not (layer2_outputs(619));
    layer3_outputs(829) <= '1';
    layer3_outputs(830) <= not(layer2_outputs(1039));
    layer3_outputs(831) <= not(layer2_outputs(1685));
    layer3_outputs(832) <= not(layer2_outputs(944)) or (layer2_outputs(2189));
    layer3_outputs(833) <= not(layer2_outputs(1826));
    layer3_outputs(834) <= not((layer2_outputs(1096)) xor (layer2_outputs(194)));
    layer3_outputs(835) <= (layer2_outputs(2394)) and (layer2_outputs(1142));
    layer3_outputs(836) <= (layer2_outputs(106)) and (layer2_outputs(1774));
    layer3_outputs(837) <= layer2_outputs(2358);
    layer3_outputs(838) <= (layer2_outputs(258)) and not (layer2_outputs(592));
    layer3_outputs(839) <= not(layer2_outputs(2552));
    layer3_outputs(840) <= '0';
    layer3_outputs(841) <= layer2_outputs(1333);
    layer3_outputs(842) <= not(layer2_outputs(312)) or (layer2_outputs(1473));
    layer3_outputs(843) <= (layer2_outputs(927)) xor (layer2_outputs(712));
    layer3_outputs(844) <= not(layer2_outputs(2207));
    layer3_outputs(845) <= not(layer2_outputs(1317));
    layer3_outputs(846) <= not(layer2_outputs(379));
    layer3_outputs(847) <= not(layer2_outputs(2431));
    layer3_outputs(848) <= (layer2_outputs(2036)) and not (layer2_outputs(1565));
    layer3_outputs(849) <= '1';
    layer3_outputs(850) <= (layer2_outputs(585)) or (layer2_outputs(1579));
    layer3_outputs(851) <= layer2_outputs(154);
    layer3_outputs(852) <= (layer2_outputs(1072)) and not (layer2_outputs(1485));
    layer3_outputs(853) <= not((layer2_outputs(1229)) or (layer2_outputs(2471)));
    layer3_outputs(854) <= not(layer2_outputs(1724));
    layer3_outputs(855) <= not(layer2_outputs(1807)) or (layer2_outputs(632));
    layer3_outputs(856) <= layer2_outputs(325);
    layer3_outputs(857) <= not((layer2_outputs(746)) or (layer2_outputs(1797)));
    layer3_outputs(858) <= not((layer2_outputs(2336)) or (layer2_outputs(1652)));
    layer3_outputs(859) <= not(layer2_outputs(691));
    layer3_outputs(860) <= not(layer2_outputs(2152));
    layer3_outputs(861) <= not(layer2_outputs(1630));
    layer3_outputs(862) <= (layer2_outputs(2436)) and not (layer2_outputs(820));
    layer3_outputs(863) <= not((layer2_outputs(1278)) xor (layer2_outputs(1768)));
    layer3_outputs(864) <= layer2_outputs(2276);
    layer3_outputs(865) <= layer2_outputs(649);
    layer3_outputs(866) <= layer2_outputs(1456);
    layer3_outputs(867) <= not(layer2_outputs(2251));
    layer3_outputs(868) <= not(layer2_outputs(1012));
    layer3_outputs(869) <= '1';
    layer3_outputs(870) <= not(layer2_outputs(1285));
    layer3_outputs(871) <= not(layer2_outputs(1826));
    layer3_outputs(872) <= layer2_outputs(1992);
    layer3_outputs(873) <= not(layer2_outputs(190));
    layer3_outputs(874) <= not(layer2_outputs(784));
    layer3_outputs(875) <= not((layer2_outputs(862)) or (layer2_outputs(1661)));
    layer3_outputs(876) <= '0';
    layer3_outputs(877) <= layer2_outputs(1517);
    layer3_outputs(878) <= not(layer2_outputs(1517));
    layer3_outputs(879) <= not((layer2_outputs(1638)) and (layer2_outputs(813)));
    layer3_outputs(880) <= not(layer2_outputs(1470)) or (layer2_outputs(152));
    layer3_outputs(881) <= '0';
    layer3_outputs(882) <= not(layer2_outputs(1819));
    layer3_outputs(883) <= not(layer2_outputs(1718)) or (layer2_outputs(2069));
    layer3_outputs(884) <= not(layer2_outputs(1135));
    layer3_outputs(885) <= layer2_outputs(2509);
    layer3_outputs(886) <= not(layer2_outputs(1876)) or (layer2_outputs(2411));
    layer3_outputs(887) <= not((layer2_outputs(1578)) or (layer2_outputs(54)));
    layer3_outputs(888) <= not(layer2_outputs(548)) or (layer2_outputs(708));
    layer3_outputs(889) <= not(layer2_outputs(203));
    layer3_outputs(890) <= not(layer2_outputs(1325));
    layer3_outputs(891) <= not(layer2_outputs(76)) or (layer2_outputs(1895));
    layer3_outputs(892) <= layer2_outputs(762);
    layer3_outputs(893) <= not(layer2_outputs(2098)) or (layer2_outputs(1024));
    layer3_outputs(894) <= '1';
    layer3_outputs(895) <= not((layer2_outputs(699)) or (layer2_outputs(2058)));
    layer3_outputs(896) <= not(layer2_outputs(93));
    layer3_outputs(897) <= not((layer2_outputs(2472)) and (layer2_outputs(744)));
    layer3_outputs(898) <= not(layer2_outputs(1741)) or (layer2_outputs(799));
    layer3_outputs(899) <= (layer2_outputs(1097)) and not (layer2_outputs(520));
    layer3_outputs(900) <= not(layer2_outputs(344)) or (layer2_outputs(617));
    layer3_outputs(901) <= not((layer2_outputs(1824)) xor (layer2_outputs(1784)));
    layer3_outputs(902) <= not(layer2_outputs(55));
    layer3_outputs(903) <= not((layer2_outputs(2203)) and (layer2_outputs(1376)));
    layer3_outputs(904) <= layer2_outputs(357);
    layer3_outputs(905) <= layer2_outputs(1131);
    layer3_outputs(906) <= not((layer2_outputs(1117)) xor (layer2_outputs(2463)));
    layer3_outputs(907) <= layer2_outputs(127);
    layer3_outputs(908) <= layer2_outputs(2259);
    layer3_outputs(909) <= '0';
    layer3_outputs(910) <= layer2_outputs(2187);
    layer3_outputs(911) <= layer2_outputs(531);
    layer3_outputs(912) <= layer2_outputs(744);
    layer3_outputs(913) <= layer2_outputs(1421);
    layer3_outputs(914) <= not(layer2_outputs(33));
    layer3_outputs(915) <= not(layer2_outputs(2279)) or (layer2_outputs(1364));
    layer3_outputs(916) <= layer2_outputs(1229);
    layer3_outputs(917) <= '1';
    layer3_outputs(918) <= not(layer2_outputs(1335)) or (layer2_outputs(1315));
    layer3_outputs(919) <= not(layer2_outputs(93)) or (layer2_outputs(179));
    layer3_outputs(920) <= (layer2_outputs(934)) and (layer2_outputs(980));
    layer3_outputs(921) <= layer2_outputs(1918);
    layer3_outputs(922) <= layer2_outputs(713);
    layer3_outputs(923) <= (layer2_outputs(2513)) and not (layer2_outputs(845));
    layer3_outputs(924) <= '0';
    layer3_outputs(925) <= not(layer2_outputs(1837)) or (layer2_outputs(851));
    layer3_outputs(926) <= (layer2_outputs(491)) or (layer2_outputs(2219));
    layer3_outputs(927) <= '1';
    layer3_outputs(928) <= layer2_outputs(759);
    layer3_outputs(929) <= (layer2_outputs(384)) xor (layer2_outputs(1754));
    layer3_outputs(930) <= layer2_outputs(1299);
    layer3_outputs(931) <= (layer2_outputs(353)) and not (layer2_outputs(1438));
    layer3_outputs(932) <= not(layer2_outputs(2540));
    layer3_outputs(933) <= not((layer2_outputs(89)) and (layer2_outputs(1971)));
    layer3_outputs(934) <= not((layer2_outputs(1737)) and (layer2_outputs(1396)));
    layer3_outputs(935) <= not(layer2_outputs(1956));
    layer3_outputs(936) <= not(layer2_outputs(1055));
    layer3_outputs(937) <= (layer2_outputs(1546)) and not (layer2_outputs(1266));
    layer3_outputs(938) <= layer2_outputs(1797);
    layer3_outputs(939) <= not(layer2_outputs(308));
    layer3_outputs(940) <= layer2_outputs(1769);
    layer3_outputs(941) <= not(layer2_outputs(34));
    layer3_outputs(942) <= not(layer2_outputs(355));
    layer3_outputs(943) <= (layer2_outputs(2450)) or (layer2_outputs(451));
    layer3_outputs(944) <= '0';
    layer3_outputs(945) <= not((layer2_outputs(1814)) or (layer2_outputs(2141)));
    layer3_outputs(946) <= not((layer2_outputs(1827)) xor (layer2_outputs(2150)));
    layer3_outputs(947) <= layer2_outputs(30);
    layer3_outputs(948) <= (layer2_outputs(607)) and (layer2_outputs(953));
    layer3_outputs(949) <= not((layer2_outputs(542)) and (layer2_outputs(378)));
    layer3_outputs(950) <= not(layer2_outputs(228)) or (layer2_outputs(1329));
    layer3_outputs(951) <= layer2_outputs(700);
    layer3_outputs(952) <= layer2_outputs(1437);
    layer3_outputs(953) <= (layer2_outputs(286)) and not (layer2_outputs(11));
    layer3_outputs(954) <= layer2_outputs(1901);
    layer3_outputs(955) <= not(layer2_outputs(2081)) or (layer2_outputs(1367));
    layer3_outputs(956) <= (layer2_outputs(1411)) and (layer2_outputs(1187));
    layer3_outputs(957) <= '0';
    layer3_outputs(958) <= '1';
    layer3_outputs(959) <= not(layer2_outputs(936));
    layer3_outputs(960) <= not(layer2_outputs(1806)) or (layer2_outputs(1423));
    layer3_outputs(961) <= not(layer2_outputs(590)) or (layer2_outputs(2051));
    layer3_outputs(962) <= layer2_outputs(1291);
    layer3_outputs(963) <= (layer2_outputs(2442)) and (layer2_outputs(1074));
    layer3_outputs(964) <= '1';
    layer3_outputs(965) <= layer2_outputs(1562);
    layer3_outputs(966) <= not(layer2_outputs(1922)) or (layer2_outputs(918));
    layer3_outputs(967) <= not(layer2_outputs(1997));
    layer3_outputs(968) <= not((layer2_outputs(420)) and (layer2_outputs(1606)));
    layer3_outputs(969) <= not(layer2_outputs(1880)) or (layer2_outputs(1109));
    layer3_outputs(970) <= layer2_outputs(1828);
    layer3_outputs(971) <= layer2_outputs(2454);
    layer3_outputs(972) <= not(layer2_outputs(1941));
    layer3_outputs(973) <= layer2_outputs(990);
    layer3_outputs(974) <= not((layer2_outputs(674)) or (layer2_outputs(1978)));
    layer3_outputs(975) <= layer2_outputs(546);
    layer3_outputs(976) <= layer2_outputs(289);
    layer3_outputs(977) <= layer2_outputs(1182);
    layer3_outputs(978) <= layer2_outputs(238);
    layer3_outputs(979) <= not(layer2_outputs(388));
    layer3_outputs(980) <= layer2_outputs(2545);
    layer3_outputs(981) <= layer2_outputs(1150);
    layer3_outputs(982) <= layer2_outputs(2233);
    layer3_outputs(983) <= layer2_outputs(678);
    layer3_outputs(984) <= not(layer2_outputs(212));
    layer3_outputs(985) <= not(layer2_outputs(686));
    layer3_outputs(986) <= (layer2_outputs(1716)) and (layer2_outputs(463));
    layer3_outputs(987) <= (layer2_outputs(883)) and not (layer2_outputs(1202));
    layer3_outputs(988) <= not(layer2_outputs(151)) or (layer2_outputs(2076));
    layer3_outputs(989) <= '0';
    layer3_outputs(990) <= not(layer2_outputs(2478));
    layer3_outputs(991) <= (layer2_outputs(687)) or (layer2_outputs(380));
    layer3_outputs(992) <= (layer2_outputs(1528)) or (layer2_outputs(1508));
    layer3_outputs(993) <= not(layer2_outputs(2000));
    layer3_outputs(994) <= not((layer2_outputs(1803)) or (layer2_outputs(1378)));
    layer3_outputs(995) <= '0';
    layer3_outputs(996) <= not(layer2_outputs(2159));
    layer3_outputs(997) <= not(layer2_outputs(1128));
    layer3_outputs(998) <= not((layer2_outputs(607)) and (layer2_outputs(1807)));
    layer3_outputs(999) <= not(layer2_outputs(2354)) or (layer2_outputs(266));
    layer3_outputs(1000) <= (layer2_outputs(2107)) and not (layer2_outputs(37));
    layer3_outputs(1001) <= not((layer2_outputs(1895)) or (layer2_outputs(900)));
    layer3_outputs(1002) <= not(layer2_outputs(324)) or (layer2_outputs(880));
    layer3_outputs(1003) <= not(layer2_outputs(562));
    layer3_outputs(1004) <= (layer2_outputs(180)) and (layer2_outputs(1996));
    layer3_outputs(1005) <= '1';
    layer3_outputs(1006) <= not(layer2_outputs(333));
    layer3_outputs(1007) <= not((layer2_outputs(1346)) and (layer2_outputs(1655)));
    layer3_outputs(1008) <= layer2_outputs(193);
    layer3_outputs(1009) <= (layer2_outputs(442)) and not (layer2_outputs(1898));
    layer3_outputs(1010) <= (layer2_outputs(1616)) and (layer2_outputs(2472));
    layer3_outputs(1011) <= (layer2_outputs(1186)) or (layer2_outputs(2048));
    layer3_outputs(1012) <= (layer2_outputs(2518)) and not (layer2_outputs(1980));
    layer3_outputs(1013) <= layer2_outputs(370);
    layer3_outputs(1014) <= layer2_outputs(822);
    layer3_outputs(1015) <= layer2_outputs(496);
    layer3_outputs(1016) <= layer2_outputs(1974);
    layer3_outputs(1017) <= layer2_outputs(608);
    layer3_outputs(1018) <= not((layer2_outputs(778)) or (layer2_outputs(807)));
    layer3_outputs(1019) <= not(layer2_outputs(874)) or (layer2_outputs(2163));
    layer3_outputs(1020) <= not(layer2_outputs(999));
    layer3_outputs(1021) <= layer2_outputs(1684);
    layer3_outputs(1022) <= (layer2_outputs(1103)) or (layer2_outputs(2053));
    layer3_outputs(1023) <= layer2_outputs(230);
    layer3_outputs(1024) <= not((layer2_outputs(1791)) xor (layer2_outputs(2099)));
    layer3_outputs(1025) <= (layer2_outputs(1106)) and not (layer2_outputs(769));
    layer3_outputs(1026) <= not(layer2_outputs(206));
    layer3_outputs(1027) <= (layer2_outputs(374)) and not (layer2_outputs(92));
    layer3_outputs(1028) <= not(layer2_outputs(1457));
    layer3_outputs(1029) <= layer2_outputs(1684);
    layer3_outputs(1030) <= layer2_outputs(437);
    layer3_outputs(1031) <= not(layer2_outputs(1509));
    layer3_outputs(1032) <= not(layer2_outputs(507));
    layer3_outputs(1033) <= not(layer2_outputs(1751)) or (layer2_outputs(923));
    layer3_outputs(1034) <= not((layer2_outputs(928)) and (layer2_outputs(1467)));
    layer3_outputs(1035) <= not(layer2_outputs(2190));
    layer3_outputs(1036) <= layer2_outputs(1476);
    layer3_outputs(1037) <= (layer2_outputs(319)) and not (layer2_outputs(890));
    layer3_outputs(1038) <= not((layer2_outputs(2031)) or (layer2_outputs(276)));
    layer3_outputs(1039) <= not(layer2_outputs(272)) or (layer2_outputs(2123));
    layer3_outputs(1040) <= not((layer2_outputs(1220)) xor (layer2_outputs(511)));
    layer3_outputs(1041) <= not((layer2_outputs(1578)) xor (layer2_outputs(1921)));
    layer3_outputs(1042) <= not(layer2_outputs(2067));
    layer3_outputs(1043) <= (layer2_outputs(1381)) and (layer2_outputs(2547));
    layer3_outputs(1044) <= (layer2_outputs(506)) or (layer2_outputs(767));
    layer3_outputs(1045) <= layer2_outputs(567);
    layer3_outputs(1046) <= not(layer2_outputs(794));
    layer3_outputs(1047) <= (layer2_outputs(1408)) and not (layer2_outputs(1513));
    layer3_outputs(1048) <= not(layer2_outputs(2160));
    layer3_outputs(1049) <= (layer2_outputs(993)) and (layer2_outputs(1376));
    layer3_outputs(1050) <= not(layer2_outputs(150));
    layer3_outputs(1051) <= not(layer2_outputs(599));
    layer3_outputs(1052) <= (layer2_outputs(1698)) and (layer2_outputs(38));
    layer3_outputs(1053) <= (layer2_outputs(1507)) or (layer2_outputs(2463));
    layer3_outputs(1054) <= not(layer2_outputs(1015)) or (layer2_outputs(2417));
    layer3_outputs(1055) <= not(layer2_outputs(1708));
    layer3_outputs(1056) <= (layer2_outputs(1454)) or (layer2_outputs(605));
    layer3_outputs(1057) <= not(layer2_outputs(950));
    layer3_outputs(1058) <= not(layer2_outputs(1496)) or (layer2_outputs(929));
    layer3_outputs(1059) <= not(layer2_outputs(162)) or (layer2_outputs(2101));
    layer3_outputs(1060) <= not(layer2_outputs(2417));
    layer3_outputs(1061) <= not(layer2_outputs(1025));
    layer3_outputs(1062) <= not(layer2_outputs(2539)) or (layer2_outputs(2403));
    layer3_outputs(1063) <= '1';
    layer3_outputs(1064) <= not(layer2_outputs(511));
    layer3_outputs(1065) <= layer2_outputs(2004);
    layer3_outputs(1066) <= (layer2_outputs(1703)) and (layer2_outputs(1810));
    layer3_outputs(1067) <= (layer2_outputs(1255)) and not (layer2_outputs(2297));
    layer3_outputs(1068) <= (layer2_outputs(907)) or (layer2_outputs(331));
    layer3_outputs(1069) <= not(layer2_outputs(2140));
    layer3_outputs(1070) <= layer2_outputs(1732);
    layer3_outputs(1071) <= layer2_outputs(299);
    layer3_outputs(1072) <= not(layer2_outputs(1098));
    layer3_outputs(1073) <= (layer2_outputs(458)) and not (layer2_outputs(1061));
    layer3_outputs(1074) <= '1';
    layer3_outputs(1075) <= not((layer2_outputs(1493)) or (layer2_outputs(2400)));
    layer3_outputs(1076) <= not(layer2_outputs(829));
    layer3_outputs(1077) <= not((layer2_outputs(1534)) or (layer2_outputs(57)));
    layer3_outputs(1078) <= not(layer2_outputs(1388));
    layer3_outputs(1079) <= not((layer2_outputs(2262)) xor (layer2_outputs(1253)));
    layer3_outputs(1080) <= (layer2_outputs(2131)) or (layer2_outputs(331));
    layer3_outputs(1081) <= not(layer2_outputs(821)) or (layer2_outputs(1696));
    layer3_outputs(1082) <= not(layer2_outputs(1188));
    layer3_outputs(1083) <= not(layer2_outputs(1040));
    layer3_outputs(1084) <= (layer2_outputs(1882)) and not (layer2_outputs(2082));
    layer3_outputs(1085) <= (layer2_outputs(1651)) or (layer2_outputs(1589));
    layer3_outputs(1086) <= (layer2_outputs(1267)) xor (layer2_outputs(2366));
    layer3_outputs(1087) <= not(layer2_outputs(2171));
    layer3_outputs(1088) <= layer2_outputs(1913);
    layer3_outputs(1089) <= not(layer2_outputs(1057)) or (layer2_outputs(1274));
    layer3_outputs(1090) <= not((layer2_outputs(1037)) or (layer2_outputs(2246)));
    layer3_outputs(1091) <= (layer2_outputs(2118)) or (layer2_outputs(2277));
    layer3_outputs(1092) <= not(layer2_outputs(1873)) or (layer2_outputs(1580));
    layer3_outputs(1093) <= '1';
    layer3_outputs(1094) <= not((layer2_outputs(1019)) and (layer2_outputs(1799)));
    layer3_outputs(1095) <= not(layer2_outputs(2203)) or (layer2_outputs(2317));
    layer3_outputs(1096) <= layer2_outputs(1839);
    layer3_outputs(1097) <= '1';
    layer3_outputs(1098) <= layer2_outputs(132);
    layer3_outputs(1099) <= not(layer2_outputs(2275));
    layer3_outputs(1100) <= (layer2_outputs(935)) and not (layer2_outputs(885));
    layer3_outputs(1101) <= not(layer2_outputs(298));
    layer3_outputs(1102) <= not(layer2_outputs(1085)) or (layer2_outputs(2222));
    layer3_outputs(1103) <= not(layer2_outputs(1514)) or (layer2_outputs(1116));
    layer3_outputs(1104) <= layer2_outputs(2291);
    layer3_outputs(1105) <= not(layer2_outputs(119));
    layer3_outputs(1106) <= '1';
    layer3_outputs(1107) <= not(layer2_outputs(236));
    layer3_outputs(1108) <= not(layer2_outputs(410)) or (layer2_outputs(60));
    layer3_outputs(1109) <= not(layer2_outputs(800)) or (layer2_outputs(729));
    layer3_outputs(1110) <= not(layer2_outputs(1104)) or (layer2_outputs(406));
    layer3_outputs(1111) <= not(layer2_outputs(966));
    layer3_outputs(1112) <= (layer2_outputs(2272)) and not (layer2_outputs(2122));
    layer3_outputs(1113) <= not((layer2_outputs(11)) or (layer2_outputs(2249)));
    layer3_outputs(1114) <= not(layer2_outputs(2367)) or (layer2_outputs(2475));
    layer3_outputs(1115) <= layer2_outputs(2505);
    layer3_outputs(1116) <= not(layer2_outputs(823));
    layer3_outputs(1117) <= not((layer2_outputs(1321)) or (layer2_outputs(47)));
    layer3_outputs(1118) <= not((layer2_outputs(754)) xor (layer2_outputs(97)));
    layer3_outputs(1119) <= not(layer2_outputs(1917));
    layer3_outputs(1120) <= (layer2_outputs(663)) and (layer2_outputs(1825));
    layer3_outputs(1121) <= (layer2_outputs(1535)) xor (layer2_outputs(514));
    layer3_outputs(1122) <= not(layer2_outputs(1183));
    layer3_outputs(1123) <= not(layer2_outputs(1952));
    layer3_outputs(1124) <= (layer2_outputs(2421)) or (layer2_outputs(1033));
    layer3_outputs(1125) <= not(layer2_outputs(870));
    layer3_outputs(1126) <= '1';
    layer3_outputs(1127) <= not((layer2_outputs(1576)) or (layer2_outputs(531)));
    layer3_outputs(1128) <= (layer2_outputs(2359)) and (layer2_outputs(1772));
    layer3_outputs(1129) <= layer2_outputs(1160);
    layer3_outputs(1130) <= not((layer2_outputs(977)) xor (layer2_outputs(1979)));
    layer3_outputs(1131) <= (layer2_outputs(1371)) and (layer2_outputs(287));
    layer3_outputs(1132) <= layer2_outputs(2432);
    layer3_outputs(1133) <= layer2_outputs(963);
    layer3_outputs(1134) <= layer2_outputs(90);
    layer3_outputs(1135) <= layer2_outputs(588);
    layer3_outputs(1136) <= not(layer2_outputs(1142));
    layer3_outputs(1137) <= not(layer2_outputs(1624));
    layer3_outputs(1138) <= (layer2_outputs(1443)) and (layer2_outputs(216));
    layer3_outputs(1139) <= not((layer2_outputs(730)) or (layer2_outputs(1264)));
    layer3_outputs(1140) <= (layer2_outputs(242)) xor (layer2_outputs(2366));
    layer3_outputs(1141) <= (layer2_outputs(438)) and not (layer2_outputs(971));
    layer3_outputs(1142) <= not((layer2_outputs(2396)) or (layer2_outputs(1151)));
    layer3_outputs(1143) <= layer2_outputs(676);
    layer3_outputs(1144) <= (layer2_outputs(2449)) or (layer2_outputs(1392));
    layer3_outputs(1145) <= layer2_outputs(2263);
    layer3_outputs(1146) <= layer2_outputs(825);
    layer3_outputs(1147) <= not((layer2_outputs(969)) and (layer2_outputs(1209)));
    layer3_outputs(1148) <= (layer2_outputs(881)) and (layer2_outputs(2236));
    layer3_outputs(1149) <= not((layer2_outputs(611)) or (layer2_outputs(1734)));
    layer3_outputs(1150) <= layer2_outputs(105);
    layer3_outputs(1151) <= (layer2_outputs(839)) and not (layer2_outputs(2084));
    layer3_outputs(1152) <= (layer2_outputs(0)) and (layer2_outputs(5));
    layer3_outputs(1153) <= not(layer2_outputs(1710));
    layer3_outputs(1154) <= not((layer2_outputs(1372)) and (layer2_outputs(456)));
    layer3_outputs(1155) <= (layer2_outputs(2496)) and not (layer2_outputs(2088));
    layer3_outputs(1156) <= layer2_outputs(1977);
    layer3_outputs(1157) <= '0';
    layer3_outputs(1158) <= layer2_outputs(55);
    layer3_outputs(1159) <= layer2_outputs(1325);
    layer3_outputs(1160) <= not((layer2_outputs(171)) or (layer2_outputs(1812)));
    layer3_outputs(1161) <= not((layer2_outputs(2124)) and (layer2_outputs(1195)));
    layer3_outputs(1162) <= not(layer2_outputs(2499));
    layer3_outputs(1163) <= not((layer2_outputs(966)) and (layer2_outputs(361)));
    layer3_outputs(1164) <= '0';
    layer3_outputs(1165) <= not(layer2_outputs(1511));
    layer3_outputs(1166) <= '1';
    layer3_outputs(1167) <= layer2_outputs(1815);
    layer3_outputs(1168) <= not(layer2_outputs(1598)) or (layer2_outputs(1089));
    layer3_outputs(1169) <= not(layer2_outputs(2162));
    layer3_outputs(1170) <= (layer2_outputs(2496)) xor (layer2_outputs(2409));
    layer3_outputs(1171) <= (layer2_outputs(40)) and not (layer2_outputs(976));
    layer3_outputs(1172) <= not(layer2_outputs(1282));
    layer3_outputs(1173) <= not(layer2_outputs(1000));
    layer3_outputs(1174) <= (layer2_outputs(1875)) and not (layer2_outputs(477));
    layer3_outputs(1175) <= not((layer2_outputs(2488)) and (layer2_outputs(658)));
    layer3_outputs(1176) <= layer2_outputs(478);
    layer3_outputs(1177) <= layer2_outputs(1286);
    layer3_outputs(1178) <= not((layer2_outputs(2495)) and (layer2_outputs(145)));
    layer3_outputs(1179) <= not(layer2_outputs(54));
    layer3_outputs(1180) <= not(layer2_outputs(1819)) or (layer2_outputs(574));
    layer3_outputs(1181) <= not(layer2_outputs(2441));
    layer3_outputs(1182) <= layer2_outputs(2468);
    layer3_outputs(1183) <= '1';
    layer3_outputs(1184) <= layer2_outputs(2310);
    layer3_outputs(1185) <= layer2_outputs(1392);
    layer3_outputs(1186) <= not(layer2_outputs(1643)) or (layer2_outputs(848));
    layer3_outputs(1187) <= '0';
    layer3_outputs(1188) <= not(layer2_outputs(1267));
    layer3_outputs(1189) <= not(layer2_outputs(95));
    layer3_outputs(1190) <= (layer2_outputs(294)) and (layer2_outputs(903));
    layer3_outputs(1191) <= not(layer2_outputs(652)) or (layer2_outputs(2288));
    layer3_outputs(1192) <= not(layer2_outputs(1322)) or (layer2_outputs(1646));
    layer3_outputs(1193) <= not(layer2_outputs(815));
    layer3_outputs(1194) <= (layer2_outputs(1541)) and (layer2_outputs(945));
    layer3_outputs(1195) <= not(layer2_outputs(1916));
    layer3_outputs(1196) <= layer2_outputs(1242);
    layer3_outputs(1197) <= not((layer2_outputs(449)) xor (layer2_outputs(2295)));
    layer3_outputs(1198) <= (layer2_outputs(1564)) or (layer2_outputs(495));
    layer3_outputs(1199) <= (layer2_outputs(849)) and not (layer2_outputs(2465));
    layer3_outputs(1200) <= not(layer2_outputs(1536));
    layer3_outputs(1201) <= not(layer2_outputs(1127));
    layer3_outputs(1202) <= '0';
    layer3_outputs(1203) <= not(layer2_outputs(861));
    layer3_outputs(1204) <= not(layer2_outputs(1459));
    layer3_outputs(1205) <= not(layer2_outputs(2040));
    layer3_outputs(1206) <= not(layer2_outputs(1737));
    layer3_outputs(1207) <= layer2_outputs(1159);
    layer3_outputs(1208) <= layer2_outputs(233);
    layer3_outputs(1209) <= not(layer2_outputs(586));
    layer3_outputs(1210) <= not(layer2_outputs(956));
    layer3_outputs(1211) <= (layer2_outputs(443)) and (layer2_outputs(500));
    layer3_outputs(1212) <= not(layer2_outputs(1464)) or (layer2_outputs(720));
    layer3_outputs(1213) <= '0';
    layer3_outputs(1214) <= '1';
    layer3_outputs(1215) <= layer2_outputs(1508);
    layer3_outputs(1216) <= (layer2_outputs(208)) and not (layer2_outputs(631));
    layer3_outputs(1217) <= '1';
    layer3_outputs(1218) <= not(layer2_outputs(1864));
    layer3_outputs(1219) <= (layer2_outputs(1559)) and (layer2_outputs(1099));
    layer3_outputs(1220) <= layer2_outputs(1759);
    layer3_outputs(1221) <= not(layer2_outputs(1111)) or (layer2_outputs(328));
    layer3_outputs(1222) <= not(layer2_outputs(940));
    layer3_outputs(1223) <= not(layer2_outputs(2104));
    layer3_outputs(1224) <= layer2_outputs(826);
    layer3_outputs(1225) <= layer2_outputs(1390);
    layer3_outputs(1226) <= (layer2_outputs(218)) and (layer2_outputs(304));
    layer3_outputs(1227) <= (layer2_outputs(348)) and (layer2_outputs(774));
    layer3_outputs(1228) <= (layer2_outputs(761)) xor (layer2_outputs(2018));
    layer3_outputs(1229) <= (layer2_outputs(581)) and not (layer2_outputs(2157));
    layer3_outputs(1230) <= (layer2_outputs(401)) xor (layer2_outputs(1058));
    layer3_outputs(1231) <= not(layer2_outputs(1845)) or (layer2_outputs(1542));
    layer3_outputs(1232) <= layer2_outputs(1301);
    layer3_outputs(1233) <= layer2_outputs(1853);
    layer3_outputs(1234) <= not(layer2_outputs(821));
    layer3_outputs(1235) <= '0';
    layer3_outputs(1236) <= layer2_outputs(1700);
    layer3_outputs(1237) <= not(layer2_outputs(393));
    layer3_outputs(1238) <= (layer2_outputs(2150)) and (layer2_outputs(1226));
    layer3_outputs(1239) <= layer2_outputs(15);
    layer3_outputs(1240) <= layer2_outputs(49);
    layer3_outputs(1241) <= (layer2_outputs(2049)) and not (layer2_outputs(1336));
    layer3_outputs(1242) <= layer2_outputs(194);
    layer3_outputs(1243) <= (layer2_outputs(2223)) and (layer2_outputs(1101));
    layer3_outputs(1244) <= (layer2_outputs(1358)) and not (layer2_outputs(764));
    layer3_outputs(1245) <= not(layer2_outputs(2335));
    layer3_outputs(1246) <= (layer2_outputs(1670)) or (layer2_outputs(1583));
    layer3_outputs(1247) <= not(layer2_outputs(286));
    layer3_outputs(1248) <= not(layer2_outputs(765));
    layer3_outputs(1249) <= not((layer2_outputs(2373)) and (layer2_outputs(669)));
    layer3_outputs(1250) <= not(layer2_outputs(1581));
    layer3_outputs(1251) <= not(layer2_outputs(322));
    layer3_outputs(1252) <= not(layer2_outputs(2389));
    layer3_outputs(1253) <= not(layer2_outputs(378)) or (layer2_outputs(2029));
    layer3_outputs(1254) <= not(layer2_outputs(1150));
    layer3_outputs(1255) <= not((layer2_outputs(1100)) and (layer2_outputs(24)));
    layer3_outputs(1256) <= not(layer2_outputs(925));
    layer3_outputs(1257) <= layer2_outputs(1605);
    layer3_outputs(1258) <= (layer2_outputs(214)) and (layer2_outputs(1728));
    layer3_outputs(1259) <= (layer2_outputs(316)) and (layer2_outputs(666));
    layer3_outputs(1260) <= not(layer2_outputs(780));
    layer3_outputs(1261) <= not(layer2_outputs(377));
    layer3_outputs(1262) <= layer2_outputs(1398);
    layer3_outputs(1263) <= (layer2_outputs(185)) xor (layer2_outputs(2136));
    layer3_outputs(1264) <= layer2_outputs(2558);
    layer3_outputs(1265) <= layer2_outputs(941);
    layer3_outputs(1266) <= layer2_outputs(268);
    layer3_outputs(1267) <= (layer2_outputs(174)) xor (layer2_outputs(1157));
    layer3_outputs(1268) <= (layer2_outputs(2103)) and not (layer2_outputs(2182));
    layer3_outputs(1269) <= not(layer2_outputs(552));
    layer3_outputs(1270) <= not(layer2_outputs(1154));
    layer3_outputs(1271) <= not(layer2_outputs(1145));
    layer3_outputs(1272) <= layer2_outputs(1860);
    layer3_outputs(1273) <= not((layer2_outputs(846)) xor (layer2_outputs(56)));
    layer3_outputs(1274) <= layer2_outputs(28);
    layer3_outputs(1275) <= not((layer2_outputs(915)) and (layer2_outputs(1869)));
    layer3_outputs(1276) <= (layer2_outputs(72)) xor (layer2_outputs(354));
    layer3_outputs(1277) <= not((layer2_outputs(857)) and (layer2_outputs(1036)));
    layer3_outputs(1278) <= not(layer2_outputs(1350)) or (layer2_outputs(2028));
    layer3_outputs(1279) <= layer2_outputs(1867);
    layer3_outputs(1280) <= not(layer2_outputs(2324)) or (layer2_outputs(1354));
    layer3_outputs(1281) <= not(layer2_outputs(1630));
    layer3_outputs(1282) <= layer2_outputs(2330);
    layer3_outputs(1283) <= layer2_outputs(271);
    layer3_outputs(1284) <= not(layer2_outputs(1474)) or (layer2_outputs(2001));
    layer3_outputs(1285) <= not(layer2_outputs(2005)) or (layer2_outputs(1164));
    layer3_outputs(1286) <= layer2_outputs(1855);
    layer3_outputs(1287) <= layer2_outputs(1768);
    layer3_outputs(1288) <= not(layer2_outputs(2369));
    layer3_outputs(1289) <= (layer2_outputs(1588)) and (layer2_outputs(706));
    layer3_outputs(1290) <= (layer2_outputs(1293)) and not (layer2_outputs(1355));
    layer3_outputs(1291) <= layer2_outputs(723);
    layer3_outputs(1292) <= not((layer2_outputs(46)) or (layer2_outputs(1892)));
    layer3_outputs(1293) <= not(layer2_outputs(672));
    layer3_outputs(1294) <= (layer2_outputs(584)) and not (layer2_outputs(1163));
    layer3_outputs(1295) <= layer2_outputs(1865);
    layer3_outputs(1296) <= not(layer2_outputs(2233));
    layer3_outputs(1297) <= not(layer2_outputs(1468)) or (layer2_outputs(186));
    layer3_outputs(1298) <= layer2_outputs(105);
    layer3_outputs(1299) <= not(layer2_outputs(920));
    layer3_outputs(1300) <= '1';
    layer3_outputs(1301) <= (layer2_outputs(1585)) or (layer2_outputs(2550));
    layer3_outputs(1302) <= not(layer2_outputs(1513));
    layer3_outputs(1303) <= (layer2_outputs(2227)) and not (layer2_outputs(1939));
    layer3_outputs(1304) <= '1';
    layer3_outputs(1305) <= layer2_outputs(468);
    layer3_outputs(1306) <= layer2_outputs(650);
    layer3_outputs(1307) <= not(layer2_outputs(1394));
    layer3_outputs(1308) <= not((layer2_outputs(143)) or (layer2_outputs(1462)));
    layer3_outputs(1309) <= layer2_outputs(618);
    layer3_outputs(1310) <= layer2_outputs(1416);
    layer3_outputs(1311) <= (layer2_outputs(1248)) xor (layer2_outputs(820));
    layer3_outputs(1312) <= not(layer2_outputs(382));
    layer3_outputs(1313) <= layer2_outputs(2239);
    layer3_outputs(1314) <= not(layer2_outputs(2199));
    layer3_outputs(1315) <= not(layer2_outputs(1494));
    layer3_outputs(1316) <= (layer2_outputs(1319)) and not (layer2_outputs(2393));
    layer3_outputs(1317) <= not((layer2_outputs(824)) xor (layer2_outputs(2229)));
    layer3_outputs(1318) <= not((layer2_outputs(498)) and (layer2_outputs(489)));
    layer3_outputs(1319) <= not(layer2_outputs(1715)) or (layer2_outputs(444));
    layer3_outputs(1320) <= (layer2_outputs(128)) and not (layer2_outputs(1258));
    layer3_outputs(1321) <= not((layer2_outputs(2185)) and (layer2_outputs(1981)));
    layer3_outputs(1322) <= layer2_outputs(2424);
    layer3_outputs(1323) <= (layer2_outputs(3)) xor (layer2_outputs(1445));
    layer3_outputs(1324) <= '0';
    layer3_outputs(1325) <= not((layer2_outputs(471)) xor (layer2_outputs(2071)));
    layer3_outputs(1326) <= not(layer2_outputs(1471));
    layer3_outputs(1327) <= not(layer2_outputs(1295)) or (layer2_outputs(884));
    layer3_outputs(1328) <= (layer2_outputs(1667)) and not (layer2_outputs(1934));
    layer3_outputs(1329) <= not(layer2_outputs(2205));
    layer3_outputs(1330) <= not(layer2_outputs(671));
    layer3_outputs(1331) <= not((layer2_outputs(17)) xor (layer2_outputs(2519)));
    layer3_outputs(1332) <= layer2_outputs(1910);
    layer3_outputs(1333) <= not(layer2_outputs(61)) or (layer2_outputs(1096));
    layer3_outputs(1334) <= not(layer2_outputs(1962));
    layer3_outputs(1335) <= (layer2_outputs(1275)) or (layer2_outputs(1841));
    layer3_outputs(1336) <= layer2_outputs(1271);
    layer3_outputs(1337) <= not(layer2_outputs(1236));
    layer3_outputs(1338) <= layer2_outputs(1992);
    layer3_outputs(1339) <= not((layer2_outputs(560)) or (layer2_outputs(1369)));
    layer3_outputs(1340) <= not(layer2_outputs(2198));
    layer3_outputs(1341) <= (layer2_outputs(1656)) and not (layer2_outputs(2381));
    layer3_outputs(1342) <= layer2_outputs(1309);
    layer3_outputs(1343) <= not(layer2_outputs(878));
    layer3_outputs(1344) <= (layer2_outputs(1269)) and not (layer2_outputs(2477));
    layer3_outputs(1345) <= not(layer2_outputs(1291));
    layer3_outputs(1346) <= (layer2_outputs(2315)) and not (layer2_outputs(1191));
    layer3_outputs(1347) <= not(layer2_outputs(1025)) or (layer2_outputs(2554));
    layer3_outputs(1348) <= not(layer2_outputs(1609)) or (layer2_outputs(1506));
    layer3_outputs(1349) <= not(layer2_outputs(853));
    layer3_outputs(1350) <= '0';
    layer3_outputs(1351) <= layer2_outputs(840);
    layer3_outputs(1352) <= layer2_outputs(83);
    layer3_outputs(1353) <= not(layer2_outputs(189));
    layer3_outputs(1354) <= layer2_outputs(1871);
    layer3_outputs(1355) <= not(layer2_outputs(2264)) or (layer2_outputs(847));
    layer3_outputs(1356) <= not(layer2_outputs(1915));
    layer3_outputs(1357) <= not(layer2_outputs(1633));
    layer3_outputs(1358) <= layer2_outputs(2479);
    layer3_outputs(1359) <= not(layer2_outputs(586));
    layer3_outputs(1360) <= (layer2_outputs(611)) and (layer2_outputs(513));
    layer3_outputs(1361) <= layer2_outputs(782);
    layer3_outputs(1362) <= (layer2_outputs(2420)) and not (layer2_outputs(2407));
    layer3_outputs(1363) <= layer2_outputs(393);
    layer3_outputs(1364) <= not(layer2_outputs(2526));
    layer3_outputs(1365) <= layer2_outputs(862);
    layer3_outputs(1366) <= not(layer2_outputs(2147));
    layer3_outputs(1367) <= layer2_outputs(2140);
    layer3_outputs(1368) <= layer2_outputs(2504);
    layer3_outputs(1369) <= not(layer2_outputs(2139));
    layer3_outputs(1370) <= (layer2_outputs(255)) and (layer2_outputs(164));
    layer3_outputs(1371) <= not(layer2_outputs(2043));
    layer3_outputs(1372) <= not((layer2_outputs(1504)) or (layer2_outputs(271)));
    layer3_outputs(1373) <= not((layer2_outputs(1320)) or (layer2_outputs(2242)));
    layer3_outputs(1374) <= not(layer2_outputs(1678));
    layer3_outputs(1375) <= layer2_outputs(625);
    layer3_outputs(1376) <= (layer2_outputs(1246)) and not (layer2_outputs(947));
    layer3_outputs(1377) <= not((layer2_outputs(2202)) and (layer2_outputs(316)));
    layer3_outputs(1378) <= '1';
    layer3_outputs(1379) <= layer2_outputs(525);
    layer3_outputs(1380) <= layer2_outputs(2422);
    layer3_outputs(1381) <= '1';
    layer3_outputs(1382) <= layer2_outputs(1760);
    layer3_outputs(1383) <= layer2_outputs(1034);
    layer3_outputs(1384) <= (layer2_outputs(2078)) xor (layer2_outputs(986));
    layer3_outputs(1385) <= not(layer2_outputs(2241)) or (layer2_outputs(808));
    layer3_outputs(1386) <= (layer2_outputs(1883)) and (layer2_outputs(398));
    layer3_outputs(1387) <= layer2_outputs(1663);
    layer3_outputs(1388) <= not((layer2_outputs(1908)) or (layer2_outputs(319)));
    layer3_outputs(1389) <= (layer2_outputs(275)) and (layer2_outputs(1635));
    layer3_outputs(1390) <= '0';
    layer3_outputs(1391) <= not((layer2_outputs(474)) or (layer2_outputs(263)));
    layer3_outputs(1392) <= layer2_outputs(685);
    layer3_outputs(1393) <= not(layer2_outputs(1623)) or (layer2_outputs(1017));
    layer3_outputs(1394) <= not(layer2_outputs(1381));
    layer3_outputs(1395) <= layer2_outputs(545);
    layer3_outputs(1396) <= not(layer2_outputs(1337)) or (layer2_outputs(2397));
    layer3_outputs(1397) <= layer2_outputs(2493);
    layer3_outputs(1398) <= not(layer2_outputs(650)) or (layer2_outputs(1912));
    layer3_outputs(1399) <= layer2_outputs(102);
    layer3_outputs(1400) <= layer2_outputs(17);
    layer3_outputs(1401) <= (layer2_outputs(1557)) and not (layer2_outputs(1002));
    layer3_outputs(1402) <= layer2_outputs(989);
    layer3_outputs(1403) <= (layer2_outputs(1618)) and not (layer2_outputs(649));
    layer3_outputs(1404) <= (layer2_outputs(1043)) and not (layer2_outputs(1443));
    layer3_outputs(1405) <= layer2_outputs(1949);
    layer3_outputs(1406) <= (layer2_outputs(521)) and (layer2_outputs(325));
    layer3_outputs(1407) <= (layer2_outputs(1010)) or (layer2_outputs(646));
    layer3_outputs(1408) <= (layer2_outputs(679)) or (layer2_outputs(2355));
    layer3_outputs(1409) <= (layer2_outputs(99)) or (layer2_outputs(930));
    layer3_outputs(1410) <= not(layer2_outputs(245)) or (layer2_outputs(1574));
    layer3_outputs(1411) <= (layer2_outputs(1623)) and not (layer2_outputs(1446));
    layer3_outputs(1412) <= not((layer2_outputs(373)) xor (layer2_outputs(1250)));
    layer3_outputs(1413) <= not(layer2_outputs(536)) or (layer2_outputs(1464));
    layer3_outputs(1414) <= layer2_outputs(1740);
    layer3_outputs(1415) <= not(layer2_outputs(2026)) or (layer2_outputs(978));
    layer3_outputs(1416) <= not(layer2_outputs(1899));
    layer3_outputs(1417) <= (layer2_outputs(1637)) and not (layer2_outputs(1626));
    layer3_outputs(1418) <= (layer2_outputs(547)) and not (layer2_outputs(1913));
    layer3_outputs(1419) <= not(layer2_outputs(1626));
    layer3_outputs(1420) <= layer2_outputs(660);
    layer3_outputs(1421) <= layer2_outputs(566);
    layer3_outputs(1422) <= not(layer2_outputs(448)) or (layer2_outputs(750));
    layer3_outputs(1423) <= not((layer2_outputs(2476)) and (layer2_outputs(1805)));
    layer3_outputs(1424) <= layer2_outputs(515);
    layer3_outputs(1425) <= (layer2_outputs(1758)) or (layer2_outputs(101));
    layer3_outputs(1426) <= not(layer2_outputs(366));
    layer3_outputs(1427) <= not((layer2_outputs(1369)) or (layer2_outputs(1422)));
    layer3_outputs(1428) <= not((layer2_outputs(1205)) xor (layer2_outputs(258)));
    layer3_outputs(1429) <= (layer2_outputs(2549)) and (layer2_outputs(465));
    layer3_outputs(1430) <= (layer2_outputs(1861)) and not (layer2_outputs(1854));
    layer3_outputs(1431) <= not(layer2_outputs(18)) or (layer2_outputs(674));
    layer3_outputs(1432) <= not(layer2_outputs(2014));
    layer3_outputs(1433) <= not((layer2_outputs(2018)) or (layer2_outputs(165)));
    layer3_outputs(1434) <= not((layer2_outputs(2083)) and (layer2_outputs(951)));
    layer3_outputs(1435) <= (layer2_outputs(1213)) and not (layer2_outputs(975));
    layer3_outputs(1436) <= (layer2_outputs(2404)) and (layer2_outputs(1610));
    layer3_outputs(1437) <= not((layer2_outputs(1940)) xor (layer2_outputs(2130)));
    layer3_outputs(1438) <= (layer2_outputs(16)) and not (layer2_outputs(64));
    layer3_outputs(1439) <= layer2_outputs(753);
    layer3_outputs(1440) <= layer2_outputs(481);
    layer3_outputs(1441) <= layer2_outputs(984);
    layer3_outputs(1442) <= (layer2_outputs(575)) and (layer2_outputs(1689));
    layer3_outputs(1443) <= not((layer2_outputs(1311)) xor (layer2_outputs(527)));
    layer3_outputs(1444) <= not(layer2_outputs(668));
    layer3_outputs(1445) <= (layer2_outputs(2504)) or (layer2_outputs(1057));
    layer3_outputs(1446) <= layer2_outputs(1729);
    layer3_outputs(1447) <= (layer2_outputs(2513)) xor (layer2_outputs(1018));
    layer3_outputs(1448) <= (layer2_outputs(893)) and not (layer2_outputs(2541));
    layer3_outputs(1449) <= layer2_outputs(337);
    layer3_outputs(1450) <= (layer2_outputs(2508)) and (layer2_outputs(1744));
    layer3_outputs(1451) <= not((layer2_outputs(1334)) or (layer2_outputs(1673)));
    layer3_outputs(1452) <= not(layer2_outputs(109));
    layer3_outputs(1453) <= not(layer2_outputs(111)) or (layer2_outputs(1091));
    layer3_outputs(1454) <= (layer2_outputs(1263)) and not (layer2_outputs(1275));
    layer3_outputs(1455) <= not(layer2_outputs(453));
    layer3_outputs(1456) <= not(layer2_outputs(2542));
    layer3_outputs(1457) <= not(layer2_outputs(1990));
    layer3_outputs(1458) <= not(layer2_outputs(2447));
    layer3_outputs(1459) <= not(layer2_outputs(2293)) or (layer2_outputs(2540));
    layer3_outputs(1460) <= not((layer2_outputs(1318)) or (layer2_outputs(1083)));
    layer3_outputs(1461) <= not((layer2_outputs(1189)) and (layer2_outputs(2453)));
    layer3_outputs(1462) <= not(layer2_outputs(630));
    layer3_outputs(1463) <= not(layer2_outputs(459));
    layer3_outputs(1464) <= not(layer2_outputs(380));
    layer3_outputs(1465) <= '1';
    layer3_outputs(1466) <= (layer2_outputs(1718)) and (layer2_outputs(2036));
    layer3_outputs(1467) <= not((layer2_outputs(755)) or (layer2_outputs(2430)));
    layer3_outputs(1468) <= not(layer2_outputs(2377));
    layer3_outputs(1469) <= (layer2_outputs(1886)) and (layer2_outputs(1706));
    layer3_outputs(1470) <= layer2_outputs(96);
    layer3_outputs(1471) <= layer2_outputs(423);
    layer3_outputs(1472) <= layer2_outputs(809);
    layer3_outputs(1473) <= not(layer2_outputs(2103));
    layer3_outputs(1474) <= not((layer2_outputs(2041)) xor (layer2_outputs(2229)));
    layer3_outputs(1475) <= not(layer2_outputs(2217)) or (layer2_outputs(2436));
    layer3_outputs(1476) <= not(layer2_outputs(2111));
    layer3_outputs(1477) <= (layer2_outputs(2007)) and (layer2_outputs(2357));
    layer3_outputs(1478) <= not(layer2_outputs(1435)) or (layer2_outputs(1));
    layer3_outputs(1479) <= not(layer2_outputs(491));
    layer3_outputs(1480) <= not(layer2_outputs(1811));
    layer3_outputs(1481) <= not((layer2_outputs(1026)) xor (layer2_outputs(1764)));
    layer3_outputs(1482) <= '0';
    layer3_outputs(1483) <= '0';
    layer3_outputs(1484) <= not(layer2_outputs(2342));
    layer3_outputs(1485) <= (layer2_outputs(1136)) or (layer2_outputs(1147));
    layer3_outputs(1486) <= (layer2_outputs(2075)) and not (layer2_outputs(1841));
    layer3_outputs(1487) <= layer2_outputs(2451);
    layer3_outputs(1488) <= not(layer2_outputs(866));
    layer3_outputs(1489) <= layer2_outputs(2299);
    layer3_outputs(1490) <= (layer2_outputs(2284)) and (layer2_outputs(334));
    layer3_outputs(1491) <= not(layer2_outputs(229)) or (layer2_outputs(1914));
    layer3_outputs(1492) <= (layer2_outputs(2296)) and not (layer2_outputs(101));
    layer3_outputs(1493) <= (layer2_outputs(2311)) and not (layer2_outputs(851));
    layer3_outputs(1494) <= not(layer2_outputs(823));
    layer3_outputs(1495) <= (layer2_outputs(56)) and (layer2_outputs(2237));
    layer3_outputs(1496) <= not(layer2_outputs(2172));
    layer3_outputs(1497) <= not(layer2_outputs(2184));
    layer3_outputs(1498) <= (layer2_outputs(1071)) or (layer2_outputs(53));
    layer3_outputs(1499) <= layer2_outputs(2074);
    layer3_outputs(1500) <= (layer2_outputs(2256)) and (layer2_outputs(2520));
    layer3_outputs(1501) <= not((layer2_outputs(1409)) and (layer2_outputs(723)));
    layer3_outputs(1502) <= '1';
    layer3_outputs(1503) <= layer2_outputs(1568);
    layer3_outputs(1504) <= not(layer2_outputs(1889));
    layer3_outputs(1505) <= not(layer2_outputs(200)) or (layer2_outputs(2442));
    layer3_outputs(1506) <= (layer2_outputs(2038)) or (layer2_outputs(1847));
    layer3_outputs(1507) <= layer2_outputs(758);
    layer3_outputs(1508) <= not(layer2_outputs(2121)) or (layer2_outputs(833));
    layer3_outputs(1509) <= (layer2_outputs(572)) xor (layer2_outputs(368));
    layer3_outputs(1510) <= (layer2_outputs(662)) and not (layer2_outputs(1165));
    layer3_outputs(1511) <= not((layer2_outputs(1490)) or (layer2_outputs(70)));
    layer3_outputs(1512) <= (layer2_outputs(1200)) or (layer2_outputs(2024));
    layer3_outputs(1513) <= layer2_outputs(2387);
    layer3_outputs(1514) <= (layer2_outputs(2265)) and not (layer2_outputs(1423));
    layer3_outputs(1515) <= not(layer2_outputs(865));
    layer3_outputs(1516) <= not(layer2_outputs(70)) or (layer2_outputs(161));
    layer3_outputs(1517) <= not(layer2_outputs(475));
    layer3_outputs(1518) <= not(layer2_outputs(173)) or (layer2_outputs(2401));
    layer3_outputs(1519) <= not(layer2_outputs(1491));
    layer3_outputs(1520) <= not(layer2_outputs(26));
    layer3_outputs(1521) <= layer2_outputs(1178);
    layer3_outputs(1522) <= not(layer2_outputs(1041));
    layer3_outputs(1523) <= not(layer2_outputs(284));
    layer3_outputs(1524) <= not(layer2_outputs(1156)) or (layer2_outputs(570));
    layer3_outputs(1525) <= layer2_outputs(698);
    layer3_outputs(1526) <= (layer2_outputs(2441)) and not (layer2_outputs(1273));
    layer3_outputs(1527) <= not(layer2_outputs(1786));
    layer3_outputs(1528) <= layer2_outputs(2362);
    layer3_outputs(1529) <= '0';
    layer3_outputs(1530) <= '1';
    layer3_outputs(1531) <= not((layer2_outputs(1489)) xor (layer2_outputs(1340)));
    layer3_outputs(1532) <= not(layer2_outputs(1884));
    layer3_outputs(1533) <= not(layer2_outputs(545));
    layer3_outputs(1534) <= not((layer2_outputs(1524)) and (layer2_outputs(1836)));
    layer3_outputs(1535) <= (layer2_outputs(1968)) and not (layer2_outputs(1400));
    layer3_outputs(1536) <= not((layer2_outputs(688)) and (layer2_outputs(1458)));
    layer3_outputs(1537) <= not((layer2_outputs(2032)) xor (layer2_outputs(771)));
    layer3_outputs(1538) <= (layer2_outputs(932)) or (layer2_outputs(2312));
    layer3_outputs(1539) <= not(layer2_outputs(1365));
    layer3_outputs(1540) <= (layer2_outputs(481)) and (layer2_outputs(2168));
    layer3_outputs(1541) <= not(layer2_outputs(1087)) or (layer2_outputs(574));
    layer3_outputs(1542) <= layer2_outputs(1424);
    layer3_outputs(1543) <= not(layer2_outputs(1990));
    layer3_outputs(1544) <= not(layer2_outputs(446)) or (layer2_outputs(515));
    layer3_outputs(1545) <= (layer2_outputs(1033)) and not (layer2_outputs(2375));
    layer3_outputs(1546) <= layer2_outputs(971);
    layer3_outputs(1547) <= (layer2_outputs(2452)) and (layer2_outputs(1821));
    layer3_outputs(1548) <= (layer2_outputs(917)) and (layer2_outputs(1817));
    layer3_outputs(1549) <= not(layer2_outputs(2087)) or (layer2_outputs(2350));
    layer3_outputs(1550) <= not((layer2_outputs(1239)) and (layer2_outputs(2279)));
    layer3_outputs(1551) <= layer2_outputs(1572);
    layer3_outputs(1552) <= not(layer2_outputs(568));
    layer3_outputs(1553) <= layer2_outputs(2259);
    layer3_outputs(1554) <= (layer2_outputs(2378)) and not (layer2_outputs(157));
    layer3_outputs(1555) <= not(layer2_outputs(1776));
    layer3_outputs(1556) <= not(layer2_outputs(667));
    layer3_outputs(1557) <= not((layer2_outputs(1700)) and (layer2_outputs(2044)));
    layer3_outputs(1558) <= not(layer2_outputs(149)) or (layer2_outputs(178));
    layer3_outputs(1559) <= layer2_outputs(396);
    layer3_outputs(1560) <= not((layer2_outputs(1353)) or (layer2_outputs(1417)));
    layer3_outputs(1561) <= layer2_outputs(2210);
    layer3_outputs(1562) <= (layer2_outputs(558)) and (layer2_outputs(1812));
    layer3_outputs(1563) <= layer2_outputs(1890);
    layer3_outputs(1564) <= (layer2_outputs(1603)) or (layer2_outputs(673));
    layer3_outputs(1565) <= layer2_outputs(1730);
    layer3_outputs(1566) <= not(layer2_outputs(1531)) or (layer2_outputs(1438));
    layer3_outputs(1567) <= (layer2_outputs(2535)) xor (layer2_outputs(1680));
    layer3_outputs(1568) <= layer2_outputs(1991);
    layer3_outputs(1569) <= (layer2_outputs(1848)) and not (layer2_outputs(1138));
    layer3_outputs(1570) <= not(layer2_outputs(524)) or (layer2_outputs(1146));
    layer3_outputs(1571) <= (layer2_outputs(1562)) xor (layer2_outputs(1222));
    layer3_outputs(1572) <= (layer2_outputs(1343)) and (layer2_outputs(1846));
    layer3_outputs(1573) <= (layer2_outputs(2044)) and not (layer2_outputs(2529));
    layer3_outputs(1574) <= not(layer2_outputs(241));
    layer3_outputs(1575) <= not(layer2_outputs(1161));
    layer3_outputs(1576) <= layer2_outputs(1838);
    layer3_outputs(1577) <= layer2_outputs(1582);
    layer3_outputs(1578) <= not((layer2_outputs(664)) xor (layer2_outputs(1391)));
    layer3_outputs(1579) <= '1';
    layer3_outputs(1580) <= not(layer2_outputs(1948)) or (layer2_outputs(540));
    layer3_outputs(1581) <= not(layer2_outputs(209)) or (layer2_outputs(961));
    layer3_outputs(1582) <= not(layer2_outputs(543));
    layer3_outputs(1583) <= layer2_outputs(2363);
    layer3_outputs(1584) <= not((layer2_outputs(439)) xor (layer2_outputs(1608)));
    layer3_outputs(1585) <= layer2_outputs(411);
    layer3_outputs(1586) <= layer2_outputs(1588);
    layer3_outputs(1587) <= not(layer2_outputs(459));
    layer3_outputs(1588) <= not(layer2_outputs(1705));
    layer3_outputs(1589) <= not(layer2_outputs(310));
    layer3_outputs(1590) <= not(layer2_outputs(2434));
    layer3_outputs(1591) <= not(layer2_outputs(1982));
    layer3_outputs(1592) <= layer2_outputs(1908);
    layer3_outputs(1593) <= not(layer2_outputs(532));
    layer3_outputs(1594) <= not((layer2_outputs(1639)) and (layer2_outputs(1506)));
    layer3_outputs(1595) <= not(layer2_outputs(251));
    layer3_outputs(1596) <= layer2_outputs(1169);
    layer3_outputs(1597) <= not(layer2_outputs(1321));
    layer3_outputs(1598) <= not((layer2_outputs(31)) xor (layer2_outputs(1401)));
    layer3_outputs(1599) <= not(layer2_outputs(403));
    layer3_outputs(1600) <= (layer2_outputs(2313)) and not (layer2_outputs(1367));
    layer3_outputs(1601) <= layer2_outputs(1813);
    layer3_outputs(1602) <= (layer2_outputs(187)) and (layer2_outputs(1604));
    layer3_outputs(1603) <= not(layer2_outputs(1673));
    layer3_outputs(1604) <= not(layer2_outputs(560));
    layer3_outputs(1605) <= layer2_outputs(244);
    layer3_outputs(1606) <= not((layer2_outputs(1622)) xor (layer2_outputs(994)));
    layer3_outputs(1607) <= (layer2_outputs(1900)) xor (layer2_outputs(2179));
    layer3_outputs(1608) <= layer2_outputs(1287);
    layer3_outputs(1609) <= not(layer2_outputs(624));
    layer3_outputs(1610) <= (layer2_outputs(2063)) and (layer2_outputs(50));
    layer3_outputs(1611) <= not(layer2_outputs(652)) or (layer2_outputs(2186));
    layer3_outputs(1612) <= layer2_outputs(1896);
    layer3_outputs(1613) <= layer2_outputs(1427);
    layer3_outputs(1614) <= not(layer2_outputs(1987));
    layer3_outputs(1615) <= (layer2_outputs(812)) and not (layer2_outputs(1387));
    layer3_outputs(1616) <= not((layer2_outputs(166)) or (layer2_outputs(643)));
    layer3_outputs(1617) <= (layer2_outputs(798)) and (layer2_outputs(1710));
    layer3_outputs(1618) <= not(layer2_outputs(1757)) or (layer2_outputs(1338));
    layer3_outputs(1619) <= layer2_outputs(175);
    layer3_outputs(1620) <= (layer2_outputs(188)) and (layer2_outputs(422));
    layer3_outputs(1621) <= (layer2_outputs(635)) and not (layer2_outputs(2026));
    layer3_outputs(1622) <= not((layer2_outputs(1185)) or (layer2_outputs(1447)));
    layer3_outputs(1623) <= not(layer2_outputs(1554)) or (layer2_outputs(2557));
    layer3_outputs(1624) <= not((layer2_outputs(1634)) or (layer2_outputs(2152)));
    layer3_outputs(1625) <= not(layer2_outputs(688));
    layer3_outputs(1626) <= not(layer2_outputs(2343)) or (layer2_outputs(1029));
    layer3_outputs(1627) <= not(layer2_outputs(1976));
    layer3_outputs(1628) <= (layer2_outputs(2412)) and not (layer2_outputs(2305));
    layer3_outputs(1629) <= '1';
    layer3_outputs(1630) <= not((layer2_outputs(551)) or (layer2_outputs(1505)));
    layer3_outputs(1631) <= not(layer2_outputs(1118));
    layer3_outputs(1632) <= layer2_outputs(1305);
    layer3_outputs(1633) <= layer2_outputs(2257);
    layer3_outputs(1634) <= not((layer2_outputs(1619)) and (layer2_outputs(1688)));
    layer3_outputs(1635) <= not(layer2_outputs(125));
    layer3_outputs(1636) <= not((layer2_outputs(1640)) and (layer2_outputs(213)));
    layer3_outputs(1637) <= layer2_outputs(1277);
    layer3_outputs(1638) <= layer2_outputs(1332);
    layer3_outputs(1639) <= layer2_outputs(640);
    layer3_outputs(1640) <= (layer2_outputs(336)) or (layer2_outputs(785));
    layer3_outputs(1641) <= layer2_outputs(239);
    layer3_outputs(1642) <= not(layer2_outputs(1384)) or (layer2_outputs(207));
    layer3_outputs(1643) <= layer2_outputs(122);
    layer3_outputs(1644) <= layer2_outputs(1774);
    layer3_outputs(1645) <= not(layer2_outputs(1865));
    layer3_outputs(1646) <= (layer2_outputs(1198)) or (layer2_outputs(1520));
    layer3_outputs(1647) <= (layer2_outputs(639)) or (layer2_outputs(1955));
    layer3_outputs(1648) <= layer2_outputs(583);
    layer3_outputs(1649) <= not(layer2_outputs(328)) or (layer2_outputs(1059));
    layer3_outputs(1650) <= layer2_outputs(50);
    layer3_outputs(1651) <= not(layer2_outputs(20));
    layer3_outputs(1652) <= '0';
    layer3_outputs(1653) <= '1';
    layer3_outputs(1654) <= not(layer2_outputs(2377));
    layer3_outputs(1655) <= '0';
    layer3_outputs(1656) <= (layer2_outputs(1918)) and not (layer2_outputs(2021));
    layer3_outputs(1657) <= layer2_outputs(2491);
    layer3_outputs(1658) <= (layer2_outputs(1559)) and not (layer2_outputs(830));
    layer3_outputs(1659) <= (layer2_outputs(1539)) or (layer2_outputs(2452));
    layer3_outputs(1660) <= not((layer2_outputs(2431)) and (layer2_outputs(2012)));
    layer3_outputs(1661) <= layer2_outputs(926);
    layer3_outputs(1662) <= not(layer2_outputs(1975));
    layer3_outputs(1663) <= not(layer2_outputs(2507));
    layer3_outputs(1664) <= not((layer2_outputs(2237)) xor (layer2_outputs(2064)));
    layer3_outputs(1665) <= not((layer2_outputs(1070)) or (layer2_outputs(634)));
    layer3_outputs(1666) <= not(layer2_outputs(2268));
    layer3_outputs(1667) <= layer2_outputs(414);
    layer3_outputs(1668) <= layer2_outputs(803);
    layer3_outputs(1669) <= (layer2_outputs(306)) and not (layer2_outputs(300));
    layer3_outputs(1670) <= '1';
    layer3_outputs(1671) <= not(layer2_outputs(1642));
    layer3_outputs(1672) <= (layer2_outputs(1301)) xor (layer2_outputs(177));
    layer3_outputs(1673) <= layer2_outputs(1782);
    layer3_outputs(1674) <= (layer2_outputs(1497)) and not (layer2_outputs(1360));
    layer3_outputs(1675) <= not((layer2_outputs(487)) and (layer2_outputs(1496)));
    layer3_outputs(1676) <= (layer2_outputs(1283)) and not (layer2_outputs(385));
    layer3_outputs(1677) <= (layer2_outputs(722)) and not (layer2_outputs(1144));
    layer3_outputs(1678) <= not(layer2_outputs(2128));
    layer3_outputs(1679) <= layer2_outputs(577);
    layer3_outputs(1680) <= not((layer2_outputs(1265)) and (layer2_outputs(1648)));
    layer3_outputs(1681) <= (layer2_outputs(727)) xor (layer2_outputs(130));
    layer3_outputs(1682) <= (layer2_outputs(382)) and (layer2_outputs(2538));
    layer3_outputs(1683) <= (layer2_outputs(1211)) or (layer2_outputs(71));
    layer3_outputs(1684) <= not(layer2_outputs(1907));
    layer3_outputs(1685) <= layer2_outputs(1786);
    layer3_outputs(1686) <= not((layer2_outputs(1421)) and (layer2_outputs(2045)));
    layer3_outputs(1687) <= (layer2_outputs(1344)) or (layer2_outputs(951));
    layer3_outputs(1688) <= (layer2_outputs(276)) and not (layer2_outputs(1656));
    layer3_outputs(1689) <= not((layer2_outputs(2002)) xor (layer2_outputs(1860)));
    layer3_outputs(1690) <= not(layer2_outputs(214));
    layer3_outputs(1691) <= not((layer2_outputs(600)) or (layer2_outputs(1567)));
    layer3_outputs(1692) <= not(layer2_outputs(87)) or (layer2_outputs(1571));
    layer3_outputs(1693) <= not(layer2_outputs(308)) or (layer2_outputs(184));
    layer3_outputs(1694) <= layer2_outputs(2006);
    layer3_outputs(1695) <= not(layer2_outputs(1988));
    layer3_outputs(1696) <= not((layer2_outputs(1410)) and (layer2_outputs(1645)));
    layer3_outputs(1697) <= not((layer2_outputs(270)) or (layer2_outputs(1235)));
    layer3_outputs(1698) <= not(layer2_outputs(2016));
    layer3_outputs(1699) <= not(layer2_outputs(2254));
    layer3_outputs(1700) <= layer2_outputs(1442);
    layer3_outputs(1701) <= (layer2_outputs(853)) and (layer2_outputs(1792));
    layer3_outputs(1702) <= not(layer2_outputs(2332));
    layer3_outputs(1703) <= layer2_outputs(845);
    layer3_outputs(1704) <= layer2_outputs(1225);
    layer3_outputs(1705) <= layer2_outputs(1527);
    layer3_outputs(1706) <= not((layer2_outputs(970)) and (layer2_outputs(1974)));
    layer3_outputs(1707) <= not(layer2_outputs(151));
    layer3_outputs(1708) <= not(layer2_outputs(2483));
    layer3_outputs(1709) <= not((layer2_outputs(1991)) and (layer2_outputs(752)));
    layer3_outputs(1710) <= (layer2_outputs(747)) and (layer2_outputs(1404));
    layer3_outputs(1711) <= (layer2_outputs(2251)) and (layer2_outputs(759));
    layer3_outputs(1712) <= not((layer2_outputs(1380)) and (layer2_outputs(2498)));
    layer3_outputs(1713) <= layer2_outputs(2543);
    layer3_outputs(1714) <= not((layer2_outputs(2070)) xor (layer2_outputs(1665)));
    layer3_outputs(1715) <= not(layer2_outputs(1598));
    layer3_outputs(1716) <= not(layer2_outputs(1594));
    layer3_outputs(1717) <= not(layer2_outputs(388));
    layer3_outputs(1718) <= not(layer2_outputs(259));
    layer3_outputs(1719) <= not(layer2_outputs(2072));
    layer3_outputs(1720) <= (layer2_outputs(407)) or (layer2_outputs(1173));
    layer3_outputs(1721) <= layer2_outputs(1731);
    layer3_outputs(1722) <= not(layer2_outputs(1830));
    layer3_outputs(1723) <= (layer2_outputs(1144)) or (layer2_outputs(961));
    layer3_outputs(1724) <= (layer2_outputs(2207)) or (layer2_outputs(2186));
    layer3_outputs(1725) <= (layer2_outputs(2062)) or (layer2_outputs(166));
    layer3_outputs(1726) <= layer2_outputs(1594);
    layer3_outputs(1727) <= not(layer2_outputs(363));
    layer3_outputs(1728) <= layer2_outputs(2545);
    layer3_outputs(1729) <= '0';
    layer3_outputs(1730) <= layer2_outputs(1140);
    layer3_outputs(1731) <= not(layer2_outputs(1237));
    layer3_outputs(1732) <= layer2_outputs(1476);
    layer3_outputs(1733) <= not(layer2_outputs(1105));
    layer3_outputs(1734) <= (layer2_outputs(1741)) xor (layer2_outputs(787));
    layer3_outputs(1735) <= layer2_outputs(2101);
    layer3_outputs(1736) <= not(layer2_outputs(2293));
    layer3_outputs(1737) <= (layer2_outputs(1176)) xor (layer2_outputs(1542));
    layer3_outputs(1738) <= '1';
    layer3_outputs(1739) <= not(layer2_outputs(113));
    layer3_outputs(1740) <= not(layer2_outputs(30));
    layer3_outputs(1741) <= not((layer2_outputs(131)) and (layer2_outputs(1790)));
    layer3_outputs(1742) <= (layer2_outputs(2503)) and not (layer2_outputs(901));
    layer3_outputs(1743) <= (layer2_outputs(198)) and (layer2_outputs(1087));
    layer3_outputs(1744) <= not((layer2_outputs(2481)) and (layer2_outputs(1021)));
    layer3_outputs(1745) <= not(layer2_outputs(1943));
    layer3_outputs(1746) <= (layer2_outputs(1616)) and (layer2_outputs(482));
    layer3_outputs(1747) <= (layer2_outputs(859)) and not (layer2_outputs(2289));
    layer3_outputs(1748) <= layer2_outputs(863);
    layer3_outputs(1749) <= (layer2_outputs(1572)) and (layer2_outputs(330));
    layer3_outputs(1750) <= not(layer2_outputs(741));
    layer3_outputs(1751) <= layer2_outputs(1152);
    layer3_outputs(1752) <= layer2_outputs(12);
    layer3_outputs(1753) <= not((layer2_outputs(1448)) and (layer2_outputs(2234)));
    layer3_outputs(1754) <= (layer2_outputs(141)) and not (layer2_outputs(832));
    layer3_outputs(1755) <= not((layer2_outputs(2138)) or (layer2_outputs(1528)));
    layer3_outputs(1756) <= (layer2_outputs(1575)) and (layer2_outputs(447));
    layer3_outputs(1757) <= not(layer2_outputs(938)) or (layer2_outputs(1682));
    layer3_outputs(1758) <= (layer2_outputs(910)) or (layer2_outputs(2529));
    layer3_outputs(1759) <= (layer2_outputs(672)) and (layer2_outputs(219));
    layer3_outputs(1760) <= layer2_outputs(733);
    layer3_outputs(1761) <= not(layer2_outputs(795));
    layer3_outputs(1762) <= not((layer2_outputs(1395)) or (layer2_outputs(167)));
    layer3_outputs(1763) <= not(layer2_outputs(1818)) or (layer2_outputs(415));
    layer3_outputs(1764) <= not(layer2_outputs(44));
    layer3_outputs(1765) <= layer2_outputs(2176);
    layer3_outputs(1766) <= (layer2_outputs(925)) and (layer2_outputs(39));
    layer3_outputs(1767) <= not(layer2_outputs(790));
    layer3_outputs(1768) <= '0';
    layer3_outputs(1769) <= (layer2_outputs(1931)) and not (layer2_outputs(1505));
    layer3_outputs(1770) <= '0';
    layer3_outputs(1771) <= not(layer2_outputs(25));
    layer3_outputs(1772) <= not(layer2_outputs(1027)) or (layer2_outputs(1328));
    layer3_outputs(1773) <= (layer2_outputs(2308)) or (layer2_outputs(703));
    layer3_outputs(1774) <= not((layer2_outputs(936)) or (layer2_outputs(86)));
    layer3_outputs(1775) <= not(layer2_outputs(1762));
    layer3_outputs(1776) <= layer2_outputs(2456);
    layer3_outputs(1777) <= layer2_outputs(2287);
    layer3_outputs(1778) <= not(layer2_outputs(2225)) or (layer2_outputs(487));
    layer3_outputs(1779) <= layer2_outputs(1692);
    layer3_outputs(1780) <= (layer2_outputs(2456)) and not (layer2_outputs(1167));
    layer3_outputs(1781) <= (layer2_outputs(1725)) or (layer2_outputs(2489));
    layer3_outputs(1782) <= not(layer2_outputs(1154)) or (layer2_outputs(2285));
    layer3_outputs(1783) <= layer2_outputs(1454);
    layer3_outputs(1784) <= not((layer2_outputs(751)) and (layer2_outputs(1852)));
    layer3_outputs(1785) <= layer2_outputs(1658);
    layer3_outputs(1786) <= layer2_outputs(181);
    layer3_outputs(1787) <= (layer2_outputs(201)) or (layer2_outputs(2499));
    layer3_outputs(1788) <= not(layer2_outputs(1198)) or (layer2_outputs(1927));
    layer3_outputs(1789) <= not(layer2_outputs(248));
    layer3_outputs(1790) <= layer2_outputs(633);
    layer3_outputs(1791) <= not(layer2_outputs(1020));
    layer3_outputs(1792) <= not(layer2_outputs(1297));
    layer3_outputs(1793) <= (layer2_outputs(2479)) and not (layer2_outputs(1994));
    layer3_outputs(1794) <= not(layer2_outputs(581));
    layer3_outputs(1795) <= not(layer2_outputs(149));
    layer3_outputs(1796) <= not((layer2_outputs(377)) xor (layer2_outputs(285)));
    layer3_outputs(1797) <= (layer2_outputs(579)) and not (layer2_outputs(2322));
    layer3_outputs(1798) <= not(layer2_outputs(160));
    layer3_outputs(1799) <= (layer2_outputs(2420)) and not (layer2_outputs(1329));
    layer3_outputs(1800) <= (layer2_outputs(190)) and not (layer2_outputs(854));
    layer3_outputs(1801) <= not(layer2_outputs(1434)) or (layer2_outputs(2193));
    layer3_outputs(1802) <= layer2_outputs(1011);
    layer3_outputs(1803) <= (layer2_outputs(238)) and not (layer2_outputs(1180));
    layer3_outputs(1804) <= layer2_outputs(87);
    layer3_outputs(1805) <= not(layer2_outputs(743));
    layer3_outputs(1806) <= not(layer2_outputs(1899));
    layer3_outputs(1807) <= (layer2_outputs(1158)) and not (layer2_outputs(620));
    layer3_outputs(1808) <= not(layer2_outputs(564));
    layer3_outputs(1809) <= not((layer2_outputs(1366)) or (layer2_outputs(608)));
    layer3_outputs(1810) <= not((layer2_outputs(1373)) or (layer2_outputs(83)));
    layer3_outputs(1811) <= not(layer2_outputs(1617));
    layer3_outputs(1812) <= not((layer2_outputs(13)) or (layer2_outputs(914)));
    layer3_outputs(1813) <= not((layer2_outputs(782)) and (layer2_outputs(927)));
    layer3_outputs(1814) <= not(layer2_outputs(1978)) or (layer2_outputs(1641));
    layer3_outputs(1815) <= not((layer2_outputs(2135)) or (layer2_outputs(2059)));
    layer3_outputs(1816) <= not((layer2_outputs(551)) or (layer2_outputs(321)));
    layer3_outputs(1817) <= (layer2_outputs(1113)) and not (layer2_outputs(973));
    layer3_outputs(1818) <= layer2_outputs(1535);
    layer3_outputs(1819) <= not(layer2_outputs(1840));
    layer3_outputs(1820) <= (layer2_outputs(1716)) or (layer2_outputs(1012));
    layer3_outputs(1821) <= not(layer2_outputs(77));
    layer3_outputs(1822) <= not(layer2_outputs(2037)) or (layer2_outputs(2369));
    layer3_outputs(1823) <= layer2_outputs(77);
    layer3_outputs(1824) <= not(layer2_outputs(132)) or (layer2_outputs(2313));
    layer3_outputs(1825) <= layer2_outputs(2009);
    layer3_outputs(1826) <= '1';
    layer3_outputs(1827) <= not(layer2_outputs(1591)) or (layer2_outputs(237));
    layer3_outputs(1828) <= not(layer2_outputs(962));
    layer3_outputs(1829) <= layer2_outputs(111);
    layer3_outputs(1830) <= not(layer2_outputs(1478)) or (layer2_outputs(953));
    layer3_outputs(1831) <= not(layer2_outputs(2443)) or (layer2_outputs(2183));
    layer3_outputs(1832) <= not((layer2_outputs(272)) or (layer2_outputs(1402)));
    layer3_outputs(1833) <= (layer2_outputs(661)) and not (layer2_outputs(1040));
    layer3_outputs(1834) <= not(layer2_outputs(1679)) or (layer2_outputs(1834));
    layer3_outputs(1835) <= layer2_outputs(1206);
    layer3_outputs(1836) <= layer2_outputs(1977);
    layer3_outputs(1837) <= layer2_outputs(1009);
    layer3_outputs(1838) <= (layer2_outputs(882)) and not (layer2_outputs(2247));
    layer3_outputs(1839) <= not(layer2_outputs(2433)) or (layer2_outputs(1629));
    layer3_outputs(1840) <= not(layer2_outputs(347));
    layer3_outputs(1841) <= (layer2_outputs(342)) or (layer2_outputs(2054));
    layer3_outputs(1842) <= (layer2_outputs(1912)) and (layer2_outputs(1926));
    layer3_outputs(1843) <= '0';
    layer3_outputs(1844) <= '1';
    layer3_outputs(1845) <= not((layer2_outputs(563)) and (layer2_outputs(590)));
    layer3_outputs(1846) <= layer2_outputs(1723);
    layer3_outputs(1847) <= (layer2_outputs(875)) and (layer2_outputs(770));
    layer3_outputs(1848) <= (layer2_outputs(663)) xor (layer2_outputs(2351));
    layer3_outputs(1849) <= not(layer2_outputs(1905));
    layer3_outputs(1850) <= (layer2_outputs(2427)) or (layer2_outputs(2185));
    layer3_outputs(1851) <= not(layer2_outputs(295)) or (layer2_outputs(2515));
    layer3_outputs(1852) <= not(layer2_outputs(91)) or (layer2_outputs(2416));
    layer3_outputs(1853) <= layer2_outputs(2090);
    layer3_outputs(1854) <= (layer2_outputs(811)) xor (layer2_outputs(2125));
    layer3_outputs(1855) <= not(layer2_outputs(619));
    layer3_outputs(1856) <= '0';
    layer3_outputs(1857) <= not(layer2_outputs(1518));
    layer3_outputs(1858) <= (layer2_outputs(1008)) or (layer2_outputs(1244));
    layer3_outputs(1859) <= not((layer2_outputs(819)) or (layer2_outputs(1252)));
    layer3_outputs(1860) <= layer2_outputs(591);
    layer3_outputs(1861) <= not(layer2_outputs(610)) or (layer2_outputs(1815));
    layer3_outputs(1862) <= '0';
    layer3_outputs(1863) <= not(layer2_outputs(640)) or (layer2_outputs(167));
    layer3_outputs(1864) <= layer2_outputs(2507);
    layer3_outputs(1865) <= layer2_outputs(818);
    layer3_outputs(1866) <= (layer2_outputs(98)) and not (layer2_outputs(1316));
    layer3_outputs(1867) <= '1';
    layer3_outputs(1868) <= not((layer2_outputs(7)) or (layer2_outputs(1961)));
    layer3_outputs(1869) <= not(layer2_outputs(1773));
    layer3_outputs(1870) <= '1';
    layer3_outputs(1871) <= not((layer2_outputs(1433)) and (layer2_outputs(324)));
    layer3_outputs(1872) <= not(layer2_outputs(1952));
    layer3_outputs(1873) <= layer2_outputs(108);
    layer3_outputs(1874) <= (layer2_outputs(1738)) and not (layer2_outputs(2304));
    layer3_outputs(1875) <= not((layer2_outputs(1740)) and (layer2_outputs(1750)));
    layer3_outputs(1876) <= not(layer2_outputs(2002));
    layer3_outputs(1877) <= layer2_outputs(1985);
    layer3_outputs(1878) <= '0';
    layer3_outputs(1879) <= (layer2_outputs(959)) or (layer2_outputs(1709));
    layer3_outputs(1880) <= layer2_outputs(741);
    layer3_outputs(1881) <= not(layer2_outputs(1172));
    layer3_outputs(1882) <= layer2_outputs(1982);
    layer3_outputs(1883) <= not(layer2_outputs(1315)) or (layer2_outputs(2386));
    layer3_outputs(1884) <= (layer2_outputs(224)) and (layer2_outputs(395));
    layer3_outputs(1885) <= layer2_outputs(1698);
    layer3_outputs(1886) <= layer2_outputs(1052);
    layer3_outputs(1887) <= not(layer2_outputs(1170));
    layer3_outputs(1888) <= (layer2_outputs(1208)) and not (layer2_outputs(1782));
    layer3_outputs(1889) <= not(layer2_outputs(1545)) or (layer2_outputs(2190));
    layer3_outputs(1890) <= (layer2_outputs(1247)) or (layer2_outputs(856));
    layer3_outputs(1891) <= '1';
    layer3_outputs(1892) <= not(layer2_outputs(513)) or (layer2_outputs(1985));
    layer3_outputs(1893) <= layer2_outputs(1779);
    layer3_outputs(1894) <= (layer2_outputs(664)) and (layer2_outputs(1056));
    layer3_outputs(1895) <= layer2_outputs(1672);
    layer3_outputs(1896) <= not(layer2_outputs(870)) or (layer2_outputs(1222));
    layer3_outputs(1897) <= not(layer2_outputs(455)) or (layer2_outputs(1429));
    layer3_outputs(1898) <= not(layer2_outputs(2455));
    layer3_outputs(1899) <= layer2_outputs(1018);
    layer3_outputs(1900) <= '1';
    layer3_outputs(1901) <= (layer2_outputs(2144)) or (layer2_outputs(168));
    layer3_outputs(1902) <= not(layer2_outputs(1016)) or (layer2_outputs(1254));
    layer3_outputs(1903) <= (layer2_outputs(868)) and not (layer2_outputs(138));
    layer3_outputs(1904) <= (layer2_outputs(2200)) and not (layer2_outputs(711));
    layer3_outputs(1905) <= layer2_outputs(1231);
    layer3_outputs(1906) <= (layer2_outputs(2197)) and not (layer2_outputs(2300));
    layer3_outputs(1907) <= layer2_outputs(2271);
    layer3_outputs(1908) <= '1';
    layer3_outputs(1909) <= (layer2_outputs(751)) or (layer2_outputs(346));
    layer3_outputs(1910) <= (layer2_outputs(208)) and (layer2_outputs(2094));
    layer3_outputs(1911) <= not(layer2_outputs(115));
    layer3_outputs(1912) <= '1';
    layer3_outputs(1913) <= not(layer2_outputs(1352));
    layer3_outputs(1914) <= '1';
    layer3_outputs(1915) <= not(layer2_outputs(1161));
    layer3_outputs(1916) <= (layer2_outputs(1805)) xor (layer2_outputs(1679));
    layer3_outputs(1917) <= not(layer2_outputs(1987));
    layer3_outputs(1918) <= not(layer2_outputs(12));
    layer3_outputs(1919) <= not(layer2_outputs(1838));
    layer3_outputs(1920) <= (layer2_outputs(117)) and (layer2_outputs(69));
    layer3_outputs(1921) <= layer2_outputs(1286);
    layer3_outputs(1922) <= (layer2_outputs(1172)) and (layer2_outputs(1511));
    layer3_outputs(1923) <= (layer2_outputs(246)) and not (layer2_outputs(444));
    layer3_outputs(1924) <= not(layer2_outputs(1550));
    layer3_outputs(1925) <= (layer2_outputs(186)) and not (layer2_outputs(2141));
    layer3_outputs(1926) <= (layer2_outputs(2438)) or (layer2_outputs(2102));
    layer3_outputs(1927) <= (layer2_outputs(326)) xor (layer2_outputs(1207));
    layer3_outputs(1928) <= layer2_outputs(507);
    layer3_outputs(1929) <= (layer2_outputs(705)) and not (layer2_outputs(1808));
    layer3_outputs(1930) <= '1';
    layer3_outputs(1931) <= '1';
    layer3_outputs(1932) <= not(layer2_outputs(2019));
    layer3_outputs(1933) <= not(layer2_outputs(575)) or (layer2_outputs(1946));
    layer3_outputs(1934) <= (layer2_outputs(1411)) and not (layer2_outputs(1212));
    layer3_outputs(1935) <= not(layer2_outputs(1460));
    layer3_outputs(1936) <= layer2_outputs(1501);
    layer3_outputs(1937) <= not(layer2_outputs(81));
    layer3_outputs(1938) <= not((layer2_outputs(2087)) or (layer2_outputs(121)));
    layer3_outputs(1939) <= layer2_outputs(1444);
    layer3_outputs(1940) <= not(layer2_outputs(512));
    layer3_outputs(1941) <= (layer2_outputs(1409)) or (layer2_outputs(94));
    layer3_outputs(1942) <= not(layer2_outputs(362));
    layer3_outputs(1943) <= (layer2_outputs(1548)) and not (layer2_outputs(1093));
    layer3_outputs(1944) <= (layer2_outputs(85)) and (layer2_outputs(464));
    layer3_outputs(1945) <= layer2_outputs(987);
    layer3_outputs(1946) <= not((layer2_outputs(832)) or (layer2_outputs(2538)));
    layer3_outputs(1947) <= not((layer2_outputs(2355)) xor (layer2_outputs(528)));
    layer3_outputs(1948) <= (layer2_outputs(1151)) or (layer2_outputs(1504));
    layer3_outputs(1949) <= not((layer2_outputs(2224)) and (layer2_outputs(662)));
    layer3_outputs(1950) <= not((layer2_outputs(1020)) and (layer2_outputs(2231)));
    layer3_outputs(1951) <= not(layer2_outputs(2534)) or (layer2_outputs(1047));
    layer3_outputs(1952) <= (layer2_outputs(2014)) and not (layer2_outputs(90));
    layer3_outputs(1953) <= not(layer2_outputs(693));
    layer3_outputs(1954) <= not((layer2_outputs(677)) and (layer2_outputs(613)));
    layer3_outputs(1955) <= not(layer2_outputs(1944));
    layer3_outputs(1956) <= not(layer2_outputs(1736));
    layer3_outputs(1957) <= (layer2_outputs(2340)) or (layer2_outputs(2276));
    layer3_outputs(1958) <= not(layer2_outputs(1800)) or (layer2_outputs(2142));
    layer3_outputs(1959) <= not(layer2_outputs(1629)) or (layer2_outputs(521));
    layer3_outputs(1960) <= not(layer2_outputs(2448)) or (layer2_outputs(601));
    layer3_outputs(1961) <= not(layer2_outputs(2062));
    layer3_outputs(1962) <= not((layer2_outputs(2250)) or (layer2_outputs(784)));
    layer3_outputs(1963) <= layer2_outputs(1747);
    layer3_outputs(1964) <= not(layer2_outputs(2348));
    layer3_outputs(1965) <= '0';
    layer3_outputs(1966) <= not(layer2_outputs(42));
    layer3_outputs(1967) <= layer2_outputs(1149);
    layer3_outputs(1968) <= not((layer2_outputs(1311)) or (layer2_outputs(1270)));
    layer3_outputs(1969) <= not(layer2_outputs(992));
    layer3_outputs(1970) <= layer2_outputs(314);
    layer3_outputs(1971) <= not(layer2_outputs(1569));
    layer3_outputs(1972) <= layer2_outputs(1446);
    layer3_outputs(1973) <= layer2_outputs(58);
    layer3_outputs(1974) <= not(layer2_outputs(806)) or (layer2_outputs(1113));
    layer3_outputs(1975) <= not(layer2_outputs(2393));
    layer3_outputs(1976) <= not((layer2_outputs(139)) or (layer2_outputs(2205)));
    layer3_outputs(1977) <= layer2_outputs(1922);
    layer3_outputs(1978) <= layer2_outputs(1076);
    layer3_outputs(1979) <= not(layer2_outputs(1422));
    layer3_outputs(1980) <= (layer2_outputs(1044)) and (layer2_outputs(1074));
    layer3_outputs(1981) <= layer2_outputs(610);
    layer3_outputs(1982) <= layer2_outputs(2414);
    layer3_outputs(1983) <= not(layer2_outputs(623)) or (layer2_outputs(1327));
    layer3_outputs(1984) <= layer2_outputs(1699);
    layer3_outputs(1985) <= not(layer2_outputs(846));
    layer3_outputs(1986) <= '0';
    layer3_outputs(1987) <= not((layer2_outputs(2270)) xor (layer2_outputs(495)));
    layer3_outputs(1988) <= (layer2_outputs(2188)) or (layer2_outputs(1481));
    layer3_outputs(1989) <= not(layer2_outputs(362));
    layer3_outputs(1990) <= (layer2_outputs(1849)) and not (layer2_outputs(1404));
    layer3_outputs(1991) <= '0';
    layer3_outputs(1992) <= '0';
    layer3_outputs(1993) <= not((layer2_outputs(2226)) or (layer2_outputs(1219)));
    layer3_outputs(1994) <= not(layer2_outputs(1168));
    layer3_outputs(1995) <= '0';
    layer3_outputs(1996) <= not((layer2_outputs(1081)) and (layer2_outputs(499)));
    layer3_outputs(1997) <= (layer2_outputs(179)) and (layer2_outputs(1322));
    layer3_outputs(1998) <= layer2_outputs(1690);
    layer3_outputs(1999) <= layer2_outputs(246);
    layer3_outputs(2000) <= (layer2_outputs(164)) and not (layer2_outputs(1359));
    layer3_outputs(2001) <= not(layer2_outputs(1625));
    layer3_outputs(2002) <= not(layer2_outputs(174)) or (layer2_outputs(828));
    layer3_outputs(2003) <= not(layer2_outputs(361));
    layer3_outputs(2004) <= (layer2_outputs(1558)) and not (layer2_outputs(924));
    layer3_outputs(2005) <= not(layer2_outputs(697));
    layer3_outputs(2006) <= not(layer2_outputs(1038)) or (layer2_outputs(767));
    layer3_outputs(2007) <= not(layer2_outputs(2405));
    layer3_outputs(2008) <= not(layer2_outputs(1211)) or (layer2_outputs(2212));
    layer3_outputs(2009) <= not(layer2_outputs(171));
    layer3_outputs(2010) <= not((layer2_outputs(1453)) xor (layer2_outputs(33)));
    layer3_outputs(2011) <= not((layer2_outputs(2023)) or (layer2_outputs(734)));
    layer3_outputs(2012) <= not(layer2_outputs(1371));
    layer3_outputs(2013) <= layer2_outputs(826);
    layer3_outputs(2014) <= (layer2_outputs(2379)) and (layer2_outputs(914));
    layer3_outputs(2015) <= layer2_outputs(1625);
    layer3_outputs(2016) <= (layer2_outputs(1004)) and (layer2_outputs(2516));
    layer3_outputs(2017) <= layer2_outputs(182);
    layer3_outputs(2018) <= (layer2_outputs(2558)) or (layer2_outputs(1383));
    layer3_outputs(2019) <= not(layer2_outputs(2528));
    layer3_outputs(2020) <= (layer2_outputs(469)) and (layer2_outputs(2487));
    layer3_outputs(2021) <= layer2_outputs(816);
    layer3_outputs(2022) <= '1';
    layer3_outputs(2023) <= layer2_outputs(1832);
    layer3_outputs(2024) <= layer2_outputs(1867);
    layer3_outputs(2025) <= (layer2_outputs(1120)) or (layer2_outputs(2484));
    layer3_outputs(2026) <= not(layer2_outputs(1449));
    layer3_outputs(2027) <= not(layer2_outputs(2137));
    layer3_outputs(2028) <= not(layer2_outputs(239)) or (layer2_outputs(2149));
    layer3_outputs(2029) <= not(layer2_outputs(302)) or (layer2_outputs(232));
    layer3_outputs(2030) <= not(layer2_outputs(248)) or (layer2_outputs(1567));
    layer3_outputs(2031) <= (layer2_outputs(143)) and not (layer2_outputs(1887));
    layer3_outputs(2032) <= not(layer2_outputs(1499));
    layer3_outputs(2033) <= layer2_outputs(905);
    layer3_outputs(2034) <= not(layer2_outputs(1664));
    layer3_outputs(2035) <= not((layer2_outputs(899)) or (layer2_outputs(2211)));
    layer3_outputs(2036) <= (layer2_outputs(775)) or (layer2_outputs(828));
    layer3_outputs(2037) <= not((layer2_outputs(1653)) and (layer2_outputs(818)));
    layer3_outputs(2038) <= not(layer2_outputs(855));
    layer3_outputs(2039) <= not((layer2_outputs(2080)) or (layer2_outputs(1837)));
    layer3_outputs(2040) <= (layer2_outputs(1773)) or (layer2_outputs(2364));
    layer3_outputs(2041) <= '0';
    layer3_outputs(2042) <= (layer2_outputs(895)) and not (layer2_outputs(2408));
    layer3_outputs(2043) <= not(layer2_outputs(1986)) or (layer2_outputs(183));
    layer3_outputs(2044) <= not((layer2_outputs(569)) or (layer2_outputs(1876)));
    layer3_outputs(2045) <= '1';
    layer3_outputs(2046) <= '0';
    layer3_outputs(2047) <= not(layer2_outputs(972));
    layer3_outputs(2048) <= (layer2_outputs(725)) and not (layer2_outputs(968));
    layer3_outputs(2049) <= layer2_outputs(789);
    layer3_outputs(2050) <= not(layer2_outputs(147)) or (layer2_outputs(618));
    layer3_outputs(2051) <= not(layer2_outputs(311));
    layer3_outputs(2052) <= layer2_outputs(2359);
    layer3_outputs(2053) <= (layer2_outputs(332)) and not (layer2_outputs(1999));
    layer3_outputs(2054) <= (layer2_outputs(1801)) or (layer2_outputs(19));
    layer3_outputs(2055) <= (layer2_outputs(2100)) xor (layer2_outputs(2085));
    layer3_outputs(2056) <= (layer2_outputs(2533)) and not (layer2_outputs(484));
    layer3_outputs(2057) <= layer2_outputs(2162);
    layer3_outputs(2058) <= not(layer2_outputs(955)) or (layer2_outputs(1035));
    layer3_outputs(2059) <= layer2_outputs(1563);
    layer3_outputs(2060) <= not((layer2_outputs(396)) or (layer2_outputs(788)));
    layer3_outputs(2061) <= (layer2_outputs(736)) or (layer2_outputs(2329));
    layer3_outputs(2062) <= layer2_outputs(1429);
    layer3_outputs(2063) <= not(layer2_outputs(2052));
    layer3_outputs(2064) <= not(layer2_outputs(264)) or (layer2_outputs(421));
    layer3_outputs(2065) <= layer2_outputs(360);
    layer3_outputs(2066) <= layer2_outputs(2265);
    layer3_outputs(2067) <= not((layer2_outputs(922)) or (layer2_outputs(1775)));
    layer3_outputs(2068) <= layer2_outputs(1481);
    layer3_outputs(2069) <= (layer2_outputs(582)) and not (layer2_outputs(930));
    layer3_outputs(2070) <= (layer2_outputs(2535)) xor (layer2_outputs(402));
    layer3_outputs(2071) <= not((layer2_outputs(940)) and (layer2_outputs(1680)));
    layer3_outputs(2072) <= layer2_outputs(667);
    layer3_outputs(2073) <= not(layer2_outputs(2327));
    layer3_outputs(2074) <= layer2_outputs(1433);
    layer3_outputs(2075) <= '1';
    layer3_outputs(2076) <= not(layer2_outputs(304)) or (layer2_outputs(1260));
    layer3_outputs(2077) <= not(layer2_outputs(2264));
    layer3_outputs(2078) <= layer2_outputs(1984);
    layer3_outputs(2079) <= (layer2_outputs(1823)) and (layer2_outputs(1969));
    layer3_outputs(2080) <= not(layer2_outputs(592));
    layer3_outputs(2081) <= not(layer2_outputs(1362));
    layer3_outputs(2082) <= not((layer2_outputs(116)) or (layer2_outputs(694)));
    layer3_outputs(2083) <= not(layer2_outputs(597));
    layer3_outputs(2084) <= not((layer2_outputs(867)) xor (layer2_outputs(854)));
    layer3_outputs(2085) <= '1';
    layer3_outputs(2086) <= not(layer2_outputs(1399));
    layer3_outputs(2087) <= layer2_outputs(1966);
    layer3_outputs(2088) <= layer2_outputs(715);
    layer3_outputs(2089) <= (layer2_outputs(1295)) and (layer2_outputs(1498));
    layer3_outputs(2090) <= not(layer2_outputs(1237)) or (layer2_outputs(1878));
    layer3_outputs(2091) <= not(layer2_outputs(2426));
    layer3_outputs(2092) <= layer2_outputs(549);
    layer3_outputs(2093) <= not((layer2_outputs(1570)) and (layer2_outputs(1031)));
    layer3_outputs(2094) <= not((layer2_outputs(142)) or (layer2_outputs(898)));
    layer3_outputs(2095) <= not(layer2_outputs(1628));
    layer3_outputs(2096) <= not(layer2_outputs(2476)) or (layer2_outputs(2166));
    layer3_outputs(2097) <= layer2_outputs(1009);
    layer3_outputs(2098) <= layer2_outputs(1327);
    layer3_outputs(2099) <= not((layer2_outputs(876)) or (layer2_outputs(1711)));
    layer3_outputs(2100) <= layer2_outputs(86);
    layer3_outputs(2101) <= (layer2_outputs(1001)) or (layer2_outputs(23));
    layer3_outputs(2102) <= (layer2_outputs(1640)) and (layer2_outputs(2069));
    layer3_outputs(2103) <= (layer2_outputs(1750)) and not (layer2_outputs(2309));
    layer3_outputs(2104) <= not(layer2_outputs(724)) or (layer2_outputs(191));
    layer3_outputs(2105) <= not(layer2_outputs(1355));
    layer3_outputs(2106) <= (layer2_outputs(412)) and not (layer2_outputs(707));
    layer3_outputs(2107) <= not(layer2_outputs(827));
    layer3_outputs(2108) <= not(layer2_outputs(2078));
    layer3_outputs(2109) <= layer2_outputs(2486);
    layer3_outputs(2110) <= not(layer2_outputs(346));
    layer3_outputs(2111) <= (layer2_outputs(1645)) or (layer2_outputs(680));
    layer3_outputs(2112) <= not(layer2_outputs(1296));
    layer3_outputs(2113) <= not(layer2_outputs(2525)) or (layer2_outputs(1822));
    layer3_outputs(2114) <= not(layer2_outputs(2310));
    layer3_outputs(2115) <= layer2_outputs(1157);
    layer3_outputs(2116) <= layer2_outputs(1658);
    layer3_outputs(2117) <= not(layer2_outputs(1016));
    layer3_outputs(2118) <= not((layer2_outputs(539)) and (layer2_outputs(2394)));
    layer3_outputs(2119) <= not(layer2_outputs(1060));
    layer3_outputs(2120) <= layer2_outputs(10);
    layer3_outputs(2121) <= (layer2_outputs(1186)) and not (layer2_outputs(2466));
    layer3_outputs(2122) <= not(layer2_outputs(290));
    layer3_outputs(2123) <= not(layer2_outputs(217));
    layer3_outputs(2124) <= not(layer2_outputs(100)) or (layer2_outputs(1461));
    layer3_outputs(2125) <= (layer2_outputs(57)) xor (layer2_outputs(114));
    layer3_outputs(2126) <= not((layer2_outputs(2448)) and (layer2_outputs(2314)));
    layer3_outputs(2127) <= '0';
    layer3_outputs(2128) <= not(layer2_outputs(277));
    layer3_outputs(2129) <= '0';
    layer3_outputs(2130) <= (layer2_outputs(39)) and (layer2_outputs(1941));
    layer3_outputs(2131) <= not(layer2_outputs(2102)) or (layer2_outputs(888));
    layer3_outputs(2132) <= (layer2_outputs(25)) and not (layer2_outputs(2059));
    layer3_outputs(2133) <= not(layer2_outputs(1870)) or (layer2_outputs(2089));
    layer3_outputs(2134) <= not(layer2_outputs(1136));
    layer3_outputs(2135) <= not(layer2_outputs(1739));
    layer3_outputs(2136) <= not(layer2_outputs(793)) or (layer2_outputs(1536));
    layer3_outputs(2137) <= not(layer2_outputs(67));
    layer3_outputs(2138) <= '0';
    layer3_outputs(2139) <= not((layer2_outputs(389)) and (layer2_outputs(837)));
    layer3_outputs(2140) <= not(layer2_outputs(842)) or (layer2_outputs(1239));
    layer3_outputs(2141) <= (layer2_outputs(2488)) and not (layer2_outputs(59));
    layer3_outputs(2142) <= (layer2_outputs(409)) and not (layer2_outputs(2223));
    layer3_outputs(2143) <= not((layer2_outputs(2316)) and (layer2_outputs(2134)));
    layer3_outputs(2144) <= not((layer2_outputs(386)) or (layer2_outputs(1184)));
    layer3_outputs(2145) <= not(layer2_outputs(1663));
    layer3_outputs(2146) <= layer2_outputs(1834);
    layer3_outputs(2147) <= not((layer2_outputs(580)) xor (layer2_outputs(2123)));
    layer3_outputs(2148) <= not(layer2_outputs(710)) or (layer2_outputs(1793));
    layer3_outputs(2149) <= (layer2_outputs(2175)) and not (layer2_outputs(62));
    layer3_outputs(2150) <= not(layer2_outputs(1395));
    layer3_outputs(2151) <= (layer2_outputs(2193)) xor (layer2_outputs(2303));
    layer3_outputs(2152) <= not((layer2_outputs(408)) and (layer2_outputs(1299)));
    layer3_outputs(2153) <= layer2_outputs(213);
    layer3_outputs(2154) <= not(layer2_outputs(1809)) or (layer2_outputs(2416));
    layer3_outputs(2155) <= layer2_outputs(1519);
    layer3_outputs(2156) <= layer2_outputs(913);
    layer3_outputs(2157) <= layer2_outputs(1108);
    layer3_outputs(2158) <= layer2_outputs(2474);
    layer3_outputs(2159) <= not(layer2_outputs(10));
    layer3_outputs(2160) <= not(layer2_outputs(1851));
    layer3_outputs(2161) <= (layer2_outputs(1251)) and not (layer2_outputs(635));
    layer3_outputs(2162) <= not(layer2_outputs(1138));
    layer3_outputs(2163) <= not((layer2_outputs(873)) and (layer2_outputs(470)));
    layer3_outputs(2164) <= (layer2_outputs(1280)) and not (layer2_outputs(446));
    layer3_outputs(2165) <= not((layer2_outputs(2138)) or (layer2_outputs(1509)));
    layer3_outputs(2166) <= (layer2_outputs(2485)) and not (layer2_outputs(394));
    layer3_outputs(2167) <= not(layer2_outputs(2446));
    layer3_outputs(2168) <= not(layer2_outputs(42));
    layer3_outputs(2169) <= not(layer2_outputs(14));
    layer3_outputs(2170) <= layer2_outputs(227);
    layer3_outputs(2171) <= (layer2_outputs(899)) xor (layer2_outputs(351));
    layer3_outputs(2172) <= (layer2_outputs(430)) or (layer2_outputs(2371));
    layer3_outputs(2173) <= not(layer2_outputs(1767));
    layer3_outputs(2174) <= not(layer2_outputs(1726));
    layer3_outputs(2175) <= not(layer2_outputs(284)) or (layer2_outputs(654));
    layer3_outputs(2176) <= layer2_outputs(1323);
    layer3_outputs(2177) <= not(layer2_outputs(1131)) or (layer2_outputs(1412));
    layer3_outputs(2178) <= not(layer2_outputs(974)) or (layer2_outputs(2039));
    layer3_outputs(2179) <= not(layer2_outputs(8));
    layer3_outputs(2180) <= layer2_outputs(1493);
    layer3_outputs(2181) <= not(layer2_outputs(1809)) or (layer2_outputs(1959));
    layer3_outputs(2182) <= layer2_outputs(760);
    layer3_outputs(2183) <= not(layer2_outputs(1001)) or (layer2_outputs(1112));
    layer3_outputs(2184) <= layer2_outputs(2490);
    layer3_outputs(2185) <= not((layer2_outputs(1889)) and (layer2_outputs(1579)));
    layer3_outputs(2186) <= not(layer2_outputs(1174));
    layer3_outputs(2187) <= not((layer2_outputs(889)) and (layer2_outputs(1079)));
    layer3_outputs(2188) <= not(layer2_outputs(1596));
    layer3_outputs(2189) <= not((layer2_outputs(2508)) or (layer2_outputs(740)));
    layer3_outputs(2190) <= not(layer2_outputs(2129));
    layer3_outputs(2191) <= layer2_outputs(1129);
    layer3_outputs(2192) <= not(layer2_outputs(2280));
    layer3_outputs(2193) <= layer2_outputs(842);
    layer3_outputs(2194) <= not(layer2_outputs(997));
    layer3_outputs(2195) <= (layer2_outputs(1435)) or (layer2_outputs(714));
    layer3_outputs(2196) <= (layer2_outputs(814)) xor (layer2_outputs(407));
    layer3_outputs(2197) <= (layer2_outputs(199)) and not (layer2_outputs(1538));
    layer3_outputs(2198) <= (layer2_outputs(1260)) and (layer2_outputs(1483));
    layer3_outputs(2199) <= not(layer2_outputs(781));
    layer3_outputs(2200) <= not(layer2_outputs(2228)) or (layer2_outputs(2517));
    layer3_outputs(2201) <= '1';
    layer3_outputs(2202) <= not(layer2_outputs(1925));
    layer3_outputs(2203) <= not(layer2_outputs(1653));
    layer3_outputs(2204) <= '0';
    layer3_outputs(2205) <= layer2_outputs(162);
    layer3_outputs(2206) <= layer2_outputs(91);
    layer3_outputs(2207) <= (layer2_outputs(1188)) and (layer2_outputs(1119));
    layer3_outputs(2208) <= layer2_outputs(1657);
    layer3_outputs(2209) <= layer2_outputs(1475);
    layer3_outputs(2210) <= '1';
    layer3_outputs(2211) <= (layer2_outputs(606)) xor (layer2_outputs(2501));
    layer3_outputs(2212) <= not(layer2_outputs(1126));
    layer3_outputs(2213) <= layer2_outputs(902);
    layer3_outputs(2214) <= (layer2_outputs(910)) and not (layer2_outputs(114));
    layer3_outputs(2215) <= not((layer2_outputs(2370)) and (layer2_outputs(2269)));
    layer3_outputs(2216) <= layer2_outputs(769);
    layer3_outputs(2217) <= layer2_outputs(2307);
    layer3_outputs(2218) <= (layer2_outputs(435)) and not (layer2_outputs(1901));
    layer3_outputs(2219) <= not(layer2_outputs(1886));
    layer3_outputs(2220) <= '1';
    layer3_outputs(2221) <= not(layer2_outputs(1997)) or (layer2_outputs(1662));
    layer3_outputs(2222) <= not((layer2_outputs(810)) or (layer2_outputs(1486)));
    layer3_outputs(2223) <= (layer2_outputs(600)) or (layer2_outputs(1039));
    layer3_outputs(2224) <= not((layer2_outputs(802)) or (layer2_outputs(1388)));
    layer3_outputs(2225) <= not(layer2_outputs(1667));
    layer3_outputs(2226) <= not((layer2_outputs(35)) and (layer2_outputs(1635)));
    layer3_outputs(2227) <= not(layer2_outputs(1021));
    layer3_outputs(2228) <= (layer2_outputs(687)) and not (layer2_outputs(2421));
    layer3_outputs(2229) <= (layer2_outputs(665)) or (layer2_outputs(1734));
    layer3_outputs(2230) <= layer2_outputs(869);
    layer3_outputs(2231) <= layer2_outputs(385);
    layer3_outputs(2232) <= not((layer2_outputs(62)) xor (layer2_outputs(523)));
    layer3_outputs(2233) <= not(layer2_outputs(905));
    layer3_outputs(2234) <= not(layer2_outputs(514)) or (layer2_outputs(2127));
    layer3_outputs(2235) <= layer2_outputs(2164);
    layer3_outputs(2236) <= (layer2_outputs(673)) or (layer2_outputs(240));
    layer3_outputs(2237) <= not(layer2_outputs(1342)) or (layer2_outputs(1413));
    layer3_outputs(2238) <= (layer2_outputs(1706)) and not (layer2_outputs(1341));
    layer3_outputs(2239) <= (layer2_outputs(1878)) and not (layer2_outputs(69));
    layer3_outputs(2240) <= (layer2_outputs(1676)) and not (layer2_outputs(755));
    layer3_outputs(2241) <= layer2_outputs(1842);
    layer3_outputs(2242) <= not(layer2_outputs(1642));
    layer3_outputs(2243) <= layer2_outputs(1526);
    layer3_outputs(2244) <= not((layer2_outputs(1586)) xor (layer2_outputs(1458)));
    layer3_outputs(2245) <= not((layer2_outputs(886)) or (layer2_outputs(359)));
    layer3_outputs(2246) <= not((layer2_outputs(2418)) or (layer2_outputs(881)));
    layer3_outputs(2247) <= not(layer2_outputs(2390));
    layer3_outputs(2248) <= (layer2_outputs(1677)) and not (layer2_outputs(1693));
    layer3_outputs(2249) <= (layer2_outputs(160)) and not (layer2_outputs(2047));
    layer3_outputs(2250) <= layer2_outputs(1049);
    layer3_outputs(2251) <= layer2_outputs(1971);
    layer3_outputs(2252) <= not(layer2_outputs(1200));
    layer3_outputs(2253) <= layer2_outputs(1980);
    layer3_outputs(2254) <= layer2_outputs(1887);
    layer3_outputs(2255) <= not((layer2_outputs(1998)) xor (layer2_outputs(2230)));
    layer3_outputs(2256) <= '1';
    layer3_outputs(2257) <= not(layer2_outputs(1044));
    layer3_outputs(2258) <= layer2_outputs(2126);
    layer3_outputs(2259) <= layer2_outputs(817);
    layer3_outputs(2260) <= not((layer2_outputs(1739)) and (layer2_outputs(85)));
    layer3_outputs(2261) <= layer2_outputs(432);
    layer3_outputs(2262) <= not(layer2_outputs(2523));
    layer3_outputs(2263) <= (layer2_outputs(1448)) xor (layer2_outputs(2212));
    layer3_outputs(2264) <= not(layer2_outputs(2012));
    layer3_outputs(2265) <= not(layer2_outputs(1225)) or (layer2_outputs(231));
    layer3_outputs(2266) <= not(layer2_outputs(833));
    layer3_outputs(2267) <= (layer2_outputs(817)) and not (layer2_outputs(1031));
    layer3_outputs(2268) <= (layer2_outputs(2195)) or (layer2_outputs(2243));
    layer3_outputs(2269) <= not((layer2_outputs(2239)) or (layer2_outputs(2071)));
    layer3_outputs(2270) <= (layer2_outputs(1386)) and not (layer2_outputs(418));
    layer3_outputs(2271) <= layer2_outputs(352);
    layer3_outputs(2272) <= not(layer2_outputs(504));
    layer3_outputs(2273) <= layer2_outputs(1840);
    layer3_outputs(2274) <= layer2_outputs(22);
    layer3_outputs(2275) <= (layer2_outputs(506)) and not (layer2_outputs(1964));
    layer3_outputs(2276) <= (layer2_outputs(485)) xor (layer2_outputs(1620));
    layer3_outputs(2277) <= (layer2_outputs(1453)) and not (layer2_outputs(1573));
    layer3_outputs(2278) <= layer2_outputs(1717);
    layer3_outputs(2279) <= layer2_outputs(329);
    layer3_outputs(2280) <= not(layer2_outputs(638));
    layer3_outputs(2281) <= not(layer2_outputs(391));
    layer3_outputs(2282) <= layer2_outputs(391);
    layer3_outputs(2283) <= (layer2_outputs(2097)) and (layer2_outputs(2243));
    layer3_outputs(2284) <= not((layer2_outputs(2045)) and (layer2_outputs(2503)));
    layer3_outputs(2285) <= '1';
    layer3_outputs(2286) <= not(layer2_outputs(2512));
    layer3_outputs(2287) <= not(layer2_outputs(1024));
    layer3_outputs(2288) <= not(layer2_outputs(193)) or (layer2_outputs(2248));
    layer3_outputs(2289) <= not(layer2_outputs(2108)) or (layer2_outputs(825));
    layer3_outputs(2290) <= not(layer2_outputs(472)) or (layer2_outputs(596));
    layer3_outputs(2291) <= '1';
    layer3_outputs(2292) <= not((layer2_outputs(1610)) xor (layer2_outputs(1894)));
    layer3_outputs(2293) <= layer2_outputs(2155);
    layer3_outputs(2294) <= not((layer2_outputs(2003)) and (layer2_outputs(1368)));
    layer3_outputs(2295) <= not(layer2_outputs(354)) or (layer2_outputs(1495));
    layer3_outputs(2296) <= not(layer2_outputs(1268));
    layer3_outputs(2297) <= not(layer2_outputs(428)) or (layer2_outputs(1946));
    layer3_outputs(2298) <= not((layer2_outputs(1139)) or (layer2_outputs(628)));
    layer3_outputs(2299) <= not(layer2_outputs(2439));
    layer3_outputs(2300) <= layer2_outputs(555);
    layer3_outputs(2301) <= (layer2_outputs(1872)) xor (layer2_outputs(372));
    layer3_outputs(2302) <= not(layer2_outputs(318)) or (layer2_outputs(658));
    layer3_outputs(2303) <= not((layer2_outputs(543)) or (layer2_outputs(2352)));
    layer3_outputs(2304) <= not((layer2_outputs(2174)) xor (layer2_outputs(764)));
    layer3_outputs(2305) <= layer2_outputs(2546);
    layer3_outputs(2306) <= not(layer2_outputs(1583)) or (layer2_outputs(1697));
    layer3_outputs(2307) <= layer2_outputs(893);
    layer3_outputs(2308) <= (layer2_outputs(2376)) and not (layer2_outputs(1115));
    layer3_outputs(2309) <= not(layer2_outputs(518)) or (layer2_outputs(1551));
    layer3_outputs(2310) <= layer2_outputs(1124);
    layer3_outputs(2311) <= not((layer2_outputs(2356)) or (layer2_outputs(1302)));
    layer3_outputs(2312) <= not(layer2_outputs(2050));
    layer3_outputs(2313) <= not(layer2_outputs(448));
    layer3_outputs(2314) <= (layer2_outputs(342)) and not (layer2_outputs(847));
    layer3_outputs(2315) <= not(layer2_outputs(1235)) or (layer2_outputs(1092));
    layer3_outputs(2316) <= (layer2_outputs(533)) and (layer2_outputs(1194));
    layer3_outputs(2317) <= not(layer2_outputs(462));
    layer3_outputs(2318) <= not(layer2_outputs(2341)) or (layer2_outputs(335));
    layer3_outputs(2319) <= not(layer2_outputs(335));
    layer3_outputs(2320) <= not(layer2_outputs(231));
    layer3_outputs(2321) <= not(layer2_outputs(2153));
    layer3_outputs(2322) <= not((layer2_outputs(1969)) and (layer2_outputs(957)));
    layer3_outputs(2323) <= layer2_outputs(1702);
    layer3_outputs(2324) <= not(layer2_outputs(1539));
    layer3_outputs(2325) <= layer2_outputs(1314);
    layer3_outputs(2326) <= layer2_outputs(137);
    layer3_outputs(2327) <= not(layer2_outputs(1885));
    layer3_outputs(2328) <= '1';
    layer3_outputs(2329) <= not(layer2_outputs(1343)) or (layer2_outputs(2371));
    layer3_outputs(2330) <= not(layer2_outputs(1379)) or (layer2_outputs(1900));
    layer3_outputs(2331) <= not(layer2_outputs(1561));
    layer3_outputs(2332) <= not(layer2_outputs(445)) or (layer2_outputs(1441));
    layer3_outputs(2333) <= layer2_outputs(638);
    layer3_outputs(2334) <= (layer2_outputs(1888)) and (layer2_outputs(2220));
    layer3_outputs(2335) <= not(layer2_outputs(2011)) or (layer2_outputs(1813));
    layer3_outputs(2336) <= not(layer2_outputs(1721));
    layer3_outputs(2337) <= not(layer2_outputs(1611)) or (layer2_outputs(1335));
    layer3_outputs(2338) <= layer2_outputs(2255);
    layer3_outputs(2339) <= layer2_outputs(1719);
    layer3_outputs(2340) <= not(layer2_outputs(498));
    layer3_outputs(2341) <= not(layer2_outputs(772)) or (layer2_outputs(1933));
    layer3_outputs(2342) <= not(layer2_outputs(776)) or (layer2_outputs(207));
    layer3_outputs(2343) <= not((layer2_outputs(2294)) or (layer2_outputs(732)));
    layer3_outputs(2344) <= layer2_outputs(368);
    layer3_outputs(2345) <= (layer2_outputs(1599)) xor (layer2_outputs(621));
    layer3_outputs(2346) <= not(layer2_outputs(2522));
    layer3_outputs(2347) <= (layer2_outputs(2425)) xor (layer2_outputs(27));
    layer3_outputs(2348) <= layer2_outputs(133);
    layer3_outputs(2349) <= (layer2_outputs(1816)) and not (layer2_outputs(1877));
    layer3_outputs(2350) <= not(layer2_outputs(995));
    layer3_outputs(2351) <= not(layer2_outputs(364));
    layer3_outputs(2352) <= (layer2_outputs(1418)) or (layer2_outputs(2246));
    layer3_outputs(2353) <= (layer2_outputs(1727)) and (layer2_outputs(416));
    layer3_outputs(2354) <= not(layer2_outputs(349));
    layer3_outputs(2355) <= (layer2_outputs(1076)) and not (layer2_outputs(2398));
    layer3_outputs(2356) <= layer2_outputs(117);
    layer3_outputs(2357) <= layer2_outputs(668);
    layer3_outputs(2358) <= (layer2_outputs(1923)) and not (layer2_outputs(2348));
    layer3_outputs(2359) <= '1';
    layer3_outputs(2360) <= not((layer2_outputs(1863)) or (layer2_outputs(2007)));
    layer3_outputs(2361) <= not((layer2_outputs(2106)) or (layer2_outputs(81)));
    layer3_outputs(2362) <= not(layer2_outputs(763));
    layer3_outputs(2363) <= not(layer2_outputs(2192));
    layer3_outputs(2364) <= layer2_outputs(1328);
    layer3_outputs(2365) <= '1';
    layer3_outputs(2366) <= '0';
    layer3_outputs(2367) <= not(layer2_outputs(1489)) or (layer2_outputs(210));
    layer3_outputs(2368) <= not(layer2_outputs(1373)) or (layer2_outputs(169));
    layer3_outputs(2369) <= layer2_outputs(1902);
    layer3_outputs(2370) <= layer2_outputs(1851);
    layer3_outputs(2371) <= layer2_outputs(301);
    layer3_outputs(2372) <= (layer2_outputs(849)) and not (layer2_outputs(2105));
    layer3_outputs(2373) <= not(layer2_outputs(2023));
    layer3_outputs(2374) <= (layer2_outputs(656)) or (layer2_outputs(240));
    layer3_outputs(2375) <= not(layer2_outputs(1390));
    layer3_outputs(2376) <= not(layer2_outputs(282)) or (layer2_outputs(1062));
    layer3_outputs(2377) <= layer2_outputs(1292);
    layer3_outputs(2378) <= layer2_outputs(692);
    layer3_outputs(2379) <= not((layer2_outputs(1474)) or (layer2_outputs(1761)));
    layer3_outputs(2380) <= (layer2_outputs(1425)) and not (layer2_outputs(2519));
    layer3_outputs(2381) <= not(layer2_outputs(2133));
    layer3_outputs(2382) <= (layer2_outputs(1621)) and (layer2_outputs(1201));
    layer3_outputs(2383) <= layer2_outputs(2539);
    layer3_outputs(2384) <= (layer2_outputs(2549)) and not (layer2_outputs(802));
    layer3_outputs(2385) <= '0';
    layer3_outputs(2386) <= not((layer2_outputs(1304)) xor (layer2_outputs(1340)));
    layer3_outputs(2387) <= layer2_outputs(509);
    layer3_outputs(2388) <= '1';
    layer3_outputs(2389) <= not((layer2_outputs(648)) and (layer2_outputs(805)));
    layer3_outputs(2390) <= layer2_outputs(2116);
    layer3_outputs(2391) <= not(layer2_outputs(202)) or (layer2_outputs(44));
    layer3_outputs(2392) <= not(layer2_outputs(1030)) or (layer2_outputs(338));
    layer3_outputs(2393) <= layer2_outputs(2267);
    layer3_outputs(2394) <= layer2_outputs(2032);
    layer3_outputs(2395) <= layer2_outputs(1428);
    layer3_outputs(2396) <= (layer2_outputs(2544)) and (layer2_outputs(1114));
    layer3_outputs(2397) <= '0';
    layer3_outputs(2398) <= not(layer2_outputs(256));
    layer3_outputs(2399) <= layer2_outputs(420);
    layer3_outputs(2400) <= layer2_outputs(1288);
    layer3_outputs(2401) <= layer2_outputs(244);
    layer3_outputs(2402) <= not(layer2_outputs(1048));
    layer3_outputs(2403) <= not(layer2_outputs(2281));
    layer3_outputs(2404) <= layer2_outputs(1103);
    layer3_outputs(2405) <= '1';
    layer3_outputs(2406) <= not(layer2_outputs(508)) or (layer2_outputs(529));
    layer3_outputs(2407) <= '1';
    layer3_outputs(2408) <= (layer2_outputs(88)) or (layer2_outputs(3));
    layer3_outputs(2409) <= (layer2_outputs(2027)) and not (layer2_outputs(1478));
    layer3_outputs(2410) <= (layer2_outputs(1770)) and (layer2_outputs(1802));
    layer3_outputs(2411) <= '0';
    layer3_outputs(2412) <= layer2_outputs(1707);
    layer3_outputs(2413) <= (layer2_outputs(1659)) or (layer2_outputs(48));
    layer3_outputs(2414) <= (layer2_outputs(1595)) and not (layer2_outputs(882));
    layer3_outputs(2415) <= not(layer2_outputs(1383)) or (layer2_outputs(1762));
    layer3_outputs(2416) <= '0';
    layer3_outputs(2417) <= not(layer2_outputs(2409));
    layer3_outputs(2418) <= layer2_outputs(1283);
    layer3_outputs(2419) <= (layer2_outputs(1444)) or (layer2_outputs(1123));
    layer3_outputs(2420) <= not((layer2_outputs(1590)) or (layer2_outputs(2263)));
    layer3_outputs(2421) <= not(layer2_outputs(34));
    layer3_outputs(2422) <= not((layer2_outputs(41)) and (layer2_outputs(1197)));
    layer3_outputs(2423) <= not((layer2_outputs(2458)) xor (layer2_outputs(493)));
    layer3_outputs(2424) <= layer2_outputs(2391);
    layer3_outputs(2425) <= not((layer2_outputs(1063)) or (layer2_outputs(931)));
    layer3_outputs(2426) <= not(layer2_outputs(332)) or (layer2_outputs(1930));
    layer3_outputs(2427) <= not(layer2_outputs(1050));
    layer3_outputs(2428) <= not(layer2_outputs(1345));
    layer3_outputs(2429) <= not(layer2_outputs(1119));
    layer3_outputs(2430) <= not((layer2_outputs(205)) and (layer2_outputs(323)));
    layer3_outputs(2431) <= (layer2_outputs(387)) or (layer2_outputs(375));
    layer3_outputs(2432) <= not(layer2_outputs(2401));
    layer3_outputs(2433) <= layer2_outputs(2058);
    layer3_outputs(2434) <= not(layer2_outputs(2268));
    layer3_outputs(2435) <= not((layer2_outputs(2167)) or (layer2_outputs(1607)));
    layer3_outputs(2436) <= layer2_outputs(1108);
    layer3_outputs(2437) <= not(layer2_outputs(211));
    layer3_outputs(2438) <= (layer2_outputs(1418)) and not (layer2_outputs(441));
    layer3_outputs(2439) <= not((layer2_outputs(561)) and (layer2_outputs(1755)));
    layer3_outputs(2440) <= not((layer2_outputs(913)) or (layer2_outputs(1501)));
    layer3_outputs(2441) <= not(layer2_outputs(330));
    layer3_outputs(2442) <= not(layer2_outputs(309));
    layer3_outputs(2443) <= layer2_outputs(135);
    layer3_outputs(2444) <= (layer2_outputs(1338)) xor (layer2_outputs(413));
    layer3_outputs(2445) <= not((layer2_outputs(988)) or (layer2_outputs(836)));
    layer3_outputs(2446) <= layer2_outputs(9);
    layer3_outputs(2447) <= layer2_outputs(1399);
    layer3_outputs(2448) <= not(layer2_outputs(1364));
    layer3_outputs(2449) <= layer2_outputs(555);
    layer3_outputs(2450) <= not(layer2_outputs(1176));
    layer3_outputs(2451) <= (layer2_outputs(1354)) or (layer2_outputs(945));
    layer3_outputs(2452) <= (layer2_outputs(1233)) and not (layer2_outputs(1344));
    layer3_outputs(2453) <= not(layer2_outputs(539));
    layer3_outputs(2454) <= (layer2_outputs(976)) and not (layer2_outputs(2385));
    layer3_outputs(2455) <= (layer2_outputs(1868)) and not (layer2_outputs(1413));
    layer3_outputs(2456) <= layer2_outputs(2379);
    layer3_outputs(2457) <= (layer2_outputs(670)) xor (layer2_outputs(251));
    layer3_outputs(2458) <= layer2_outputs(2347);
    layer3_outputs(2459) <= '1';
    layer3_outputs(2460) <= (layer2_outputs(1436)) and (layer2_outputs(2081));
    layer3_outputs(2461) <= (layer2_outputs(2177)) and (layer2_outputs(8));
    layer3_outputs(2462) <= (layer2_outputs(360)) and (layer2_outputs(1993));
    layer3_outputs(2463) <= not(layer2_outputs(2089));
    layer3_outputs(2464) <= (layer2_outputs(259)) or (layer2_outputs(372));
    layer3_outputs(2465) <= not(layer2_outputs(353));
    layer3_outputs(2466) <= '1';
    layer3_outputs(2467) <= not((layer2_outputs(6)) xor (layer2_outputs(2003)));
    layer3_outputs(2468) <= layer2_outputs(1724);
    layer3_outputs(2469) <= layer2_outputs(2210);
    layer3_outputs(2470) <= '1';
    layer3_outputs(2471) <= not(layer2_outputs(2248));
    layer3_outputs(2472) <= (layer2_outputs(1305)) and (layer2_outputs(2095));
    layer3_outputs(2473) <= layer2_outputs(798);
    layer3_outputs(2474) <= layer2_outputs(395);
    layer3_outputs(2475) <= not(layer2_outputs(2451));
    layer3_outputs(2476) <= layer2_outputs(1347);
    layer3_outputs(2477) <= (layer2_outputs(850)) or (layer2_outputs(1585));
    layer3_outputs(2478) <= '1';
    layer3_outputs(2479) <= layer2_outputs(2067);
    layer3_outputs(2480) <= not(layer2_outputs(381));
    layer3_outputs(2481) <= not(layer2_outputs(333));
    layer3_outputs(2482) <= not((layer2_outputs(1414)) or (layer2_outputs(956)));
    layer3_outputs(2483) <= not(layer2_outputs(2475));
    layer3_outputs(2484) <= layer2_outputs(230);
    layer3_outputs(2485) <= layer2_outputs(1864);
    layer3_outputs(2486) <= '1';
    layer3_outputs(2487) <= (layer2_outputs(522)) and not (layer2_outputs(604));
    layer3_outputs(2488) <= not(layer2_outputs(1027)) or (layer2_outputs(1368));
    layer3_outputs(2489) <= not((layer2_outputs(1303)) or (layer2_outputs(1491)));
    layer3_outputs(2490) <= layer2_outputs(2464);
    layer3_outputs(2491) <= not(layer2_outputs(88));
    layer3_outputs(2492) <= layer2_outputs(2177);
    layer3_outputs(2493) <= not(layer2_outputs(195));
    layer3_outputs(2494) <= layer2_outputs(1238);
    layer3_outputs(2495) <= not(layer2_outputs(1780));
    layer3_outputs(2496) <= not(layer2_outputs(1330)) or (layer2_outputs(1822));
    layer3_outputs(2497) <= (layer2_outputs(1082)) and not (layer2_outputs(1253));
    layer3_outputs(2498) <= not(layer2_outputs(243));
    layer3_outputs(2499) <= (layer2_outputs(1412)) and (layer2_outputs(232));
    layer3_outputs(2500) <= layer2_outputs(1573);
    layer3_outputs(2501) <= not(layer2_outputs(99));
    layer3_outputs(2502) <= layer2_outputs(1788);
    layer3_outputs(2503) <= layer2_outputs(1234);
    layer3_outputs(2504) <= layer2_outputs(809);
    layer3_outputs(2505) <= not(layer2_outputs(127));
    layer3_outputs(2506) <= not(layer2_outputs(1926));
    layer3_outputs(2507) <= (layer2_outputs(584)) and (layer2_outputs(1345));
    layer3_outputs(2508) <= not(layer2_outputs(1924));
    layer3_outputs(2509) <= not(layer2_outputs(478));
    layer3_outputs(2510) <= not(layer2_outputs(1733));
    layer3_outputs(2511) <= not(layer2_outputs(1185)) or (layer2_outputs(413));
    layer3_outputs(2512) <= layer2_outputs(1880);
    layer3_outputs(2513) <= not((layer2_outputs(301)) or (layer2_outputs(2473)));
    layer3_outputs(2514) <= (layer2_outputs(960)) or (layer2_outputs(510));
    layer3_outputs(2515) <= not((layer2_outputs(470)) xor (layer2_outputs(1770)));
    layer3_outputs(2516) <= not(layer2_outputs(315));
    layer3_outputs(2517) <= not((layer2_outputs(884)) or (layer2_outputs(1516)));
    layer3_outputs(2518) <= '1';
    layer3_outputs(2519) <= '0';
    layer3_outputs(2520) <= not(layer2_outputs(1155)) or (layer2_outputs(1784));
    layer3_outputs(2521) <= (layer2_outputs(250)) and not (layer2_outputs(2232));
    layer3_outputs(2522) <= (layer2_outputs(1863)) xor (layer2_outputs(417));
    layer3_outputs(2523) <= layer2_outputs(136);
    layer3_outputs(2524) <= (layer2_outputs(577)) and (layer2_outputs(904));
    layer3_outputs(2525) <= not(layer2_outputs(1760));
    layer3_outputs(2526) <= (layer2_outputs(1897)) and not (layer2_outputs(2387));
    layer3_outputs(2527) <= '1';
    layer3_outputs(2528) <= layer2_outputs(1215);
    layer3_outputs(2529) <= not((layer2_outputs(1257)) and (layer2_outputs(1045)));
    layer3_outputs(2530) <= not(layer2_outputs(13));
    layer3_outputs(2531) <= layer2_outputs(866);
    layer3_outputs(2532) <= (layer2_outputs(1232)) or (layer2_outputs(1638));
    layer3_outputs(2533) <= layer2_outputs(2542);
    layer3_outputs(2534) <= (layer2_outputs(647)) or (layer2_outputs(126));
    layer3_outputs(2535) <= '1';
    layer3_outputs(2536) <= not(layer2_outputs(1252));
    layer3_outputs(2537) <= (layer2_outputs(922)) and not (layer2_outputs(2261));
    layer3_outputs(2538) <= not(layer2_outputs(2199));
    layer3_outputs(2539) <= not((layer2_outputs(1945)) or (layer2_outputs(1465)));
    layer3_outputs(2540) <= '1';
    layer3_outputs(2541) <= (layer2_outputs(501)) or (layer2_outputs(49));
    layer3_outputs(2542) <= layer2_outputs(903);
    layer3_outputs(2543) <= not(layer2_outputs(680));
    layer3_outputs(2544) <= not(layer2_outputs(2051));
    layer3_outputs(2545) <= layer2_outputs(1920);
    layer3_outputs(2546) <= '1';
    layer3_outputs(2547) <= layer2_outputs(1691);
    layer3_outputs(2548) <= not(layer2_outputs(172));
    layer3_outputs(2549) <= not(layer2_outputs(1967));
    layer3_outputs(2550) <= layer2_outputs(1601);
    layer3_outputs(2551) <= not(layer2_outputs(1177));
    layer3_outputs(2552) <= not(layer2_outputs(2454));
    layer3_outputs(2553) <= not(layer2_outputs(400));
    layer3_outputs(2554) <= layer2_outputs(691);
    layer3_outputs(2555) <= (layer2_outputs(1451)) or (layer2_outputs(2290));
    layer3_outputs(2556) <= layer2_outputs(754);
    layer3_outputs(2557) <= not(layer2_outputs(197));
    layer3_outputs(2558) <= (layer2_outputs(1587)) xor (layer2_outputs(1571));
    layer3_outputs(2559) <= not(layer2_outputs(170));
    layer4_outputs(0) <= layer3_outputs(1302);
    layer4_outputs(1) <= not(layer3_outputs(1103));
    layer4_outputs(2) <= '1';
    layer4_outputs(3) <= layer3_outputs(2050);
    layer4_outputs(4) <= not(layer3_outputs(428)) or (layer3_outputs(154));
    layer4_outputs(5) <= layer3_outputs(324);
    layer4_outputs(6) <= layer3_outputs(672);
    layer4_outputs(7) <= not(layer3_outputs(1109)) or (layer3_outputs(2499));
    layer4_outputs(8) <= not(layer3_outputs(340));
    layer4_outputs(9) <= not(layer3_outputs(2102));
    layer4_outputs(10) <= (layer3_outputs(2534)) or (layer3_outputs(1352));
    layer4_outputs(11) <= (layer3_outputs(753)) and (layer3_outputs(915));
    layer4_outputs(12) <= not(layer3_outputs(1375));
    layer4_outputs(13) <= (layer3_outputs(914)) or (layer3_outputs(132));
    layer4_outputs(14) <= not(layer3_outputs(711));
    layer4_outputs(15) <= '0';
    layer4_outputs(16) <= layer3_outputs(223);
    layer4_outputs(17) <= (layer3_outputs(694)) and not (layer3_outputs(203));
    layer4_outputs(18) <= not((layer3_outputs(896)) and (layer3_outputs(2021)));
    layer4_outputs(19) <= (layer3_outputs(1395)) xor (layer3_outputs(669));
    layer4_outputs(20) <= not(layer3_outputs(1392)) or (layer3_outputs(1293));
    layer4_outputs(21) <= (layer3_outputs(1634)) or (layer3_outputs(1192));
    layer4_outputs(22) <= not(layer3_outputs(78));
    layer4_outputs(23) <= not((layer3_outputs(322)) or (layer3_outputs(517)));
    layer4_outputs(24) <= not((layer3_outputs(536)) or (layer3_outputs(309)));
    layer4_outputs(25) <= '1';
    layer4_outputs(26) <= layer3_outputs(2034);
    layer4_outputs(27) <= (layer3_outputs(660)) and not (layer3_outputs(2214));
    layer4_outputs(28) <= (layer3_outputs(90)) xor (layer3_outputs(1062));
    layer4_outputs(29) <= (layer3_outputs(1728)) and not (layer3_outputs(1032));
    layer4_outputs(30) <= not((layer3_outputs(2474)) or (layer3_outputs(620)));
    layer4_outputs(31) <= layer3_outputs(2531);
    layer4_outputs(32) <= not(layer3_outputs(1260)) or (layer3_outputs(349));
    layer4_outputs(33) <= not(layer3_outputs(2213)) or (layer3_outputs(1287));
    layer4_outputs(34) <= not(layer3_outputs(2120));
    layer4_outputs(35) <= not((layer3_outputs(802)) xor (layer3_outputs(1794)));
    layer4_outputs(36) <= not((layer3_outputs(1204)) or (layer3_outputs(307)));
    layer4_outputs(37) <= not(layer3_outputs(837));
    layer4_outputs(38) <= not(layer3_outputs(495));
    layer4_outputs(39) <= layer3_outputs(1915);
    layer4_outputs(40) <= not((layer3_outputs(1171)) and (layer3_outputs(1722)));
    layer4_outputs(41) <= not(layer3_outputs(1913));
    layer4_outputs(42) <= layer3_outputs(1276);
    layer4_outputs(43) <= (layer3_outputs(1328)) and not (layer3_outputs(1246));
    layer4_outputs(44) <= not(layer3_outputs(936));
    layer4_outputs(45) <= layer3_outputs(706);
    layer4_outputs(46) <= not(layer3_outputs(2316));
    layer4_outputs(47) <= layer3_outputs(1427);
    layer4_outputs(48) <= not(layer3_outputs(2104)) or (layer3_outputs(2409));
    layer4_outputs(49) <= not((layer3_outputs(1796)) xor (layer3_outputs(1796)));
    layer4_outputs(50) <= not(layer3_outputs(1638));
    layer4_outputs(51) <= layer3_outputs(2055);
    layer4_outputs(52) <= layer3_outputs(2108);
    layer4_outputs(53) <= '0';
    layer4_outputs(54) <= layer3_outputs(772);
    layer4_outputs(55) <= (layer3_outputs(247)) and not (layer3_outputs(2173));
    layer4_outputs(56) <= not(layer3_outputs(841));
    layer4_outputs(57) <= (layer3_outputs(1190)) and not (layer3_outputs(823));
    layer4_outputs(58) <= not(layer3_outputs(448)) or (layer3_outputs(2454));
    layer4_outputs(59) <= (layer3_outputs(759)) and (layer3_outputs(39));
    layer4_outputs(60) <= not(layer3_outputs(1331)) or (layer3_outputs(1145));
    layer4_outputs(61) <= not(layer3_outputs(765)) or (layer3_outputs(1009));
    layer4_outputs(62) <= not((layer3_outputs(698)) or (layer3_outputs(2042)));
    layer4_outputs(63) <= layer3_outputs(983);
    layer4_outputs(64) <= (layer3_outputs(1058)) and not (layer3_outputs(832));
    layer4_outputs(65) <= (layer3_outputs(1497)) and (layer3_outputs(1505));
    layer4_outputs(66) <= not(layer3_outputs(596));
    layer4_outputs(67) <= not((layer3_outputs(2331)) or (layer3_outputs(1097)));
    layer4_outputs(68) <= layer3_outputs(2272);
    layer4_outputs(69) <= layer3_outputs(217);
    layer4_outputs(70) <= (layer3_outputs(761)) and not (layer3_outputs(2412));
    layer4_outputs(71) <= not(layer3_outputs(1455));
    layer4_outputs(72) <= layer3_outputs(431);
    layer4_outputs(73) <= (layer3_outputs(1883)) and not (layer3_outputs(1166));
    layer4_outputs(74) <= not(layer3_outputs(502));
    layer4_outputs(75) <= not(layer3_outputs(894));
    layer4_outputs(76) <= (layer3_outputs(734)) and not (layer3_outputs(2431));
    layer4_outputs(77) <= not(layer3_outputs(2516));
    layer4_outputs(78) <= not(layer3_outputs(1005));
    layer4_outputs(79) <= not(layer3_outputs(311));
    layer4_outputs(80) <= not((layer3_outputs(1582)) and (layer3_outputs(583)));
    layer4_outputs(81) <= not((layer3_outputs(2073)) and (layer3_outputs(1135)));
    layer4_outputs(82) <= not(layer3_outputs(1635));
    layer4_outputs(83) <= (layer3_outputs(2491)) and not (layer3_outputs(52));
    layer4_outputs(84) <= layer3_outputs(1347);
    layer4_outputs(85) <= not(layer3_outputs(1203));
    layer4_outputs(86) <= not(layer3_outputs(1312));
    layer4_outputs(87) <= not(layer3_outputs(383));
    layer4_outputs(88) <= not((layer3_outputs(144)) or (layer3_outputs(354)));
    layer4_outputs(89) <= not(layer3_outputs(948));
    layer4_outputs(90) <= not((layer3_outputs(225)) xor (layer3_outputs(1434)));
    layer4_outputs(91) <= (layer3_outputs(1674)) or (layer3_outputs(1964));
    layer4_outputs(92) <= not(layer3_outputs(37));
    layer4_outputs(93) <= not((layer3_outputs(14)) xor (layer3_outputs(1337)));
    layer4_outputs(94) <= '1';
    layer4_outputs(95) <= layer3_outputs(609);
    layer4_outputs(96) <= not(layer3_outputs(2006)) or (layer3_outputs(1250));
    layer4_outputs(97) <= not(layer3_outputs(1556)) or (layer3_outputs(1295));
    layer4_outputs(98) <= '0';
    layer4_outputs(99) <= (layer3_outputs(420)) and not (layer3_outputs(1977));
    layer4_outputs(100) <= layer3_outputs(892);
    layer4_outputs(101) <= (layer3_outputs(1330)) xor (layer3_outputs(769));
    layer4_outputs(102) <= not(layer3_outputs(1820));
    layer4_outputs(103) <= not(layer3_outputs(2469));
    layer4_outputs(104) <= layer3_outputs(2558);
    layer4_outputs(105) <= not((layer3_outputs(1946)) xor (layer3_outputs(1298)));
    layer4_outputs(106) <= not(layer3_outputs(873)) or (layer3_outputs(1472));
    layer4_outputs(107) <= not((layer3_outputs(2085)) and (layer3_outputs(1506)));
    layer4_outputs(108) <= (layer3_outputs(1983)) or (layer3_outputs(1415));
    layer4_outputs(109) <= not(layer3_outputs(1810));
    layer4_outputs(110) <= (layer3_outputs(1924)) and not (layer3_outputs(1533));
    layer4_outputs(111) <= (layer3_outputs(2217)) and not (layer3_outputs(303));
    layer4_outputs(112) <= not(layer3_outputs(2317));
    layer4_outputs(113) <= (layer3_outputs(1701)) and not (layer3_outputs(261));
    layer4_outputs(114) <= layer3_outputs(1951);
    layer4_outputs(115) <= '1';
    layer4_outputs(116) <= layer3_outputs(1134);
    layer4_outputs(117) <= not(layer3_outputs(2009));
    layer4_outputs(118) <= not(layer3_outputs(101)) or (layer3_outputs(1584));
    layer4_outputs(119) <= not(layer3_outputs(1693));
    layer4_outputs(120) <= (layer3_outputs(340)) or (layer3_outputs(1271));
    layer4_outputs(121) <= not(layer3_outputs(186));
    layer4_outputs(122) <= not((layer3_outputs(2123)) xor (layer3_outputs(1473)));
    layer4_outputs(123) <= (layer3_outputs(975)) and not (layer3_outputs(1605));
    layer4_outputs(124) <= (layer3_outputs(178)) and not (layer3_outputs(698));
    layer4_outputs(125) <= '1';
    layer4_outputs(126) <= not(layer3_outputs(1216));
    layer4_outputs(127) <= (layer3_outputs(424)) and not (layer3_outputs(334));
    layer4_outputs(128) <= not(layer3_outputs(1026));
    layer4_outputs(129) <= layer3_outputs(362);
    layer4_outputs(130) <= not(layer3_outputs(1631));
    layer4_outputs(131) <= not(layer3_outputs(744));
    layer4_outputs(132) <= layer3_outputs(1336);
    layer4_outputs(133) <= not(layer3_outputs(1647));
    layer4_outputs(134) <= not(layer3_outputs(2162)) or (layer3_outputs(2197));
    layer4_outputs(135) <= layer3_outputs(2349);
    layer4_outputs(136) <= (layer3_outputs(1848)) or (layer3_outputs(2267));
    layer4_outputs(137) <= (layer3_outputs(1288)) and not (layer3_outputs(1002));
    layer4_outputs(138) <= (layer3_outputs(754)) and not (layer3_outputs(4));
    layer4_outputs(139) <= layer3_outputs(1403);
    layer4_outputs(140) <= not(layer3_outputs(2099));
    layer4_outputs(141) <= not(layer3_outputs(1606));
    layer4_outputs(142) <= not(layer3_outputs(2135));
    layer4_outputs(143) <= layer3_outputs(347);
    layer4_outputs(144) <= layer3_outputs(1905);
    layer4_outputs(145) <= layer3_outputs(181);
    layer4_outputs(146) <= not(layer3_outputs(244));
    layer4_outputs(147) <= (layer3_outputs(1962)) or (layer3_outputs(1069));
    layer4_outputs(148) <= layer3_outputs(10);
    layer4_outputs(149) <= not(layer3_outputs(407));
    layer4_outputs(150) <= layer3_outputs(1045);
    layer4_outputs(151) <= (layer3_outputs(588)) and not (layer3_outputs(1872));
    layer4_outputs(152) <= (layer3_outputs(2280)) or (layer3_outputs(520));
    layer4_outputs(153) <= layer3_outputs(140);
    layer4_outputs(154) <= layer3_outputs(1354);
    layer4_outputs(155) <= not(layer3_outputs(2273));
    layer4_outputs(156) <= not(layer3_outputs(160));
    layer4_outputs(157) <= (layer3_outputs(2126)) xor (layer3_outputs(2253));
    layer4_outputs(158) <= not((layer3_outputs(755)) or (layer3_outputs(2232)));
    layer4_outputs(159) <= (layer3_outputs(67)) or (layer3_outputs(1949));
    layer4_outputs(160) <= layer3_outputs(2156);
    layer4_outputs(161) <= not(layer3_outputs(1835));
    layer4_outputs(162) <= layer3_outputs(206);
    layer4_outputs(163) <= layer3_outputs(2405);
    layer4_outputs(164) <= not((layer3_outputs(1033)) and (layer3_outputs(1169)));
    layer4_outputs(165) <= (layer3_outputs(995)) and not (layer3_outputs(1814));
    layer4_outputs(166) <= layer3_outputs(371);
    layer4_outputs(167) <= (layer3_outputs(871)) and not (layer3_outputs(2542));
    layer4_outputs(168) <= not((layer3_outputs(2435)) xor (layer3_outputs(1275)));
    layer4_outputs(169) <= '1';
    layer4_outputs(170) <= layer3_outputs(1808);
    layer4_outputs(171) <= not((layer3_outputs(2107)) and (layer3_outputs(2196)));
    layer4_outputs(172) <= (layer3_outputs(1720)) and not (layer3_outputs(1748));
    layer4_outputs(173) <= not((layer3_outputs(1143)) or (layer3_outputs(322)));
    layer4_outputs(174) <= not(layer3_outputs(946)) or (layer3_outputs(2477));
    layer4_outputs(175) <= layer3_outputs(2465);
    layer4_outputs(176) <= not((layer3_outputs(2492)) xor (layer3_outputs(988)));
    layer4_outputs(177) <= (layer3_outputs(2100)) xor (layer3_outputs(1562));
    layer4_outputs(178) <= not((layer3_outputs(1878)) xor (layer3_outputs(1813)));
    layer4_outputs(179) <= (layer3_outputs(1595)) and (layer3_outputs(1069));
    layer4_outputs(180) <= not((layer3_outputs(1367)) or (layer3_outputs(109)));
    layer4_outputs(181) <= layer3_outputs(380);
    layer4_outputs(182) <= not(layer3_outputs(947));
    layer4_outputs(183) <= (layer3_outputs(221)) and not (layer3_outputs(839));
    layer4_outputs(184) <= layer3_outputs(2373);
    layer4_outputs(185) <= layer3_outputs(333);
    layer4_outputs(186) <= not((layer3_outputs(1447)) xor (layer3_outputs(1421)));
    layer4_outputs(187) <= not(layer3_outputs(1379));
    layer4_outputs(188) <= (layer3_outputs(2187)) and (layer3_outputs(150));
    layer4_outputs(189) <= (layer3_outputs(1650)) and not (layer3_outputs(2165));
    layer4_outputs(190) <= layer3_outputs(2137);
    layer4_outputs(191) <= (layer3_outputs(709)) and (layer3_outputs(260));
    layer4_outputs(192) <= layer3_outputs(1576);
    layer4_outputs(193) <= (layer3_outputs(2157)) or (layer3_outputs(532));
    layer4_outputs(194) <= not(layer3_outputs(1470));
    layer4_outputs(195) <= layer3_outputs(1257);
    layer4_outputs(196) <= layer3_outputs(2310);
    layer4_outputs(197) <= layer3_outputs(1242);
    layer4_outputs(198) <= layer3_outputs(1804);
    layer4_outputs(199) <= not(layer3_outputs(1578));
    layer4_outputs(200) <= not(layer3_outputs(1037));
    layer4_outputs(201) <= not(layer3_outputs(2065)) or (layer3_outputs(1091));
    layer4_outputs(202) <= layer3_outputs(227);
    layer4_outputs(203) <= '1';
    layer4_outputs(204) <= layer3_outputs(197);
    layer4_outputs(205) <= (layer3_outputs(414)) xor (layer3_outputs(1228));
    layer4_outputs(206) <= layer3_outputs(415);
    layer4_outputs(207) <= not(layer3_outputs(2495));
    layer4_outputs(208) <= not((layer3_outputs(1928)) xor (layer3_outputs(202)));
    layer4_outputs(209) <= (layer3_outputs(855)) and not (layer3_outputs(1752));
    layer4_outputs(210) <= not(layer3_outputs(2068));
    layer4_outputs(211) <= (layer3_outputs(270)) and not (layer3_outputs(1816));
    layer4_outputs(212) <= (layer3_outputs(717)) xor (layer3_outputs(1725));
    layer4_outputs(213) <= not((layer3_outputs(129)) and (layer3_outputs(1142)));
    layer4_outputs(214) <= layer3_outputs(1078);
    layer4_outputs(215) <= layer3_outputs(807);
    layer4_outputs(216) <= (layer3_outputs(729)) and not (layer3_outputs(1161));
    layer4_outputs(217) <= layer3_outputs(2186);
    layer4_outputs(218) <= not((layer3_outputs(317)) and (layer3_outputs(971)));
    layer4_outputs(219) <= not(layer3_outputs(222));
    layer4_outputs(220) <= (layer3_outputs(401)) xor (layer3_outputs(282));
    layer4_outputs(221) <= not(layer3_outputs(1685));
    layer4_outputs(222) <= (layer3_outputs(2122)) and not (layer3_outputs(766));
    layer4_outputs(223) <= (layer3_outputs(293)) or (layer3_outputs(124));
    layer4_outputs(224) <= not(layer3_outputs(1165));
    layer4_outputs(225) <= layer3_outputs(2049);
    layer4_outputs(226) <= not(layer3_outputs(62));
    layer4_outputs(227) <= layer3_outputs(208);
    layer4_outputs(228) <= (layer3_outputs(5)) or (layer3_outputs(2512));
    layer4_outputs(229) <= not((layer3_outputs(864)) or (layer3_outputs(1836)));
    layer4_outputs(230) <= (layer3_outputs(673)) and not (layer3_outputs(2334));
    layer4_outputs(231) <= not(layer3_outputs(110)) or (layer3_outputs(1693));
    layer4_outputs(232) <= (layer3_outputs(1230)) and (layer3_outputs(2369));
    layer4_outputs(233) <= not(layer3_outputs(684));
    layer4_outputs(234) <= not(layer3_outputs(1592));
    layer4_outputs(235) <= not((layer3_outputs(1438)) or (layer3_outputs(1261)));
    layer4_outputs(236) <= not(layer3_outputs(2021)) or (layer3_outputs(1736));
    layer4_outputs(237) <= not(layer3_outputs(797));
    layer4_outputs(238) <= (layer3_outputs(2555)) and (layer3_outputs(1526));
    layer4_outputs(239) <= not((layer3_outputs(2073)) and (layer3_outputs(1430)));
    layer4_outputs(240) <= not(layer3_outputs(2133)) or (layer3_outputs(2444));
    layer4_outputs(241) <= not(layer3_outputs(2081));
    layer4_outputs(242) <= not(layer3_outputs(56)) or (layer3_outputs(689));
    layer4_outputs(243) <= layer3_outputs(1200);
    layer4_outputs(244) <= layer3_outputs(1563);
    layer4_outputs(245) <= not(layer3_outputs(2004)) or (layer3_outputs(1815));
    layer4_outputs(246) <= (layer3_outputs(87)) xor (layer3_outputs(1456));
    layer4_outputs(247) <= not(layer3_outputs(1940));
    layer4_outputs(248) <= not(layer3_outputs(494));
    layer4_outputs(249) <= layer3_outputs(2059);
    layer4_outputs(250) <= not(layer3_outputs(211));
    layer4_outputs(251) <= not(layer3_outputs(1985));
    layer4_outputs(252) <= '1';
    layer4_outputs(253) <= not(layer3_outputs(1101)) or (layer3_outputs(1782));
    layer4_outputs(254) <= not(layer3_outputs(1208));
    layer4_outputs(255) <= not(layer3_outputs(619));
    layer4_outputs(256) <= layer3_outputs(148);
    layer4_outputs(257) <= (layer3_outputs(847)) and (layer3_outputs(1014));
    layer4_outputs(258) <= (layer3_outputs(649)) or (layer3_outputs(439));
    layer4_outputs(259) <= not(layer3_outputs(1981));
    layer4_outputs(260) <= not(layer3_outputs(1448));
    layer4_outputs(261) <= not(layer3_outputs(61)) or (layer3_outputs(2216));
    layer4_outputs(262) <= (layer3_outputs(283)) xor (layer3_outputs(291));
    layer4_outputs(263) <= not(layer3_outputs(2337));
    layer4_outputs(264) <= not(layer3_outputs(1774)) or (layer3_outputs(1087));
    layer4_outputs(265) <= not((layer3_outputs(1350)) xor (layer3_outputs(1993)));
    layer4_outputs(266) <= (layer3_outputs(1888)) xor (layer3_outputs(993));
    layer4_outputs(267) <= not(layer3_outputs(2114)) or (layer3_outputs(179));
    layer4_outputs(268) <= (layer3_outputs(1958)) and not (layer3_outputs(1683));
    layer4_outputs(269) <= not(layer3_outputs(1461));
    layer4_outputs(270) <= not(layer3_outputs(2378)) or (layer3_outputs(1372));
    layer4_outputs(271) <= layer3_outputs(2475);
    layer4_outputs(272) <= not(layer3_outputs(1444)) or (layer3_outputs(670));
    layer4_outputs(273) <= (layer3_outputs(970)) and not (layer3_outputs(2090));
    layer4_outputs(274) <= layer3_outputs(445);
    layer4_outputs(275) <= (layer3_outputs(1412)) and (layer3_outputs(1971));
    layer4_outputs(276) <= layer3_outputs(9);
    layer4_outputs(277) <= not(layer3_outputs(1950)) or (layer3_outputs(944));
    layer4_outputs(278) <= '0';
    layer4_outputs(279) <= layer3_outputs(2145);
    layer4_outputs(280) <= layer3_outputs(1846);
    layer4_outputs(281) <= not(layer3_outputs(2355));
    layer4_outputs(282) <= not(layer3_outputs(197));
    layer4_outputs(283) <= (layer3_outputs(1792)) and not (layer3_outputs(851));
    layer4_outputs(284) <= (layer3_outputs(2226)) xor (layer3_outputs(1355));
    layer4_outputs(285) <= not(layer3_outputs(2539));
    layer4_outputs(286) <= not(layer3_outputs(877));
    layer4_outputs(287) <= layer3_outputs(38);
    layer4_outputs(288) <= (layer3_outputs(514)) and not (layer3_outputs(2018));
    layer4_outputs(289) <= not(layer3_outputs(551));
    layer4_outputs(290) <= (layer3_outputs(2543)) xor (layer3_outputs(434));
    layer4_outputs(291) <= (layer3_outputs(751)) or (layer3_outputs(2279));
    layer4_outputs(292) <= layer3_outputs(1790);
    layer4_outputs(293) <= not(layer3_outputs(1994));
    layer4_outputs(294) <= (layer3_outputs(1191)) and (layer3_outputs(1845));
    layer4_outputs(295) <= not((layer3_outputs(2027)) and (layer3_outputs(788)));
    layer4_outputs(296) <= not(layer3_outputs(1316));
    layer4_outputs(297) <= layer3_outputs(688);
    layer4_outputs(298) <= not(layer3_outputs(1840)) or (layer3_outputs(933));
    layer4_outputs(299) <= layer3_outputs(1000);
    layer4_outputs(300) <= (layer3_outputs(408)) and (layer3_outputs(1493));
    layer4_outputs(301) <= '1';
    layer4_outputs(302) <= not(layer3_outputs(2130)) or (layer3_outputs(1647));
    layer4_outputs(303) <= not(layer3_outputs(1921));
    layer4_outputs(304) <= layer3_outputs(274);
    layer4_outputs(305) <= layer3_outputs(1388);
    layer4_outputs(306) <= layer3_outputs(844);
    layer4_outputs(307) <= (layer3_outputs(1743)) and not (layer3_outputs(2425));
    layer4_outputs(308) <= not(layer3_outputs(1315));
    layer4_outputs(309) <= (layer3_outputs(1886)) xor (layer3_outputs(191));
    layer4_outputs(310) <= layer3_outputs(804);
    layer4_outputs(311) <= layer3_outputs(171);
    layer4_outputs(312) <= layer3_outputs(1596);
    layer4_outputs(313) <= not((layer3_outputs(2459)) or (layer3_outputs(1858)));
    layer4_outputs(314) <= (layer3_outputs(1709)) and not (layer3_outputs(1041));
    layer4_outputs(315) <= not(layer3_outputs(235));
    layer4_outputs(316) <= (layer3_outputs(422)) xor (layer3_outputs(1891));
    layer4_outputs(317) <= not(layer3_outputs(2446));
    layer4_outputs(318) <= not(layer3_outputs(1800));
    layer4_outputs(319) <= layer3_outputs(1307);
    layer4_outputs(320) <= not(layer3_outputs(2284));
    layer4_outputs(321) <= layer3_outputs(961);
    layer4_outputs(322) <= layer3_outputs(1262);
    layer4_outputs(323) <= layer3_outputs(2223);
    layer4_outputs(324) <= layer3_outputs(1976);
    layer4_outputs(325) <= not((layer3_outputs(800)) or (layer3_outputs(1537)));
    layer4_outputs(326) <= not(layer3_outputs(1490)) or (layer3_outputs(2538));
    layer4_outputs(327) <= not(layer3_outputs(871)) or (layer3_outputs(1215));
    layer4_outputs(328) <= not((layer3_outputs(2038)) or (layer3_outputs(903)));
    layer4_outputs(329) <= not((layer3_outputs(1095)) or (layer3_outputs(918)));
    layer4_outputs(330) <= layer3_outputs(2281);
    layer4_outputs(331) <= (layer3_outputs(1616)) and (layer3_outputs(546));
    layer4_outputs(332) <= (layer3_outputs(868)) xor (layer3_outputs(829));
    layer4_outputs(333) <= layer3_outputs(24);
    layer4_outputs(334) <= not((layer3_outputs(2226)) and (layer3_outputs(2229)));
    layer4_outputs(335) <= (layer3_outputs(1129)) and (layer3_outputs(436));
    layer4_outputs(336) <= not((layer3_outputs(2265)) xor (layer3_outputs(1531)));
    layer4_outputs(337) <= (layer3_outputs(1192)) and not (layer3_outputs(1418));
    layer4_outputs(338) <= layer3_outputs(1131);
    layer4_outputs(339) <= (layer3_outputs(1093)) xor (layer3_outputs(2153));
    layer4_outputs(340) <= layer3_outputs(830);
    layer4_outputs(341) <= layer3_outputs(665);
    layer4_outputs(342) <= not(layer3_outputs(1838));
    layer4_outputs(343) <= (layer3_outputs(663)) and not (layer3_outputs(1733));
    layer4_outputs(344) <= not(layer3_outputs(7));
    layer4_outputs(345) <= not(layer3_outputs(1224));
    layer4_outputs(346) <= (layer3_outputs(2478)) xor (layer3_outputs(2151));
    layer4_outputs(347) <= not((layer3_outputs(492)) or (layer3_outputs(2105)));
    layer4_outputs(348) <= not(layer3_outputs(2245)) or (layer3_outputs(1805));
    layer4_outputs(349) <= layer3_outputs(756);
    layer4_outputs(350) <= layer3_outputs(1955);
    layer4_outputs(351) <= not(layer3_outputs(1681));
    layer4_outputs(352) <= layer3_outputs(1668);
    layer4_outputs(353) <= layer3_outputs(2434);
    layer4_outputs(354) <= (layer3_outputs(1084)) or (layer3_outputs(455));
    layer4_outputs(355) <= layer3_outputs(168);
    layer4_outputs(356) <= not(layer3_outputs(2440));
    layer4_outputs(357) <= not(layer3_outputs(750));
    layer4_outputs(358) <= (layer3_outputs(1422)) or (layer3_outputs(2003));
    layer4_outputs(359) <= not(layer3_outputs(916));
    layer4_outputs(360) <= (layer3_outputs(1151)) and (layer3_outputs(732));
    layer4_outputs(361) <= (layer3_outputs(1969)) xor (layer3_outputs(1897));
    layer4_outputs(362) <= not((layer3_outputs(927)) xor (layer3_outputs(2056)));
    layer4_outputs(363) <= not((layer3_outputs(1708)) or (layer3_outputs(1525)));
    layer4_outputs(364) <= not(layer3_outputs(1454)) or (layer3_outputs(1539));
    layer4_outputs(365) <= not((layer3_outputs(226)) or (layer3_outputs(460)));
    layer4_outputs(366) <= layer3_outputs(1821);
    layer4_outputs(367) <= (layer3_outputs(2426)) or (layer3_outputs(1637));
    layer4_outputs(368) <= not((layer3_outputs(2362)) xor (layer3_outputs(2514)));
    layer4_outputs(369) <= layer3_outputs(667);
    layer4_outputs(370) <= not(layer3_outputs(1011)) or (layer3_outputs(606));
    layer4_outputs(371) <= (layer3_outputs(2211)) and not (layer3_outputs(2171));
    layer4_outputs(372) <= (layer3_outputs(83)) and not (layer3_outputs(1576));
    layer4_outputs(373) <= not(layer3_outputs(1212)) or (layer3_outputs(1252));
    layer4_outputs(374) <= not((layer3_outputs(599)) and (layer3_outputs(1624)));
    layer4_outputs(375) <= layer3_outputs(1437);
    layer4_outputs(376) <= (layer3_outputs(2051)) xor (layer3_outputs(2497));
    layer4_outputs(377) <= not(layer3_outputs(2423));
    layer4_outputs(378) <= (layer3_outputs(845)) xor (layer3_outputs(1496));
    layer4_outputs(379) <= not(layer3_outputs(2361));
    layer4_outputs(380) <= not((layer3_outputs(981)) or (layer3_outputs(1253)));
    layer4_outputs(381) <= (layer3_outputs(484)) and not (layer3_outputs(1786));
    layer4_outputs(382) <= not(layer3_outputs(676)) or (layer3_outputs(1832));
    layer4_outputs(383) <= layer3_outputs(2165);
    layer4_outputs(384) <= not(layer3_outputs(2534));
    layer4_outputs(385) <= not(layer3_outputs(1215));
    layer4_outputs(386) <= not(layer3_outputs(644));
    layer4_outputs(387) <= not(layer3_outputs(429));
    layer4_outputs(388) <= (layer3_outputs(2012)) and (layer3_outputs(2058));
    layer4_outputs(389) <= layer3_outputs(1397);
    layer4_outputs(390) <= not((layer3_outputs(943)) xor (layer3_outputs(857)));
    layer4_outputs(391) <= (layer3_outputs(1117)) and not (layer3_outputs(207));
    layer4_outputs(392) <= not(layer3_outputs(1051));
    layer4_outputs(393) <= layer3_outputs(2053);
    layer4_outputs(394) <= (layer3_outputs(2530)) and not (layer3_outputs(1676));
    layer4_outputs(395) <= layer3_outputs(2425);
    layer4_outputs(396) <= not((layer3_outputs(946)) or (layer3_outputs(872)));
    layer4_outputs(397) <= layer3_outputs(1464);
    layer4_outputs(398) <= layer3_outputs(2078);
    layer4_outputs(399) <= not((layer3_outputs(1390)) or (layer3_outputs(1054)));
    layer4_outputs(400) <= not(layer3_outputs(1574));
    layer4_outputs(401) <= not(layer3_outputs(499));
    layer4_outputs(402) <= layer3_outputs(709);
    layer4_outputs(403) <= not(layer3_outputs(1784)) or (layer3_outputs(1764));
    layer4_outputs(404) <= layer3_outputs(2377);
    layer4_outputs(405) <= not(layer3_outputs(1758)) or (layer3_outputs(2418));
    layer4_outputs(406) <= not((layer3_outputs(627)) and (layer3_outputs(583)));
    layer4_outputs(407) <= not(layer3_outputs(1400)) or (layer3_outputs(1811));
    layer4_outputs(408) <= not(layer3_outputs(2220)) or (layer3_outputs(1954));
    layer4_outputs(409) <= layer3_outputs(2303);
    layer4_outputs(410) <= layer3_outputs(40);
    layer4_outputs(411) <= layer3_outputs(189);
    layer4_outputs(412) <= layer3_outputs(2554);
    layer4_outputs(413) <= (layer3_outputs(696)) and not (layer3_outputs(795));
    layer4_outputs(414) <= not(layer3_outputs(254));
    layer4_outputs(415) <= layer3_outputs(1283);
    layer4_outputs(416) <= not(layer3_outputs(1446));
    layer4_outputs(417) <= layer3_outputs(1510);
    layer4_outputs(418) <= (layer3_outputs(1285)) and not (layer3_outputs(980));
    layer4_outputs(419) <= not(layer3_outputs(639));
    layer4_outputs(420) <= (layer3_outputs(1465)) and not (layer3_outputs(1167));
    layer4_outputs(421) <= not(layer3_outputs(2392)) or (layer3_outputs(1257));
    layer4_outputs(422) <= not((layer3_outputs(2134)) and (layer3_outputs(2244)));
    layer4_outputs(423) <= (layer3_outputs(419)) and not (layer3_outputs(915));
    layer4_outputs(424) <= layer3_outputs(957);
    layer4_outputs(425) <= layer3_outputs(2235);
    layer4_outputs(426) <= not(layer3_outputs(1476));
    layer4_outputs(427) <= layer3_outputs(1436);
    layer4_outputs(428) <= not(layer3_outputs(2066));
    layer4_outputs(429) <= not((layer3_outputs(222)) or (layer3_outputs(972)));
    layer4_outputs(430) <= not(layer3_outputs(2230));
    layer4_outputs(431) <= not(layer3_outputs(2509)) or (layer3_outputs(615));
    layer4_outputs(432) <= layer3_outputs(1189);
    layer4_outputs(433) <= not((layer3_outputs(612)) or (layer3_outputs(2122)));
    layer4_outputs(434) <= not((layer3_outputs(2278)) xor (layer3_outputs(1806)));
    layer4_outputs(435) <= (layer3_outputs(836)) and not (layer3_outputs(1930));
    layer4_outputs(436) <= not(layer3_outputs(1225)) or (layer3_outputs(874));
    layer4_outputs(437) <= layer3_outputs(964);
    layer4_outputs(438) <= layer3_outputs(2507);
    layer4_outputs(439) <= layer3_outputs(693);
    layer4_outputs(440) <= (layer3_outputs(266)) and not (layer3_outputs(2493));
    layer4_outputs(441) <= not(layer3_outputs(458));
    layer4_outputs(442) <= not(layer3_outputs(1782));
    layer4_outputs(443) <= not(layer3_outputs(438));
    layer4_outputs(444) <= layer3_outputs(1850);
    layer4_outputs(445) <= not((layer3_outputs(1050)) and (layer3_outputs(1632)));
    layer4_outputs(446) <= not(layer3_outputs(2379));
    layer4_outputs(447) <= not(layer3_outputs(216));
    layer4_outputs(448) <= layer3_outputs(99);
    layer4_outputs(449) <= not(layer3_outputs(1482));
    layer4_outputs(450) <= layer3_outputs(2511);
    layer4_outputs(451) <= '1';
    layer4_outputs(452) <= (layer3_outputs(1345)) and not (layer3_outputs(160));
    layer4_outputs(453) <= layer3_outputs(573);
    layer4_outputs(454) <= not(layer3_outputs(2512));
    layer4_outputs(455) <= (layer3_outputs(2107)) and not (layer3_outputs(1929));
    layer4_outputs(456) <= '1';
    layer4_outputs(457) <= layer3_outputs(741);
    layer4_outputs(458) <= not((layer3_outputs(1262)) xor (layer3_outputs(2257)));
    layer4_outputs(459) <= not(layer3_outputs(449));
    layer4_outputs(460) <= (layer3_outputs(1993)) and (layer3_outputs(1712));
    layer4_outputs(461) <= not(layer3_outputs(17));
    layer4_outputs(462) <= (layer3_outputs(1724)) or (layer3_outputs(970));
    layer4_outputs(463) <= (layer3_outputs(426)) and not (layer3_outputs(65));
    layer4_outputs(464) <= layer3_outputs(1992);
    layer4_outputs(465) <= not(layer3_outputs(2030));
    layer4_outputs(466) <= not(layer3_outputs(2203));
    layer4_outputs(467) <= layer3_outputs(542);
    layer4_outputs(468) <= layer3_outputs(759);
    layer4_outputs(469) <= not(layer3_outputs(563));
    layer4_outputs(470) <= (layer3_outputs(2342)) and not (layer3_outputs(628));
    layer4_outputs(471) <= not(layer3_outputs(528));
    layer4_outputs(472) <= layer3_outputs(161);
    layer4_outputs(473) <= (layer3_outputs(1826)) and not (layer3_outputs(1414));
    layer4_outputs(474) <= not(layer3_outputs(2408)) or (layer3_outputs(2482));
    layer4_outputs(475) <= not(layer3_outputs(1684));
    layer4_outputs(476) <= not(layer3_outputs(328));
    layer4_outputs(477) <= not(layer3_outputs(810));
    layer4_outputs(478) <= layer3_outputs(1353);
    layer4_outputs(479) <= layer3_outputs(2421);
    layer4_outputs(480) <= not(layer3_outputs(2185));
    layer4_outputs(481) <= not(layer3_outputs(789));
    layer4_outputs(482) <= (layer3_outputs(1129)) and not (layer3_outputs(1361));
    layer4_outputs(483) <= not(layer3_outputs(1893));
    layer4_outputs(484) <= not(layer3_outputs(2268));
    layer4_outputs(485) <= not(layer3_outputs(2277));
    layer4_outputs(486) <= (layer3_outputs(229)) xor (layer3_outputs(973));
    layer4_outputs(487) <= not((layer3_outputs(35)) and (layer3_outputs(917)));
    layer4_outputs(488) <= layer3_outputs(2341);
    layer4_outputs(489) <= (layer3_outputs(885)) xor (layer3_outputs(1124));
    layer4_outputs(490) <= (layer3_outputs(2497)) and not (layer3_outputs(672));
    layer4_outputs(491) <= layer3_outputs(2442);
    layer4_outputs(492) <= layer3_outputs(563);
    layer4_outputs(493) <= not(layer3_outputs(1343));
    layer4_outputs(494) <= not((layer3_outputs(1619)) xor (layer3_outputs(2335)));
    layer4_outputs(495) <= layer3_outputs(8);
    layer4_outputs(496) <= layer3_outputs(1795);
    layer4_outputs(497) <= layer3_outputs(1216);
    layer4_outputs(498) <= layer3_outputs(760);
    layer4_outputs(499) <= not((layer3_outputs(975)) xor (layer3_outputs(2427)));
    layer4_outputs(500) <= (layer3_outputs(2108)) or (layer3_outputs(49));
    layer4_outputs(501) <= not(layer3_outputs(1036));
    layer4_outputs(502) <= layer3_outputs(2327);
    layer4_outputs(503) <= layer3_outputs(448);
    layer4_outputs(504) <= not((layer3_outputs(1718)) xor (layer3_outputs(622)));
    layer4_outputs(505) <= not(layer3_outputs(2206)) or (layer3_outputs(412));
    layer4_outputs(506) <= layer3_outputs(1875);
    layer4_outputs(507) <= (layer3_outputs(685)) or (layer3_outputs(1970));
    layer4_outputs(508) <= layer3_outputs(301);
    layer4_outputs(509) <= (layer3_outputs(891)) xor (layer3_outputs(1326));
    layer4_outputs(510) <= not(layer3_outputs(1978));
    layer4_outputs(511) <= layer3_outputs(1321);
    layer4_outputs(512) <= layer3_outputs(2120);
    layer4_outputs(513) <= not(layer3_outputs(1133));
    layer4_outputs(514) <= layer3_outputs(577);
    layer4_outputs(515) <= layer3_outputs(2408);
    layer4_outputs(516) <= not(layer3_outputs(1997));
    layer4_outputs(517) <= layer3_outputs(1515);
    layer4_outputs(518) <= (layer3_outputs(1465)) and not (layer3_outputs(2443));
    layer4_outputs(519) <= not(layer3_outputs(748));
    layer4_outputs(520) <= '1';
    layer4_outputs(521) <= layer3_outputs(294);
    layer4_outputs(522) <= layer3_outputs(1780);
    layer4_outputs(523) <= not(layer3_outputs(2214));
    layer4_outputs(524) <= not(layer3_outputs(589));
    layer4_outputs(525) <= layer3_outputs(1898);
    layer4_outputs(526) <= layer3_outputs(730);
    layer4_outputs(527) <= not(layer3_outputs(2146));
    layer4_outputs(528) <= not((layer3_outputs(2180)) or (layer3_outputs(454)));
    layer4_outputs(529) <= not(layer3_outputs(1340)) or (layer3_outputs(1818));
    layer4_outputs(530) <= not(layer3_outputs(1488));
    layer4_outputs(531) <= (layer3_outputs(1453)) and not (layer3_outputs(1471));
    layer4_outputs(532) <= '1';
    layer4_outputs(533) <= (layer3_outputs(1096)) xor (layer3_outputs(436));
    layer4_outputs(534) <= layer3_outputs(1562);
    layer4_outputs(535) <= not(layer3_outputs(189));
    layer4_outputs(536) <= layer3_outputs(1356);
    layer4_outputs(537) <= (layer3_outputs(2450)) or (layer3_outputs(1263));
    layer4_outputs(538) <= layer3_outputs(866);
    layer4_outputs(539) <= not(layer3_outputs(1199));
    layer4_outputs(540) <= (layer3_outputs(482)) and not (layer3_outputs(1196));
    layer4_outputs(541) <= not((layer3_outputs(2245)) xor (layer3_outputs(906)));
    layer4_outputs(542) <= not((layer3_outputs(1349)) or (layer3_outputs(747)));
    layer4_outputs(543) <= layer3_outputs(1512);
    layer4_outputs(544) <= not(layer3_outputs(237));
    layer4_outputs(545) <= not(layer3_outputs(1681));
    layer4_outputs(546) <= not(layer3_outputs(1679));
    layer4_outputs(547) <= layer3_outputs(2421);
    layer4_outputs(548) <= not(layer3_outputs(737));
    layer4_outputs(549) <= not(layer3_outputs(1691));
    layer4_outputs(550) <= not(layer3_outputs(472));
    layer4_outputs(551) <= not(layer3_outputs(1182));
    layer4_outputs(552) <= not(layer3_outputs(1045));
    layer4_outputs(553) <= layer3_outputs(699);
    layer4_outputs(554) <= not(layer3_outputs(842));
    layer4_outputs(555) <= (layer3_outputs(1053)) or (layer3_outputs(865));
    layer4_outputs(556) <= not(layer3_outputs(990));
    layer4_outputs(557) <= not(layer3_outputs(2437));
    layer4_outputs(558) <= not(layer3_outputs(1750));
    layer4_outputs(559) <= not(layer3_outputs(357));
    layer4_outputs(560) <= (layer3_outputs(895)) or (layer3_outputs(1487));
    layer4_outputs(561) <= layer3_outputs(2247);
    layer4_outputs(562) <= not(layer3_outputs(2520)) or (layer3_outputs(1627));
    layer4_outputs(563) <= layer3_outputs(150);
    layer4_outputs(564) <= (layer3_outputs(2188)) and not (layer3_outputs(635));
    layer4_outputs(565) <= not((layer3_outputs(1797)) and (layer3_outputs(671)));
    layer4_outputs(566) <= layer3_outputs(1739);
    layer4_outputs(567) <= (layer3_outputs(809)) xor (layer3_outputs(2134));
    layer4_outputs(568) <= layer3_outputs(574);
    layer4_outputs(569) <= not(layer3_outputs(485));
    layer4_outputs(570) <= not((layer3_outputs(2375)) and (layer3_outputs(1026)));
    layer4_outputs(571) <= not(layer3_outputs(2211));
    layer4_outputs(572) <= (layer3_outputs(60)) and not (layer3_outputs(1162));
    layer4_outputs(573) <= not(layer3_outputs(1450)) or (layer3_outputs(268));
    layer4_outputs(574) <= layer3_outputs(1551);
    layer4_outputs(575) <= layer3_outputs(1760);
    layer4_outputs(576) <= not((layer3_outputs(1442)) xor (layer3_outputs(1355)));
    layer4_outputs(577) <= (layer3_outputs(1489)) and not (layer3_outputs(238));
    layer4_outputs(578) <= not(layer3_outputs(1616));
    layer4_outputs(579) <= layer3_outputs(134);
    layer4_outputs(580) <= (layer3_outputs(2422)) and (layer3_outputs(1012));
    layer4_outputs(581) <= '1';
    layer4_outputs(582) <= not(layer3_outputs(2062));
    layer4_outputs(583) <= layer3_outputs(1888);
    layer4_outputs(584) <= not(layer3_outputs(687));
    layer4_outputs(585) <= (layer3_outputs(2544)) and not (layer3_outputs(496));
    layer4_outputs(586) <= (layer3_outputs(1322)) and (layer3_outputs(1455));
    layer4_outputs(587) <= not((layer3_outputs(663)) or (layer3_outputs(1320)));
    layer4_outputs(588) <= not(layer3_outputs(126));
    layer4_outputs(589) <= layer3_outputs(1672);
    layer4_outputs(590) <= layer3_outputs(1879);
    layer4_outputs(591) <= '1';
    layer4_outputs(592) <= (layer3_outputs(441)) and not (layer3_outputs(1845));
    layer4_outputs(593) <= not(layer3_outputs(1081));
    layer4_outputs(594) <= (layer3_outputs(2041)) xor (layer3_outputs(600));
    layer4_outputs(595) <= not(layer3_outputs(2234));
    layer4_outputs(596) <= layer3_outputs(1890);
    layer4_outputs(597) <= not((layer3_outputs(1199)) and (layer3_outputs(2210)));
    layer4_outputs(598) <= (layer3_outputs(473)) or (layer3_outputs(134));
    layer4_outputs(599) <= layer3_outputs(266);
    layer4_outputs(600) <= (layer3_outputs(572)) or (layer3_outputs(735));
    layer4_outputs(601) <= (layer3_outputs(1488)) and (layer3_outputs(1942));
    layer4_outputs(602) <= not((layer3_outputs(751)) and (layer3_outputs(713)));
    layer4_outputs(603) <= not((layer3_outputs(165)) xor (layer3_outputs(1305)));
    layer4_outputs(604) <= (layer3_outputs(492)) or (layer3_outputs(320));
    layer4_outputs(605) <= (layer3_outputs(2124)) and (layer3_outputs(1813));
    layer4_outputs(606) <= not(layer3_outputs(1394)) or (layer3_outputs(1878));
    layer4_outputs(607) <= not(layer3_outputs(2205));
    layer4_outputs(608) <= layer3_outputs(816);
    layer4_outputs(609) <= not(layer3_outputs(86));
    layer4_outputs(610) <= not(layer3_outputs(2494));
    layer4_outputs(611) <= not(layer3_outputs(2209));
    layer4_outputs(612) <= not(layer3_outputs(1531));
    layer4_outputs(613) <= (layer3_outputs(951)) or (layer3_outputs(781));
    layer4_outputs(614) <= not(layer3_outputs(1072)) or (layer3_outputs(1723));
    layer4_outputs(615) <= layer3_outputs(1754);
    layer4_outputs(616) <= not((layer3_outputs(2181)) xor (layer3_outputs(2110)));
    layer4_outputs(617) <= '0';
    layer4_outputs(618) <= not(layer3_outputs(239));
    layer4_outputs(619) <= (layer3_outputs(1364)) and (layer3_outputs(2181));
    layer4_outputs(620) <= not(layer3_outputs(2213)) or (layer3_outputs(1264));
    layer4_outputs(621) <= layer3_outputs(1559);
    layer4_outputs(622) <= layer3_outputs(1198);
    layer4_outputs(623) <= layer3_outputs(2190);
    layer4_outputs(624) <= layer3_outputs(865);
    layer4_outputs(625) <= not(layer3_outputs(2191));
    layer4_outputs(626) <= not((layer3_outputs(157)) or (layer3_outputs(1899)));
    layer4_outputs(627) <= not(layer3_outputs(560));
    layer4_outputs(628) <= not(layer3_outputs(1550));
    layer4_outputs(629) <= (layer3_outputs(2363)) and not (layer3_outputs(909));
    layer4_outputs(630) <= not((layer3_outputs(2302)) and (layer3_outputs(2037)));
    layer4_outputs(631) <= (layer3_outputs(1718)) or (layer3_outputs(984));
    layer4_outputs(632) <= not(layer3_outputs(628)) or (layer3_outputs(1613));
    layer4_outputs(633) <= layer3_outputs(779);
    layer4_outputs(634) <= not(layer3_outputs(1380));
    layer4_outputs(635) <= not(layer3_outputs(1132));
    layer4_outputs(636) <= (layer3_outputs(824)) xor (layer3_outputs(512));
    layer4_outputs(637) <= not((layer3_outputs(1042)) or (layer3_outputs(1686)));
    layer4_outputs(638) <= layer3_outputs(2376);
    layer4_outputs(639) <= layer3_outputs(1310);
    layer4_outputs(640) <= '0';
    layer4_outputs(641) <= layer3_outputs(610);
    layer4_outputs(642) <= (layer3_outputs(1166)) and (layer3_outputs(447));
    layer4_outputs(643) <= not(layer3_outputs(2328));
    layer4_outputs(644) <= not((layer3_outputs(1998)) or (layer3_outputs(133)));
    layer4_outputs(645) <= layer3_outputs(1184);
    layer4_outputs(646) <= layer3_outputs(1452);
    layer4_outputs(647) <= (layer3_outputs(2143)) and not (layer3_outputs(522));
    layer4_outputs(648) <= (layer3_outputs(864)) and (layer3_outputs(1121));
    layer4_outputs(649) <= layer3_outputs(1104);
    layer4_outputs(650) <= not((layer3_outputs(926)) or (layer3_outputs(1097)));
    layer4_outputs(651) <= (layer3_outputs(1148)) or (layer3_outputs(1948));
    layer4_outputs(652) <= (layer3_outputs(1480)) xor (layer3_outputs(1976));
    layer4_outputs(653) <= not((layer3_outputs(2046)) xor (layer3_outputs(2249)));
    layer4_outputs(654) <= not(layer3_outputs(573)) or (layer3_outputs(450));
    layer4_outputs(655) <= (layer3_outputs(198)) and not (layer3_outputs(2516));
    layer4_outputs(656) <= layer3_outputs(439);
    layer4_outputs(657) <= not((layer3_outputs(149)) and (layer3_outputs(2299)));
    layer4_outputs(658) <= not((layer3_outputs(1272)) xor (layer3_outputs(253)));
    layer4_outputs(659) <= not((layer3_outputs(272)) and (layer3_outputs(860)));
    layer4_outputs(660) <= '1';
    layer4_outputs(661) <= (layer3_outputs(1825)) and not (layer3_outputs(1917));
    layer4_outputs(662) <= layer3_outputs(1812);
    layer4_outputs(663) <= not((layer3_outputs(1866)) xor (layer3_outputs(1386)));
    layer4_outputs(664) <= layer3_outputs(2052);
    layer4_outputs(665) <= (layer3_outputs(2057)) xor (layer3_outputs(1147));
    layer4_outputs(666) <= not(layer3_outputs(1898));
    layer4_outputs(667) <= layer3_outputs(662);
    layer4_outputs(668) <= not(layer3_outputs(2436));
    layer4_outputs(669) <= not((layer3_outputs(363)) xor (layer3_outputs(526)));
    layer4_outputs(670) <= layer3_outputs(2128);
    layer4_outputs(671) <= not(layer3_outputs(1925));
    layer4_outputs(672) <= not(layer3_outputs(2259));
    layer4_outputs(673) <= (layer3_outputs(2081)) or (layer3_outputs(510));
    layer4_outputs(674) <= layer3_outputs(79);
    layer4_outputs(675) <= (layer3_outputs(188)) xor (layer3_outputs(416));
    layer4_outputs(676) <= '1';
    layer4_outputs(677) <= (layer3_outputs(1421)) and not (layer3_outputs(1528));
    layer4_outputs(678) <= not((layer3_outputs(384)) or (layer3_outputs(124)));
    layer4_outputs(679) <= layer3_outputs(1723);
    layer4_outputs(680) <= not(layer3_outputs(1258));
    layer4_outputs(681) <= layer3_outputs(1344);
    layer4_outputs(682) <= layer3_outputs(2194);
    layer4_outputs(683) <= (layer3_outputs(670)) xor (layer3_outputs(1391));
    layer4_outputs(684) <= not(layer3_outputs(1218)) or (layer3_outputs(2208));
    layer4_outputs(685) <= not(layer3_outputs(996)) or (layer3_outputs(1780));
    layer4_outputs(686) <= not((layer3_outputs(224)) xor (layer3_outputs(2458)));
    layer4_outputs(687) <= layer3_outputs(1156);
    layer4_outputs(688) <= (layer3_outputs(2432)) and not (layer3_outputs(400));
    layer4_outputs(689) <= layer3_outputs(1947);
    layer4_outputs(690) <= layer3_outputs(1052);
    layer4_outputs(691) <= layer3_outputs(342);
    layer4_outputs(692) <= (layer3_outputs(1945)) xor (layer3_outputs(1009));
    layer4_outputs(693) <= not((layer3_outputs(535)) or (layer3_outputs(982)));
    layer4_outputs(694) <= (layer3_outputs(2224)) and (layer3_outputs(88));
    layer4_outputs(695) <= not(layer3_outputs(2531));
    layer4_outputs(696) <= not(layer3_outputs(826));
    layer4_outputs(697) <= layer3_outputs(1354);
    layer4_outputs(698) <= not(layer3_outputs(2048)) or (layer3_outputs(745));
    layer4_outputs(699) <= not((layer3_outputs(2127)) xor (layer3_outputs(481)));
    layer4_outputs(700) <= (layer3_outputs(1824)) and not (layer3_outputs(1842));
    layer4_outputs(701) <= not((layer3_outputs(2216)) and (layer3_outputs(1677)));
    layer4_outputs(702) <= not(layer3_outputs(2174));
    layer4_outputs(703) <= (layer3_outputs(2391)) and (layer3_outputs(205));
    layer4_outputs(704) <= not(layer3_outputs(2500));
    layer4_outputs(705) <= (layer3_outputs(143)) or (layer3_outputs(261));
    layer4_outputs(706) <= not(layer3_outputs(1824)) or (layer3_outputs(38));
    layer4_outputs(707) <= not(layer3_outputs(1828));
    layer4_outputs(708) <= layer3_outputs(2192);
    layer4_outputs(709) <= layer3_outputs(128);
    layer4_outputs(710) <= not((layer3_outputs(2129)) or (layer3_outputs(416)));
    layer4_outputs(711) <= not((layer3_outputs(2043)) or (layer3_outputs(142)));
    layer4_outputs(712) <= not((layer3_outputs(199)) xor (layer3_outputs(1991)));
    layer4_outputs(713) <= not(layer3_outputs(2280));
    layer4_outputs(714) <= layer3_outputs(2177);
    layer4_outputs(715) <= not((layer3_outputs(433)) and (layer3_outputs(1155)));
    layer4_outputs(716) <= (layer3_outputs(1644)) and not (layer3_outputs(1731));
    layer4_outputs(717) <= (layer3_outputs(323)) and not (layer3_outputs(757));
    layer4_outputs(718) <= not(layer3_outputs(2223));
    layer4_outputs(719) <= layer3_outputs(730);
    layer4_outputs(720) <= not(layer3_outputs(912));
    layer4_outputs(721) <= not(layer3_outputs(1365));
    layer4_outputs(722) <= not(layer3_outputs(226));
    layer4_outputs(723) <= not((layer3_outputs(2031)) and (layer3_outputs(2196)));
    layer4_outputs(724) <= layer3_outputs(2119);
    layer4_outputs(725) <= not((layer3_outputs(547)) or (layer3_outputs(1368)));
    layer4_outputs(726) <= layer3_outputs(445);
    layer4_outputs(727) <= layer3_outputs(2413);
    layer4_outputs(728) <= not((layer3_outputs(722)) and (layer3_outputs(675)));
    layer4_outputs(729) <= '0';
    layer4_outputs(730) <= (layer3_outputs(2544)) or (layer3_outputs(474));
    layer4_outputs(731) <= layer3_outputs(314);
    layer4_outputs(732) <= not(layer3_outputs(1568));
    layer4_outputs(733) <= not((layer3_outputs(1433)) or (layer3_outputs(1948)));
    layer4_outputs(734) <= not(layer3_outputs(2150)) or (layer3_outputs(1662));
    layer4_outputs(735) <= not(layer3_outputs(2043)) or (layer3_outputs(2231));
    layer4_outputs(736) <= not(layer3_outputs(1293));
    layer4_outputs(737) <= (layer3_outputs(533)) and not (layer3_outputs(746));
    layer4_outputs(738) <= layer3_outputs(141);
    layer4_outputs(739) <= (layer3_outputs(1366)) xor (layer3_outputs(2144));
    layer4_outputs(740) <= not(layer3_outputs(1546)) or (layer3_outputs(2248));
    layer4_outputs(741) <= not(layer3_outputs(1873));
    layer4_outputs(742) <= not((layer3_outputs(1558)) or (layer3_outputs(1405)));
    layer4_outputs(743) <= not(layer3_outputs(2436));
    layer4_outputs(744) <= not(layer3_outputs(756));
    layer4_outputs(745) <= layer3_outputs(432);
    layer4_outputs(746) <= layer3_outputs(1150);
    layer4_outputs(747) <= layer3_outputs(1613);
    layer4_outputs(748) <= (layer3_outputs(1379)) and not (layer3_outputs(461));
    layer4_outputs(749) <= not(layer3_outputs(867));
    layer4_outputs(750) <= not((layer3_outputs(1286)) xor (layer3_outputs(1061)));
    layer4_outputs(751) <= not(layer3_outputs(1255));
    layer4_outputs(752) <= layer3_outputs(1420);
    layer4_outputs(753) <= layer3_outputs(777);
    layer4_outputs(754) <= layer3_outputs(2351);
    layer4_outputs(755) <= not(layer3_outputs(608)) or (layer3_outputs(1908));
    layer4_outputs(756) <= (layer3_outputs(1580)) and (layer3_outputs(2272));
    layer4_outputs(757) <= layer3_outputs(1467);
    layer4_outputs(758) <= (layer3_outputs(1214)) or (layer3_outputs(749));
    layer4_outputs(759) <= not(layer3_outputs(2254));
    layer4_outputs(760) <= not(layer3_outputs(798));
    layer4_outputs(761) <= (layer3_outputs(280)) and (layer3_outputs(280));
    layer4_outputs(762) <= (layer3_outputs(1203)) or (layer3_outputs(193));
    layer4_outputs(763) <= layer3_outputs(1091);
    layer4_outputs(764) <= layer3_outputs(494);
    layer4_outputs(765) <= layer3_outputs(1593);
    layer4_outputs(766) <= not((layer3_outputs(743)) xor (layer3_outputs(695)));
    layer4_outputs(767) <= layer3_outputs(1252);
    layer4_outputs(768) <= not((layer3_outputs(713)) xor (layer3_outputs(565)));
    layer4_outputs(769) <= not(layer3_outputs(1781));
    layer4_outputs(770) <= layer3_outputs(1851);
    layer4_outputs(771) <= not((layer3_outputs(714)) xor (layer3_outputs(882)));
    layer4_outputs(772) <= not(layer3_outputs(544));
    layer4_outputs(773) <= not(layer3_outputs(82));
    layer4_outputs(774) <= (layer3_outputs(1559)) or (layer3_outputs(1198));
    layer4_outputs(775) <= (layer3_outputs(1877)) xor (layer3_outputs(1159));
    layer4_outputs(776) <= not(layer3_outputs(2307));
    layer4_outputs(777) <= not(layer3_outputs(1882));
    layer4_outputs(778) <= not((layer3_outputs(576)) xor (layer3_outputs(2205)));
    layer4_outputs(779) <= layer3_outputs(2069);
    layer4_outputs(780) <= (layer3_outputs(2220)) xor (layer3_outputs(2557));
    layer4_outputs(781) <= not(layer3_outputs(411));
    layer4_outputs(782) <= (layer3_outputs(2175)) and (layer3_outputs(271));
    layer4_outputs(783) <= layer3_outputs(252);
    layer4_outputs(784) <= (layer3_outputs(605)) xor (layer3_outputs(2001));
    layer4_outputs(785) <= (layer3_outputs(2198)) and (layer3_outputs(1341));
    layer4_outputs(786) <= layer3_outputs(1789);
    layer4_outputs(787) <= layer3_outputs(1517);
    layer4_outputs(788) <= (layer3_outputs(1552)) xor (layer3_outputs(1569));
    layer4_outputs(789) <= not((layer3_outputs(243)) or (layer3_outputs(1265)));
    layer4_outputs(790) <= '1';
    layer4_outputs(791) <= not(layer3_outputs(1065));
    layer4_outputs(792) <= not((layer3_outputs(1629)) xor (layer3_outputs(1892)));
    layer4_outputs(793) <= layer3_outputs(1116);
    layer4_outputs(794) <= layer3_outputs(620);
    layer4_outputs(795) <= not((layer3_outputs(183)) xor (layer3_outputs(368)));
    layer4_outputs(796) <= not(layer3_outputs(51));
    layer4_outputs(797) <= not(layer3_outputs(723)) or (layer3_outputs(218));
    layer4_outputs(798) <= layer3_outputs(1233);
    layer4_outputs(799) <= (layer3_outputs(575)) and not (layer3_outputs(1876));
    layer4_outputs(800) <= layer3_outputs(1035);
    layer4_outputs(801) <= layer3_outputs(71);
    layer4_outputs(802) <= layer3_outputs(1513);
    layer4_outputs(803) <= layer3_outputs(1953);
    layer4_outputs(804) <= not((layer3_outputs(642)) and (layer3_outputs(1370)));
    layer4_outputs(805) <= not((layer3_outputs(2373)) or (layer3_outputs(937)));
    layer4_outputs(806) <= (layer3_outputs(605)) and not (layer3_outputs(929));
    layer4_outputs(807) <= (layer3_outputs(2423)) xor (layer3_outputs(612));
    layer4_outputs(808) <= not(layer3_outputs(2150));
    layer4_outputs(809) <= (layer3_outputs(1498)) and not (layer3_outputs(1443));
    layer4_outputs(810) <= layer3_outputs(2301);
    layer4_outputs(811) <= (layer3_outputs(155)) and not (layer3_outputs(69));
    layer4_outputs(812) <= layer3_outputs(2333);
    layer4_outputs(813) <= layer3_outputs(2260);
    layer4_outputs(814) <= not(layer3_outputs(26));
    layer4_outputs(815) <= not(layer3_outputs(390)) or (layer3_outputs(1376));
    layer4_outputs(816) <= '0';
    layer4_outputs(817) <= not((layer3_outputs(557)) or (layer3_outputs(1496)));
    layer4_outputs(818) <= not(layer3_outputs(1136)) or (layer3_outputs(262));
    layer4_outputs(819) <= not((layer3_outputs(304)) or (layer3_outputs(1523)));
    layer4_outputs(820) <= layer3_outputs(2114);
    layer4_outputs(821) <= not((layer3_outputs(2471)) or (layer3_outputs(1143)));
    layer4_outputs(822) <= not(layer3_outputs(321));
    layer4_outputs(823) <= (layer3_outputs(486)) and not (layer3_outputs(590));
    layer4_outputs(824) <= not(layer3_outputs(446)) or (layer3_outputs(1753));
    layer4_outputs(825) <= '0';
    layer4_outputs(826) <= not(layer3_outputs(681));
    layer4_outputs(827) <= not(layer3_outputs(2453));
    layer4_outputs(828) <= not(layer3_outputs(59));
    layer4_outputs(829) <= (layer3_outputs(595)) xor (layer3_outputs(1389));
    layer4_outputs(830) <= (layer3_outputs(1425)) and not (layer3_outputs(885));
    layer4_outputs(831) <= (layer3_outputs(2155)) and (layer3_outputs(1570));
    layer4_outputs(832) <= layer3_outputs(941);
    layer4_outputs(833) <= not(layer3_outputs(326));
    layer4_outputs(834) <= not(layer3_outputs(233)) or (layer3_outputs(513));
    layer4_outputs(835) <= (layer3_outputs(1934)) and not (layer3_outputs(295));
    layer4_outputs(836) <= not((layer3_outputs(2058)) xor (layer3_outputs(1020)));
    layer4_outputs(837) <= layer3_outputs(144);
    layer4_outputs(838) <= not(layer3_outputs(2167)) or (layer3_outputs(1417));
    layer4_outputs(839) <= layer3_outputs(857);
    layer4_outputs(840) <= not(layer3_outputs(1419));
    layer4_outputs(841) <= layer3_outputs(820);
    layer4_outputs(842) <= not(layer3_outputs(417));
    layer4_outputs(843) <= not(layer3_outputs(754));
    layer4_outputs(844) <= not((layer3_outputs(2424)) or (layer3_outputs(1901)));
    layer4_outputs(845) <= not(layer3_outputs(1819));
    layer4_outputs(846) <= not(layer3_outputs(1684));
    layer4_outputs(847) <= layer3_outputs(24);
    layer4_outputs(848) <= not((layer3_outputs(1160)) and (layer3_outputs(1209)));
    layer4_outputs(849) <= layer3_outputs(2080);
    layer4_outputs(850) <= not(layer3_outputs(350)) or (layer3_outputs(1396));
    layer4_outputs(851) <= layer3_outputs(2491);
    layer4_outputs(852) <= not((layer3_outputs(108)) and (layer3_outputs(1986)));
    layer4_outputs(853) <= not(layer3_outputs(2522));
    layer4_outputs(854) <= (layer3_outputs(1333)) and (layer3_outputs(468));
    layer4_outputs(855) <= not(layer3_outputs(64)) or (layer3_outputs(96));
    layer4_outputs(856) <= not(layer3_outputs(2362));
    layer4_outputs(857) <= not(layer3_outputs(1791));
    layer4_outputs(858) <= (layer3_outputs(1063)) xor (layer3_outputs(2218));
    layer4_outputs(859) <= not(layer3_outputs(2445));
    layer4_outputs(860) <= not(layer3_outputs(1532));
    layer4_outputs(861) <= layer3_outputs(2393);
    layer4_outputs(862) <= (layer3_outputs(2348)) and not (layer3_outputs(424));
    layer4_outputs(863) <= (layer3_outputs(1949)) and not (layer3_outputs(1701));
    layer4_outputs(864) <= not(layer3_outputs(2403));
    layer4_outputs(865) <= (layer3_outputs(1362)) and (layer3_outputs(1560));
    layer4_outputs(866) <= not(layer3_outputs(1961));
    layer4_outputs(867) <= not(layer3_outputs(1413));
    layer4_outputs(868) <= layer3_outputs(2467);
    layer4_outputs(869) <= layer3_outputs(2311);
    layer4_outputs(870) <= (layer3_outputs(2424)) and not (layer3_outputs(1485));
    layer4_outputs(871) <= (layer3_outputs(1765)) and (layer3_outputs(943));
    layer4_outputs(872) <= (layer3_outputs(478)) xor (layer3_outputs(1389));
    layer4_outputs(873) <= not((layer3_outputs(2045)) xor (layer3_outputs(702)));
    layer4_outputs(874) <= not(layer3_outputs(363));
    layer4_outputs(875) <= (layer3_outputs(2222)) and not (layer3_outputs(1329));
    layer4_outputs(876) <= not(layer3_outputs(859));
    layer4_outputs(877) <= not((layer3_outputs(342)) or (layer3_outputs(735)));
    layer4_outputs(878) <= (layer3_outputs(1910)) and not (layer3_outputs(1011));
    layer4_outputs(879) <= not((layer3_outputs(100)) and (layer3_outputs(138)));
    layer4_outputs(880) <= layer3_outputs(2500);
    layer4_outputs(881) <= not(layer3_outputs(2199));
    layer4_outputs(882) <= not((layer3_outputs(708)) or (layer3_outputs(2429)));
    layer4_outputs(883) <= layer3_outputs(913);
    layer4_outputs(884) <= layer3_outputs(1522);
    layer4_outputs(885) <= not((layer3_outputs(1625)) or (layer3_outputs(777)));
    layer4_outputs(886) <= (layer3_outputs(1606)) and (layer3_outputs(111));
    layer4_outputs(887) <= not(layer3_outputs(2332));
    layer4_outputs(888) <= '1';
    layer4_outputs(889) <= not((layer3_outputs(1746)) or (layer3_outputs(1066)));
    layer4_outputs(890) <= not((layer3_outputs(968)) xor (layer3_outputs(393)));
    layer4_outputs(891) <= not(layer3_outputs(686));
    layer4_outputs(892) <= not(layer3_outputs(55));
    layer4_outputs(893) <= not(layer3_outputs(525)) or (layer3_outputs(1347));
    layer4_outputs(894) <= (layer3_outputs(1350)) xor (layer3_outputs(33));
    layer4_outputs(895) <= layer3_outputs(1394);
    layer4_outputs(896) <= not((layer3_outputs(2341)) xor (layer3_outputs(1118)));
    layer4_outputs(897) <= not(layer3_outputs(597));
    layer4_outputs(898) <= not((layer3_outputs(1182)) xor (layer3_outputs(332)));
    layer4_outputs(899) <= not(layer3_outputs(1115));
    layer4_outputs(900) <= not(layer3_outputs(750));
    layer4_outputs(901) <= not(layer3_outputs(1515));
    layer4_outputs(902) <= not(layer3_outputs(571));
    layer4_outputs(903) <= (layer3_outputs(2143)) xor (layer3_outputs(1566));
    layer4_outputs(904) <= layer3_outputs(2457);
    layer4_outputs(905) <= '1';
    layer4_outputs(906) <= (layer3_outputs(1371)) and not (layer3_outputs(1549));
    layer4_outputs(907) <= not((layer3_outputs(2309)) and (layer3_outputs(774)));
    layer4_outputs(908) <= layer3_outputs(523);
    layer4_outputs(909) <= not((layer3_outputs(1500)) or (layer3_outputs(1134)));
    layer4_outputs(910) <= (layer3_outputs(1247)) and (layer3_outputs(355));
    layer4_outputs(911) <= layer3_outputs(210);
    layer4_outputs(912) <= not(layer3_outputs(2433)) or (layer3_outputs(1990));
    layer4_outputs(913) <= not(layer3_outputs(63));
    layer4_outputs(914) <= not((layer3_outputs(690)) or (layer3_outputs(2123)));
    layer4_outputs(915) <= (layer3_outputs(2559)) xor (layer3_outputs(1999));
    layer4_outputs(916) <= not(layer3_outputs(1639));
    layer4_outputs(917) <= not(layer3_outputs(1495));
    layer4_outputs(918) <= (layer3_outputs(2012)) and not (layer3_outputs(1378));
    layer4_outputs(919) <= not((layer3_outputs(2546)) xor (layer3_outputs(1811)));
    layer4_outputs(920) <= not(layer3_outputs(2091));
    layer4_outputs(921) <= not(layer3_outputs(561));
    layer4_outputs(922) <= not(layer3_outputs(2419));
    layer4_outputs(923) <= layer3_outputs(42);
    layer4_outputs(924) <= (layer3_outputs(548)) and not (layer3_outputs(1339));
    layer4_outputs(925) <= not(layer3_outputs(121));
    layer4_outputs(926) <= not(layer3_outputs(437));
    layer4_outputs(927) <= (layer3_outputs(1665)) or (layer3_outputs(1906));
    layer4_outputs(928) <= not(layer3_outputs(2365));
    layer4_outputs(929) <= not(layer3_outputs(538));
    layer4_outputs(930) <= not(layer3_outputs(1676));
    layer4_outputs(931) <= not((layer3_outputs(982)) and (layer3_outputs(1649)));
    layer4_outputs(932) <= (layer3_outputs(1374)) or (layer3_outputs(1236));
    layer4_outputs(933) <= layer3_outputs(388);
    layer4_outputs(934) <= not(layer3_outputs(859)) or (layer3_outputs(702));
    layer4_outputs(935) <= layer3_outputs(749);
    layer4_outputs(936) <= (layer3_outputs(2286)) and not (layer3_outputs(1833));
    layer4_outputs(937) <= layer3_outputs(1322);
    layer4_outputs(938) <= not((layer3_outputs(2399)) and (layer3_outputs(889)));
    layer4_outputs(939) <= not(layer3_outputs(1426)) or (layer3_outputs(955));
    layer4_outputs(940) <= '0';
    layer4_outputs(941) <= layer3_outputs(590);
    layer4_outputs(942) <= not(layer3_outputs(1730));
    layer4_outputs(943) <= (layer3_outputs(1622)) and not (layer3_outputs(163));
    layer4_outputs(944) <= not((layer3_outputs(470)) and (layer3_outputs(111)));
    layer4_outputs(945) <= not(layer3_outputs(2357));
    layer4_outputs(946) <= '0';
    layer4_outputs(947) <= (layer3_outputs(1121)) and not (layer3_outputs(1989));
    layer4_outputs(948) <= not(layer3_outputs(2305));
    layer4_outputs(949) <= not((layer3_outputs(2354)) or (layer3_outputs(1587)));
    layer4_outputs(950) <= (layer3_outputs(2079)) or (layer3_outputs(75));
    layer4_outputs(951) <= not((layer3_outputs(2044)) or (layer3_outputs(1493)));
    layer4_outputs(952) <= '1';
    layer4_outputs(953) <= layer3_outputs(403);
    layer4_outputs(954) <= not(layer3_outputs(2490)) or (layer3_outputs(1460));
    layer4_outputs(955) <= not(layer3_outputs(922));
    layer4_outputs(956) <= not(layer3_outputs(344)) or (layer3_outputs(1735));
    layer4_outputs(957) <= not((layer3_outputs(1319)) and (layer3_outputs(1095)));
    layer4_outputs(958) <= layer3_outputs(2040);
    layer4_outputs(959) <= not(layer3_outputs(1149)) or (layer3_outputs(170));
    layer4_outputs(960) <= layer3_outputs(1602);
    layer4_outputs(961) <= not(layer3_outputs(1997));
    layer4_outputs(962) <= layer3_outputs(691);
    layer4_outputs(963) <= (layer3_outputs(450)) or (layer3_outputs(1342));
    layer4_outputs(964) <= not(layer3_outputs(57));
    layer4_outputs(965) <= (layer3_outputs(905)) and not (layer3_outputs(848));
    layer4_outputs(966) <= not((layer3_outputs(1028)) xor (layer3_outputs(1035)));
    layer4_outputs(967) <= layer3_outputs(572);
    layer4_outputs(968) <= not((layer3_outputs(1411)) and (layer3_outputs(1096)));
    layer4_outputs(969) <= not((layer3_outputs(2517)) and (layer3_outputs(2414)));
    layer4_outputs(970) <= not((layer3_outputs(131)) and (layer3_outputs(166)));
    layer4_outputs(971) <= layer3_outputs(41);
    layer4_outputs(972) <= (layer3_outputs(167)) or (layer3_outputs(986));
    layer4_outputs(973) <= layer3_outputs(2003);
    layer4_outputs(974) <= not((layer3_outputs(468)) and (layer3_outputs(58)));
    layer4_outputs(975) <= not(layer3_outputs(173));
    layer4_outputs(976) <= layer3_outputs(1696);
    layer4_outputs(977) <= layer3_outputs(1959);
    layer4_outputs(978) <= '0';
    layer4_outputs(979) <= (layer3_outputs(1775)) and not (layer3_outputs(1186));
    layer4_outputs(980) <= not(layer3_outputs(1572)) or (layer3_outputs(1757));
    layer4_outputs(981) <= not((layer3_outputs(296)) xor (layer3_outputs(2480)));
    layer4_outputs(982) <= layer3_outputs(2498);
    layer4_outputs(983) <= '1';
    layer4_outputs(984) <= layer3_outputs(596);
    layer4_outputs(985) <= not(layer3_outputs(762));
    layer4_outputs(986) <= not((layer3_outputs(1348)) or (layer3_outputs(159)));
    layer4_outputs(987) <= (layer3_outputs(1666)) xor (layer3_outputs(1534));
    layer4_outputs(988) <= not(layer3_outputs(1569));
    layer4_outputs(989) <= '0';
    layer4_outputs(990) <= not((layer3_outputs(409)) xor (layer3_outputs(2537)));
    layer4_outputs(991) <= not((layer3_outputs(2338)) and (layer3_outputs(508)));
    layer4_outputs(992) <= not(layer3_outputs(1049));
    layer4_outputs(993) <= not(layer3_outputs(1929));
    layer4_outputs(994) <= (layer3_outputs(2328)) xor (layer3_outputs(1127));
    layer4_outputs(995) <= not(layer3_outputs(1391));
    layer4_outputs(996) <= (layer3_outputs(2402)) or (layer3_outputs(2394));
    layer4_outputs(997) <= layer3_outputs(707);
    layer4_outputs(998) <= (layer3_outputs(2526)) and (layer3_outputs(902));
    layer4_outputs(999) <= not(layer3_outputs(116)) or (layer3_outputs(853));
    layer4_outputs(1000) <= not(layer3_outputs(1561)) or (layer3_outputs(22));
    layer4_outputs(1001) <= not(layer3_outputs(2293));
    layer4_outputs(1002) <= (layer3_outputs(1092)) and not (layer3_outputs(366));
    layer4_outputs(1003) <= (layer3_outputs(1909)) and not (layer3_outputs(1237));
    layer4_outputs(1004) <= not(layer3_outputs(2457));
    layer4_outputs(1005) <= not((layer3_outputs(1453)) and (layer3_outputs(1538)));
    layer4_outputs(1006) <= (layer3_outputs(501)) and not (layer3_outputs(1303));
    layer4_outputs(1007) <= layer3_outputs(119);
    layer4_outputs(1008) <= (layer3_outputs(2087)) xor (layer3_outputs(2448));
    layer4_outputs(1009) <= (layer3_outputs(1235)) and not (layer3_outputs(2536));
    layer4_outputs(1010) <= not((layer3_outputs(2399)) xor (layer3_outputs(1834)));
    layer4_outputs(1011) <= layer3_outputs(30);
    layer4_outputs(1012) <= layer3_outputs(616);
    layer4_outputs(1013) <= (layer3_outputs(59)) xor (layer3_outputs(1874));
    layer4_outputs(1014) <= not(layer3_outputs(211));
    layer4_outputs(1015) <= not(layer3_outputs(587));
    layer4_outputs(1016) <= (layer3_outputs(2519)) and (layer3_outputs(1341));
    layer4_outputs(1017) <= not(layer3_outputs(387));
    layer4_outputs(1018) <= (layer3_outputs(1575)) and not (layer3_outputs(983));
    layer4_outputs(1019) <= layer3_outputs(103);
    layer4_outputs(1020) <= layer3_outputs(1671);
    layer4_outputs(1021) <= not(layer3_outputs(2267));
    layer4_outputs(1022) <= '0';
    layer4_outputs(1023) <= layer3_outputs(1188);
    layer4_outputs(1024) <= (layer3_outputs(357)) xor (layer3_outputs(910));
    layer4_outputs(1025) <= layer3_outputs(104);
    layer4_outputs(1026) <= (layer3_outputs(2052)) and (layer3_outputs(1699));
    layer4_outputs(1027) <= (layer3_outputs(681)) xor (layer3_outputs(1429));
    layer4_outputs(1028) <= not(layer3_outputs(1861));
    layer4_outputs(1029) <= not((layer3_outputs(2468)) xor (layer3_outputs(666)));
    layer4_outputs(1030) <= (layer3_outputs(930)) and not (layer3_outputs(2161));
    layer4_outputs(1031) <= not((layer3_outputs(314)) and (layer3_outputs(1895)));
    layer4_outputs(1032) <= not(layer3_outputs(1979));
    layer4_outputs(1033) <= not((layer3_outputs(1273)) and (layer3_outputs(1281)));
    layer4_outputs(1034) <= layer3_outputs(377);
    layer4_outputs(1035) <= not(layer3_outputs(2319));
    layer4_outputs(1036) <= not(layer3_outputs(1808));
    layer4_outputs(1037) <= not(layer3_outputs(215));
    layer4_outputs(1038) <= not((layer3_outputs(110)) and (layer3_outputs(1525)));
    layer4_outputs(1039) <= not(layer3_outputs(2030));
    layer4_outputs(1040) <= layer3_outputs(655);
    layer4_outputs(1041) <= (layer3_outputs(359)) xor (layer3_outputs(940));
    layer4_outputs(1042) <= (layer3_outputs(525)) and not (layer3_outputs(888));
    layer4_outputs(1043) <= layer3_outputs(127);
    layer4_outputs(1044) <= not(layer3_outputs(427));
    layer4_outputs(1045) <= layer3_outputs(2252);
    layer4_outputs(1046) <= not(layer3_outputs(539));
    layer4_outputs(1047) <= not(layer3_outputs(1709)) or (layer3_outputs(980));
    layer4_outputs(1048) <= not(layer3_outputs(978));
    layer4_outputs(1049) <= (layer3_outputs(2100)) and not (layer3_outputs(2229));
    layer4_outputs(1050) <= (layer3_outputs(2339)) and not (layer3_outputs(2338));
    layer4_outputs(1051) <= layer3_outputs(827);
    layer4_outputs(1052) <= not((layer3_outputs(904)) xor (layer3_outputs(1268)));
    layer4_outputs(1053) <= not((layer3_outputs(1007)) and (layer3_outputs(1800)));
    layer4_outputs(1054) <= (layer3_outputs(1029)) xor (layer3_outputs(267));
    layer4_outputs(1055) <= layer3_outputs(1607);
    layer4_outputs(1056) <= (layer3_outputs(2249)) and not (layer3_outputs(1778));
    layer4_outputs(1057) <= '0';
    layer4_outputs(1058) <= layer3_outputs(958);
    layer4_outputs(1059) <= not(layer3_outputs(1073)) or (layer3_outputs(1980));
    layer4_outputs(1060) <= not(layer3_outputs(242));
    layer4_outputs(1061) <= (layer3_outputs(2300)) and not (layer3_outputs(976));
    layer4_outputs(1062) <= not(layer3_outputs(44));
    layer4_outputs(1063) <= layer3_outputs(232);
    layer4_outputs(1064) <= (layer3_outputs(1237)) and not (layer3_outputs(502));
    layer4_outputs(1065) <= not(layer3_outputs(1));
    layer4_outputs(1066) <= layer3_outputs(325);
    layer4_outputs(1067) <= layer3_outputs(680);
    layer4_outputs(1068) <= not(layer3_outputs(2467));
    layer4_outputs(1069) <= not(layer3_outputs(1243)) or (layer3_outputs(683));
    layer4_outputs(1070) <= not(layer3_outputs(1936));
    layer4_outputs(1071) <= not(layer3_outputs(2233));
    layer4_outputs(1072) <= layer3_outputs(1604);
    layer4_outputs(1073) <= not(layer3_outputs(2112)) or (layer3_outputs(95));
    layer4_outputs(1074) <= layer3_outputs(1659);
    layer4_outputs(1075) <= not((layer3_outputs(948)) and (layer3_outputs(617)));
    layer4_outputs(1076) <= not((layer3_outputs(499)) or (layer3_outputs(1317)));
    layer4_outputs(1077) <= not(layer3_outputs(843));
    layer4_outputs(1078) <= not(layer3_outputs(1881));
    layer4_outputs(1079) <= (layer3_outputs(1165)) xor (layer3_outputs(1291));
    layer4_outputs(1080) <= not((layer3_outputs(2346)) and (layer3_outputs(897)));
    layer4_outputs(1081) <= layer3_outputs(2404);
    layer4_outputs(1082) <= layer3_outputs(928);
    layer4_outputs(1083) <= (layer3_outputs(577)) xor (layer3_outputs(1498));
    layer4_outputs(1084) <= not((layer3_outputs(674)) and (layer3_outputs(2208)));
    layer4_outputs(1085) <= layer3_outputs(1056);
    layer4_outputs(1086) <= '0';
    layer4_outputs(1087) <= layer3_outputs(108);
    layer4_outputs(1088) <= not(layer3_outputs(138));
    layer4_outputs(1089) <= (layer3_outputs(312)) xor (layer3_outputs(95));
    layer4_outputs(1090) <= (layer3_outputs(715)) and not (layer3_outputs(2400));
    layer4_outputs(1091) <= not((layer3_outputs(1139)) xor (layer3_outputs(1390)));
    layer4_outputs(1092) <= layer3_outputs(1577);
    layer4_outputs(1093) <= layer3_outputs(1196);
    layer4_outputs(1094) <= (layer3_outputs(716)) and not (layer3_outputs(629));
    layer4_outputs(1095) <= not(layer3_outputs(2231));
    layer4_outputs(1096) <= not(layer3_outputs(1115));
    layer4_outputs(1097) <= layer3_outputs(2290);
    layer4_outputs(1098) <= layer3_outputs(873);
    layer4_outputs(1099) <= not(layer3_outputs(658));
    layer4_outputs(1100) <= layer3_outputs(1521);
    layer4_outputs(1101) <= (layer3_outputs(2086)) and (layer3_outputs(1603));
    layer4_outputs(1102) <= (layer3_outputs(1854)) xor (layer3_outputs(1107));
    layer4_outputs(1103) <= layer3_outputs(790);
    layer4_outputs(1104) <= layer3_outputs(0);
    layer4_outputs(1105) <= not(layer3_outputs(817));
    layer4_outputs(1106) <= (layer3_outputs(2375)) and not (layer3_outputs(862));
    layer4_outputs(1107) <= layer3_outputs(1218);
    layer4_outputs(1108) <= not(layer3_outputs(2558));
    layer4_outputs(1109) <= not((layer3_outputs(2317)) or (layer3_outputs(487)));
    layer4_outputs(1110) <= not(layer3_outputs(1597));
    layer4_outputs(1111) <= not(layer3_outputs(1851)) or (layer3_outputs(2217));
    layer4_outputs(1112) <= (layer3_outputs(2378)) and (layer3_outputs(1542));
    layer4_outputs(1113) <= not(layer3_outputs(153)) or (layer3_outputs(1087));
    layer4_outputs(1114) <= layer3_outputs(2380);
    layer4_outputs(1115) <= not(layer3_outputs(2278));
    layer4_outputs(1116) <= layer3_outputs(35);
    layer4_outputs(1117) <= layer3_outputs(2506);
    layer4_outputs(1118) <= not(layer3_outputs(1988)) or (layer3_outputs(2484));
    layer4_outputs(1119) <= '1';
    layer4_outputs(1120) <= (layer3_outputs(1769)) and (layer3_outputs(1812));
    layer4_outputs(1121) <= not((layer3_outputs(1269)) or (layer3_outputs(344)));
    layer4_outputs(1122) <= layer3_outputs(539);
    layer4_outputs(1123) <= not((layer3_outputs(952)) and (layer3_outputs(457)));
    layer4_outputs(1124) <= not(layer3_outputs(973)) or (layer3_outputs(229));
    layer4_outputs(1125) <= not(layer3_outputs(29));
    layer4_outputs(1126) <= layer3_outputs(1499);
    layer4_outputs(1127) <= layer3_outputs(719);
    layer4_outputs(1128) <= not(layer3_outputs(405));
    layer4_outputs(1129) <= not(layer3_outputs(235));
    layer4_outputs(1130) <= not(layer3_outputs(2542));
    layer4_outputs(1131) <= (layer3_outputs(2142)) or (layer3_outputs(1853));
    layer4_outputs(1132) <= not(layer3_outputs(1703)) or (layer3_outputs(1860));
    layer4_outputs(1133) <= not(layer3_outputs(2462));
    layer4_outputs(1134) <= not(layer3_outputs(861));
    layer4_outputs(1135) <= not(layer3_outputs(803)) or (layer3_outputs(1609));
    layer4_outputs(1136) <= not(layer3_outputs(1979)) or (layer3_outputs(1144));
    layer4_outputs(1137) <= not(layer3_outputs(1554));
    layer4_outputs(1138) <= layer3_outputs(512);
    layer4_outputs(1139) <= (layer3_outputs(1181)) and (layer3_outputs(2339));
    layer4_outputs(1140) <= not(layer3_outputs(1618));
    layer4_outputs(1141) <= layer3_outputs(2106);
    layer4_outputs(1142) <= not(layer3_outputs(1365));
    layer4_outputs(1143) <= not(layer3_outputs(1773)) or (layer3_outputs(302));
    layer4_outputs(1144) <= not((layer3_outputs(879)) and (layer3_outputs(1752)));
    layer4_outputs(1145) <= not((layer3_outputs(696)) and (layer3_outputs(740)));
    layer4_outputs(1146) <= not(layer3_outputs(1177));
    layer4_outputs(1147) <= (layer3_outputs(465)) and not (layer3_outputs(1219));
    layer4_outputs(1148) <= layer3_outputs(299);
    layer4_outputs(1149) <= (layer3_outputs(1486)) xor (layer3_outputs(28));
    layer4_outputs(1150) <= not(layer3_outputs(1514));
    layer4_outputs(1151) <= (layer3_outputs(209)) and (layer3_outputs(1335));
    layer4_outputs(1152) <= not(layer3_outputs(2200));
    layer4_outputs(1153) <= not(layer3_outputs(123));
    layer4_outputs(1154) <= not(layer3_outputs(758)) or (layer3_outputs(2102));
    layer4_outputs(1155) <= not(layer3_outputs(1642));
    layer4_outputs(1156) <= not(layer3_outputs(1274));
    layer4_outputs(1157) <= layer3_outputs(172);
    layer4_outputs(1158) <= not(layer3_outputs(1714));
    layer4_outputs(1159) <= (layer3_outputs(402)) xor (layer3_outputs(1108));
    layer4_outputs(1160) <= layer3_outputs(2330);
    layer4_outputs(1161) <= '0';
    layer4_outputs(1162) <= (layer3_outputs(1286)) and not (layer3_outputs(748));
    layer4_outputs(1163) <= layer3_outputs(1682);
    layer4_outputs(1164) <= (layer3_outputs(2383)) xor (layer3_outputs(2189));
    layer4_outputs(1165) <= not(layer3_outputs(1516));
    layer4_outputs(1166) <= not(layer3_outputs(1171));
    layer4_outputs(1167) <= not(layer3_outputs(2335));
    layer4_outputs(1168) <= not(layer3_outputs(1163));
    layer4_outputs(1169) <= (layer3_outputs(2265)) and not (layer3_outputs(2041));
    layer4_outputs(1170) <= layer3_outputs(2443);
    layer4_outputs(1171) <= not((layer3_outputs(1520)) xor (layer3_outputs(2131)));
    layer4_outputs(1172) <= not(layer3_outputs(353));
    layer4_outputs(1173) <= not(layer3_outputs(2455)) or (layer3_outputs(2344));
    layer4_outputs(1174) <= not(layer3_outputs(1975));
    layer4_outputs(1175) <= '1';
    layer4_outputs(1176) <= layer3_outputs(1904);
    layer4_outputs(1177) <= layer3_outputs(2301);
    layer4_outputs(1178) <= not(layer3_outputs(2472));
    layer4_outputs(1179) <= not((layer3_outputs(1705)) and (layer3_outputs(105)));
    layer4_outputs(1180) <= not(layer3_outputs(1747));
    layer4_outputs(1181) <= (layer3_outputs(2417)) and not (layer3_outputs(406));
    layer4_outputs(1182) <= not((layer3_outputs(2488)) and (layer3_outputs(286)));
    layer4_outputs(1183) <= not(layer3_outputs(1751));
    layer4_outputs(1184) <= not((layer3_outputs(907)) and (layer3_outputs(1056)));
    layer4_outputs(1185) <= not((layer3_outputs(2237)) or (layer3_outputs(102)));
    layer4_outputs(1186) <= (layer3_outputs(1086)) and not (layer3_outputs(1621));
    layer4_outputs(1187) <= (layer3_outputs(640)) and not (layer3_outputs(2420));
    layer4_outputs(1188) <= not((layer3_outputs(279)) xor (layer3_outputs(1195)));
    layer4_outputs(1189) <= not(layer3_outputs(257)) or (layer3_outputs(1395));
    layer4_outputs(1190) <= not((layer3_outputs(1000)) or (layer3_outputs(1589)));
    layer4_outputs(1191) <= (layer3_outputs(45)) or (layer3_outputs(1474));
    layer4_outputs(1192) <= not(layer3_outputs(1585)) or (layer3_outputs(825));
    layer4_outputs(1193) <= not(layer3_outputs(1029)) or (layer3_outputs(1548));
    layer4_outputs(1194) <= not(layer3_outputs(548)) or (layer3_outputs(1435));
    layer4_outputs(1195) <= (layer3_outputs(2286)) and not (layer3_outputs(1571));
    layer4_outputs(1196) <= not((layer3_outputs(745)) and (layer3_outputs(360)));
    layer4_outputs(1197) <= not((layer3_outputs(1207)) xor (layer3_outputs(373)));
    layer4_outputs(1198) <= not(layer3_outputs(2382));
    layer4_outputs(1199) <= (layer3_outputs(742)) or (layer3_outputs(330));
    layer4_outputs(1200) <= (layer3_outputs(300)) xor (layer3_outputs(368));
    layer4_outputs(1201) <= not(layer3_outputs(2345));
    layer4_outputs(1202) <= not(layer3_outputs(1060));
    layer4_outputs(1203) <= not((layer3_outputs(2264)) xor (layer3_outputs(2046)));
    layer4_outputs(1204) <= layer3_outputs(1802);
    layer4_outputs(1205) <= (layer3_outputs(1038)) and not (layer3_outputs(839));
    layer4_outputs(1206) <= '1';
    layer4_outputs(1207) <= not(layer3_outputs(1288));
    layer4_outputs(1208) <= layer3_outputs(306);
    layer4_outputs(1209) <= not(layer3_outputs(119));
    layer4_outputs(1210) <= layer3_outputs(1608);
    layer4_outputs(1211) <= layer3_outputs(234);
    layer4_outputs(1212) <= (layer3_outputs(2409)) and not (layer3_outputs(510));
    layer4_outputs(1213) <= (layer3_outputs(490)) and not (layer3_outputs(724));
    layer4_outputs(1214) <= not((layer3_outputs(1210)) or (layer3_outputs(148)));
    layer4_outputs(1215) <= layer3_outputs(2083);
    layer4_outputs(1216) <= layer3_outputs(1698);
    layer4_outputs(1217) <= (layer3_outputs(227)) xor (layer3_outputs(1457));
    layer4_outputs(1218) <= not(layer3_outputs(372)) or (layer3_outputs(2482));
    layer4_outputs(1219) <= '1';
    layer4_outputs(1220) <= layer3_outputs(42);
    layer4_outputs(1221) <= layer3_outputs(2068);
    layer4_outputs(1222) <= layer3_outputs(1014);
    layer4_outputs(1223) <= layer3_outputs(808);
    layer4_outputs(1224) <= not(layer3_outputs(1761));
    layer4_outputs(1225) <= not(layer3_outputs(2479));
    layer4_outputs(1226) <= layer3_outputs(2275);
    layer4_outputs(1227) <= layer3_outputs(1695);
    layer4_outputs(1228) <= (layer3_outputs(1417)) xor (layer3_outputs(849));
    layer4_outputs(1229) <= layer3_outputs(28);
    layer4_outputs(1230) <= layer3_outputs(1980);
    layer4_outputs(1231) <= layer3_outputs(1716);
    layer4_outputs(1232) <= (layer3_outputs(1271)) and not (layer3_outputs(2014));
    layer4_outputs(1233) <= not(layer3_outputs(1563));
    layer4_outputs(1234) <= (layer3_outputs(244)) and not (layer3_outputs(2315));
    layer4_outputs(1235) <= (layer3_outputs(781)) xor (layer3_outputs(2259));
    layer4_outputs(1236) <= layer3_outputs(2282);
    layer4_outputs(1237) <= not(layer3_outputs(1623));
    layer4_outputs(1238) <= (layer3_outputs(2140)) and not (layer3_outputs(1967));
    layer4_outputs(1239) <= not(layer3_outputs(1107)) or (layer3_outputs(964));
    layer4_outputs(1240) <= layer3_outputs(1076);
    layer4_outputs(1241) <= layer3_outputs(462);
    layer4_outputs(1242) <= (layer3_outputs(1457)) and not (layer3_outputs(1383));
    layer4_outputs(1243) <= layer3_outputs(1896);
    layer4_outputs(1244) <= not(layer3_outputs(582));
    layer4_outputs(1245) <= (layer3_outputs(1705)) or (layer3_outputs(530));
    layer4_outputs(1246) <= (layer3_outputs(11)) and not (layer3_outputs(385));
    layer4_outputs(1247) <= not((layer3_outputs(755)) or (layer3_outputs(786)));
    layer4_outputs(1248) <= layer3_outputs(2238);
    layer4_outputs(1249) <= (layer3_outputs(2283)) or (layer3_outputs(2524));
    layer4_outputs(1250) <= (layer3_outputs(47)) and not (layer3_outputs(2489));
    layer4_outputs(1251) <= (layer3_outputs(903)) and not (layer3_outputs(838));
    layer4_outputs(1252) <= (layer3_outputs(1088)) xor (layer3_outputs(985));
    layer4_outputs(1253) <= not(layer3_outputs(1013));
    layer4_outputs(1254) <= not(layer3_outputs(2538));
    layer4_outputs(1255) <= (layer3_outputs(1969)) and (layer3_outputs(1624));
    layer4_outputs(1256) <= not(layer3_outputs(212)) or (layer3_outputs(1856));
    layer4_outputs(1257) <= '0';
    layer4_outputs(1258) <= layer3_outputs(1917);
    layer4_outputs(1259) <= (layer3_outputs(737)) or (layer3_outputs(1497));
    layer4_outputs(1260) <= not(layer3_outputs(1575));
    layer4_outputs(1261) <= not(layer3_outputs(645)) or (layer3_outputs(2227));
    layer4_outputs(1262) <= not(layer3_outputs(18));
    layer4_outputs(1263) <= layer3_outputs(1018);
    layer4_outputs(1264) <= (layer3_outputs(994)) and not (layer3_outputs(1669));
    layer4_outputs(1265) <= (layer3_outputs(345)) and (layer3_outputs(827));
    layer4_outputs(1266) <= (layer3_outputs(1374)) and (layer3_outputs(1290));
    layer4_outputs(1267) <= not(layer3_outputs(84));
    layer4_outputs(1268) <= (layer3_outputs(1598)) and (layer3_outputs(2368));
    layer4_outputs(1269) <= not(layer3_outputs(1957));
    layer4_outputs(1270) <= (layer3_outputs(886)) and not (layer3_outputs(914));
    layer4_outputs(1271) <= (layer3_outputs(647)) and not (layer3_outputs(2183));
    layer4_outputs(1272) <= not(layer3_outputs(1222));
    layer4_outputs(1273) <= (layer3_outputs(668)) and not (layer3_outputs(1746));
    layer4_outputs(1274) <= not(layer3_outputs(629));
    layer4_outputs(1275) <= layer3_outputs(1597);
    layer4_outputs(1276) <= (layer3_outputs(277)) or (layer3_outputs(356));
    layer4_outputs(1277) <= layer3_outputs(117);
    layer4_outputs(1278) <= not((layer3_outputs(972)) xor (layer3_outputs(1212)));
    layer4_outputs(1279) <= not(layer3_outputs(58));
    layer4_outputs(1280) <= (layer3_outputs(1768)) xor (layer3_outputs(565));
    layer4_outputs(1281) <= not(layer3_outputs(1397));
    layer4_outputs(1282) <= not((layer3_outputs(741)) or (layer3_outputs(743)));
    layer4_outputs(1283) <= not(layer3_outputs(2523)) or (layer3_outputs(1255));
    layer4_outputs(1284) <= (layer3_outputs(1600)) or (layer3_outputs(120));
    layer4_outputs(1285) <= layer3_outputs(1021);
    layer4_outputs(1286) <= layer3_outputs(1123);
    layer4_outputs(1287) <= not(layer3_outputs(1864));
    layer4_outputs(1288) <= layer3_outputs(1537);
    layer4_outputs(1289) <= (layer3_outputs(618)) and not (layer3_outputs(804));
    layer4_outputs(1290) <= not(layer3_outputs(1193));
    layer4_outputs(1291) <= layer3_outputs(641);
    layer4_outputs(1292) <= layer3_outputs(2025);
    layer4_outputs(1293) <= layer3_outputs(2242);
    layer4_outputs(1294) <= not(layer3_outputs(2126)) or (layer3_outputs(1592));
    layer4_outputs(1295) <= layer3_outputs(415);
    layer4_outputs(1296) <= not(layer3_outputs(476));
    layer4_outputs(1297) <= not(layer3_outputs(1145));
    layer4_outputs(1298) <= layer3_outputs(1033);
    layer4_outputs(1299) <= layer3_outputs(1149);
    layer4_outputs(1300) <= not(layer3_outputs(426)) or (layer3_outputs(788));
    layer4_outputs(1301) <= layer3_outputs(2149);
    layer4_outputs(1302) <= not(layer3_outputs(1744));
    layer4_outputs(1303) <= (layer3_outputs(29)) and not (layer3_outputs(1722));
    layer4_outputs(1304) <= not(layer3_outputs(528)) or (layer3_outputs(1688));
    layer4_outputs(1305) <= not(layer3_outputs(803));
    layer4_outputs(1306) <= layer3_outputs(787);
    layer4_outputs(1307) <= not(layer3_outputs(1343));
    layer4_outputs(1308) <= '0';
    layer4_outputs(1309) <= not(layer3_outputs(1187)) or (layer3_outputs(887));
    layer4_outputs(1310) <= (layer3_outputs(1884)) and not (layer3_outputs(921));
    layer4_outputs(1311) <= layer3_outputs(1120);
    layer4_outputs(1312) <= not(layer3_outputs(784));
    layer4_outputs(1313) <= layer3_outputs(1725);
    layer4_outputs(1314) <= not(layer3_outputs(1049));
    layer4_outputs(1315) <= layer3_outputs(621);
    layer4_outputs(1316) <= layer3_outputs(752);
    layer4_outputs(1317) <= (layer3_outputs(2246)) or (layer3_outputs(1278));
    layer4_outputs(1318) <= not(layer3_outputs(2553));
    layer4_outputs(1319) <= not((layer3_outputs(161)) and (layer3_outputs(1046)));
    layer4_outputs(1320) <= layer3_outputs(407);
    layer4_outputs(1321) <= not((layer3_outputs(92)) or (layer3_outputs(1944)));
    layer4_outputs(1322) <= not(layer3_outputs(2366)) or (layer3_outputs(805));
    layer4_outputs(1323) <= layer3_outputs(2307);
    layer4_outputs(1324) <= layer3_outputs(2503);
    layer4_outputs(1325) <= not((layer3_outputs(1210)) or (layer3_outputs(440)));
    layer4_outputs(1326) <= (layer3_outputs(34)) and not (layer3_outputs(503));
    layer4_outputs(1327) <= not(layer3_outputs(1221)) or (layer3_outputs(70));
    layer4_outputs(1328) <= not(layer3_outputs(1755));
    layer4_outputs(1329) <= not(layer3_outputs(1407));
    layer4_outputs(1330) <= (layer3_outputs(856)) and not (layer3_outputs(1721));
    layer4_outputs(1331) <= (layer3_outputs(1500)) or (layer3_outputs(866));
    layer4_outputs(1332) <= (layer3_outputs(352)) and not (layer3_outputs(2305));
    layer4_outputs(1333) <= not(layer3_outputs(2297));
    layer4_outputs(1334) <= (layer3_outputs(2016)) and (layer3_outputs(1771));
    layer4_outputs(1335) <= not((layer3_outputs(1844)) xor (layer3_outputs(251)));
    layer4_outputs(1336) <= layer3_outputs(480);
    layer4_outputs(1337) <= (layer3_outputs(912)) and not (layer3_outputs(195));
    layer4_outputs(1338) <= not(layer3_outputs(2454));
    layer4_outputs(1339) <= (layer3_outputs(1118)) and not (layer3_outputs(843));
    layer4_outputs(1340) <= not(layer3_outputs(657)) or (layer3_outputs(531));
    layer4_outputs(1341) <= not(layer3_outputs(2087));
    layer4_outputs(1342) <= (layer3_outputs(1443)) or (layer3_outputs(1415));
    layer4_outputs(1343) <= layer3_outputs(343);
    layer4_outputs(1344) <= not(layer3_outputs(680)) or (layer3_outputs(2479));
    layer4_outputs(1345) <= not(layer3_outputs(487));
    layer4_outputs(1346) <= not(layer3_outputs(498));
    layer4_outputs(1347) <= not(layer3_outputs(1490)) or (layer3_outputs(243));
    layer4_outputs(1348) <= not((layer3_outputs(899)) or (layer3_outputs(2157)));
    layer4_outputs(1349) <= not(layer3_outputs(299)) or (layer3_outputs(2273));
    layer4_outputs(1350) <= not(layer3_outputs(1828));
    layer4_outputs(1351) <= not(layer3_outputs(1316));
    layer4_outputs(1352) <= layer3_outputs(872);
    layer4_outputs(1353) <= layer3_outputs(2255);
    layer4_outputs(1354) <= (layer3_outputs(1544)) and (layer3_outputs(1239));
    layer4_outputs(1355) <= not(layer3_outputs(78));
    layer4_outputs(1356) <= not(layer3_outputs(1654));
    layer4_outputs(1357) <= not(layer3_outputs(1082)) or (layer3_outputs(125));
    layer4_outputs(1358) <= not(layer3_outputs(248));
    layer4_outputs(1359) <= layer3_outputs(2361);
    layer4_outputs(1360) <= (layer3_outputs(1689)) and not (layer3_outputs(1245));
    layer4_outputs(1361) <= not(layer3_outputs(2224));
    layer4_outputs(1362) <= layer3_outputs(246);
    layer4_outputs(1363) <= layer3_outputs(2412);
    layer4_outputs(1364) <= not(layer3_outputs(2549));
    layer4_outputs(1365) <= not((layer3_outputs(879)) xor (layer3_outputs(71)));
    layer4_outputs(1366) <= not((layer3_outputs(2117)) or (layer3_outputs(195)));
    layer4_outputs(1367) <= layer3_outputs(1849);
    layer4_outputs(1368) <= not(layer3_outputs(186));
    layer4_outputs(1369) <= not((layer3_outputs(1193)) xor (layer3_outputs(480)));
    layer4_outputs(1370) <= not((layer3_outputs(37)) and (layer3_outputs(483)));
    layer4_outputs(1371) <= not(layer3_outputs(180));
    layer4_outputs(1372) <= layer3_outputs(51);
    layer4_outputs(1373) <= '1';
    layer4_outputs(1374) <= not(layer3_outputs(2296));
    layer4_outputs(1375) <= not(layer3_outputs(947));
    layer4_outputs(1376) <= not((layer3_outputs(1795)) and (layer3_outputs(1167)));
    layer4_outputs(1377) <= layer3_outputs(1785);
    layer4_outputs(1378) <= layer3_outputs(2084);
    layer4_outputs(1379) <= (layer3_outputs(437)) and not (layer3_outputs(48));
    layer4_outputs(1380) <= not(layer3_outputs(783));
    layer4_outputs(1381) <= not((layer3_outputs(1022)) and (layer3_outputs(410)));
    layer4_outputs(1382) <= not(layer3_outputs(671));
    layer4_outputs(1383) <= not(layer3_outputs(23));
    layer4_outputs(1384) <= not((layer3_outputs(540)) or (layer3_outputs(1753)));
    layer4_outputs(1385) <= not(layer3_outputs(951));
    layer4_outputs(1386) <= not((layer3_outputs(504)) xor (layer3_outputs(880)));
    layer4_outputs(1387) <= not(layer3_outputs(1050));
    layer4_outputs(1388) <= (layer3_outputs(2314)) xor (layer3_outputs(1032));
    layer4_outputs(1389) <= layer3_outputs(556);
    layer4_outputs(1390) <= not((layer3_outputs(2295)) xor (layer3_outputs(1429)));
    layer4_outputs(1391) <= not(layer3_outputs(801));
    layer4_outputs(1392) <= not(layer3_outputs(1393));
    layer4_outputs(1393) <= (layer3_outputs(684)) and not (layer3_outputs(163));
    layer4_outputs(1394) <= layer3_outputs(1449);
    layer4_outputs(1395) <= layer3_outputs(1798);
    layer4_outputs(1396) <= layer3_outputs(2067);
    layer4_outputs(1397) <= (layer3_outputs(1814)) and not (layer3_outputs(1801));
    layer4_outputs(1398) <= not(layer3_outputs(1363));
    layer4_outputs(1399) <= not(layer3_outputs(2032));
    layer4_outputs(1400) <= layer3_outputs(806);
    layer4_outputs(1401) <= layer3_outputs(765);
    layer4_outputs(1402) <= layer3_outputs(2156);
    layer4_outputs(1403) <= not(layer3_outputs(281));
    layer4_outputs(1404) <= not(layer3_outputs(2074));
    layer4_outputs(1405) <= layer3_outputs(2007);
    layer4_outputs(1406) <= not(layer3_outputs(50));
    layer4_outputs(1407) <= not((layer3_outputs(256)) xor (layer3_outputs(2312)));
    layer4_outputs(1408) <= not(layer3_outputs(183));
    layer4_outputs(1409) <= layer3_outputs(1323);
    layer4_outputs(1410) <= layer3_outputs(2485);
    layer4_outputs(1411) <= layer3_outputs(832);
    layer4_outputs(1412) <= (layer3_outputs(93)) xor (layer3_outputs(305));
    layer4_outputs(1413) <= not(layer3_outputs(1849));
    layer4_outputs(1414) <= not((layer3_outputs(2415)) or (layer3_outputs(1231)));
    layer4_outputs(1415) <= (layer3_outputs(338)) xor (layer3_outputs(501));
    layer4_outputs(1416) <= not(layer3_outputs(2192));
    layer4_outputs(1417) <= layer3_outputs(897);
    layer4_outputs(1418) <= not(layer3_outputs(2481));
    layer4_outputs(1419) <= (layer3_outputs(2313)) or (layer3_outputs(1942));
    layer4_outputs(1420) <= layer3_outputs(2066);
    layer4_outputs(1421) <= (layer3_outputs(1296)) or (layer3_outputs(399));
    layer4_outputs(1422) <= not(layer3_outputs(1327));
    layer4_outputs(1423) <= (layer3_outputs(932)) and (layer3_outputs(580));
    layer4_outputs(1424) <= not(layer3_outputs(688));
    layer4_outputs(1425) <= layer3_outputs(1405);
    layer4_outputs(1426) <= layer3_outputs(120);
    layer4_outputs(1427) <= not(layer3_outputs(1040));
    layer4_outputs(1428) <= layer3_outputs(1170);
    layer4_outputs(1429) <= layer3_outputs(1740);
    layer4_outputs(1430) <= not(layer3_outputs(1063));
    layer4_outputs(1431) <= (layer3_outputs(0)) and (layer3_outputs(246));
    layer4_outputs(1432) <= not(layer3_outputs(2296));
    layer4_outputs(1433) <= (layer3_outputs(112)) and not (layer3_outputs(1855));
    layer4_outputs(1434) <= not((layer3_outputs(97)) or (layer3_outputs(1088)));
    layer4_outputs(1435) <= layer3_outputs(2487);
    layer4_outputs(1436) <= not((layer3_outputs(718)) and (layer3_outputs(1892)));
    layer4_outputs(1437) <= layer3_outputs(1044);
    layer4_outputs(1438) <= layer3_outputs(192);
    layer4_outputs(1439) <= not(layer3_outputs(1479)) or (layer3_outputs(1206));
    layer4_outputs(1440) <= not(layer3_outputs(2193));
    layer4_outputs(1441) <= layer3_outputs(979);
    layer4_outputs(1442) <= layer3_outputs(34);
    layer4_outputs(1443) <= layer3_outputs(825);
    layer4_outputs(1444) <= not((layer3_outputs(325)) xor (layer3_outputs(1242)));
    layer4_outputs(1445) <= layer3_outputs(1139);
    layer4_outputs(1446) <= layer3_outputs(2236);
    layer4_outputs(1447) <= (layer3_outputs(293)) xor (layer3_outputs(513));
    layer4_outputs(1448) <= not((layer3_outputs(2322)) and (layer3_outputs(599)));
    layer4_outputs(1449) <= not((layer3_outputs(691)) and (layer3_outputs(831)));
    layer4_outputs(1450) <= layer3_outputs(255);
    layer4_outputs(1451) <= not(layer3_outputs(1636)) or (layer3_outputs(2327));
    layer4_outputs(1452) <= not(layer3_outputs(780));
    layer4_outputs(1453) <= layer3_outputs(516);
    layer4_outputs(1454) <= (layer3_outputs(776)) and not (layer3_outputs(1924));
    layer4_outputs(1455) <= not(layer3_outputs(2514));
    layer4_outputs(1456) <= (layer3_outputs(1822)) and not (layer3_outputs(1256));
    layer4_outputs(1457) <= not((layer3_outputs(586)) or (layer3_outputs(1346)));
    layer4_outputs(1458) <= (layer3_outputs(1550)) and not (layer3_outputs(2435));
    layer4_outputs(1459) <= layer3_outputs(1992);
    layer4_outputs(1460) <= not(layer3_outputs(1937)) or (layer3_outputs(656));
    layer4_outputs(1461) <= not(layer3_outputs(1920));
    layer4_outputs(1462) <= (layer3_outputs(761)) or (layer3_outputs(942));
    layer4_outputs(1463) <= not(layer3_outputs(53));
    layer4_outputs(1464) <= not((layer3_outputs(474)) or (layer3_outputs(1186)));
    layer4_outputs(1465) <= not(layer3_outputs(1830));
    layer4_outputs(1466) <= not(layer3_outputs(158));
    layer4_outputs(1467) <= layer3_outputs(1416);
    layer4_outputs(1468) <= layer3_outputs(893);
    layer4_outputs(1469) <= (layer3_outputs(901)) and not (layer3_outputs(657));
    layer4_outputs(1470) <= not(layer3_outputs(944));
    layer4_outputs(1471) <= not(layer3_outputs(622)) or (layer3_outputs(1962));
    layer4_outputs(1472) <= not((layer3_outputs(2430)) or (layer3_outputs(1944)));
    layer4_outputs(1473) <= (layer3_outputs(542)) or (layer3_outputs(392));
    layer4_outputs(1474) <= not(layer3_outputs(218));
    layer4_outputs(1475) <= layer3_outputs(406);
    layer4_outputs(1476) <= (layer3_outputs(1468)) or (layer3_outputs(171));
    layer4_outputs(1477) <= not((layer3_outputs(2127)) xor (layer3_outputs(1274)));
    layer4_outputs(1478) <= (layer3_outputs(19)) and (layer3_outputs(1848));
    layer4_outputs(1479) <= layer3_outputs(1102);
    layer4_outputs(1480) <= (layer3_outputs(1213)) xor (layer3_outputs(1792));
    layer4_outputs(1481) <= not((layer3_outputs(792)) or (layer3_outputs(1187)));
    layer4_outputs(1482) <= layer3_outputs(2384);
    layer4_outputs(1483) <= layer3_outputs(1779);
    layer4_outputs(1484) <= not(layer3_outputs(1831));
    layer4_outputs(1485) <= not(layer3_outputs(2172));
    layer4_outputs(1486) <= layer3_outputs(1651);
    layer4_outputs(1487) <= not(layer3_outputs(841));
    layer4_outputs(1488) <= (layer3_outputs(2308)) and not (layer3_outputs(25));
    layer4_outputs(1489) <= layer3_outputs(1439);
    layer4_outputs(1490) <= (layer3_outputs(1658)) xor (layer3_outputs(1535));
    layer4_outputs(1491) <= not(layer3_outputs(453)) or (layer3_outputs(1799));
    layer4_outputs(1492) <= layer3_outputs(1590);
    layer4_outputs(1493) <= not(layer3_outputs(2513));
    layer4_outputs(1494) <= layer3_outputs(1809);
    layer4_outputs(1495) <= (layer3_outputs(337)) and not (layer3_outputs(1546));
    layer4_outputs(1496) <= not(layer3_outputs(2174)) or (layer3_outputs(1424));
    layer4_outputs(1497) <= (layer3_outputs(397)) and (layer3_outputs(1090));
    layer4_outputs(1498) <= layer3_outputs(1116);
    layer4_outputs(1499) <= (layer3_outputs(1972)) and not (layer3_outputs(67));
    layer4_outputs(1500) <= (layer3_outputs(1450)) and (layer3_outputs(2528));
    layer4_outputs(1501) <= not(layer3_outputs(2398));
    layer4_outputs(1502) <= not(layer3_outputs(911));
    layer4_outputs(1503) <= layer3_outputs(2061);
    layer4_outputs(1504) <= (layer3_outputs(2020)) and (layer3_outputs(1326));
    layer4_outputs(1505) <= not(layer3_outputs(2103)) or (layer3_outputs(2396));
    layer4_outputs(1506) <= not((layer3_outputs(2397)) or (layer3_outputs(633)));
    layer4_outputs(1507) <= not(layer3_outputs(693)) or (layer3_outputs(318));
    layer4_outputs(1508) <= layer3_outputs(1176);
    layer4_outputs(1509) <= not(layer3_outputs(378)) or (layer3_outputs(389));
    layer4_outputs(1510) <= not(layer3_outputs(2261));
    layer4_outputs(1511) <= not((layer3_outputs(1741)) or (layer3_outputs(1071)));
    layer4_outputs(1512) <= layer3_outputs(2266);
    layer4_outputs(1513) <= layer3_outputs(1329);
    layer4_outputs(1514) <= not(layer3_outputs(1692)) or (layer3_outputs(1057));
    layer4_outputs(1515) <= not(layer3_outputs(2179));
    layer4_outputs(1516) <= layer3_outputs(404);
    layer4_outputs(1517) <= (layer3_outputs(1225)) and (layer3_outputs(867));
    layer4_outputs(1518) <= (layer3_outputs(118)) and not (layer3_outputs(85));
    layer4_outputs(1519) <= not(layer3_outputs(441));
    layer4_outputs(1520) <= not(layer3_outputs(656));
    layer4_outputs(1521) <= (layer3_outputs(1030)) and (layer3_outputs(828));
    layer4_outputs(1522) <= not(layer3_outputs(162));
    layer4_outputs(1523) <= layer3_outputs(826);
    layer4_outputs(1524) <= not((layer3_outputs(2287)) and (layer3_outputs(1702)));
    layer4_outputs(1525) <= not(layer3_outputs(1251)) or (layer3_outputs(2414));
    layer4_outputs(1526) <= '0';
    layer4_outputs(1527) <= not((layer3_outputs(2289)) xor (layer3_outputs(2185)));
    layer4_outputs(1528) <= layer3_outputs(2556);
    layer4_outputs(1529) <= not((layer3_outputs(126)) or (layer3_outputs(725)));
    layer4_outputs(1530) <= (layer3_outputs(2498)) or (layer3_outputs(925));
    layer4_outputs(1531) <= not((layer3_outputs(164)) xor (layer3_outputs(679)));
    layer4_outputs(1532) <= not(layer3_outputs(1727));
    layer4_outputs(1533) <= not((layer3_outputs(1607)) and (layer3_outputs(2008)));
    layer4_outputs(1534) <= not(layer3_outputs(212));
    layer4_outputs(1535) <= not(layer3_outputs(1886));
    layer4_outputs(1536) <= layer3_outputs(2473);
    layer4_outputs(1537) <= not(layer3_outputs(2330));
    layer4_outputs(1538) <= layer3_outputs(169);
    layer4_outputs(1539) <= layer3_outputs(1113);
    layer4_outputs(1540) <= not((layer3_outputs(1841)) or (layer3_outputs(579)));
    layer4_outputs(1541) <= not((layer3_outputs(2356)) xor (layer3_outputs(1912)));
    layer4_outputs(1542) <= (layer3_outputs(2326)) and not (layer3_outputs(1781));
    layer4_outputs(1543) <= layer3_outputs(1400);
    layer4_outputs(1544) <= not(layer3_outputs(515));
    layer4_outputs(1545) <= not(layer3_outputs(694));
    layer4_outputs(1546) <= layer3_outputs(692);
    layer4_outputs(1547) <= not(layer3_outputs(328));
    layer4_outputs(1548) <= layer3_outputs(833);
    layer4_outputs(1549) <= (layer3_outputs(2417)) and not (layer3_outputs(1601));
    layer4_outputs(1550) <= not(layer3_outputs(251));
    layer4_outputs(1551) <= not(layer3_outputs(860)) or (layer3_outputs(2202));
    layer4_outputs(1552) <= not(layer3_outputs(198));
    layer4_outputs(1553) <= layer3_outputs(1220);
    layer4_outputs(1554) <= not(layer3_outputs(1963));
    layer4_outputs(1555) <= layer3_outputs(1907);
    layer4_outputs(1556) <= '0';
    layer4_outputs(1557) <= (layer3_outputs(869)) and (layer3_outputs(308));
    layer4_outputs(1558) <= layer3_outputs(341);
    layer4_outputs(1559) <= layer3_outputs(2067);
    layer4_outputs(1560) <= (layer3_outputs(495)) and (layer3_outputs(2369));
    layer4_outputs(1561) <= not(layer3_outputs(1603));
    layer4_outputs(1562) <= layer3_outputs(1356);
    layer4_outputs(1563) <= not(layer3_outputs(399)) or (layer3_outputs(370));
    layer4_outputs(1564) <= (layer3_outputs(853)) and not (layer3_outputs(549));
    layer4_outputs(1565) <= layer3_outputs(2433);
    layer4_outputs(1566) <= layer3_outputs(801);
    layer4_outputs(1567) <= not(layer3_outputs(237)) or (layer3_outputs(324));
    layer4_outputs(1568) <= not((layer3_outputs(1183)) xor (layer3_outputs(1234)));
    layer4_outputs(1569) <= not((layer3_outputs(2314)) and (layer3_outputs(172)));
    layer4_outputs(1570) <= not(layer3_outputs(2251));
    layer4_outputs(1571) <= layer3_outputs(1680);
    layer4_outputs(1572) <= layer3_outputs(2268);
    layer4_outputs(1573) <= (layer3_outputs(1783)) or (layer3_outputs(1825));
    layer4_outputs(1574) <= not((layer3_outputs(1661)) or (layer3_outputs(94)));
    layer4_outputs(1575) <= (layer3_outputs(2456)) and (layer3_outputs(388));
    layer4_outputs(1576) <= not(layer3_outputs(1711));
    layer4_outputs(1577) <= not((layer3_outputs(1100)) or (layer3_outputs(1267)));
    layer4_outputs(1578) <= not(layer3_outputs(2523));
    layer4_outputs(1579) <= layer3_outputs(545);
    layer4_outputs(1580) <= layer3_outputs(391);
    layer4_outputs(1581) <= layer3_outputs(68);
    layer4_outputs(1582) <= not((layer3_outputs(1079)) or (layer3_outputs(2162)));
    layer4_outputs(1583) <= not(layer3_outputs(883));
    layer4_outputs(1584) <= not(layer3_outputs(1542));
    layer4_outputs(1585) <= (layer3_outputs(2464)) and (layer3_outputs(1627));
    layer4_outputs(1586) <= not(layer3_outputs(630));
    layer4_outputs(1587) <= not(layer3_outputs(2310));
    layer4_outputs(1588) <= not(layer3_outputs(1633)) or (layer3_outputs(1696));
    layer4_outputs(1589) <= (layer3_outputs(1154)) and not (layer3_outputs(500));
    layer4_outputs(1590) <= not(layer3_outputs(2191)) or (layer3_outputs(2168));
    layer4_outputs(1591) <= not((layer3_outputs(1923)) or (layer3_outputs(2525)));
    layer4_outputs(1592) <= not((layer3_outputs(634)) and (layer3_outputs(2136)));
    layer4_outputs(1593) <= (layer3_outputs(123)) xor (layer3_outputs(2040));
    layer4_outputs(1594) <= not((layer3_outputs(2406)) xor (layer3_outputs(327)));
    layer4_outputs(1595) <= not(layer3_outputs(1553)) or (layer3_outputs(1547));
    layer4_outputs(1596) <= not(layer3_outputs(2152)) or (layer3_outputs(2250));
    layer4_outputs(1597) <= not(layer3_outputs(156));
    layer4_outputs(1598) <= not(layer3_outputs(2242));
    layer4_outputs(1599) <= (layer3_outputs(551)) and (layer3_outputs(260));
    layer4_outputs(1600) <= not(layer3_outputs(1524)) or (layer3_outputs(2502));
    layer4_outputs(1601) <= not((layer3_outputs(2149)) or (layer3_outputs(54)));
    layer4_outputs(1602) <= not((layer3_outputs(2309)) xor (layer3_outputs(854)));
    layer4_outputs(1603) <= (layer3_outputs(1857)) and (layer3_outputs(587));
    layer4_outputs(1604) <= layer3_outputs(1762);
    layer4_outputs(1605) <= (layer3_outputs(896)) or (layer3_outputs(870));
    layer4_outputs(1606) <= layer3_outputs(2347);
    layer4_outputs(1607) <= (layer3_outputs(1048)) and not (layer3_outputs(2360));
    layer4_outputs(1608) <= not(layer3_outputs(1666));
    layer4_outputs(1609) <= not(layer3_outputs(1754));
    layer4_outputs(1610) <= layer3_outputs(1582);
    layer4_outputs(1611) <= (layer3_outputs(1999)) and not (layer3_outputs(1181));
    layer4_outputs(1612) <= not(layer3_outputs(1734));
    layer4_outputs(1613) <= not(layer3_outputs(2264));
    layer4_outputs(1614) <= not(layer3_outputs(1059)) or (layer3_outputs(794));
    layer4_outputs(1615) <= (layer3_outputs(2154)) xor (layer3_outputs(2113));
    layer4_outputs(1616) <= (layer3_outputs(491)) xor (layer3_outputs(928));
    layer4_outputs(1617) <= not(layer3_outputs(1079));
    layer4_outputs(1618) <= not((layer3_outputs(432)) xor (layer3_outputs(2548)));
    layer4_outputs(1619) <= not(layer3_outputs(767));
    layer4_outputs(1620) <= not(layer3_outputs(852));
    layer4_outputs(1621) <= not((layer3_outputs(362)) and (layer3_outputs(950)));
    layer4_outputs(1622) <= (layer3_outputs(1017)) and not (layer3_outputs(369));
    layer4_outputs(1623) <= not(layer3_outputs(1947));
    layer4_outputs(1624) <= not((layer3_outputs(1916)) and (layer3_outputs(2502)));
    layer4_outputs(1625) <= (layer3_outputs(2366)) and not (layer3_outputs(2406));
    layer4_outputs(1626) <= not(layer3_outputs(1538));
    layer4_outputs(1627) <= not(layer3_outputs(2541)) or (layer3_outputs(1599));
    layer4_outputs(1628) <= layer3_outputs(1102);
    layer4_outputs(1629) <= layer3_outputs(687);
    layer4_outputs(1630) <= not(layer3_outputs(435)) or (layer3_outputs(1220));
    layer4_outputs(1631) <= not(layer3_outputs(497));
    layer4_outputs(1632) <= not((layer3_outputs(814)) and (layer3_outputs(678)));
    layer4_outputs(1633) <= not(layer3_outputs(2326)) or (layer3_outputs(821));
    layer4_outputs(1634) <= not(layer3_outputs(1357));
    layer4_outputs(1635) <= layer3_outputs(1830);
    layer4_outputs(1636) <= '1';
    layer4_outputs(1637) <= not(layer3_outputs(375));
    layer4_outputs(1638) <= not((layer3_outputs(2221)) or (layer3_outputs(2551)));
    layer4_outputs(1639) <= not((layer3_outputs(1112)) or (layer3_outputs(1325)));
    layer4_outputs(1640) <= (layer3_outputs(2212)) and not (layer3_outputs(2271));
    layer4_outputs(1641) <= layer3_outputs(278);
    layer4_outputs(1642) <= not(layer3_outputs(2180));
    layer4_outputs(1643) <= (layer3_outputs(721)) or (layer3_outputs(2446));
    layer4_outputs(1644) <= not((layer3_outputs(275)) or (layer3_outputs(742)));
    layer4_outputs(1645) <= (layer3_outputs(2533)) or (layer3_outputs(145));
    layer4_outputs(1646) <= layer3_outputs(1776);
    layer4_outputs(1647) <= not((layer3_outputs(118)) and (layer3_outputs(2532)));
    layer4_outputs(1648) <= not(layer3_outputs(1424));
    layer4_outputs(1649) <= not((layer3_outputs(637)) and (layer3_outputs(2348)));
    layer4_outputs(1650) <= not(layer3_outputs(527));
    layer4_outputs(1651) <= layer3_outputs(2130);
    layer4_outputs(1652) <= not(layer3_outputs(559));
    layer4_outputs(1653) <= not(layer3_outputs(1385));
    layer4_outputs(1654) <= not(layer3_outputs(1158)) or (layer3_outputs(974));
    layer4_outputs(1655) <= (layer3_outputs(1086)) and (layer3_outputs(2147));
    layer4_outputs(1656) <= not(layer3_outputs(1863));
    layer4_outputs(1657) <= layer3_outputs(1628);
    layer4_outputs(1658) <= not((layer3_outputs(1148)) xor (layer3_outputs(1137)));
    layer4_outputs(1659) <= not(layer3_outputs(1678));
    layer4_outputs(1660) <= not(layer3_outputs(2550));
    layer4_outputs(1661) <= layer3_outputs(1311);
    layer4_outputs(1662) <= (layer3_outputs(1636)) and not (layer3_outputs(2019));
    layer4_outputs(1663) <= not(layer3_outputs(655));
    layer4_outputs(1664) <= layer3_outputs(570);
    layer4_outputs(1665) <= layer3_outputs(1766);
    layer4_outputs(1666) <= (layer3_outputs(386)) and not (layer3_outputs(1428));
    layer4_outputs(1667) <= not((layer3_outputs(231)) or (layer3_outputs(910)));
    layer4_outputs(1668) <= not((layer3_outputs(1568)) xor (layer3_outputs(1431)));
    layer4_outputs(1669) <= not((layer3_outputs(1657)) xor (layer3_outputs(2480)));
    layer4_outputs(1670) <= layer3_outputs(2029);
    layer4_outputs(1671) <= (layer3_outputs(2010)) and not (layer3_outputs(376));
    layer4_outputs(1672) <= (layer3_outputs(2381)) and not (layer3_outputs(805));
    layer4_outputs(1673) <= not(layer3_outputs(393));
    layer4_outputs(1674) <= layer3_outputs(345);
    layer4_outputs(1675) <= layer3_outputs(1984);
    layer4_outputs(1676) <= not(layer3_outputs(2495)) or (layer3_outputs(1153));
    layer4_outputs(1677) <= not((layer3_outputs(854)) xor (layer3_outputs(451)));
    layer4_outputs(1678) <= not((layer3_outputs(2017)) xor (layer3_outputs(1914)));
    layer4_outputs(1679) <= not(layer3_outputs(2274));
    layer4_outputs(1680) <= not(layer3_outputs(1247)) or (layer3_outputs(522));
    layer4_outputs(1681) <= layer3_outputs(292);
    layer4_outputs(1682) <= layer3_outputs(264);
    layer4_outputs(1683) <= (layer3_outputs(950)) and (layer3_outputs(1161));
    layer4_outputs(1684) <= layer3_outputs(2450);
    layer4_outputs(1685) <= layer3_outputs(106);
    layer4_outputs(1686) <= (layer3_outputs(2275)) and (layer3_outputs(2391));
    layer4_outputs(1687) <= not(layer3_outputs(467));
    layer4_outputs(1688) <= (layer3_outputs(794)) and not (layer3_outputs(297));
    layer4_outputs(1689) <= (layer3_outputs(607)) or (layer3_outputs(269));
    layer4_outputs(1690) <= not(layer3_outputs(147));
    layer4_outputs(1691) <= not(layer3_outputs(1234));
    layer4_outputs(1692) <= (layer3_outputs(1526)) and (layer3_outputs(1377));
    layer4_outputs(1693) <= not((layer3_outputs(32)) or (layer3_outputs(2354)));
    layer4_outputs(1694) <= layer3_outputs(2386);
    layer4_outputs(1695) <= not(layer3_outputs(2508));
    layer4_outputs(1696) <= (layer3_outputs(1448)) and not (layer3_outputs(1687));
    layer4_outputs(1697) <= not(layer3_outputs(1558));
    layer4_outputs(1698) <= layer3_outputs(316);
    layer4_outputs(1699) <= not(layer3_outputs(537)) or (layer3_outputs(376));
    layer4_outputs(1700) <= not(layer3_outputs(1015));
    layer4_outputs(1701) <= not(layer3_outputs(1553));
    layer4_outputs(1702) <= not(layer3_outputs(603));
    layer4_outputs(1703) <= not(layer3_outputs(1658));
    layer4_outputs(1704) <= not(layer3_outputs(329));
    layer4_outputs(1705) <= not(layer3_outputs(752));
    layer4_outputs(1706) <= layer3_outputs(316);
    layer4_outputs(1707) <= not(layer3_outputs(550));
    layer4_outputs(1708) <= layer3_outputs(818);
    layer4_outputs(1709) <= layer3_outputs(73);
    layer4_outputs(1710) <= layer3_outputs(1100);
    layer4_outputs(1711) <= not(layer3_outputs(1065));
    layer4_outputs(1712) <= layer3_outputs(1481);
    layer4_outputs(1713) <= not(layer3_outputs(651));
    layer4_outputs(1714) <= not((layer3_outputs(1407)) and (layer3_outputs(2503)));
    layer4_outputs(1715) <= (layer3_outputs(1177)) and not (layer3_outputs(420));
    layer4_outputs(1716) <= not((layer3_outputs(475)) or (layer3_outputs(1484)));
    layer4_outputs(1717) <= layer3_outputs(1180);
    layer4_outputs(1718) <= not(layer3_outputs(2088));
    layer4_outputs(1719) <= not(layer3_outputs(2318));
    layer4_outputs(1720) <= layer3_outputs(236);
    layer4_outputs(1721) <= layer3_outputs(985);
    layer4_outputs(1722) <= not(layer3_outputs(2400));
    layer4_outputs(1723) <= layer3_outputs(1765);
    layer4_outputs(1724) <= not(layer3_outputs(2319)) or (layer3_outputs(1432));
    layer4_outputs(1725) <= (layer3_outputs(137)) and not (layer3_outputs(2469));
    layer4_outputs(1726) <= not((layer3_outputs(2306)) or (layer3_outputs(1818)));
    layer4_outputs(1727) <= not(layer3_outputs(585));
    layer4_outputs(1728) <= layer3_outputs(1144);
    layer4_outputs(1729) <= layer3_outputs(286);
    layer4_outputs(1730) <= not((layer3_outputs(1710)) xor (layer3_outputs(1772)));
    layer4_outputs(1731) <= not(layer3_outputs(616)) or (layer3_outputs(1952));
    layer4_outputs(1732) <= layer3_outputs(206);
    layer4_outputs(1733) <= not((layer3_outputs(1535)) xor (layer3_outputs(16)));
    layer4_outputs(1734) <= (layer3_outputs(479)) and not (layer3_outputs(190));
    layer4_outputs(1735) <= not(layer3_outputs(1119));
    layer4_outputs(1736) <= not(layer3_outputs(204));
    layer4_outputs(1737) <= not(layer3_outputs(178));
    layer4_outputs(1738) <= not((layer3_outputs(1319)) and (layer3_outputs(1599)));
    layer4_outputs(1739) <= not(layer3_outputs(147));
    layer4_outputs(1740) <= layer3_outputs(1543);
    layer4_outputs(1741) <= layer3_outputs(1708);
    layer4_outputs(1742) <= layer3_outputs(2132);
    layer4_outputs(1743) <= (layer3_outputs(1223)) and not (layer3_outputs(1965));
    layer4_outputs(1744) <= not((layer3_outputs(710)) and (layer3_outputs(1001)));
    layer4_outputs(1745) <= (layer3_outputs(177)) and (layer3_outputs(1406));
    layer4_outputs(1746) <= layer3_outputs(2083);
    layer4_outputs(1747) <= layer3_outputs(711);
    layer4_outputs(1748) <= (layer3_outputs(726)) and (layer3_outputs(1903));
    layer4_outputs(1749) <= not(layer3_outputs(1184));
    layer4_outputs(1750) <= layer3_outputs(994);
    layer4_outputs(1751) <= layer3_outputs(386);
    layer4_outputs(1752) <= (layer3_outputs(1932)) and not (layer3_outputs(575));
    layer4_outputs(1753) <= not(layer3_outputs(1246));
    layer4_outputs(1754) <= layer3_outputs(2034);
    layer4_outputs(1755) <= layer3_outputs(953);
    layer4_outputs(1756) <= layer3_outputs(560);
    layer4_outputs(1757) <= not((layer3_outputs(1823)) or (layer3_outputs(1268)));
    layer4_outputs(1758) <= (layer3_outputs(1598)) and not (layer3_outputs(1351));
    layer4_outputs(1759) <= layer3_outputs(1309);
    layer4_outputs(1760) <= not(layer3_outputs(651));
    layer4_outputs(1761) <= not(layer3_outputs(453)) or (layer3_outputs(49));
    layer4_outputs(1762) <= (layer3_outputs(544)) or (layer3_outputs(1698));
    layer4_outputs(1763) <= layer3_outputs(2458);
    layer4_outputs(1764) <= layer3_outputs(2011);
    layer4_outputs(1765) <= not(layer3_outputs(2063));
    layer4_outputs(1766) <= not(layer3_outputs(2055));
    layer4_outputs(1767) <= layer3_outputs(2080);
    layer4_outputs(1768) <= layer3_outputs(1922);
    layer4_outputs(1769) <= (layer3_outputs(1168)) and not (layer3_outputs(1756));
    layer4_outputs(1770) <= layer3_outputs(107);
    layer4_outputs(1771) <= (layer3_outputs(1879)) and not (layer3_outputs(1282));
    layer4_outputs(1772) <= not((layer3_outputs(2365)) xor (layer3_outputs(242)));
    layer4_outputs(1773) <= not(layer3_outputs(1667));
    layer4_outputs(1774) <= layer3_outputs(2440);
    layer4_outputs(1775) <= layer3_outputs(1730);
    layer4_outputs(1776) <= (layer3_outputs(1950)) and not (layer3_outputs(1205));
    layer4_outputs(1777) <= (layer3_outputs(780)) and not (layer3_outputs(2051));
    layer4_outputs(1778) <= not(layer3_outputs(875)) or (layer3_outputs(1180));
    layer4_outputs(1779) <= not((layer3_outputs(1174)) and (layer3_outputs(726)));
    layer4_outputs(1780) <= layer3_outputs(1726);
    layer4_outputs(1781) <= not(layer3_outputs(2395));
    layer4_outputs(1782) <= not(layer3_outputs(831)) or (layer3_outputs(1070));
    layer4_outputs(1783) <= layer3_outputs(2420);
    layer4_outputs(1784) <= not((layer3_outputs(1715)) or (layer3_outputs(1833)));
    layer4_outputs(1785) <= layer3_outputs(579);
    layer4_outputs(1786) <= not(layer3_outputs(2061));
    layer4_outputs(1787) <= layer3_outputs(1914);
    layer4_outputs(1788) <= not(layer3_outputs(1643));
    layer4_outputs(1789) <= layer3_outputs(1463);
    layer4_outputs(1790) <= layer3_outputs(1010);
    layer4_outputs(1791) <= (layer3_outputs(270)) or (layer3_outputs(2094));
    layer4_outputs(1792) <= not(layer3_outputs(2096)) or (layer3_outputs(1002));
    layer4_outputs(1793) <= not(layer3_outputs(2320));
    layer4_outputs(1794) <= layer3_outputs(2364);
    layer4_outputs(1795) <= not((layer3_outputs(541)) or (layer3_outputs(2427)));
    layer4_outputs(1796) <= not(layer3_outputs(2139));
    layer4_outputs(1797) <= not(layer3_outputs(1881)) or (layer3_outputs(934));
    layer4_outputs(1798) <= (layer3_outputs(1945)) and not (layer3_outputs(1441));
    layer4_outputs(1799) <= not(layer3_outputs(2345));
    layer4_outputs(1800) <= layer3_outputs(1970);
    layer4_outputs(1801) <= layer3_outputs(1172);
    layer4_outputs(1802) <= layer3_outputs(1127);
    layer4_outputs(1803) <= not((layer3_outputs(768)) xor (layer3_outputs(1548)));
    layer4_outputs(1804) <= not(layer3_outputs(2115)) or (layer3_outputs(351));
    layer4_outputs(1805) <= not(layer3_outputs(861));
    layer4_outputs(1806) <= not(layer3_outputs(278));
    layer4_outputs(1807) <= not((layer3_outputs(175)) and (layer3_outputs(1816)));
    layer4_outputs(1808) <= not(layer3_outputs(1918)) or (layer3_outputs(2292));
    layer4_outputs(1809) <= not(layer3_outputs(66)) or (layer3_outputs(1244));
    layer4_outputs(1810) <= layer3_outputs(967);
    layer4_outputs(1811) <= not((layer3_outputs(818)) and (layer3_outputs(1082)));
    layer4_outputs(1812) <= (layer3_outputs(1690)) or (layer3_outputs(1003));
    layer4_outputs(1813) <= not(layer3_outputs(905));
    layer4_outputs(1814) <= (layer3_outputs(1839)) or (layer3_outputs(493));
    layer4_outputs(1815) <= not((layer3_outputs(187)) and (layer3_outputs(1266)));
    layer4_outputs(1816) <= not(layer3_outputs(555)) or (layer3_outputs(1128));
    layer4_outputs(1817) <= not(layer3_outputs(1583));
    layer4_outputs(1818) <= layer3_outputs(1943);
    layer4_outputs(1819) <= not(layer3_outputs(1523));
    layer4_outputs(1820) <= not((layer3_outputs(133)) xor (layer3_outputs(812)));
    layer4_outputs(1821) <= not(layer3_outputs(956));
    layer4_outputs(1822) <= not((layer3_outputs(182)) and (layer3_outputs(1866)));
    layer4_outputs(1823) <= layer3_outputs(1549);
    layer4_outputs(1824) <= (layer3_outputs(1076)) and not (layer3_outputs(800));
    layer4_outputs(1825) <= layer3_outputs(1470);
    layer4_outputs(1826) <= not((layer3_outputs(1690)) and (layer3_outputs(1476)));
    layer4_outputs(1827) <= not((layer3_outputs(1545)) and (layer3_outputs(989)));
    layer4_outputs(1828) <= not(layer3_outputs(1870)) or (layer3_outputs(1111));
    layer4_outputs(1829) <= layer3_outputs(46);
    layer4_outputs(1830) <= (layer3_outputs(2372)) and not (layer3_outputs(1573));
    layer4_outputs(1831) <= layer3_outputs(2283);
    layer4_outputs(1832) <= (layer3_outputs(1420)) and (layer3_outputs(736));
    layer4_outputs(1833) <= (layer3_outputs(2418)) and (layer3_outputs(1333));
    layer4_outputs(1834) <= not(layer3_outputs(1519));
    layer4_outputs(1835) <= not(layer3_outputs(925)) or (layer3_outputs(220));
    layer4_outputs(1836) <= layer3_outputs(2203);
    layer4_outputs(1837) <= not(layer3_outputs(1527));
    layer4_outputs(1838) <= layer3_outputs(1158);
    layer4_outputs(1839) <= not(layer3_outputs(1870)) or (layer3_outputs(1265));
    layer4_outputs(1840) <= not((layer3_outputs(1868)) xor (layer3_outputs(2064)));
    layer4_outputs(1841) <= not((layer3_outputs(394)) xor (layer3_outputs(762)));
    layer4_outputs(1842) <= (layer3_outputs(2530)) and not (layer3_outputs(1105));
    layer4_outputs(1843) <= not(layer3_outputs(81));
    layer4_outputs(1844) <= not((layer3_outputs(2461)) or (layer3_outputs(1202)));
    layer4_outputs(1845) <= not((layer3_outputs(396)) or (layer3_outputs(648)));
    layer4_outputs(1846) <= not(layer3_outputs(2151));
    layer4_outputs(1847) <= layer3_outputs(1188);
    layer4_outputs(1848) <= not(layer3_outputs(381)) or (layer3_outputs(1555));
    layer4_outputs(1849) <= layer3_outputs(1611);
    layer4_outputs(1850) <= not(layer3_outputs(1325));
    layer4_outputs(1851) <= not(layer3_outputs(1194));
    layer4_outputs(1852) <= layer3_outputs(1820);
    layer4_outputs(1853) <= not((layer3_outputs(640)) and (layer3_outputs(489)));
    layer4_outputs(1854) <= not(layer3_outputs(1806));
    layer4_outputs(1855) <= (layer3_outputs(621)) and (layer3_outputs(1711));
    layer4_outputs(1856) <= (layer3_outputs(812)) xor (layer3_outputs(1074));
    layer4_outputs(1857) <= (layer3_outputs(1889)) and (layer3_outputs(1514));
    layer4_outputs(1858) <= not(layer3_outputs(1543));
    layer4_outputs(1859) <= layer3_outputs(1864);
    layer4_outputs(1860) <= (layer3_outputs(1197)) and (layer3_outputs(2475));
    layer4_outputs(1861) <= (layer3_outputs(1819)) and not (layer3_outputs(899));
    layer4_outputs(1862) <= not(layer3_outputs(766));
    layer4_outputs(1863) <= layer3_outputs(997);
    layer4_outputs(1864) <= (layer3_outputs(1713)) and not (layer3_outputs(1259));
    layer4_outputs(1865) <= layer3_outputs(290);
    layer4_outputs(1866) <= not(layer3_outputs(1630)) or (layer3_outputs(1226));
    layer4_outputs(1867) <= not(layer3_outputs(1963)) or (layer3_outputs(1669));
    layer4_outputs(1868) <= not((layer3_outputs(1652)) and (layer3_outputs(624)));
    layer4_outputs(1869) <= not(layer3_outputs(356));
    layer4_outputs(1870) <= (layer3_outputs(107)) and not (layer3_outputs(923));
    layer4_outputs(1871) <= not((layer3_outputs(1985)) or (layer3_outputs(1617)));
    layer4_outputs(1872) <= not(layer3_outputs(963));
    layer4_outputs(1873) <= (layer3_outputs(850)) or (layer3_outputs(203));
    layer4_outputs(1874) <= (layer3_outputs(908)) and (layer3_outputs(1377));
    layer4_outputs(1875) <= '1';
    layer4_outputs(1876) <= (layer3_outputs(753)) and not (layer3_outputs(1375));
    layer4_outputs(1877) <= not(layer3_outputs(1089));
    layer4_outputs(1878) <= layer3_outputs(2474);
    layer4_outputs(1879) <= not(layer3_outputs(1663));
    layer4_outputs(1880) <= layer3_outputs(113);
    layer4_outputs(1881) <= layer3_outputs(1919);
    layer4_outputs(1882) <= (layer3_outputs(403)) xor (layer3_outputs(1677));
    layer4_outputs(1883) <= not(layer3_outputs(2367));
    layer4_outputs(1884) <= not((layer3_outputs(838)) and (layer3_outputs(2545)));
    layer4_outputs(1885) <= not((layer3_outputs(1791)) or (layer3_outputs(2129)));
    layer4_outputs(1886) <= (layer3_outputs(1499)) or (layer3_outputs(2206));
    layer4_outputs(1887) <= not(layer3_outputs(848));
    layer4_outputs(1888) <= not((layer3_outputs(2270)) or (layer3_outputs(1644)));
    layer4_outputs(1889) <= not(layer3_outputs(319));
    layer4_outputs(1890) <= not((layer3_outputs(1308)) and (layer3_outputs(1734)));
    layer4_outputs(1891) <= not((layer3_outputs(258)) or (layer3_outputs(808)));
    layer4_outputs(1892) <= not(layer3_outputs(2145));
    layer4_outputs(1893) <= not(layer3_outputs(1591)) or (layer3_outputs(423));
    layer4_outputs(1894) <= '0';
    layer4_outputs(1895) <= layer3_outputs(2357);
    layer4_outputs(1896) <= not((layer3_outputs(1847)) or (layer3_outputs(1437)));
    layer4_outputs(1897) <= not(layer3_outputs(471)) or (layer3_outputs(214));
    layer4_outputs(1898) <= not((layer3_outputs(282)) xor (layer3_outputs(1414)));
    layer4_outputs(1899) <= not(layer3_outputs(1494));
    layer4_outputs(1900) <= not(layer3_outputs(2047));
    layer4_outputs(1901) <= not(layer3_outputs(2026));
    layer4_outputs(1902) <= not(layer3_outputs(760));
    layer4_outputs(1903) <= not(layer3_outputs(790));
    layer4_outputs(1904) <= '1';
    layer4_outputs(1905) <= layer3_outputs(1369);
    layer4_outputs(1906) <= layer3_outputs(1909);
    layer4_outputs(1907) <= not((layer3_outputs(2398)) and (layer3_outputs(151)));
    layer4_outputs(1908) <= not(layer3_outputs(1745));
    layer4_outputs(1909) <= (layer3_outputs(1207)) and not (layer3_outputs(717));
    layer4_outputs(1910) <= not(layer3_outputs(1635));
    layer4_outputs(1911) <= (layer3_outputs(80)) and (layer3_outputs(2451));
    layer4_outputs(1912) <= '0';
    layer4_outputs(1913) <= not((layer3_outputs(1675)) xor (layer3_outputs(466)));
    layer4_outputs(1914) <= not(layer3_outputs(1564));
    layer4_outputs(1915) <= not((layer3_outputs(1891)) or (layer3_outputs(2250)));
    layer4_outputs(1916) <= layer3_outputs(105);
    layer4_outputs(1917) <= (layer3_outputs(647)) and (layer3_outputs(2449));
    layer4_outputs(1918) <= (layer3_outputs(1098)) and not (layer3_outputs(1412));
    layer4_outputs(1919) <= not((layer3_outputs(701)) or (layer3_outputs(2470)));
    layer4_outputs(1920) <= layer3_outputs(991);
    layer4_outputs(1921) <= layer3_outputs(1835);
    layer4_outputs(1922) <= not(layer3_outputs(782));
    layer4_outputs(1923) <= (layer3_outputs(1933)) xor (layer3_outputs(1452));
    layer4_outputs(1924) <= (layer3_outputs(296)) or (layer3_outputs(190));
    layer4_outputs(1925) <= not(layer3_outputs(2118));
    layer4_outputs(1926) <= (layer3_outputs(569)) and (layer3_outputs(1313));
    layer4_outputs(1927) <= not(layer3_outputs(2000)) or (layer3_outputs(1915));
    layer4_outputs(1928) <= '0';
    layer4_outputs(1929) <= (layer3_outputs(2298)) or (layer3_outputs(1522));
    layer4_outputs(1930) <= not((layer3_outputs(254)) and (layer3_outputs(1610)));
    layer4_outputs(1931) <= (layer3_outputs(1019)) and (layer3_outputs(1671));
    layer4_outputs(1932) <= layer3_outputs(1006);
    layer4_outputs(1933) <= layer3_outputs(1504);
    layer4_outputs(1934) <= layer3_outputs(8);
    layer4_outputs(1935) <= not(layer3_outputs(2430));
    layer4_outputs(1936) <= (layer3_outputs(2023)) or (layer3_outputs(987));
    layer4_outputs(1937) <= not(layer3_outputs(132));
    layer4_outputs(1938) <= not(layer3_outputs(554));
    layer4_outputs(1939) <= layer3_outputs(658);
    layer4_outputs(1940) <= not((layer3_outputs(76)) and (layer3_outputs(876)));
    layer4_outputs(1941) <= not(layer3_outputs(2047));
    layer4_outputs(1942) <= layer3_outputs(606);
    layer4_outputs(1943) <= layer3_outputs(1628);
    layer4_outputs(1944) <= not(layer3_outputs(1052)) or (layer3_outputs(2251));
    layer4_outputs(1945) <= not((layer3_outputs(1614)) xor (layer3_outputs(2221)));
    layer4_outputs(1946) <= layer3_outputs(401);
    layer4_outputs(1947) <= not(layer3_outputs(1771));
    layer4_outputs(1948) <= layer3_outputs(1307);
    layer4_outputs(1949) <= not(layer3_outputs(2554));
    layer4_outputs(1950) <= not(layer3_outputs(1738));
    layer4_outputs(1951) <= not(layer3_outputs(715));
    layer4_outputs(1952) <= (layer3_outputs(2109)) or (layer3_outputs(834));
    layer4_outputs(1953) <= layer3_outputs(2441);
    layer4_outputs(1954) <= not((layer3_outputs(900)) xor (layer3_outputs(1048)));
    layer4_outputs(1955) <= layer3_outputs(1040);
    layer4_outputs(1956) <= not(layer3_outputs(16)) or (layer3_outputs(127));
    layer4_outputs(1957) <= layer3_outputs(1822);
    layer4_outputs(1958) <= '1';
    layer4_outputs(1959) <= layer3_outputs(2340);
    layer4_outputs(1960) <= not((layer3_outputs(524)) xor (layer3_outputs(1959)));
    layer4_outputs(1961) <= not((layer3_outputs(2460)) xor (layer3_outputs(1626)));
    layer4_outputs(1962) <= (layer3_outputs(2104)) and not (layer3_outputs(2094));
    layer4_outputs(1963) <= '0';
    layer4_outputs(1964) <= layer3_outputs(1578);
    layer4_outputs(1965) <= not(layer3_outputs(1986)) or (layer3_outputs(442));
    layer4_outputs(1966) <= not(layer3_outputs(1871)) or (layer3_outputs(2277));
    layer4_outputs(1967) <= layer3_outputs(884);
    layer4_outputs(1968) <= not(layer3_outputs(2057));
    layer4_outputs(1969) <= layer3_outputs(810);
    layer4_outputs(1970) <= not((layer3_outputs(109)) xor (layer3_outputs(710)));
    layer4_outputs(1971) <= not((layer3_outputs(259)) and (layer3_outputs(1964)));
    layer4_outputs(1972) <= (layer3_outputs(335)) and not (layer3_outputs(1314));
    layer4_outputs(1973) <= (layer3_outputs(1804)) and (layer3_outputs(2163));
    layer4_outputs(1974) <= layer3_outputs(594);
    layer4_outputs(1975) <= layer3_outputs(519);
    layer4_outputs(1976) <= not(layer3_outputs(30));
    layer4_outputs(1977) <= layer3_outputs(937);
    layer4_outputs(1978) <= layer3_outputs(1533);
    layer4_outputs(1979) <= (layer3_outputs(1966)) and not (layer3_outputs(1164));
    layer4_outputs(1980) <= not((layer3_outputs(2195)) xor (layer3_outputs(62)));
    layer4_outputs(1981) <= not(layer3_outputs(2302));
    layer4_outputs(1982) <= not(layer3_outputs(1910)) or (layer3_outputs(2164));
    layer4_outputs(1983) <= layer3_outputs(2109);
    layer4_outputs(1984) <= (layer3_outputs(926)) xor (layer3_outputs(862));
    layer4_outputs(1985) <= not(layer3_outputs(1456));
    layer4_outputs(1986) <= not(layer3_outputs(1401));
    layer4_outputs(1987) <= not(layer3_outputs(323)) or (layer3_outputs(1132));
    layer4_outputs(1988) <= (layer3_outputs(2287)) and not (layer3_outputs(503));
    layer4_outputs(1989) <= (layer3_outputs(644)) or (layer3_outputs(523));
    layer4_outputs(1990) <= (layer3_outputs(106)) and not (layer3_outputs(75));
    layer4_outputs(1991) <= not(layer3_outputs(1209));
    layer4_outputs(1992) <= (layer3_outputs(856)) and not (layer3_outputs(1399));
    layer4_outputs(1993) <= not((layer3_outputs(2263)) and (layer3_outputs(354)));
    layer4_outputs(1994) <= not(layer3_outputs(736));
    layer4_outputs(1995) <= (layer3_outputs(1310)) and not (layer3_outputs(1590));
    layer4_outputs(1996) <= layer3_outputs(792);
    layer4_outputs(1997) <= not(layer3_outputs(1974));
    layer4_outputs(1998) <= (layer3_outputs(85)) and (layer3_outputs(2212));
    layer4_outputs(1999) <= not((layer3_outputs(1827)) xor (layer3_outputs(1587)));
    layer4_outputs(2000) <= not(layer3_outputs(2374)) or (layer3_outputs(1802));
    layer4_outputs(2001) <= not((layer3_outputs(1772)) xor (layer3_outputs(53)));
    layer4_outputs(2002) <= not(layer3_outputs(2071)) or (layer3_outputs(154));
    layer4_outputs(2003) <= not((layer3_outputs(1843)) or (layer3_outputs(1057)));
    layer4_outputs(2004) <= not(layer3_outputs(185));
    layer4_outputs(2005) <= (layer3_outputs(433)) and not (layer3_outputs(2044));
    layer4_outputs(2006) <= (layer3_outputs(2032)) and not (layer3_outputs(408));
    layer4_outputs(2007) <= (layer3_outputs(2198)) xor (layer3_outputs(318));
    layer4_outputs(2008) <= layer3_outputs(1439);
    layer4_outputs(2009) <= (layer3_outputs(999)) and (layer3_outputs(774));
    layer4_outputs(2010) <= (layer3_outputs(213)) or (layer3_outputs(2509));
    layer4_outputs(2011) <= (layer3_outputs(1566)) xor (layer3_outputs(2023));
    layer4_outputs(2012) <= (layer3_outputs(2528)) and (layer3_outputs(74));
    layer4_outputs(2013) <= layer3_outputs(697);
    layer4_outputs(2014) <= layer3_outputs(1445);
    layer4_outputs(2015) <= not(layer3_outputs(413));
    layer4_outputs(2016) <= not((layer3_outputs(1054)) and (layer3_outputs(1458)));
    layer4_outputs(2017) <= layer3_outputs(2325);
    layer4_outputs(2018) <= not(layer3_outputs(1596)) or (layer3_outputs(1867));
    layer4_outputs(2019) <= not(layer3_outputs(1682));
    layer4_outputs(2020) <= layer3_outputs(728);
    layer4_outputs(2021) <= not((layer3_outputs(842)) or (layer3_outputs(1077)));
    layer4_outputs(2022) <= not(layer3_outputs(2085));
    layer4_outputs(2023) <= layer3_outputs(1494);
    layer4_outputs(2024) <= (layer3_outputs(1419)) and not (layer3_outputs(1342));
    layer4_outputs(2025) <= layer3_outputs(1683);
    layer4_outputs(2026) <= layer3_outputs(380);
    layer4_outputs(2027) <= layer3_outputs(343);
    layer4_outputs(2028) <= not(layer3_outputs(2360));
    layer4_outputs(2029) <= not((layer3_outputs(1043)) xor (layer3_outputs(1194)));
    layer4_outputs(2030) <= (layer3_outputs(1788)) and (layer3_outputs(400));
    layer4_outputs(2031) <= layer3_outputs(1401);
    layer4_outputs(2032) <= not(layer3_outputs(2288));
    layer4_outputs(2033) <= (layer3_outputs(373)) and not (layer3_outputs(1445));
    layer4_outputs(2034) <= layer3_outputs(541);
    layer4_outputs(2035) <= layer3_outputs(615);
    layer4_outputs(2036) <= not(layer3_outputs(603)) or (layer3_outputs(464));
    layer4_outputs(2037) <= (layer3_outputs(2526)) and not (layer3_outputs(1085));
    layer4_outputs(2038) <= not(layer3_outputs(959)) or (layer3_outputs(1777));
    layer4_outputs(2039) <= (layer3_outputs(739)) xor (layer3_outputs(315));
    layer4_outputs(2040) <= (layer3_outputs(2282)) and (layer3_outputs(274));
    layer4_outputs(2041) <= not(layer3_outputs(1978));
    layer4_outputs(2042) <= not(layer3_outputs(1973));
    layer4_outputs(2043) <= layer3_outputs(775);
    layer4_outputs(2044) <= layer3_outputs(1280);
    layer4_outputs(2045) <= not((layer3_outputs(636)) or (layer3_outputs(516)));
    layer4_outputs(2046) <= layer3_outputs(1618);
    layer4_outputs(2047) <= (layer3_outputs(336)) or (layer3_outputs(770));
    layer4_outputs(2048) <= not(layer3_outputs(1506)) or (layer3_outputs(2095));
    layer4_outputs(2049) <= not(layer3_outputs(1359));
    layer4_outputs(2050) <= not(layer3_outputs(2403)) or (layer3_outputs(2105));
    layer4_outputs(2051) <= (layer3_outputs(1642)) and not (layer3_outputs(1385));
    layer4_outputs(2052) <= (layer3_outputs(2089)) xor (layer3_outputs(418));
    layer4_outputs(2053) <= (layer3_outputs(2329)) and not (layer3_outputs(1905));
    layer4_outputs(2054) <= layer3_outputs(1762);
    layer4_outputs(2055) <= not(layer3_outputs(114));
    layer4_outputs(2056) <= (layer3_outputs(288)) and not (layer3_outputs(689));
    layer4_outputs(2057) <= (layer3_outputs(465)) and (layer3_outputs(1292));
    layer4_outputs(2058) <= layer3_outputs(706);
    layer4_outputs(2059) <= not((layer3_outputs(668)) or (layer3_outputs(2049)));
    layer4_outputs(2060) <= (layer3_outputs(292)) and not (layer3_outputs(1823));
    layer4_outputs(2061) <= layer3_outputs(1266);
    layer4_outputs(2062) <= layer3_outputs(922);
    layer4_outputs(2063) <= not((layer3_outputs(1475)) and (layer3_outputs(634)));
    layer4_outputs(2064) <= '0';
    layer4_outputs(2065) <= not(layer3_outputs(2199)) or (layer3_outputs(2334));
    layer4_outputs(2066) <= (layer3_outputs(2276)) and (layer3_outputs(2381));
    layer4_outputs(2067) <= layer3_outputs(87);
    layer4_outputs(2068) <= not(layer3_outputs(1173)) or (layer3_outputs(1124));
    layer4_outputs(2069) <= (layer3_outputs(724)) and not (layer3_outputs(1454));
    layer4_outputs(2070) <= layer3_outputs(1767);
    layer4_outputs(2071) <= not(layer3_outputs(1409));
    layer4_outputs(2072) <= (layer3_outputs(2204)) and not (layer3_outputs(1668));
    layer4_outputs(2073) <= not(layer3_outputs(954));
    layer4_outputs(2074) <= not(layer3_outputs(1586)) or (layer3_outputs(1351));
    layer4_outputs(2075) <= layer3_outputs(1836);
    layer4_outputs(2076) <= (layer3_outputs(2077)) or (layer3_outputs(1880));
    layer4_outputs(2077) <= not(layer3_outputs(1646));
    layer4_outputs(2078) <= '1';
    layer4_outputs(2079) <= layer3_outputs(1920);
    layer4_outputs(2080) <= not(layer3_outputs(1240));
    layer4_outputs(2081) <= not((layer3_outputs(733)) or (layer3_outputs(69)));
    layer4_outputs(2082) <= (layer3_outputs(130)) or (layer3_outputs(20));
    layer4_outputs(2083) <= not(layer3_outputs(799));
    layer4_outputs(2084) <= layer3_outputs(520);
    layer4_outputs(2085) <= not(layer3_outputs(17));
    layer4_outputs(2086) <= not(layer3_outputs(1556));
    layer4_outputs(2087) <= not(layer3_outputs(1093)) or (layer3_outputs(2549));
    layer4_outputs(2088) <= not(layer3_outputs(423));
    layer4_outputs(2089) <= layer3_outputs(2036);
    layer4_outputs(2090) <= (layer3_outputs(1757)) or (layer3_outputs(659));
    layer4_outputs(2091) <= (layer3_outputs(1847)) and not (layer3_outputs(546));
    layer4_outputs(2092) <= layer3_outputs(2321);
    layer4_outputs(2093) <= not(layer3_outputs(1224));
    layer4_outputs(2094) <= not((layer3_outputs(2350)) xor (layer3_outputs(2501)));
    layer4_outputs(2095) <= '0';
    layer4_outputs(2096) <= (layer3_outputs(2254)) and (layer3_outputs(1444));
    layer4_outputs(2097) <= not((layer3_outputs(1858)) and (layer3_outputs(1750)));
    layer4_outputs(2098) <= not(layer3_outputs(1513)) or (layer3_outputs(819));
    layer4_outputs(2099) <= layer3_outputs(213);
    layer4_outputs(2100) <= layer3_outputs(1435);
    layer4_outputs(2101) <= (layer3_outputs(1790)) and not (layer3_outputs(256));
    layer4_outputs(2102) <= layer3_outputs(1700);
    layer4_outputs(2103) <= layer3_outputs(351);
    layer4_outputs(2104) <= '1';
    layer4_outputs(2105) <= layer3_outputs(1850);
    layer4_outputs(2106) <= not(layer3_outputs(2088));
    layer4_outputs(2107) <= (layer3_outputs(419)) and (layer3_outputs(1738));
    layer4_outputs(2108) <= not((layer3_outputs(1640)) or (layer3_outputs(2308)));
    layer4_outputs(2109) <= (layer3_outputs(1788)) or (layer3_outputs(1951));
    layer4_outputs(2110) <= not(layer3_outputs(1528)) or (layer3_outputs(568));
    layer4_outputs(2111) <= layer3_outputs(417);
    layer4_outputs(2112) <= (layer3_outputs(113)) and not (layer3_outputs(1743));
    layer4_outputs(2113) <= not(layer3_outputs(1422));
    layer4_outputs(2114) <= not(layer3_outputs(1937));
    layer4_outputs(2115) <= not(layer3_outputs(1931)) or (layer3_outputs(1315));
    layer4_outputs(2116) <= not(layer3_outputs(367));
    layer4_outputs(2117) <= not(layer3_outputs(547));
    layer4_outputs(2118) <= layer3_outputs(1041);
    layer4_outputs(2119) <= not((layer3_outputs(934)) and (layer3_outputs(2101)));
    layer4_outputs(2120) <= (layer3_outputs(661)) and not (layer3_outputs(1827));
    layer4_outputs(2121) <= not(layer3_outputs(32));
    layer4_outputs(2122) <= (layer3_outputs(1799)) and not (layer3_outputs(552));
    layer4_outputs(2123) <= layer3_outputs(1719);
    layer4_outputs(2124) <= not(layer3_outputs(473));
    layer4_outputs(2125) <= (layer3_outputs(1075)) and (layer3_outputs(100));
    layer4_outputs(2126) <= not(layer3_outputs(591));
    layer4_outputs(2127) <= not(layer3_outputs(236));
    layer4_outputs(2128) <= not(layer3_outputs(1232));
    layer4_outputs(2129) <= not(layer3_outputs(2266));
    layer4_outputs(2130) <= (layer3_outputs(608)) and not (layer3_outputs(623));
    layer4_outputs(2131) <= (layer3_outputs(902)) or (layer3_outputs(1229));
    layer4_outputs(2132) <= not(layer3_outputs(149)) or (layer3_outputs(811));
    layer4_outputs(2133) <= layer3_outputs(82);
    layer4_outputs(2134) <= not(layer3_outputs(939)) or (layer3_outputs(2008));
    layer4_outputs(2135) <= layer3_outputs(1660);
    layer4_outputs(2136) <= layer3_outputs(1146);
    layer4_outputs(2137) <= (layer3_outputs(1106)) xor (layer3_outputs(1885));
    layer4_outputs(2138) <= layer3_outputs(787);
    layer4_outputs(2139) <= layer3_outputs(1728);
    layer4_outputs(2140) <= not((layer3_outputs(1704)) or (layer3_outputs(2062)));
    layer4_outputs(2141) <= not((layer3_outputs(919)) xor (layer3_outputs(174)));
    layer4_outputs(2142) <= layer3_outputs(529);
    layer4_outputs(2143) <= not(layer3_outputs(346));
    layer4_outputs(2144) <= not(layer3_outputs(936));
    layer4_outputs(2145) <= not(layer3_outputs(2201));
    layer4_outputs(2146) <= (layer3_outputs(1540)) xor (layer3_outputs(2228));
    layer4_outputs(2147) <= '0';
    layer4_outputs(2148) <= not((layer3_outputs(969)) and (layer3_outputs(2556)));
    layer4_outputs(2149) <= not(layer3_outputs(1678));
    layer4_outputs(2150) <= not((layer3_outputs(757)) xor (layer3_outputs(1689)));
    layer4_outputs(2151) <= layer3_outputs(1064);
    layer4_outputs(2152) <= (layer3_outputs(793)) or (layer3_outputs(6));
    layer4_outputs(2153) <= '0';
    layer4_outputs(2154) <= (layer3_outputs(153)) and (layer3_outputs(273));
    layer4_outputs(2155) <= not(layer3_outputs(1783)) or (layer3_outputs(115));
    layer4_outputs(2156) <= not(layer3_outputs(833)) or (layer3_outputs(876));
    layer4_outputs(2157) <= (layer3_outputs(1620)) and not (layer3_outputs(1025));
    layer4_outputs(2158) <= layer3_outputs(491);
    layer4_outputs(2159) <= layer3_outputs(2371);
    layer4_outputs(2160) <= not((layer3_outputs(719)) or (layer3_outputs(182)));
    layer4_outputs(2161) <= (layer3_outputs(2318)) and (layer3_outputs(1794));
    layer4_outputs(2162) <= not(layer3_outputs(1901)) or (layer3_outputs(976));
    layer4_outputs(2163) <= not((layer3_outputs(1441)) or (layer3_outputs(571)));
    layer4_outputs(2164) <= not(layer3_outputs(2476)) or (layer3_outputs(1518));
    layer4_outputs(2165) <= not(layer3_outputs(2376));
    layer4_outputs(2166) <= not((layer3_outputs(1103)) and (layer3_outputs(2358)));
    layer4_outputs(2167) <= (layer3_outputs(2505)) and not (layer3_outputs(2344));
    layer4_outputs(2168) <= not(layer3_outputs(962));
    layer4_outputs(2169) <= layer3_outputs(1231);
    layer4_outputs(2170) <= layer3_outputs(1741);
    layer4_outputs(2171) <= (layer3_outputs(2352)) and (layer3_outputs(1270));
    layer4_outputs(2172) <= not((layer3_outputs(690)) or (layer3_outputs(471)));
    layer4_outputs(2173) <= not(layer3_outputs(553)) or (layer3_outputs(637));
    layer4_outputs(2174) <= layer3_outputs(738);
    layer4_outputs(2175) <= not(layer3_outputs(92));
    layer4_outputs(2176) <= (layer3_outputs(230)) and (layer3_outputs(1570));
    layer4_outputs(2177) <= not(layer3_outputs(2197));
    layer4_outputs(2178) <= not(layer3_outputs(185));
    layer4_outputs(2179) <= layer3_outputs(771);
    layer4_outputs(2180) <= layer3_outputs(1777);
    layer4_outputs(2181) <= (layer3_outputs(2045)) xor (layer3_outputs(1451));
    layer4_outputs(2182) <= layer3_outputs(2387);
    layer4_outputs(2183) <= '0';
    layer4_outputs(2184) <= not((layer3_outputs(1467)) and (layer3_outputs(2082)));
    layer4_outputs(2185) <= layer3_outputs(2358);
    layer4_outputs(2186) <= not(layer3_outputs(1581)) or (layer3_outputs(2079));
    layer4_outputs(2187) <= layer3_outputs(2496);
    layer4_outputs(2188) <= not((layer3_outputs(1793)) or (layer3_outputs(2261)));
    layer4_outputs(2189) <= layer3_outputs(1426);
    layer4_outputs(2190) <= (layer3_outputs(712)) and not (layer3_outputs(992));
    layer4_outputs(2191) <= layer3_outputs(2056);
    layer4_outputs(2192) <= not(layer3_outputs(1789)) or (layer3_outputs(1588));
    layer4_outputs(2193) <= not(layer3_outputs(2139));
    layer4_outputs(2194) <= not(layer3_outputs(475));
    layer4_outputs(2195) <= not(layer3_outputs(1302)) or (layer3_outputs(677));
    layer4_outputs(2196) <= (layer3_outputs(20)) or (layer3_outputs(1732));
    layer4_outputs(2197) <= not(layer3_outputs(1785));
    layer4_outputs(2198) <= not(layer3_outputs(1561));
    layer4_outputs(2199) <= not(layer3_outputs(1784));
    layer4_outputs(2200) <= layer3_outputs(1489);
    layer4_outputs(2201) <= not(layer3_outputs(2320)) or (layer3_outputs(712));
    layer4_outputs(2202) <= not(layer3_outputs(1140));
    layer4_outputs(2203) <= layer3_outputs(858);
    layer4_outputs(2204) <= (layer3_outputs(2016)) and not (layer3_outputs(2451));
    layer4_outputs(2205) <= not(layer3_outputs(747));
    layer4_outputs(2206) <= not(layer3_outputs(9));
    layer4_outputs(2207) <= not(layer3_outputs(22));
    layer4_outputs(2208) <= '1';
    layer4_outputs(2209) <= (layer3_outputs(2207)) or (layer3_outputs(676));
    layer4_outputs(2210) <= (layer3_outputs(2036)) and (layer3_outputs(2552));
    layer4_outputs(2211) <= layer3_outputs(2054);
    layer4_outputs(2212) <= (layer3_outputs(128)) or (layer3_outputs(779));
    layer4_outputs(2213) <= not((layer3_outputs(2363)) or (layer3_outputs(435)));
    layer4_outputs(2214) <= (layer3_outputs(1239)) and not (layer3_outputs(2382));
    layer4_outputs(2215) <= not((layer3_outputs(1364)) or (layer3_outputs(666)));
    layer4_outputs(2216) <= not(layer3_outputs(1099));
    layer4_outputs(2217) <= layer3_outputs(898);
    layer4_outputs(2218) <= layer3_outputs(2492);
    layer4_outputs(2219) <= layer3_outputs(2401);
    layer4_outputs(2220) <= not((layer3_outputs(2359)) xor (layer3_outputs(654)));
    layer4_outputs(2221) <= (layer3_outputs(2035)) or (layer3_outputs(1605));
    layer4_outputs(2222) <= not(layer3_outputs(1645));
    layer4_outputs(2223) <= not((layer3_outputs(2024)) or (layer3_outputs(1191)));
    layer4_outputs(2224) <= (layer3_outputs(2219)) and not (layer3_outputs(21));
    layer4_outputs(2225) <= layer3_outputs(518);
    layer4_outputs(2226) <= not((layer3_outputs(2158)) xor (layer3_outputs(2323)));
    layer4_outputs(2227) <= not((layer3_outputs(2269)) or (layer3_outputs(1869)));
    layer4_outputs(2228) <= layer3_outputs(767);
    layer4_outputs(2229) <= not(layer3_outputs(1172)) or (layer3_outputs(2447));
    layer4_outputs(2230) <= not(layer3_outputs(1968));
    layer4_outputs(2231) <= layer3_outputs(72);
    layer4_outputs(2232) <= layer3_outputs(346);
    layer4_outputs(2233) <= not(layer3_outputs(1664));
    layer4_outputs(2234) <= not(layer3_outputs(2179));
    layer4_outputs(2235) <= (layer3_outputs(632)) and not (layer3_outputs(1321));
    layer4_outputs(2236) <= layer3_outputs(52);
    layer4_outputs(2237) <= layer3_outputs(452);
    layer4_outputs(2238) <= not((layer3_outputs(1477)) or (layer3_outputs(63)));
    layer4_outputs(2239) <= (layer3_outputs(2155)) and not (layer3_outputs(705));
    layer4_outputs(2240) <= not(layer3_outputs(1366)) or (layer3_outputs(564));
    layer4_outputs(2241) <= not(layer3_outputs(310)) or (layer3_outputs(1089));
    layer4_outputs(2242) <= not(layer3_outputs(844));
    layer4_outputs(2243) <= (layer3_outputs(768)) or (layer3_outputs(1254));
    layer4_outputs(2244) <= layer3_outputs(1842);
    layer4_outputs(2245) <= not((layer3_outputs(971)) and (layer3_outputs(449)));
    layer4_outputs(2246) <= not((layer3_outputs(559)) or (layer3_outputs(2160)));
    layer4_outputs(2247) <= not((layer3_outputs(460)) xor (layer3_outputs(1927)));
    layer4_outputs(2248) <= layer3_outputs(479);
    layer4_outputs(2249) <= not((layer3_outputs(1034)) xor (layer3_outputs(1345)));
    layer4_outputs(2250) <= (layer3_outputs(412)) and (layer3_outputs(1114));
    layer4_outputs(2251) <= not(layer3_outputs(1719));
    layer4_outputs(2252) <= not(layer3_outputs(1071));
    layer4_outputs(2253) <= (layer3_outputs(1303)) or (layer3_outputs(2323));
    layer4_outputs(2254) <= not(layer3_outputs(907)) or (layer3_outputs(2233));
    layer4_outputs(2255) <= not(layer3_outputs(1243));
    layer4_outputs(2256) <= '1';
    layer4_outputs(2257) <= not(layer3_outputs(1078));
    layer4_outputs(2258) <= not(layer3_outputs(1382));
    layer4_outputs(2259) <= layer3_outputs(1253);
    layer4_outputs(2260) <= (layer3_outputs(27)) and not (layer3_outputs(23));
    layer4_outputs(2261) <= not(layer3_outputs(940)) or (layer3_outputs(2353));
    layer4_outputs(2262) <= layer3_outputs(2300);
    layer4_outputs(2263) <= (layer3_outputs(1921)) or (layer3_outputs(1984));
    layer4_outputs(2264) <= layer3_outputs(117);
    layer4_outputs(2265) <= not(layer3_outputs(1585));
    layer4_outputs(2266) <= not(layer3_outputs(887));
    layer4_outputs(2267) <= not((layer3_outputs(2209)) xor (layer3_outputs(215)));
    layer4_outputs(2268) <= '1';
    layer4_outputs(2269) <= (layer3_outputs(686)) and not (layer3_outputs(1279));
    layer4_outputs(2270) <= not(layer3_outputs(1016));
    layer4_outputs(2271) <= layer3_outputs(1179);
    layer4_outputs(2272) <= not(layer3_outputs(1248));
    layer4_outputs(2273) <= not(layer3_outputs(2336));
    layer4_outputs(2274) <= layer3_outputs(1507);
    layer4_outputs(2275) <= (layer3_outputs(257)) and not (layer3_outputs(2506));
    layer4_outputs(2276) <= layer3_outputs(14);
    layer4_outputs(2277) <= not(layer3_outputs(1536));
    layer4_outputs(2278) <= not(layer3_outputs(488));
    layer4_outputs(2279) <= not(layer3_outputs(552));
    layer4_outputs(2280) <= layer3_outputs(1433);
    layer4_outputs(2281) <= not(layer3_outputs(962));
    layer4_outputs(2282) <= (layer3_outputs(1436)) and (layer3_outputs(319));
    layer4_outputs(2283) <= (layer3_outputs(5)) and not (layer3_outputs(358));
    layer4_outputs(2284) <= not(layer3_outputs(1278)) or (layer3_outputs(2160));
    layer4_outputs(2285) <= not(layer3_outputs(2370));
    layer4_outputs(2286) <= not(layer3_outputs(447));
    layer4_outputs(2287) <= (layer3_outputs(929)) and (layer3_outputs(1739));
    layer4_outputs(2288) <= (layer3_outputs(1023)) or (layer3_outputs(2269));
    layer4_outputs(2289) <= not(layer3_outputs(1280));
    layer4_outputs(2290) <= not(layer3_outputs(1829)) or (layer3_outputs(1529));
    layer4_outputs(2291) <= (layer3_outputs(101)) and not (layer3_outputs(2210));
    layer4_outputs(2292) <= not(layer3_outputs(678));
    layer4_outputs(2293) <= not(layer3_outputs(1258));
    layer4_outputs(2294) <= (layer3_outputs(2207)) or (layer3_outputs(697));
    layer4_outputs(2295) <= layer3_outputs(2184);
    layer4_outputs(2296) <= not(layer3_outputs(1645));
    layer4_outputs(2297) <= (layer3_outputs(692)) and not (layer3_outputs(675));
    layer4_outputs(2298) <= not((layer3_outputs(562)) and (layer3_outputs(2462)));
    layer4_outputs(2299) <= not(layer3_outputs(1484)) or (layer3_outputs(1941));
    layer4_outputs(2300) <= (layer3_outputs(1560)) or (layer3_outputs(955));
    layer4_outputs(2301) <= (layer3_outputs(456)) and not (layer3_outputs(727));
    layer4_outputs(2302) <= not((layer3_outputs(2007)) xor (layer3_outputs(597)));
    layer4_outputs(2303) <= layer3_outputs(1545);
    layer4_outputs(2304) <= (layer3_outputs(1517)) and not (layer3_outputs(2117));
    layer4_outputs(2305) <= not(layer3_outputs(1622));
    layer4_outputs(2306) <= not(layer3_outputs(567));
    layer4_outputs(2307) <= (layer3_outputs(196)) and (layer3_outputs(91));
    layer4_outputs(2308) <= not((layer3_outputs(370)) and (layer3_outputs(434)));
    layer4_outputs(2309) <= not(layer3_outputs(1142));
    layer4_outputs(2310) <= layer3_outputs(2037);
    layer4_outputs(2311) <= not((layer3_outputs(457)) or (layer3_outputs(1442)));
    layer4_outputs(2312) <= (layer3_outputs(1897)) xor (layer3_outputs(265));
    layer4_outputs(2313) <= not((layer3_outputs(61)) xor (layer3_outputs(2510)));
    layer4_outputs(2314) <= (layer3_outputs(2527)) and not (layer3_outputs(1200));
    layer4_outputs(2315) <= layer3_outputs(310);
    layer4_outputs(2316) <= layer3_outputs(1175);
    layer4_outputs(2317) <= (layer3_outputs(2075)) and not (layer3_outputs(1604));
    layer4_outputs(2318) <= layer3_outputs(430);
    layer4_outputs(2319) <= not(layer3_outputs(2426)) or (layer3_outputs(2293));
    layer4_outputs(2320) <= layer3_outputs(2009);
    layer4_outputs(2321) <= (layer3_outputs(1977)) and (layer3_outputs(220));
    layer4_outputs(2322) <= (layer3_outputs(1108)) and not (layer3_outputs(1289));
    layer4_outputs(2323) <= (layer3_outputs(2002)) xor (layer3_outputs(2035));
    layer4_outputs(2324) <= layer3_outputs(1031);
    layer4_outputs(2325) <= not(layer3_outputs(891));
    layer4_outputs(2326) <= (layer3_outputs(1084)) and not (layer3_outputs(2324));
    layer4_outputs(2327) <= not(layer3_outputs(2172)) or (layer3_outputs(653));
    layer4_outputs(2328) <= (layer3_outputs(1431)) xor (layer3_outputs(2060));
    layer4_outputs(2329) <= layer3_outputs(673);
    layer4_outputs(2330) <= (layer3_outputs(1334)) xor (layer3_outputs(720));
    layer4_outputs(2331) <= (layer3_outputs(2063)) or (layer3_outputs(444));
    layer4_outputs(2332) <= not(layer3_outputs(2395));
    layer4_outputs(2333) <= not(layer3_outputs(1853)) or (layer3_outputs(701));
    layer4_outputs(2334) <= layer3_outputs(2434);
    layer4_outputs(2335) <= not(layer3_outputs(2390));
    layer4_outputs(2336) <= (layer3_outputs(791)) xor (layer3_outputs(2175));
    layer4_outputs(2337) <= layer3_outputs(1241);
    layer4_outputs(2338) <= layer3_outputs(2356);
    layer4_outputs(2339) <= not(layer3_outputs(2033));
    layer4_outputs(2340) <= layer3_outputs(11);
    layer4_outputs(2341) <= not(layer3_outputs(1279)) or (layer3_outputs(255));
    layer4_outputs(2342) <= not(layer3_outputs(15));
    layer4_outputs(2343) <= layer3_outputs(920);
    layer4_outputs(2344) <= layer3_outputs(1875);
    layer4_outputs(2345) <= not((layer3_outputs(505)) and (layer3_outputs(2524)));
    layer4_outputs(2346) <= (layer3_outputs(301)) and not (layer3_outputs(738));
    layer4_outputs(2347) <= not(layer3_outputs(1038)) or (layer3_outputs(1801));
    layer4_outputs(2348) <= not((layer3_outputs(2547)) or (layer3_outputs(1298)));
    layer4_outputs(2349) <= not(layer3_outputs(582));
    layer4_outputs(2350) <= not(layer3_outputs(1090));
    layer4_outputs(2351) <= not(layer3_outputs(1501));
    layer4_outputs(2352) <= (layer3_outputs(919)) and not (layer3_outputs(1988));
    layer4_outputs(2353) <= not(layer3_outputs(326)) or (layer3_outputs(1859));
    layer4_outputs(2354) <= not(layer3_outputs(307)) or (layer3_outputs(146));
    layer4_outputs(2355) <= layer3_outputs(2183);
    layer4_outputs(2356) <= not(layer3_outputs(2324));
    layer4_outputs(2357) <= not(layer3_outputs(2187)) or (layer3_outputs(2428));
    layer4_outputs(2358) <= layer3_outputs(1702);
    layer4_outputs(2359) <= (layer3_outputs(2333)) and not (layer3_outputs(535));
    layer4_outputs(2360) <= layer3_outputs(1081);
    layer4_outputs(2361) <= (layer3_outputs(2027)) and not (layer3_outputs(935));
    layer4_outputs(2362) <= not(layer3_outputs(430));
    layer4_outputs(2363) <= not(layer3_outputs(1527)) or (layer3_outputs(901));
    layer4_outputs(2364) <= not((layer3_outputs(604)) xor (layer3_outputs(1114)));
    layer4_outputs(2365) <= not((layer3_outputs(366)) and (layer3_outputs(847)));
    layer4_outputs(2366) <= layer3_outputs(73);
    layer4_outputs(2367) <= not((layer3_outputs(1961)) xor (layer3_outputs(1995)));
    layer4_outputs(2368) <= not(layer3_outputs(1859));
    layer4_outputs(2369) <= (layer3_outputs(2390)) xor (layer3_outputs(1282));
    layer4_outputs(2370) <= (layer3_outputs(878)) and not (layer3_outputs(176));
    layer4_outputs(2371) <= not(layer3_outputs(1650));
    layer4_outputs(2372) <= not(layer3_outputs(1630));
    layer4_outputs(2373) <= not((layer3_outputs(2336)) xor (layer3_outputs(1991)));
    layer4_outputs(2374) <= (layer3_outputs(1047)) xor (layer3_outputs(2355));
    layer4_outputs(2375) <= (layer3_outputs(1368)) and not (layer3_outputs(835));
    layer4_outputs(2376) <= not((layer3_outputs(578)) or (layer3_outputs(2258)));
    layer4_outputs(2377) <= not(layer3_outputs(598));
    layer4_outputs(2378) <= layer3_outputs(1277);
    layer4_outputs(2379) <= (layer3_outputs(2006)) and (layer3_outputs(1294));
    layer4_outputs(2380) <= (layer3_outputs(1540)) or (layer3_outputs(581));
    layer4_outputs(2381) <= not(layer3_outputs(524));
    layer4_outputs(2382) <= not((layer3_outputs(200)) xor (layer3_outputs(965)));
    layer4_outputs(2383) <= not(layer3_outputs(1922));
    layer4_outputs(2384) <= not(layer3_outputs(223)) or (layer3_outputs(1362));
    layer4_outputs(2385) <= (layer3_outputs(413)) and not (layer3_outputs(2464));
    layer4_outputs(2386) <= not(layer3_outputs(398));
    layer4_outputs(2387) <= not(layer3_outputs(611));
    layer4_outputs(2388) <= not(layer3_outputs(56)) or (layer3_outputs(1179));
    layer4_outputs(2389) <= '1';
    layer4_outputs(2390) <= not(layer3_outputs(2137));
    layer4_outputs(2391) <= not((layer3_outputs(2059)) and (layer3_outputs(2136)));
    layer4_outputs(2392) <= layer3_outputs(2393);
    layer4_outputs(2393) <= not(layer3_outputs(1662)) or (layer3_outputs(641));
    layer4_outputs(2394) <= not((layer3_outputs(168)) xor (layer3_outputs(1459)));
    layer4_outputs(2395) <= not(layer3_outputs(602));
    layer4_outputs(2396) <= layer3_outputs(2504);
    layer4_outputs(2397) <= layer3_outputs(782);
    layer4_outputs(2398) <= (layer3_outputs(1837)) and (layer3_outputs(1983));
    layer4_outputs(2399) <= not(layer3_outputs(784));
    layer4_outputs(2400) <= layer3_outputs(2193);
    layer4_outputs(2401) <= not(layer3_outputs(2527)) or (layer3_outputs(1189));
    layer4_outputs(2402) <= not((layer3_outputs(778)) or (layer3_outputs(181)));
    layer4_outputs(2403) <= layer3_outputs(923);
    layer4_outputs(2404) <= not(layer3_outputs(1284)) or (layer3_outputs(329));
    layer4_outputs(2405) <= not(layer3_outputs(734)) or (layer3_outputs(2483));
    layer4_outputs(2406) <= not((layer3_outputs(36)) or (layer3_outputs(303)));
    layer4_outputs(2407) <= layer3_outputs(1406);
    layer4_outputs(2408) <= (layer3_outputs(909)) xor (layer3_outputs(1679));
    layer4_outputs(2409) <= not(layer3_outputs(570));
    layer4_outputs(2410) <= not(layer3_outputs(1085));
    layer4_outputs(2411) <= not(layer3_outputs(1335));
    layer4_outputs(2412) <= (layer3_outputs(1930)) and not (layer3_outputs(1773));
    layer4_outputs(2413) <= not(layer3_outputs(2159)) or (layer3_outputs(2288));
    layer4_outputs(2414) <= not((layer3_outputs(938)) or (layer3_outputs(155)));
    layer4_outputs(2415) <= not(layer3_outputs(1487));
    layer4_outputs(2416) <= not((layer3_outputs(507)) or (layer3_outputs(1492)));
    layer4_outputs(2417) <= layer3_outputs(1989);
    layer4_outputs(2418) <= not(layer3_outputs(191));
    layer4_outputs(2419) <= not(layer3_outputs(773));
    layer4_outputs(2420) <= (layer3_outputs(377)) and (layer3_outputs(10));
    layer4_outputs(2421) <= layer3_outputs(2505);
    layer4_outputs(2422) <= layer3_outputs(1292);
    layer4_outputs(2423) <= not((layer3_outputs(1747)) and (layer3_outputs(139)));
    layer4_outputs(2424) <= not((layer3_outputs(1384)) or (layer3_outputs(1044)));
    layer4_outputs(2425) <= layer3_outputs(802);
    layer4_outputs(2426) <= not(layer3_outputs(464));
    layer4_outputs(2427) <= not(layer3_outputs(46));
    layer4_outputs(2428) <= not(layer3_outputs(1332)) or (layer3_outputs(2263));
    layer4_outputs(2429) <= layer3_outputs(1297);
    layer4_outputs(2430) <= not(layer3_outputs(2089));
    layer4_outputs(2431) <= (layer3_outputs(1111)) or (layer3_outputs(1839));
    layer4_outputs(2432) <= layer3_outputs(1297);
    layer4_outputs(2433) <= layer3_outputs(1027);
    layer4_outputs(2434) <= not(layer3_outputs(931)) or (layer3_outputs(1037));
    layer4_outputs(2435) <= not(layer3_outputs(604));
    layer4_outputs(2436) <= not(layer3_outputs(1334));
    layer4_outputs(2437) <= layer3_outputs(869);
    layer4_outputs(2438) <= layer3_outputs(209);
    layer4_outputs(2439) <= not(layer3_outputs(1064)) or (layer3_outputs(2529));
    layer4_outputs(2440) <= not(layer3_outputs(614));
    layer4_outputs(2441) <= (layer3_outputs(1157)) and not (layer3_outputs(466));
    layer4_outputs(2442) <= layer3_outputs(2386);
    layer4_outputs(2443) <= (layer3_outputs(1055)) and not (layer3_outputs(425));
    layer4_outputs(2444) <= layer3_outputs(289);
    layer4_outputs(2445) <= (layer3_outputs(1641)) or (layer3_outputs(511));
    layer4_outputs(2446) <= not(layer3_outputs(2077)) or (layer3_outputs(289));
    layer4_outputs(2447) <= not(layer3_outputs(1015));
    layer4_outputs(2448) <= '1';
    layer4_outputs(2449) <= layer3_outputs(2461);
    layer4_outputs(2450) <= not(layer3_outputs(1895)) or (layer3_outputs(1313));
    layer4_outputs(2451) <= layer3_outputs(361);
    layer4_outputs(2452) <= not(layer3_outputs(1185));
    layer4_outputs(2453) <= (layer3_outputs(440)) xor (layer3_outputs(1281));
    layer4_outputs(2454) <= not(layer3_outputs(1130));
    layer4_outputs(2455) <= layer3_outputs(1797);
    layer4_outputs(2456) <= (layer3_outputs(799)) and not (layer3_outputs(2010));
    layer4_outputs(2457) <= layer3_outputs(2359);
    layer4_outputs(2458) <= not(layer3_outputs(1717));
    layer4_outputs(2459) <= not(layer3_outputs(68));
    layer4_outputs(2460) <= (layer3_outputs(364)) or (layer3_outputs(2377));
    layer4_outputs(2461) <= not(layer3_outputs(661));
    layer4_outputs(2462) <= layer3_outputs(789);
    layer4_outputs(2463) <= layer3_outputs(2404);
    layer4_outputs(2464) <= (layer3_outputs(558)) and (layer3_outputs(1306));
    layer4_outputs(2465) <= layer3_outputs(580);
    layer4_outputs(2466) <= layer3_outputs(878);
    layer4_outputs(2467) <= not(layer3_outputs(2060));
    layer4_outputs(2468) <= layer3_outputs(167);
    layer4_outputs(2469) <= not(layer3_outputs(1787));
    layer4_outputs(2470) <= (layer3_outputs(1152)) xor (layer3_outputs(993));
    layer4_outputs(2471) <= not(layer3_outputs(1904)) or (layer3_outputs(1150));
    layer4_outputs(2472) <= layer3_outputs(2225);
    layer4_outputs(2473) <= not(layer3_outputs(2487));
    layer4_outputs(2474) <= not(layer3_outputs(157));
    layer4_outputs(2475) <= not(layer3_outputs(44));
    layer4_outputs(2476) <= not((layer3_outputs(115)) and (layer3_outputs(594)));
    layer4_outputs(2477) <= layer3_outputs(642);
    layer4_outputs(2478) <= not((layer3_outputs(1010)) or (layer3_outputs(796)));
    layer4_outputs(2479) <= not(layer3_outputs(1852)) or (layer3_outputs(1761));
    layer4_outputs(2480) <= not((layer3_outputs(1153)) or (layer3_outputs(1176)));
    layer4_outputs(2481) <= not(layer3_outputs(205));
    layer4_outputs(2482) <= not(layer3_outputs(648)) or (layer3_outputs(481));
    layer4_outputs(2483) <= not((layer3_outputs(241)) or (layer3_outputs(1524)));
    layer4_outputs(2484) <= (layer3_outputs(2138)) and not (layer3_outputs(497));
    layer4_outputs(2485) <= layer3_outputs(2419);
    layer4_outputs(2486) <= not(layer3_outputs(431));
    layer4_outputs(2487) <= (layer3_outputs(1902)) xor (layer3_outputs(558));
    layer4_outputs(2488) <= (layer3_outputs(965)) and not (layer3_outputs(1440));
    layer4_outputs(2489) <= not(layer3_outputs(1600));
    layer4_outputs(2490) <= layer3_outputs(179);
    layer4_outputs(2491) <= '0';
    layer4_outputs(2492) <= not((layer3_outputs(2248)) or (layer3_outputs(1477)));
    layer4_outputs(2493) <= not(layer3_outputs(2086));
    layer4_outputs(2494) <= layer3_outputs(3);
    layer4_outputs(2495) <= not((layer3_outputs(2048)) xor (layer3_outputs(631)));
    layer4_outputs(2496) <= not(layer3_outputs(1778)) or (layer3_outputs(2241));
    layer4_outputs(2497) <= not(layer3_outputs(2387));
    layer4_outputs(2498) <= layer3_outputs(619);
    layer4_outputs(2499) <= not(layer3_outputs(822));
    layer4_outputs(2500) <= not((layer3_outputs(1138)) or (layer3_outputs(2483)));
    layer4_outputs(2501) <= not((layer3_outputs(1675)) or (layer3_outputs(1416)));
    layer4_outputs(2502) <= not(layer3_outputs(511));
    layer4_outputs(2503) <= not(layer3_outputs(2017)) or (layer3_outputs(1998));
    layer4_outputs(2504) <= not(layer3_outputs(396)) or (layer3_outputs(2106));
    layer4_outputs(2505) <= not(layer3_outputs(1208));
    layer4_outputs(2506) <= layer3_outputs(954);
    layer4_outputs(2507) <= not(layer3_outputs(653));
    layer4_outputs(2508) <= not(layer3_outputs(1957));
    layer4_outputs(2509) <= layer3_outputs(505);
    layer4_outputs(2510) <= not(layer3_outputs(1882)) or (layer3_outputs(1099));
    layer4_outputs(2511) <= (layer3_outputs(2090)) or (layer3_outputs(2298));
    layer4_outputs(2512) <= not(layer3_outputs(1565));
    layer4_outputs(2513) <= not(layer3_outputs(1595));
    layer4_outputs(2514) <= not((layer3_outputs(1233)) and (layer3_outputs(540)));
    layer4_outputs(2515) <= not(layer3_outputs(1760));
    layer4_outputs(2516) <= layer3_outputs(2456);
    layer4_outputs(2517) <= not(layer3_outputs(2389));
    layer4_outputs(2518) <= not((layer3_outputs(2241)) or (layer3_outputs(1648)));
    layer4_outputs(2519) <= layer3_outputs(383);
    layer4_outputs(2520) <= layer3_outputs(821);
    layer4_outputs(2521) <= not((layer3_outputs(2135)) or (layer3_outputs(152)));
    layer4_outputs(2522) <= not(layer3_outputs(1940)) or (layer3_outputs(2383));
    layer4_outputs(2523) <= (layer3_outputs(313)) and (layer3_outputs(2513));
    layer4_outputs(2524) <= (layer3_outputs(1926)) xor (layer3_outputs(1122));
    layer4_outputs(2525) <= not(layer3_outputs(900));
    layer4_outputs(2526) <= layer3_outputs(414);
    layer4_outputs(2527) <= not((layer3_outputs(335)) and (layer3_outputs(238)));
    layer4_outputs(2528) <= layer3_outputs(1446);
    layer4_outputs(2529) <= not(layer3_outputs(1053)) or (layer3_outputs(12));
    layer4_outputs(2530) <= not((layer3_outputs(588)) and (layer3_outputs(2092)));
    layer4_outputs(2531) <= layer3_outputs(429);
    layer4_outputs(2532) <= not((layer3_outputs(130)) or (layer3_outputs(1338)));
    layer4_outputs(2533) <= not(layer3_outputs(1338));
    layer4_outputs(2534) <= (layer3_outputs(829)) and not (layer3_outputs(581));
    layer4_outputs(2535) <= not(layer3_outputs(2541));
    layer4_outputs(2536) <= layer3_outputs(2153);
    layer4_outputs(2537) <= not(layer3_outputs(509)) or (layer3_outputs(250));
    layer4_outputs(2538) <= layer3_outputs(1609);
    layer4_outputs(2539) <= not(layer3_outputs(731));
    layer4_outputs(2540) <= (layer3_outputs(2410)) and not (layer3_outputs(2099));
    layer4_outputs(2541) <= not(layer3_outputs(966));
    layer4_outputs(2542) <= '1';
    layer4_outputs(2543) <= not(layer3_outputs(1403));
    layer4_outputs(2544) <= (layer3_outputs(1055)) or (layer3_outputs(151));
    layer4_outputs(2545) <= (layer3_outputs(112)) and not (layer3_outputs(1554));
    layer4_outputs(2546) <= (layer3_outputs(1486)) xor (layer3_outputs(247));
    layer4_outputs(2547) <= not((layer3_outputs(1694)) or (layer3_outputs(43)));
    layer4_outputs(2548) <= (layer3_outputs(2141)) and not (layer3_outputs(233));
    layer4_outputs(2549) <= layer3_outputs(1821);
    layer4_outputs(2550) <= not(layer3_outputs(514));
    layer4_outputs(2551) <= (layer3_outputs(284)) and (layer3_outputs(1913));
    layer4_outputs(2552) <= (layer3_outputs(27)) or (layer3_outputs(315));
    layer4_outputs(2553) <= not(layer3_outputs(234));
    layer4_outputs(2554) <= layer3_outputs(1885);
    layer4_outputs(2555) <= not(layer3_outputs(2128)) or (layer3_outputs(1291));
    layer4_outputs(2556) <= not((layer3_outputs(1008)) and (layer3_outputs(367)));
    layer4_outputs(2557) <= (layer3_outputs(2235)) and (layer3_outputs(184));
    layer4_outputs(2558) <= not(layer3_outputs(1023));
    layer4_outputs(2559) <= (layer3_outputs(486)) and not (layer3_outputs(2015));
    outputs(0) <= not(layer4_outputs(1547));
    outputs(1) <= (layer4_outputs(2293)) and (layer4_outputs(1418));
    outputs(2) <= layer4_outputs(635);
    outputs(3) <= (layer4_outputs(54)) and not (layer4_outputs(1507));
    outputs(4) <= layer4_outputs(1942);
    outputs(5) <= not((layer4_outputs(1219)) xor (layer4_outputs(326)));
    outputs(6) <= (layer4_outputs(1903)) and not (layer4_outputs(247));
    outputs(7) <= not(layer4_outputs(1216));
    outputs(8) <= (layer4_outputs(1059)) and not (layer4_outputs(1770));
    outputs(9) <= (layer4_outputs(1680)) and not (layer4_outputs(2099));
    outputs(10) <= not(layer4_outputs(2058));
    outputs(11) <= layer4_outputs(694);
    outputs(12) <= layer4_outputs(1040);
    outputs(13) <= layer4_outputs(1229);
    outputs(14) <= not((layer4_outputs(981)) xor (layer4_outputs(1016)));
    outputs(15) <= layer4_outputs(2232);
    outputs(16) <= layer4_outputs(1892);
    outputs(17) <= (layer4_outputs(1246)) and not (layer4_outputs(252));
    outputs(18) <= not(layer4_outputs(1757));
    outputs(19) <= (layer4_outputs(488)) and not (layer4_outputs(266));
    outputs(20) <= (layer4_outputs(449)) and (layer4_outputs(761));
    outputs(21) <= (layer4_outputs(1017)) and (layer4_outputs(265));
    outputs(22) <= not(layer4_outputs(1141));
    outputs(23) <= not(layer4_outputs(1298));
    outputs(24) <= (layer4_outputs(894)) and (layer4_outputs(2191));
    outputs(25) <= (layer4_outputs(2124)) and not (layer4_outputs(487));
    outputs(26) <= not((layer4_outputs(1136)) and (layer4_outputs(673)));
    outputs(27) <= layer4_outputs(1463);
    outputs(28) <= not(layer4_outputs(2504));
    outputs(29) <= layer4_outputs(176);
    outputs(30) <= not(layer4_outputs(1790));
    outputs(31) <= not(layer4_outputs(616));
    outputs(32) <= not(layer4_outputs(590));
    outputs(33) <= (layer4_outputs(1347)) and not (layer4_outputs(2024));
    outputs(34) <= (layer4_outputs(797)) xor (layer4_outputs(730));
    outputs(35) <= layer4_outputs(1885);
    outputs(36) <= not((layer4_outputs(686)) xor (layer4_outputs(2284)));
    outputs(37) <= not(layer4_outputs(1181));
    outputs(38) <= layer4_outputs(289);
    outputs(39) <= (layer4_outputs(2020)) and not (layer4_outputs(1916));
    outputs(40) <= (layer4_outputs(488)) and not (layer4_outputs(936));
    outputs(41) <= (layer4_outputs(2068)) and not (layer4_outputs(1618));
    outputs(42) <= not((layer4_outputs(2089)) xor (layer4_outputs(1100)));
    outputs(43) <= layer4_outputs(550);
    outputs(44) <= layer4_outputs(776);
    outputs(45) <= (layer4_outputs(1734)) and not (layer4_outputs(1379));
    outputs(46) <= layer4_outputs(2328);
    outputs(47) <= (layer4_outputs(2389)) and (layer4_outputs(137));
    outputs(48) <= layer4_outputs(1417);
    outputs(49) <= not(layer4_outputs(1567));
    outputs(50) <= not(layer4_outputs(530));
    outputs(51) <= not((layer4_outputs(1514)) xor (layer4_outputs(1787)));
    outputs(52) <= not((layer4_outputs(1798)) or (layer4_outputs(1088)));
    outputs(53) <= not(layer4_outputs(1177));
    outputs(54) <= not((layer4_outputs(1588)) xor (layer4_outputs(2248)));
    outputs(55) <= (layer4_outputs(1135)) and not (layer4_outputs(1144));
    outputs(56) <= layer4_outputs(2402);
    outputs(57) <= not(layer4_outputs(2527)) or (layer4_outputs(402));
    outputs(58) <= layer4_outputs(1608);
    outputs(59) <= (layer4_outputs(1079)) xor (layer4_outputs(1603));
    outputs(60) <= layer4_outputs(2296);
    outputs(61) <= (layer4_outputs(876)) and not (layer4_outputs(1200));
    outputs(62) <= not((layer4_outputs(1553)) and (layer4_outputs(2313)));
    outputs(63) <= not((layer4_outputs(1854)) or (layer4_outputs(1962)));
    outputs(64) <= (layer4_outputs(75)) or (layer4_outputs(2440));
    outputs(65) <= not((layer4_outputs(1287)) xor (layer4_outputs(2527)));
    outputs(66) <= layer4_outputs(1125);
    outputs(67) <= not(layer4_outputs(713));
    outputs(68) <= not((layer4_outputs(287)) or (layer4_outputs(1943)));
    outputs(69) <= layer4_outputs(1036);
    outputs(70) <= layer4_outputs(1869);
    outputs(71) <= (layer4_outputs(321)) and not (layer4_outputs(316));
    outputs(72) <= not(layer4_outputs(924));
    outputs(73) <= layer4_outputs(2319);
    outputs(74) <= layer4_outputs(2295);
    outputs(75) <= (layer4_outputs(214)) and not (layer4_outputs(616));
    outputs(76) <= not(layer4_outputs(46));
    outputs(77) <= not((layer4_outputs(464)) xor (layer4_outputs(1231)));
    outputs(78) <= not(layer4_outputs(1870));
    outputs(79) <= (layer4_outputs(675)) and not (layer4_outputs(837));
    outputs(80) <= not(layer4_outputs(2465));
    outputs(81) <= not(layer4_outputs(847));
    outputs(82) <= (layer4_outputs(461)) and not (layer4_outputs(2474));
    outputs(83) <= (layer4_outputs(199)) xor (layer4_outputs(1239));
    outputs(84) <= (layer4_outputs(1469)) xor (layer4_outputs(729));
    outputs(85) <= (layer4_outputs(439)) xor (layer4_outputs(2438));
    outputs(86) <= layer4_outputs(275);
    outputs(87) <= (layer4_outputs(2212)) and (layer4_outputs(1998));
    outputs(88) <= (layer4_outputs(2551)) or (layer4_outputs(2080));
    outputs(89) <= layer4_outputs(2029);
    outputs(90) <= layer4_outputs(2352);
    outputs(91) <= not((layer4_outputs(937)) or (layer4_outputs(1092)));
    outputs(92) <= layer4_outputs(162);
    outputs(93) <= not(layer4_outputs(345));
    outputs(94) <= (layer4_outputs(425)) and not (layer4_outputs(535));
    outputs(95) <= not(layer4_outputs(981));
    outputs(96) <= (layer4_outputs(1137)) or (layer4_outputs(460));
    outputs(97) <= (layer4_outputs(242)) and not (layer4_outputs(1527));
    outputs(98) <= not(layer4_outputs(2386));
    outputs(99) <= not(layer4_outputs(1914));
    outputs(100) <= not(layer4_outputs(2073));
    outputs(101) <= layer4_outputs(512);
    outputs(102) <= layer4_outputs(1482);
    outputs(103) <= layer4_outputs(2530);
    outputs(104) <= layer4_outputs(1858);
    outputs(105) <= not((layer4_outputs(1975)) xor (layer4_outputs(1093)));
    outputs(106) <= layer4_outputs(2523);
    outputs(107) <= (layer4_outputs(1443)) and (layer4_outputs(204));
    outputs(108) <= not((layer4_outputs(1089)) or (layer4_outputs(1985)));
    outputs(109) <= not(layer4_outputs(604));
    outputs(110) <= not(layer4_outputs(2177));
    outputs(111) <= not((layer4_outputs(801)) or (layer4_outputs(2432)));
    outputs(112) <= not(layer4_outputs(1080));
    outputs(113) <= not(layer4_outputs(187));
    outputs(114) <= (layer4_outputs(1695)) xor (layer4_outputs(155));
    outputs(115) <= layer4_outputs(1491);
    outputs(116) <= not(layer4_outputs(921));
    outputs(117) <= layer4_outputs(277);
    outputs(118) <= layer4_outputs(547);
    outputs(119) <= not(layer4_outputs(2181));
    outputs(120) <= not(layer4_outputs(2254));
    outputs(121) <= (layer4_outputs(2348)) or (layer4_outputs(1704));
    outputs(122) <= layer4_outputs(1126);
    outputs(123) <= layer4_outputs(414);
    outputs(124) <= (layer4_outputs(1884)) xor (layer4_outputs(513));
    outputs(125) <= not(layer4_outputs(2058));
    outputs(126) <= (layer4_outputs(2268)) and not (layer4_outputs(1164));
    outputs(127) <= (layer4_outputs(406)) and not (layer4_outputs(1465));
    outputs(128) <= layer4_outputs(1888);
    outputs(129) <= (layer4_outputs(148)) and not (layer4_outputs(133));
    outputs(130) <= layer4_outputs(1125);
    outputs(131) <= not(layer4_outputs(2522));
    outputs(132) <= not((layer4_outputs(2445)) xor (layer4_outputs(2299)));
    outputs(133) <= (layer4_outputs(280)) xor (layer4_outputs(991));
    outputs(134) <= (layer4_outputs(539)) and (layer4_outputs(97));
    outputs(135) <= layer4_outputs(327);
    outputs(136) <= (layer4_outputs(307)) and not (layer4_outputs(329));
    outputs(137) <= not(layer4_outputs(2195));
    outputs(138) <= layer4_outputs(310);
    outputs(139) <= not((layer4_outputs(1796)) or (layer4_outputs(798)));
    outputs(140) <= not(layer4_outputs(354));
    outputs(141) <= not(layer4_outputs(2399));
    outputs(142) <= not(layer4_outputs(147));
    outputs(143) <= not(layer4_outputs(2432));
    outputs(144) <= not(layer4_outputs(1838));
    outputs(145) <= (layer4_outputs(1284)) and not (layer4_outputs(306));
    outputs(146) <= not((layer4_outputs(1119)) and (layer4_outputs(646)));
    outputs(147) <= not(layer4_outputs(128));
    outputs(148) <= (layer4_outputs(68)) and not (layer4_outputs(884));
    outputs(149) <= not(layer4_outputs(856));
    outputs(150) <= (layer4_outputs(422)) and not (layer4_outputs(2513));
    outputs(151) <= not((layer4_outputs(1750)) or (layer4_outputs(333)));
    outputs(152) <= (layer4_outputs(1737)) and not (layer4_outputs(35));
    outputs(153) <= not(layer4_outputs(839));
    outputs(154) <= not(layer4_outputs(2112));
    outputs(155) <= layer4_outputs(1898);
    outputs(156) <= not(layer4_outputs(365));
    outputs(157) <= not(layer4_outputs(2004));
    outputs(158) <= layer4_outputs(868);
    outputs(159) <= not(layer4_outputs(1565)) or (layer4_outputs(869));
    outputs(160) <= not(layer4_outputs(2335));
    outputs(161) <= (layer4_outputs(749)) and not (layer4_outputs(1131));
    outputs(162) <= layer4_outputs(957);
    outputs(163) <= not(layer4_outputs(1920));
    outputs(164) <= not(layer4_outputs(202)) or (layer4_outputs(2517));
    outputs(165) <= layer4_outputs(2417);
    outputs(166) <= (layer4_outputs(815)) xor (layer4_outputs(1884));
    outputs(167) <= layer4_outputs(1407);
    outputs(168) <= not(layer4_outputs(1144));
    outputs(169) <= (layer4_outputs(859)) and (layer4_outputs(546));
    outputs(170) <= layer4_outputs(726);
    outputs(171) <= not((layer4_outputs(847)) or (layer4_outputs(1771)));
    outputs(172) <= not(layer4_outputs(2148));
    outputs(173) <= (layer4_outputs(1536)) and not (layer4_outputs(1578));
    outputs(174) <= not(layer4_outputs(961));
    outputs(175) <= not(layer4_outputs(3));
    outputs(176) <= not((layer4_outputs(732)) or (layer4_outputs(974)));
    outputs(177) <= layer4_outputs(275);
    outputs(178) <= layer4_outputs(63);
    outputs(179) <= (layer4_outputs(976)) xor (layer4_outputs(1529));
    outputs(180) <= not((layer4_outputs(1177)) or (layer4_outputs(1183)));
    outputs(181) <= layer4_outputs(137);
    outputs(182) <= (layer4_outputs(74)) and not (layer4_outputs(478));
    outputs(183) <= layer4_outputs(1675);
    outputs(184) <= not(layer4_outputs(95));
    outputs(185) <= not((layer4_outputs(781)) and (layer4_outputs(2230)));
    outputs(186) <= layer4_outputs(1521);
    outputs(187) <= layer4_outputs(864);
    outputs(188) <= layer4_outputs(235);
    outputs(189) <= not(layer4_outputs(1924));
    outputs(190) <= not(layer4_outputs(2373));
    outputs(191) <= not((layer4_outputs(999)) and (layer4_outputs(1683)));
    outputs(192) <= (layer4_outputs(2357)) and not (layer4_outputs(194));
    outputs(193) <= not(layer4_outputs(2336));
    outputs(194) <= (layer4_outputs(633)) xor (layer4_outputs(1653));
    outputs(195) <= not(layer4_outputs(1875)) or (layer4_outputs(1205));
    outputs(196) <= layer4_outputs(523);
    outputs(197) <= not(layer4_outputs(938)) or (layer4_outputs(1621));
    outputs(198) <= (layer4_outputs(693)) and (layer4_outputs(2184));
    outputs(199) <= layer4_outputs(47);
    outputs(200) <= (layer4_outputs(2324)) and not (layer4_outputs(692));
    outputs(201) <= layer4_outputs(892);
    outputs(202) <= layer4_outputs(1360);
    outputs(203) <= layer4_outputs(256);
    outputs(204) <= not((layer4_outputs(269)) xor (layer4_outputs(907)));
    outputs(205) <= not(layer4_outputs(316)) or (layer4_outputs(113));
    outputs(206) <= layer4_outputs(678);
    outputs(207) <= not(layer4_outputs(685));
    outputs(208) <= (layer4_outputs(977)) and not (layer4_outputs(5));
    outputs(209) <= layer4_outputs(348);
    outputs(210) <= layer4_outputs(249);
    outputs(211) <= layer4_outputs(1408);
    outputs(212) <= layer4_outputs(143);
    outputs(213) <= not(layer4_outputs(709));
    outputs(214) <= layer4_outputs(554);
    outputs(215) <= not((layer4_outputs(1946)) or (layer4_outputs(1736)));
    outputs(216) <= (layer4_outputs(2213)) xor (layer4_outputs(594));
    outputs(217) <= (layer4_outputs(601)) and not (layer4_outputs(2153));
    outputs(218) <= not(layer4_outputs(1074));
    outputs(219) <= (layer4_outputs(1868)) and (layer4_outputs(1998));
    outputs(220) <= (layer4_outputs(2202)) and (layer4_outputs(461));
    outputs(221) <= layer4_outputs(1973);
    outputs(222) <= not(layer4_outputs(2097));
    outputs(223) <= not((layer4_outputs(283)) or (layer4_outputs(432)));
    outputs(224) <= (layer4_outputs(146)) and (layer4_outputs(1138));
    outputs(225) <= not((layer4_outputs(579)) or (layer4_outputs(925)));
    outputs(226) <= (layer4_outputs(250)) and not (layer4_outputs(2549));
    outputs(227) <= not(layer4_outputs(1321));
    outputs(228) <= not((layer4_outputs(1668)) xor (layer4_outputs(169)));
    outputs(229) <= not(layer4_outputs(170));
    outputs(230) <= not(layer4_outputs(366));
    outputs(231) <= layer4_outputs(1427);
    outputs(232) <= layer4_outputs(1662);
    outputs(233) <= layer4_outputs(2045);
    outputs(234) <= (layer4_outputs(1922)) and not (layer4_outputs(1324));
    outputs(235) <= layer4_outputs(1469);
    outputs(236) <= (layer4_outputs(1878)) and not (layer4_outputs(608));
    outputs(237) <= layer4_outputs(766);
    outputs(238) <= not((layer4_outputs(115)) xor (layer4_outputs(1552)));
    outputs(239) <= not(layer4_outputs(1614));
    outputs(240) <= layer4_outputs(2114);
    outputs(241) <= layer4_outputs(397);
    outputs(242) <= (layer4_outputs(2330)) and not (layer4_outputs(1134));
    outputs(243) <= not(layer4_outputs(649));
    outputs(244) <= layer4_outputs(1983);
    outputs(245) <= not(layer4_outputs(1447));
    outputs(246) <= (layer4_outputs(2131)) and not (layer4_outputs(1770));
    outputs(247) <= not(layer4_outputs(2430));
    outputs(248) <= not(layer4_outputs(1271));
    outputs(249) <= not(layer4_outputs(929));
    outputs(250) <= not((layer4_outputs(671)) xor (layer4_outputs(82)));
    outputs(251) <= layer4_outputs(486);
    outputs(252) <= layer4_outputs(1273);
    outputs(253) <= (layer4_outputs(2245)) xor (layer4_outputs(25));
    outputs(254) <= layer4_outputs(1969);
    outputs(255) <= layer4_outputs(600);
    outputs(256) <= not(layer4_outputs(1782));
    outputs(257) <= not(layer4_outputs(1402));
    outputs(258) <= layer4_outputs(1423);
    outputs(259) <= (layer4_outputs(1141)) and not (layer4_outputs(1460));
    outputs(260) <= not(layer4_outputs(949));
    outputs(261) <= (layer4_outputs(1182)) and not (layer4_outputs(2053));
    outputs(262) <= layer4_outputs(1830);
    outputs(263) <= not((layer4_outputs(348)) or (layer4_outputs(1896)));
    outputs(264) <= (layer4_outputs(814)) and (layer4_outputs(318));
    outputs(265) <= layer4_outputs(1049);
    outputs(266) <= not(layer4_outputs(369)) or (layer4_outputs(2167));
    outputs(267) <= not(layer4_outputs(160));
    outputs(268) <= layer4_outputs(1210);
    outputs(269) <= (layer4_outputs(129)) and not (layer4_outputs(2192));
    outputs(270) <= not((layer4_outputs(1376)) or (layer4_outputs(1227)));
    outputs(271) <= (layer4_outputs(536)) and (layer4_outputs(2337));
    outputs(272) <= (layer4_outputs(2361)) and not (layer4_outputs(2082));
    outputs(273) <= layer4_outputs(1040);
    outputs(274) <= not((layer4_outputs(1398)) or (layer4_outputs(909)));
    outputs(275) <= layer4_outputs(1171);
    outputs(276) <= (layer4_outputs(476)) and not (layer4_outputs(868));
    outputs(277) <= not(layer4_outputs(2170));
    outputs(278) <= not(layer4_outputs(1006));
    outputs(279) <= layer4_outputs(392);
    outputs(280) <= (layer4_outputs(569)) and not (layer4_outputs(791));
    outputs(281) <= (layer4_outputs(2199)) and not (layer4_outputs(1025));
    outputs(282) <= layer4_outputs(151);
    outputs(283) <= layer4_outputs(1315);
    outputs(284) <= layer4_outputs(1555);
    outputs(285) <= not(layer4_outputs(1127));
    outputs(286) <= not(layer4_outputs(374));
    outputs(287) <= (layer4_outputs(95)) and (layer4_outputs(2313));
    outputs(288) <= layer4_outputs(2287);
    outputs(289) <= (layer4_outputs(438)) xor (layer4_outputs(2511));
    outputs(290) <= layer4_outputs(365);
    outputs(291) <= not((layer4_outputs(94)) xor (layer4_outputs(402)));
    outputs(292) <= (layer4_outputs(2300)) and (layer4_outputs(1289));
    outputs(293) <= layer4_outputs(8);
    outputs(294) <= (layer4_outputs(962)) and not (layer4_outputs(1156));
    outputs(295) <= (layer4_outputs(1589)) and not (layer4_outputs(916));
    outputs(296) <= layer4_outputs(1686);
    outputs(297) <= layer4_outputs(2269);
    outputs(298) <= layer4_outputs(2012);
    outputs(299) <= (layer4_outputs(2536)) and (layer4_outputs(238));
    outputs(300) <= layer4_outputs(1661);
    outputs(301) <= layer4_outputs(2260);
    outputs(302) <= (layer4_outputs(1058)) and not (layer4_outputs(762));
    outputs(303) <= not(layer4_outputs(415));
    outputs(304) <= layer4_outputs(1142);
    outputs(305) <= layer4_outputs(1532);
    outputs(306) <= not(layer4_outputs(1927));
    outputs(307) <= (layer4_outputs(2157)) and (layer4_outputs(1343));
    outputs(308) <= layer4_outputs(1056);
    outputs(309) <= (layer4_outputs(1877)) and not (layer4_outputs(253));
    outputs(310) <= layer4_outputs(432);
    outputs(311) <= not((layer4_outputs(530)) xor (layer4_outputs(1101)));
    outputs(312) <= not((layer4_outputs(1632)) or (layer4_outputs(1889)));
    outputs(313) <= not((layer4_outputs(2044)) or (layer4_outputs(1973)));
    outputs(314) <= not(layer4_outputs(1319));
    outputs(315) <= (layer4_outputs(1450)) and (layer4_outputs(1044));
    outputs(316) <= not((layer4_outputs(1458)) or (layer4_outputs(2304)));
    outputs(317) <= not(layer4_outputs(493));
    outputs(318) <= layer4_outputs(1147);
    outputs(319) <= (layer4_outputs(2447)) and not (layer4_outputs(1855));
    outputs(320) <= layer4_outputs(501);
    outputs(321) <= not(layer4_outputs(1778));
    outputs(322) <= (layer4_outputs(2476)) and not (layer4_outputs(2387));
    outputs(323) <= not(layer4_outputs(2299));
    outputs(324) <= (layer4_outputs(1157)) and not (layer4_outputs(1463));
    outputs(325) <= layer4_outputs(2207);
    outputs(326) <= (layer4_outputs(1940)) and not (layer4_outputs(774));
    outputs(327) <= (layer4_outputs(1067)) and (layer4_outputs(314));
    outputs(328) <= not(layer4_outputs(1989));
    outputs(329) <= (layer4_outputs(2200)) and not (layer4_outputs(302));
    outputs(330) <= layer4_outputs(2282);
    outputs(331) <= not((layer4_outputs(656)) or (layer4_outputs(697)));
    outputs(332) <= layer4_outputs(1788);
    outputs(333) <= not((layer4_outputs(1220)) or (layer4_outputs(140)));
    outputs(334) <= layer4_outputs(427);
    outputs(335) <= layer4_outputs(429);
    outputs(336) <= layer4_outputs(1383);
    outputs(337) <= layer4_outputs(957);
    outputs(338) <= not(layer4_outputs(1370));
    outputs(339) <= not((layer4_outputs(1030)) or (layer4_outputs(1716)));
    outputs(340) <= (layer4_outputs(1601)) and not (layer4_outputs(1952));
    outputs(341) <= layer4_outputs(2148);
    outputs(342) <= not((layer4_outputs(160)) or (layer4_outputs(1460)));
    outputs(343) <= (layer4_outputs(2223)) or (layer4_outputs(138));
    outputs(344) <= not(layer4_outputs(2211));
    outputs(345) <= layer4_outputs(1736);
    outputs(346) <= not(layer4_outputs(806));
    outputs(347) <= (layer4_outputs(116)) and (layer4_outputs(1324));
    outputs(348) <= not(layer4_outputs(702));
    outputs(349) <= (layer4_outputs(757)) and not (layer4_outputs(1477));
    outputs(350) <= (layer4_outputs(1184)) and (layer4_outputs(1692));
    outputs(351) <= layer4_outputs(745);
    outputs(352) <= (layer4_outputs(238)) and not (layer4_outputs(1286));
    outputs(353) <= layer4_outputs(1165);
    outputs(354) <= not(layer4_outputs(1804));
    outputs(355) <= (layer4_outputs(1781)) and (layer4_outputs(99));
    outputs(356) <= not(layer4_outputs(1580));
    outputs(357) <= not(layer4_outputs(1592));
    outputs(358) <= (layer4_outputs(231)) and not (layer4_outputs(2103));
    outputs(359) <= (layer4_outputs(2522)) and (layer4_outputs(2367));
    outputs(360) <= (layer4_outputs(596)) and not (layer4_outputs(2255));
    outputs(361) <= not((layer4_outputs(1382)) or (layer4_outputs(2044)));
    outputs(362) <= not(layer4_outputs(1501));
    outputs(363) <= layer4_outputs(1832);
    outputs(364) <= not((layer4_outputs(1118)) or (layer4_outputs(1432)));
    outputs(365) <= not((layer4_outputs(2107)) or (layer4_outputs(2494)));
    outputs(366) <= layer4_outputs(1891);
    outputs(367) <= (layer4_outputs(300)) or (layer4_outputs(1656));
    outputs(368) <= (layer4_outputs(1313)) and not (layer4_outputs(2322));
    outputs(369) <= (layer4_outputs(1726)) and (layer4_outputs(2090));
    outputs(370) <= (layer4_outputs(2433)) and not (layer4_outputs(1733));
    outputs(371) <= layer4_outputs(85);
    outputs(372) <= (layer4_outputs(33)) and not (layer4_outputs(2467));
    outputs(373) <= not(layer4_outputs(1150)) or (layer4_outputs(1777));
    outputs(374) <= layer4_outputs(811);
    outputs(375) <= layer4_outputs(2275);
    outputs(376) <= (layer4_outputs(2013)) and not (layer4_outputs(1413));
    outputs(377) <= not(layer4_outputs(249));
    outputs(378) <= layer4_outputs(2209);
    outputs(379) <= not(layer4_outputs(2131));
    outputs(380) <= layer4_outputs(548);
    outputs(381) <= (layer4_outputs(1836)) xor (layer4_outputs(283));
    outputs(382) <= layer4_outputs(2410);
    outputs(383) <= (layer4_outputs(2521)) and not (layer4_outputs(404));
    outputs(384) <= layer4_outputs(1103);
    outputs(385) <= not(layer4_outputs(1386));
    outputs(386) <= not(layer4_outputs(1530));
    outputs(387) <= not(layer4_outputs(1678)) or (layer4_outputs(1684));
    outputs(388) <= not((layer4_outputs(2137)) or (layer4_outputs(968)));
    outputs(389) <= not(layer4_outputs(632));
    outputs(390) <= (layer4_outputs(1593)) and not (layer4_outputs(1449));
    outputs(391) <= not(layer4_outputs(1799));
    outputs(392) <= (layer4_outputs(468)) and not (layer4_outputs(1848));
    outputs(393) <= (layer4_outputs(798)) or (layer4_outputs(579));
    outputs(394) <= not(layer4_outputs(838)) or (layer4_outputs(1833));
    outputs(395) <= (layer4_outputs(1816)) and not (layer4_outputs(2428));
    outputs(396) <= layer4_outputs(2167);
    outputs(397) <= layer4_outputs(177);
    outputs(398) <= (layer4_outputs(1381)) and not (layer4_outputs(2205));
    outputs(399) <= not(layer4_outputs(2530));
    outputs(400) <= layer4_outputs(2060);
    outputs(401) <= (layer4_outputs(637)) and (layer4_outputs(873));
    outputs(402) <= not((layer4_outputs(1883)) xor (layer4_outputs(1941)));
    outputs(403) <= not((layer4_outputs(1730)) or (layer4_outputs(932)));
    outputs(404) <= not(layer4_outputs(1737));
    outputs(405) <= layer4_outputs(232);
    outputs(406) <= layer4_outputs(2346);
    outputs(407) <= not(layer4_outputs(1608));
    outputs(408) <= (layer4_outputs(1017)) and (layer4_outputs(1670));
    outputs(409) <= not(layer4_outputs(582));
    outputs(410) <= not((layer4_outputs(341)) or (layer4_outputs(1989)));
    outputs(411) <= layer4_outputs(1457);
    outputs(412) <= not((layer4_outputs(2084)) or (layer4_outputs(1913)));
    outputs(413) <= not(layer4_outputs(2168));
    outputs(414) <= (layer4_outputs(1866)) and not (layer4_outputs(1952));
    outputs(415) <= (layer4_outputs(508)) and not (layer4_outputs(384));
    outputs(416) <= layer4_outputs(1271);
    outputs(417) <= not((layer4_outputs(1320)) or (layer4_outputs(367)));
    outputs(418) <= layer4_outputs(429);
    outputs(419) <= (layer4_outputs(1967)) and (layer4_outputs(1844));
    outputs(420) <= layer4_outputs(1);
    outputs(421) <= not(layer4_outputs(184));
    outputs(422) <= (layer4_outputs(1379)) and not (layer4_outputs(1192));
    outputs(423) <= not((layer4_outputs(1741)) or (layer4_outputs(872)));
    outputs(424) <= (layer4_outputs(2129)) and not (layer4_outputs(339));
    outputs(425) <= layer4_outputs(1604);
    outputs(426) <= not(layer4_outputs(2395));
    outputs(427) <= (layer4_outputs(2013)) and not (layer4_outputs(2098));
    outputs(428) <= not(layer4_outputs(136));
    outputs(429) <= layer4_outputs(1155);
    outputs(430) <= (layer4_outputs(2406)) and not (layer4_outputs(2135));
    outputs(431) <= layer4_outputs(1043);
    outputs(432) <= not(layer4_outputs(1322)) or (layer4_outputs(574));
    outputs(433) <= not(layer4_outputs(689));
    outputs(434) <= not((layer4_outputs(172)) or (layer4_outputs(1015)));
    outputs(435) <= not(layer4_outputs(84));
    outputs(436) <= layer4_outputs(1626);
    outputs(437) <= (layer4_outputs(152)) and not (layer4_outputs(1819));
    outputs(438) <= layer4_outputs(1003);
    outputs(439) <= not((layer4_outputs(2284)) xor (layer4_outputs(17)));
    outputs(440) <= (layer4_outputs(2499)) and not (layer4_outputs(2028));
    outputs(441) <= not(layer4_outputs(797)) or (layer4_outputs(2149));
    outputs(442) <= not((layer4_outputs(1939)) xor (layer4_outputs(1262)));
    outputs(443) <= not((layer4_outputs(331)) or (layer4_outputs(951)));
    outputs(444) <= layer4_outputs(141);
    outputs(445) <= not(layer4_outputs(1496));
    outputs(446) <= layer4_outputs(328);
    outputs(447) <= not((layer4_outputs(1605)) or (layer4_outputs(2264)));
    outputs(448) <= (layer4_outputs(2238)) and not (layer4_outputs(2239));
    outputs(449) <= layer4_outputs(1946);
    outputs(450) <= (layer4_outputs(2193)) and not (layer4_outputs(1325));
    outputs(451) <= not(layer4_outputs(2208)) or (layer4_outputs(2370));
    outputs(452) <= not((layer4_outputs(307)) or (layer4_outputs(774)));
    outputs(453) <= (layer4_outputs(477)) and not (layer4_outputs(2229));
    outputs(454) <= (layer4_outputs(1721)) and not (layer4_outputs(111));
    outputs(455) <= (layer4_outputs(672)) and not (layer4_outputs(716));
    outputs(456) <= (layer4_outputs(1842)) and (layer4_outputs(1252));
    outputs(457) <= (layer4_outputs(1686)) and not (layer4_outputs(992));
    outputs(458) <= not(layer4_outputs(471));
    outputs(459) <= not(layer4_outputs(370));
    outputs(460) <= layer4_outputs(400);
    outputs(461) <= (layer4_outputs(803)) and not (layer4_outputs(2452));
    outputs(462) <= not(layer4_outputs(930));
    outputs(463) <= not(layer4_outputs(1717));
    outputs(464) <= (layer4_outputs(2516)) and not (layer4_outputs(287));
    outputs(465) <= not((layer4_outputs(2005)) or (layer4_outputs(1336)));
    outputs(466) <= (layer4_outputs(925)) and not (layer4_outputs(2352));
    outputs(467) <= layer4_outputs(121);
    outputs(468) <= not((layer4_outputs(444)) xor (layer4_outputs(985)));
    outputs(469) <= layer4_outputs(1093);
    outputs(470) <= layer4_outputs(290);
    outputs(471) <= not((layer4_outputs(1226)) xor (layer4_outputs(1821)));
    outputs(472) <= (layer4_outputs(1359)) and (layer4_outputs(1629));
    outputs(473) <= (layer4_outputs(1676)) and (layer4_outputs(1490));
    outputs(474) <= not((layer4_outputs(1174)) or (layer4_outputs(593)));
    outputs(475) <= (layer4_outputs(667)) and (layer4_outputs(1453));
    outputs(476) <= layer4_outputs(222);
    outputs(477) <= layer4_outputs(719);
    outputs(478) <= not(layer4_outputs(1208));
    outputs(479) <= not(layer4_outputs(2192));
    outputs(480) <= (layer4_outputs(225)) and not (layer4_outputs(1314));
    outputs(481) <= not(layer4_outputs(2233));
    outputs(482) <= not((layer4_outputs(2424)) xor (layer4_outputs(820)));
    outputs(483) <= layer4_outputs(123);
    outputs(484) <= not((layer4_outputs(479)) xor (layer4_outputs(816)));
    outputs(485) <= (layer4_outputs(1003)) and not (layer4_outputs(356));
    outputs(486) <= not((layer4_outputs(1633)) or (layer4_outputs(991)));
    outputs(487) <= (layer4_outputs(1551)) and (layer4_outputs(1250));
    outputs(488) <= (layer4_outputs(528)) xor (layer4_outputs(1806));
    outputs(489) <= not(layer4_outputs(697));
    outputs(490) <= (layer4_outputs(1679)) and not (layer4_outputs(642));
    outputs(491) <= (layer4_outputs(1033)) and (layer4_outputs(1935));
    outputs(492) <= not(layer4_outputs(1663));
    outputs(493) <= layer4_outputs(1504);
    outputs(494) <= not(layer4_outputs(2378)) or (layer4_outputs(897));
    outputs(495) <= not(layer4_outputs(804));
    outputs(496) <= not((layer4_outputs(224)) or (layer4_outputs(362)));
    outputs(497) <= (layer4_outputs(1250)) and (layer4_outputs(2035));
    outputs(498) <= not((layer4_outputs(1008)) or (layer4_outputs(0)));
    outputs(499) <= layer4_outputs(1153);
    outputs(500) <= not(layer4_outputs(1069));
    outputs(501) <= layer4_outputs(586);
    outputs(502) <= layer4_outputs(1393);
    outputs(503) <= (layer4_outputs(169)) xor (layer4_outputs(2196));
    outputs(504) <= layer4_outputs(2054);
    outputs(505) <= layer4_outputs(121);
    outputs(506) <= not(layer4_outputs(258));
    outputs(507) <= layer4_outputs(1049);
    outputs(508) <= not((layer4_outputs(517)) xor (layer4_outputs(1606)));
    outputs(509) <= not((layer4_outputs(1217)) or (layer4_outputs(465)));
    outputs(510) <= layer4_outputs(70);
    outputs(511) <= (layer4_outputs(2496)) and (layer4_outputs(767));
    outputs(512) <= not(layer4_outputs(2503)) or (layer4_outputs(2540));
    outputs(513) <= not(layer4_outputs(2273));
    outputs(514) <= layer4_outputs(341);
    outputs(515) <= layer4_outputs(1650);
    outputs(516) <= not(layer4_outputs(419));
    outputs(517) <= not(layer4_outputs(828));
    outputs(518) <= (layer4_outputs(1297)) and (layer4_outputs(492));
    outputs(519) <= not((layer4_outputs(524)) xor (layer4_outputs(560)));
    outputs(520) <= layer4_outputs(497);
    outputs(521) <= not(layer4_outputs(813));
    outputs(522) <= not((layer4_outputs(1955)) xor (layer4_outputs(2201)));
    outputs(523) <= (layer4_outputs(738)) and not (layer4_outputs(1850));
    outputs(524) <= not(layer4_outputs(1982));
    outputs(525) <= (layer4_outputs(942)) and (layer4_outputs(990));
    outputs(526) <= not((layer4_outputs(1748)) xor (layer4_outputs(2475)));
    outputs(527) <= (layer4_outputs(1588)) xor (layer4_outputs(1380));
    outputs(528) <= not(layer4_outputs(949));
    outputs(529) <= not(layer4_outputs(2353));
    outputs(530) <= (layer4_outputs(851)) and (layer4_outputs(1300));
    outputs(531) <= not(layer4_outputs(2118));
    outputs(532) <= not(layer4_outputs(659));
    outputs(533) <= layer4_outputs(2460);
    outputs(534) <= layer4_outputs(1717);
    outputs(535) <= (layer4_outputs(2463)) xor (layer4_outputs(37));
    outputs(536) <= layer4_outputs(1936);
    outputs(537) <= layer4_outputs(625);
    outputs(538) <= layer4_outputs(281);
    outputs(539) <= not((layer4_outputs(2091)) xor (layer4_outputs(1517)));
    outputs(540) <= layer4_outputs(1122);
    outputs(541) <= layer4_outputs(297);
    outputs(542) <= not(layer4_outputs(1791));
    outputs(543) <= not(layer4_outputs(1648)) or (layer4_outputs(534));
    outputs(544) <= (layer4_outputs(2184)) xor (layer4_outputs(294));
    outputs(545) <= layer4_outputs(1711);
    outputs(546) <= not(layer4_outputs(2448)) or (layer4_outputs(2466));
    outputs(547) <= not(layer4_outputs(711));
    outputs(548) <= not(layer4_outputs(1187));
    outputs(549) <= (layer4_outputs(1526)) xor (layer4_outputs(373));
    outputs(550) <= layer4_outputs(1749);
    outputs(551) <= not(layer4_outputs(527));
    outputs(552) <= not(layer4_outputs(2185));
    outputs(553) <= not(layer4_outputs(2366));
    outputs(554) <= not(layer4_outputs(1182)) or (layer4_outputs(1432));
    outputs(555) <= not((layer4_outputs(1626)) xor (layer4_outputs(2104)));
    outputs(556) <= not(layer4_outputs(1269));
    outputs(557) <= not(layer4_outputs(1544)) or (layer4_outputs(412));
    outputs(558) <= layer4_outputs(1984);
    outputs(559) <= not(layer4_outputs(1012));
    outputs(560) <= not(layer4_outputs(2249));
    outputs(561) <= not(layer4_outputs(2056));
    outputs(562) <= not(layer4_outputs(2170));
    outputs(563) <= not(layer4_outputs(2176));
    outputs(564) <= layer4_outputs(1684);
    outputs(565) <= not(layer4_outputs(2162)) or (layer4_outputs(1607));
    outputs(566) <= not(layer4_outputs(2393));
    outputs(567) <= layer4_outputs(1829);
    outputs(568) <= layer4_outputs(1461);
    outputs(569) <= not(layer4_outputs(2338));
    outputs(570) <= not(layer4_outputs(444));
    outputs(571) <= not((layer4_outputs(398)) and (layer4_outputs(1245)));
    outputs(572) <= not(layer4_outputs(741));
    outputs(573) <= not(layer4_outputs(2494));
    outputs(574) <= not(layer4_outputs(1569));
    outputs(575) <= not((layer4_outputs(331)) xor (layer4_outputs(570)));
    outputs(576) <= layer4_outputs(2286);
    outputs(577) <= not((layer4_outputs(470)) or (layer4_outputs(2056)));
    outputs(578) <= not((layer4_outputs(1424)) and (layer4_outputs(653)));
    outputs(579) <= layer4_outputs(1238);
    outputs(580) <= layer4_outputs(1710);
    outputs(581) <= (layer4_outputs(2500)) or (layer4_outputs(210));
    outputs(582) <= layer4_outputs(877);
    outputs(583) <= layer4_outputs(415);
    outputs(584) <= not(layer4_outputs(288));
    outputs(585) <= (layer4_outputs(938)) and (layer4_outputs(2068));
    outputs(586) <= (layer4_outputs(865)) or (layer4_outputs(93));
    outputs(587) <= not(layer4_outputs(143));
    outputs(588) <= not(layer4_outputs(184));
    outputs(589) <= layer4_outputs(841);
    outputs(590) <= layer4_outputs(271);
    outputs(591) <= not(layer4_outputs(2467));
    outputs(592) <= layer4_outputs(2460);
    outputs(593) <= not(layer4_outputs(575));
    outputs(594) <= not(layer4_outputs(28));
    outputs(595) <= not(layer4_outputs(1241));
    outputs(596) <= layer4_outputs(942);
    outputs(597) <= (layer4_outputs(1511)) or (layer4_outputs(2163));
    outputs(598) <= (layer4_outputs(552)) and not (layer4_outputs(919));
    outputs(599) <= not(layer4_outputs(960));
    outputs(600) <= not(layer4_outputs(1569));
    outputs(601) <= layer4_outputs(1859);
    outputs(602) <= layer4_outputs(1783);
    outputs(603) <= not(layer4_outputs(378));
    outputs(604) <= layer4_outputs(2165);
    outputs(605) <= not(layer4_outputs(2350)) or (layer4_outputs(2035));
    outputs(606) <= layer4_outputs(212);
    outputs(607) <= (layer4_outputs(1667)) and (layer4_outputs(2262));
    outputs(608) <= not(layer4_outputs(1073)) or (layer4_outputs(1258));
    outputs(609) <= (layer4_outputs(714)) and not (layer4_outputs(1142));
    outputs(610) <= not(layer4_outputs(1676));
    outputs(611) <= (layer4_outputs(2505)) or (layer4_outputs(1925));
    outputs(612) <= layer4_outputs(547);
    outputs(613) <= (layer4_outputs(1649)) and not (layer4_outputs(1559));
    outputs(614) <= not(layer4_outputs(724));
    outputs(615) <= not(layer4_outputs(1228));
    outputs(616) <= not(layer4_outputs(2511));
    outputs(617) <= not((layer4_outputs(2300)) xor (layer4_outputs(420)));
    outputs(618) <= layer4_outputs(542);
    outputs(619) <= (layer4_outputs(1869)) xor (layer4_outputs(2069));
    outputs(620) <= layer4_outputs(431);
    outputs(621) <= not(layer4_outputs(338));
    outputs(622) <= not(layer4_outputs(505));
    outputs(623) <= not(layer4_outputs(1032));
    outputs(624) <= layer4_outputs(1111);
    outputs(625) <= not(layer4_outputs(1994));
    outputs(626) <= not(layer4_outputs(392));
    outputs(627) <= layer4_outputs(1355);
    outputs(628) <= (layer4_outputs(930)) and not (layer4_outputs(126));
    outputs(629) <= not(layer4_outputs(1514));
    outputs(630) <= layer4_outputs(1272);
    outputs(631) <= layer4_outputs(572);
    outputs(632) <= layer4_outputs(192);
    outputs(633) <= not(layer4_outputs(355)) or (layer4_outputs(343));
    outputs(634) <= not(layer4_outputs(1675));
    outputs(635) <= not((layer4_outputs(346)) or (layer4_outputs(2531)));
    outputs(636) <= '1';
    outputs(637) <= layer4_outputs(954);
    outputs(638) <= layer4_outputs(1020);
    outputs(639) <= not(layer4_outputs(1264));
    outputs(640) <= (layer4_outputs(592)) or (layer4_outputs(1696));
    outputs(641) <= not((layer4_outputs(1817)) xor (layer4_outputs(1918)));
    outputs(642) <= not(layer4_outputs(752));
    outputs(643) <= not(layer4_outputs(2556));
    outputs(644) <= not(layer4_outputs(621));
    outputs(645) <= not((layer4_outputs(1573)) and (layer4_outputs(1387)));
    outputs(646) <= not((layer4_outputs(460)) xor (layer4_outputs(1446)));
    outputs(647) <= layer4_outputs(23);
    outputs(648) <= layer4_outputs(384);
    outputs(649) <= not(layer4_outputs(2243));
    outputs(650) <= layer4_outputs(827);
    outputs(651) <= not(layer4_outputs(2065));
    outputs(652) <= not(layer4_outputs(614)) or (layer4_outputs(877));
    outputs(653) <= (layer4_outputs(1195)) xor (layer4_outputs(223));
    outputs(654) <= (layer4_outputs(1215)) xor (layer4_outputs(285));
    outputs(655) <= not(layer4_outputs(840));
    outputs(656) <= (layer4_outputs(640)) or (layer4_outputs(156));
    outputs(657) <= not(layer4_outputs(61));
    outputs(658) <= layer4_outputs(2174);
    outputs(659) <= layer4_outputs(535);
    outputs(660) <= (layer4_outputs(2368)) and not (layer4_outputs(1776));
    outputs(661) <= not((layer4_outputs(1772)) or (layer4_outputs(2318)));
    outputs(662) <= not(layer4_outputs(267)) or (layer4_outputs(2344));
    outputs(663) <= (layer4_outputs(2469)) xor (layer4_outputs(763));
    outputs(664) <= not((layer4_outputs(969)) xor (layer4_outputs(955)));
    outputs(665) <= (layer4_outputs(286)) and not (layer4_outputs(2062));
    outputs(666) <= not(layer4_outputs(1046));
    outputs(667) <= layer4_outputs(2124);
    outputs(668) <= not((layer4_outputs(2294)) and (layer4_outputs(519)));
    outputs(669) <= layer4_outputs(2016);
    outputs(670) <= not(layer4_outputs(260));
    outputs(671) <= not(layer4_outputs(1961));
    outputs(672) <= layer4_outputs(1354);
    outputs(673) <= not(layer4_outputs(2132));
    outputs(674) <= not(layer4_outputs(927));
    outputs(675) <= (layer4_outputs(496)) and not (layer4_outputs(808));
    outputs(676) <= not(layer4_outputs(1805));
    outputs(677) <= (layer4_outputs(1479)) xor (layer4_outputs(2196));
    outputs(678) <= not(layer4_outputs(1709));
    outputs(679) <= layer4_outputs(1401);
    outputs(680) <= (layer4_outputs(1233)) and (layer4_outputs(1475));
    outputs(681) <= not((layer4_outputs(612)) xor (layer4_outputs(135)));
    outputs(682) <= layer4_outputs(289);
    outputs(683) <= not(layer4_outputs(2261));
    outputs(684) <= not(layer4_outputs(204));
    outputs(685) <= not(layer4_outputs(507));
    outputs(686) <= not(layer4_outputs(610));
    outputs(687) <= not(layer4_outputs(1554));
    outputs(688) <= (layer4_outputs(1193)) xor (layer4_outputs(1468));
    outputs(689) <= not(layer4_outputs(1306));
    outputs(690) <= layer4_outputs(637);
    outputs(691) <= not((layer4_outputs(2084)) or (layer4_outputs(1681)));
    outputs(692) <= (layer4_outputs(2422)) or (layer4_outputs(110));
    outputs(693) <= not(layer4_outputs(845)) or (layer4_outputs(2142));
    outputs(694) <= layer4_outputs(2403);
    outputs(695) <= (layer4_outputs(1047)) and not (layer4_outputs(764));
    outputs(696) <= not((layer4_outputs(1525)) xor (layer4_outputs(1232)));
    outputs(697) <= not(layer4_outputs(2427)) or (layer4_outputs(1441));
    outputs(698) <= not(layer4_outputs(2355));
    outputs(699) <= layer4_outputs(192);
    outputs(700) <= not(layer4_outputs(1754));
    outputs(701) <= not((layer4_outputs(503)) xor (layer4_outputs(678)));
    outputs(702) <= (layer4_outputs(805)) and not (layer4_outputs(43));
    outputs(703) <= not(layer4_outputs(200));
    outputs(704) <= layer4_outputs(841);
    outputs(705) <= layer4_outputs(2280);
    outputs(706) <= (layer4_outputs(1120)) or (layer4_outputs(124));
    outputs(707) <= layer4_outputs(2016);
    outputs(708) <= not(layer4_outputs(848));
    outputs(709) <= not((layer4_outputs(2022)) xor (layer4_outputs(1910)));
    outputs(710) <= not(layer4_outputs(1969));
    outputs(711) <= (layer4_outputs(1877)) and not (layer4_outputs(1167));
    outputs(712) <= not(layer4_outputs(782));
    outputs(713) <= not(layer4_outputs(207));
    outputs(714) <= not(layer4_outputs(344));
    outputs(715) <= not((layer4_outputs(366)) and (layer4_outputs(2178)));
    outputs(716) <= not(layer4_outputs(2250));
    outputs(717) <= layer4_outputs(1729);
    outputs(718) <= not(layer4_outputs(2160));
    outputs(719) <= layer4_outputs(1323);
    outputs(720) <= not((layer4_outputs(79)) and (layer4_outputs(1630)));
    outputs(721) <= (layer4_outputs(2477)) and not (layer4_outputs(712));
    outputs(722) <= layer4_outputs(1397);
    outputs(723) <= not(layer4_outputs(1347));
    outputs(724) <= not(layer4_outputs(566));
    outputs(725) <= not(layer4_outputs(1599));
    outputs(726) <= not(layer4_outputs(2206));
    outputs(727) <= (layer4_outputs(609)) and not (layer4_outputs(2478));
    outputs(728) <= not(layer4_outputs(1425));
    outputs(729) <= layer4_outputs(1558);
    outputs(730) <= not(layer4_outputs(1368));
    outputs(731) <= not(layer4_outputs(1978));
    outputs(732) <= layer4_outputs(1550);
    outputs(733) <= not((layer4_outputs(1022)) or (layer4_outputs(1128)));
    outputs(734) <= not(layer4_outputs(2327));
    outputs(735) <= layer4_outputs(769);
    outputs(736) <= layer4_outputs(2529);
    outputs(737) <= (layer4_outputs(1756)) and not (layer4_outputs(146));
    outputs(738) <= (layer4_outputs(67)) xor (layer4_outputs(896));
    outputs(739) <= layer4_outputs(1786);
    outputs(740) <= (layer4_outputs(1880)) xor (layer4_outputs(1755));
    outputs(741) <= layer4_outputs(1107);
    outputs(742) <= layer4_outputs(1011);
    outputs(743) <= not(layer4_outputs(505));
    outputs(744) <= not(layer4_outputs(264));
    outputs(745) <= layer4_outputs(2158);
    outputs(746) <= not((layer4_outputs(1819)) and (layer4_outputs(1873)));
    outputs(747) <= not((layer4_outputs(310)) or (layer4_outputs(1094)));
    outputs(748) <= (layer4_outputs(262)) or (layer4_outputs(1555));
    outputs(749) <= not(layer4_outputs(2533));
    outputs(750) <= layer4_outputs(1088);
    outputs(751) <= not(layer4_outputs(1380));
    outputs(752) <= (layer4_outputs(2266)) and not (layer4_outputs(536));
    outputs(753) <= (layer4_outputs(210)) or (layer4_outputs(69));
    outputs(754) <= (layer4_outputs(698)) and (layer4_outputs(2075));
    outputs(755) <= not(layer4_outputs(831));
    outputs(756) <= not(layer4_outputs(1288));
    outputs(757) <= layer4_outputs(1711);
    outputs(758) <= not(layer4_outputs(2121)) or (layer4_outputs(2081));
    outputs(759) <= not(layer4_outputs(197));
    outputs(760) <= (layer4_outputs(400)) and not (layer4_outputs(2492));
    outputs(761) <= layer4_outputs(1731);
    outputs(762) <= layer4_outputs(22);
    outputs(763) <= not(layer4_outputs(1240));
    outputs(764) <= not(layer4_outputs(1706));
    outputs(765) <= layer4_outputs(1350);
    outputs(766) <= layer4_outputs(2283);
    outputs(767) <= layer4_outputs(1294);
    outputs(768) <= layer4_outputs(1205);
    outputs(769) <= layer4_outputs(340);
    outputs(770) <= not((layer4_outputs(587)) or (layer4_outputs(885)));
    outputs(771) <= (layer4_outputs(1911)) and not (layer4_outputs(363));
    outputs(772) <= layer4_outputs(161);
    outputs(773) <= layer4_outputs(950);
    outputs(774) <= layer4_outputs(696);
    outputs(775) <= layer4_outputs(558);
    outputs(776) <= layer4_outputs(79);
    outputs(777) <= (layer4_outputs(843)) or (layer4_outputs(1094));
    outputs(778) <= not(layer4_outputs(652));
    outputs(779) <= not((layer4_outputs(707)) and (layer4_outputs(1462)));
    outputs(780) <= (layer4_outputs(2186)) and not (layer4_outputs(2440));
    outputs(781) <= not((layer4_outputs(1702)) or (layer4_outputs(585)));
    outputs(782) <= not((layer4_outputs(1501)) or (layer4_outputs(339)));
    outputs(783) <= not(layer4_outputs(1456));
    outputs(784) <= not(layer4_outputs(81));
    outputs(785) <= (layer4_outputs(2135)) or (layer4_outputs(1912));
    outputs(786) <= not(layer4_outputs(1394));
    outputs(787) <= layer4_outputs(1914);
    outputs(788) <= layer4_outputs(183);
    outputs(789) <= layer4_outputs(1900);
    outputs(790) <= (layer4_outputs(1402)) and not (layer4_outputs(772));
    outputs(791) <= not(layer4_outputs(2227));
    outputs(792) <= not(layer4_outputs(1439));
    outputs(793) <= layer4_outputs(1311);
    outputs(794) <= not(layer4_outputs(915));
    outputs(795) <= not(layer4_outputs(881));
    outputs(796) <= not(layer4_outputs(1326));
    outputs(797) <= (layer4_outputs(164)) xor (layer4_outputs(1609));
    outputs(798) <= layer4_outputs(1305);
    outputs(799) <= layer4_outputs(1160);
    outputs(800) <= not(layer4_outputs(1562));
    outputs(801) <= not(layer4_outputs(701));
    outputs(802) <= layer4_outputs(883);
    outputs(803) <= not((layer4_outputs(940)) xor (layer4_outputs(606)));
    outputs(804) <= not(layer4_outputs(1253));
    outputs(805) <= not(layer4_outputs(1335));
    outputs(806) <= layer4_outputs(639);
    outputs(807) <= layer4_outputs(1348);
    outputs(808) <= layer4_outputs(1520);
    outputs(809) <= layer4_outputs(1330);
    outputs(810) <= layer4_outputs(746);
    outputs(811) <= not(layer4_outputs(2328));
    outputs(812) <= not(layer4_outputs(722));
    outputs(813) <= not((layer4_outputs(1826)) or (layer4_outputs(1939)));
    outputs(814) <= not(layer4_outputs(1138));
    outputs(815) <= not(layer4_outputs(2439));
    outputs(816) <= not(layer4_outputs(37));
    outputs(817) <= layer4_outputs(2429);
    outputs(818) <= not(layer4_outputs(1340));
    outputs(819) <= (layer4_outputs(793)) and not (layer4_outputs(540));
    outputs(820) <= layer4_outputs(1836);
    outputs(821) <= layer4_outputs(2004);
    outputs(822) <= (layer4_outputs(2134)) and (layer4_outputs(1591));
    outputs(823) <= not(layer4_outputs(1697));
    outputs(824) <= not(layer4_outputs(1503));
    outputs(825) <= layer4_outputs(2283);
    outputs(826) <= layer4_outputs(2309);
    outputs(827) <= not(layer4_outputs(900));
    outputs(828) <= layer4_outputs(3);
    outputs(829) <= not((layer4_outputs(1651)) xor (layer4_outputs(280)));
    outputs(830) <= layer4_outputs(2151);
    outputs(831) <= not((layer4_outputs(875)) and (layer4_outputs(1609)));
    outputs(832) <= not(layer4_outputs(1879));
    outputs(833) <= not((layer4_outputs(867)) and (layer4_outputs(1456)));
    outputs(834) <= (layer4_outputs(514)) xor (layer4_outputs(1161));
    outputs(835) <= not((layer4_outputs(1201)) and (layer4_outputs(107)));
    outputs(836) <= not(layer4_outputs(141)) or (layer4_outputs(1745));
    outputs(837) <= not(layer4_outputs(2347));
    outputs(838) <= not(layer4_outputs(1576));
    outputs(839) <= layer4_outputs(1062);
    outputs(840) <= not((layer4_outputs(55)) xor (layer4_outputs(1441)));
    outputs(841) <= not(layer4_outputs(1948));
    outputs(842) <= not(layer4_outputs(131));
    outputs(843) <= (layer4_outputs(1718)) and not (layer4_outputs(744));
    outputs(844) <= layer4_outputs(179);
    outputs(845) <= not((layer4_outputs(988)) or (layer4_outputs(917)));
    outputs(846) <= layer4_outputs(274);
    outputs(847) <= layer4_outputs(627);
    outputs(848) <= layer4_outputs(998);
    outputs(849) <= not(layer4_outputs(1417));
    outputs(850) <= not(layer4_outputs(1528));
    outputs(851) <= not(layer4_outputs(1377));
    outputs(852) <= layer4_outputs(1772);
    outputs(853) <= not((layer4_outputs(1789)) or (layer4_outputs(1023)));
    outputs(854) <= (layer4_outputs(2415)) xor (layer4_outputs(1722));
    outputs(855) <= not(layer4_outputs(822));
    outputs(856) <= layer4_outputs(1964);
    outputs(857) <= layer4_outputs(1109);
    outputs(858) <= not(layer4_outputs(2331));
    outputs(859) <= layer4_outputs(597);
    outputs(860) <= (layer4_outputs(2458)) and not (layer4_outputs(1487));
    outputs(861) <= not((layer4_outputs(2258)) or (layer4_outputs(854)));
    outputs(862) <= not(layer4_outputs(2360));
    outputs(863) <= not((layer4_outputs(1661)) xor (layer4_outputs(875)));
    outputs(864) <= layer4_outputs(1574);
    outputs(865) <= layer4_outputs(1480);
    outputs(866) <= layer4_outputs(92);
    outputs(867) <= layer4_outputs(1242);
    outputs(868) <= layer4_outputs(1433);
    outputs(869) <= (layer4_outputs(1502)) and (layer4_outputs(483));
    outputs(870) <= not((layer4_outputs(71)) or (layer4_outputs(2107)));
    outputs(871) <= layer4_outputs(1007);
    outputs(872) <= layer4_outputs(454);
    outputs(873) <= not((layer4_outputs(632)) or (layer4_outputs(1719)));
    outputs(874) <= (layer4_outputs(14)) and not (layer4_outputs(1898));
    outputs(875) <= (layer4_outputs(66)) and not (layer4_outputs(1174));
    outputs(876) <= not(layer4_outputs(2259));
    outputs(877) <= not(layer4_outputs(789)) or (layer4_outputs(2370));
    outputs(878) <= layer4_outputs(767);
    outputs(879) <= layer4_outputs(1151);
    outputs(880) <= layer4_outputs(281);
    outputs(881) <= layer4_outputs(830);
    outputs(882) <= not(layer4_outputs(2450));
    outputs(883) <= not(layer4_outputs(846));
    outputs(884) <= not(layer4_outputs(1808));
    outputs(885) <= (layer4_outputs(347)) and not (layer4_outputs(139));
    outputs(886) <= layer4_outputs(2231);
    outputs(887) <= (layer4_outputs(895)) and not (layer4_outputs(1867));
    outputs(888) <= not((layer4_outputs(677)) or (layer4_outputs(1568)));
    outputs(889) <= not(layer4_outputs(642));
    outputs(890) <= layer4_outputs(2359);
    outputs(891) <= not(layer4_outputs(2554));
    outputs(892) <= (layer4_outputs(297)) and not (layer4_outputs(1999));
    outputs(893) <= (layer4_outputs(2077)) xor (layer4_outputs(465));
    outputs(894) <= layer4_outputs(257);
    outputs(895) <= (layer4_outputs(2333)) and not (layer4_outputs(1207));
    outputs(896) <= not(layer4_outputs(1751));
    outputs(897) <= (layer4_outputs(936)) and not (layer4_outputs(1846));
    outputs(898) <= (layer4_outputs(458)) and not (layer4_outputs(885));
    outputs(899) <= layer4_outputs(2383);
    outputs(900) <= not(layer4_outputs(584));
    outputs(901) <= not(layer4_outputs(846));
    outputs(902) <= (layer4_outputs(2421)) and (layer4_outputs(2380));
    outputs(903) <= not(layer4_outputs(1097));
    outputs(904) <= not(layer4_outputs(674));
    outputs(905) <= (layer4_outputs(1742)) and not (layer4_outputs(2073));
    outputs(906) <= layer4_outputs(2507);
    outputs(907) <= layer4_outputs(72);
    outputs(908) <= not(layer4_outputs(2252));
    outputs(909) <= not(layer4_outputs(1687));
    outputs(910) <= not(layer4_outputs(1687));
    outputs(911) <= layer4_outputs(1028);
    outputs(912) <= not((layer4_outputs(1512)) xor (layer4_outputs(1415)));
    outputs(913) <= not(layer4_outputs(1327));
    outputs(914) <= not(layer4_outputs(1646)) or (layer4_outputs(1052));
    outputs(915) <= not(layer4_outputs(2218));
    outputs(916) <= (layer4_outputs(989)) xor (layer4_outputs(1905));
    outputs(917) <= layer4_outputs(1006);
    outputs(918) <= not((layer4_outputs(1124)) or (layer4_outputs(2521)));
    outputs(919) <= layer4_outputs(648);
    outputs(920) <= layer4_outputs(577);
    outputs(921) <= not(layer4_outputs(2156));
    outputs(922) <= not(layer4_outputs(1400));
    outputs(923) <= layer4_outputs(904);
    outputs(924) <= layer4_outputs(1041);
    outputs(925) <= not(layer4_outputs(1198));
    outputs(926) <= (layer4_outputs(2261)) and not (layer4_outputs(1813));
    outputs(927) <= layer4_outputs(920);
    outputs(928) <= not(layer4_outputs(903));
    outputs(929) <= layer4_outputs(1655);
    outputs(930) <= not(layer4_outputs(1124));
    outputs(931) <= not(layer4_outputs(2194));
    outputs(932) <= layer4_outputs(1312);
    outputs(933) <= not(layer4_outputs(2442));
    outputs(934) <= layer4_outputs(1202);
    outputs(935) <= layer4_outputs(2312);
    outputs(936) <= not(layer4_outputs(2187));
    outputs(937) <= not((layer4_outputs(720)) or (layer4_outputs(2110)));
    outputs(938) <= (layer4_outputs(27)) xor (layer4_outputs(799));
    outputs(939) <= layer4_outputs(1951);
    outputs(940) <= layer4_outputs(2512);
    outputs(941) <= (layer4_outputs(2251)) and not (layer4_outputs(512));
    outputs(942) <= (layer4_outputs(1167)) and not (layer4_outputs(721));
    outputs(943) <= not(layer4_outputs(1277));
    outputs(944) <= not(layer4_outputs(2007));
    outputs(945) <= (layer4_outputs(961)) xor (layer4_outputs(897));
    outputs(946) <= (layer4_outputs(516)) and not (layer4_outputs(2474));
    outputs(947) <= not(layer4_outputs(722));
    outputs(948) <= (layer4_outputs(2153)) xor (layer4_outputs(96));
    outputs(949) <= (layer4_outputs(445)) and (layer4_outputs(1450));
    outputs(950) <= layer4_outputs(910);
    outputs(951) <= (layer4_outputs(58)) and not (layer4_outputs(1743));
    outputs(952) <= not(layer4_outputs(1528));
    outputs(953) <= not((layer4_outputs(710)) and (layer4_outputs(1236)));
    outputs(954) <= (layer4_outputs(1316)) and (layer4_outputs(2233));
    outputs(955) <= (layer4_outputs(659)) and (layer4_outputs(2310));
    outputs(956) <= layer4_outputs(1398);
    outputs(957) <= layer4_outputs(982);
    outputs(958) <= (layer4_outputs(1303)) or (layer4_outputs(2066));
    outputs(959) <= not((layer4_outputs(965)) xor (layer4_outputs(1787)));
    outputs(960) <= layer4_outputs(77);
    outputs(961) <= (layer4_outputs(73)) xor (layer4_outputs(489));
    outputs(962) <= layer4_outputs(2001);
    outputs(963) <= not(layer4_outputs(2486)) or (layer4_outputs(1519));
    outputs(964) <= not(layer4_outputs(2455));
    outputs(965) <= (layer4_outputs(2011)) and not (layer4_outputs(1732));
    outputs(966) <= layer4_outputs(1633);
    outputs(967) <= (layer4_outputs(1013)) and (layer4_outputs(1486));
    outputs(968) <= (layer4_outputs(1673)) and not (layer4_outputs(2032));
    outputs(969) <= layer4_outputs(1931);
    outputs(970) <= (layer4_outputs(1333)) xor (layer4_outputs(1139));
    outputs(971) <= (layer4_outputs(347)) and not (layer4_outputs(1878));
    outputs(972) <= not(layer4_outputs(1173));
    outputs(973) <= layer4_outputs(1062);
    outputs(974) <= not(layer4_outputs(299));
    outputs(975) <= layer4_outputs(2451);
    outputs(976) <= layer4_outputs(688);
    outputs(977) <= layer4_outputs(648);
    outputs(978) <= (layer4_outputs(1011)) and not (layer4_outputs(446));
    outputs(979) <= layer4_outputs(1499);
    outputs(980) <= layer4_outputs(380);
    outputs(981) <= not((layer4_outputs(39)) xor (layer4_outputs(1353)));
    outputs(982) <= not(layer4_outputs(1511));
    outputs(983) <= not((layer4_outputs(390)) and (layer4_outputs(104)));
    outputs(984) <= (layer4_outputs(1941)) and (layer4_outputs(1746));
    outputs(985) <= (layer4_outputs(1063)) and not (layer4_outputs(1255));
    outputs(986) <= not(layer4_outputs(1209));
    outputs(987) <= layer4_outputs(1543);
    outputs(988) <= not(layer4_outputs(1));
    outputs(989) <= not(layer4_outputs(2453));
    outputs(990) <= layer4_outputs(968);
    outputs(991) <= (layer4_outputs(1897)) and (layer4_outputs(2516));
    outputs(992) <= not((layer4_outputs(1112)) or (layer4_outputs(1750)));
    outputs(993) <= layer4_outputs(1232);
    outputs(994) <= layer4_outputs(2092);
    outputs(995) <= not((layer4_outputs(1871)) or (layer4_outputs(2481)));
    outputs(996) <= not(layer4_outputs(479));
    outputs(997) <= not(layer4_outputs(788));
    outputs(998) <= not(layer4_outputs(1664));
    outputs(999) <= layer4_outputs(1996);
    outputs(1000) <= layer4_outputs(211);
    outputs(1001) <= not(layer4_outputs(56));
    outputs(1002) <= (layer4_outputs(709)) and not (layer4_outputs(943));
    outputs(1003) <= not(layer4_outputs(592));
    outputs(1004) <= (layer4_outputs(1084)) and not (layer4_outputs(2158));
    outputs(1005) <= layer4_outputs(945);
    outputs(1006) <= (layer4_outputs(2473)) and (layer4_outputs(665));
    outputs(1007) <= not((layer4_outputs(63)) or (layer4_outputs(2375)));
    outputs(1008) <= layer4_outputs(237);
    outputs(1009) <= (layer4_outputs(206)) xor (layer4_outputs(2501));
    outputs(1010) <= not(layer4_outputs(1235));
    outputs(1011) <= (layer4_outputs(1128)) and (layer4_outputs(1496));
    outputs(1012) <= (layer4_outputs(158)) xor (layer4_outputs(59));
    outputs(1013) <= not((layer4_outputs(2085)) and (layer4_outputs(970)));
    outputs(1014) <= not(layer4_outputs(1666));
    outputs(1015) <= layer4_outputs(330);
    outputs(1016) <= layer4_outputs(1917);
    outputs(1017) <= layer4_outputs(862);
    outputs(1018) <= layer4_outputs(1640);
    outputs(1019) <= not(layer4_outputs(2063));
    outputs(1020) <= layer4_outputs(72);
    outputs(1021) <= (layer4_outputs(2119)) and (layer4_outputs(2139));
    outputs(1022) <= not((layer4_outputs(682)) or (layer4_outputs(2314)));
    outputs(1023) <= not((layer4_outputs(358)) xor (layer4_outputs(1762)));
    outputs(1024) <= (layer4_outputs(338)) and not (layer4_outputs(88));
    outputs(1025) <= not(layer4_outputs(379));
    outputs(1026) <= layer4_outputs(2356);
    outputs(1027) <= layer4_outputs(241);
    outputs(1028) <= not(layer4_outputs(2384));
    outputs(1029) <= (layer4_outputs(1483)) or (layer4_outputs(1540));
    outputs(1030) <= layer4_outputs(1064);
    outputs(1031) <= (layer4_outputs(2039)) and not (layer4_outputs(2322));
    outputs(1032) <= not(layer4_outputs(1852));
    outputs(1033) <= not(layer4_outputs(2401));
    outputs(1034) <= layer4_outputs(2143);
    outputs(1035) <= not((layer4_outputs(2390)) and (layer4_outputs(202)));
    outputs(1036) <= layer4_outputs(1214);
    outputs(1037) <= layer4_outputs(1553);
    outputs(1038) <= layer4_outputs(1774);
    outputs(1039) <= layer4_outputs(2528);
    outputs(1040) <= (layer4_outputs(420)) xor (layer4_outputs(1307));
    outputs(1041) <= not((layer4_outputs(2189)) xor (layer4_outputs(1623)));
    outputs(1042) <= not(layer4_outputs(576));
    outputs(1043) <= (layer4_outputs(2553)) or (layer4_outputs(1582));
    outputs(1044) <= not(layer4_outputs(1784));
    outputs(1045) <= (layer4_outputs(1027)) and not (layer4_outputs(1639));
    outputs(1046) <= layer4_outputs(708);
    outputs(1047) <= layer4_outputs(182);
    outputs(1048) <= layer4_outputs(2398);
    outputs(1049) <= (layer4_outputs(107)) and not (layer4_outputs(1408));
    outputs(1050) <= not(layer4_outputs(680));
    outputs(1051) <= not(layer4_outputs(1602));
    outputs(1052) <= layer4_outputs(1949);
    outputs(1053) <= layer4_outputs(409);
    outputs(1054) <= not(layer4_outputs(980)) or (layer4_outputs(336));
    outputs(1055) <= not(layer4_outputs(361));
    outputs(1056) <= not(layer4_outputs(582));
    outputs(1057) <= not((layer4_outputs(2125)) xor (layer4_outputs(2137)));
    outputs(1058) <= layer4_outputs(1986);
    outputs(1059) <= (layer4_outputs(1078)) and not (layer4_outputs(1426));
    outputs(1060) <= (layer4_outputs(401)) and (layer4_outputs(2391));
    outputs(1061) <= not(layer4_outputs(2363));
    outputs(1062) <= layer4_outputs(1871);
    outputs(1063) <= not(layer4_outputs(1031));
    outputs(1064) <= not(layer4_outputs(1344)) or (layer4_outputs(1861));
    outputs(1065) <= not(layer4_outputs(462)) or (layer4_outputs(1042));
    outputs(1066) <= not((layer4_outputs(883)) or (layer4_outputs(1163)));
    outputs(1067) <= layer4_outputs(1587);
    outputs(1068) <= layer4_outputs(1796);
    outputs(1069) <= layer4_outputs(1114);
    outputs(1070) <= not(layer4_outputs(2315));
    outputs(1071) <= not(layer4_outputs(183));
    outputs(1072) <= not((layer4_outputs(1440)) or (layer4_outputs(1153)));
    outputs(1073) <= layer4_outputs(2094);
    outputs(1074) <= not(layer4_outputs(246));
    outputs(1075) <= (layer4_outputs(155)) and not (layer4_outputs(168));
    outputs(1076) <= layer4_outputs(1481);
    outputs(1077) <= not(layer4_outputs(2248));
    outputs(1078) <= not((layer4_outputs(2276)) or (layer4_outputs(358)));
    outputs(1079) <= layer4_outputs(1359);
    outputs(1080) <= not(layer4_outputs(2031));
    outputs(1081) <= not(layer4_outputs(863));
    outputs(1082) <= layer4_outputs(1846);
    outputs(1083) <= (layer4_outputs(929)) and not (layer4_outputs(2422));
    outputs(1084) <= layer4_outputs(2339);
    outputs(1085) <= not(layer4_outputs(2388));
    outputs(1086) <= not(layer4_outputs(1283));
    outputs(1087) <= layer4_outputs(8);
    outputs(1088) <= layer4_outputs(1363);
    outputs(1089) <= layer4_outputs(1291);
    outputs(1090) <= layer4_outputs(858);
    outputs(1091) <= layer4_outputs(1209);
    outputs(1092) <= layer4_outputs(1328);
    outputs(1093) <= not(layer4_outputs(1145));
    outputs(1094) <= (layer4_outputs(118)) and not (layer4_outputs(40));
    outputs(1095) <= layer4_outputs(2127);
    outputs(1096) <= not((layer4_outputs(2420)) or (layer4_outputs(64)));
    outputs(1097) <= (layer4_outputs(2394)) and not (layer4_outputs(1688));
    outputs(1098) <= not(layer4_outputs(198));
    outputs(1099) <= layer4_outputs(571);
    outputs(1100) <= layer4_outputs(538);
    outputs(1101) <= (layer4_outputs(758)) and not (layer4_outputs(1279));
    outputs(1102) <= (layer4_outputs(837)) and not (layer4_outputs(1293));
    outputs(1103) <= not(layer4_outputs(2358));
    outputs(1104) <= (layer4_outputs(739)) xor (layer4_outputs(1980));
    outputs(1105) <= layer4_outputs(700);
    outputs(1106) <= not(layer4_outputs(1126));
    outputs(1107) <= layer4_outputs(1945);
    outputs(1108) <= layer4_outputs(1429);
    outputs(1109) <= not(layer4_outputs(1116));
    outputs(1110) <= not(layer4_outputs(2083));
    outputs(1111) <= not((layer4_outputs(312)) xor (layer4_outputs(1668)));
    outputs(1112) <= (layer4_outputs(810)) and (layer4_outputs(1114));
    outputs(1113) <= layer4_outputs(1210);
    outputs(1114) <= layer4_outputs(1235);
    outputs(1115) <= not(layer4_outputs(1056));
    outputs(1116) <= (layer4_outputs(824)) and not (layer4_outputs(246));
    outputs(1117) <= (layer4_outputs(2371)) xor (layer4_outputs(2183));
    outputs(1118) <= layer4_outputs(1121);
    outputs(1119) <= not(layer4_outputs(1319));
    outputs(1120) <= layer4_outputs(1410);
    outputs(1121) <= not(layer4_outputs(2099));
    outputs(1122) <= layer4_outputs(413);
    outputs(1123) <= not(layer4_outputs(6));
    outputs(1124) <= not((layer4_outputs(261)) xor (layer4_outputs(1455)));
    outputs(1125) <= not(layer4_outputs(30));
    outputs(1126) <= layer4_outputs(1976);
    outputs(1127) <= layer4_outputs(1032);
    outputs(1128) <= (layer4_outputs(1997)) and not (layer4_outputs(511));
    outputs(1129) <= (layer4_outputs(1582)) or (layer4_outputs(1494));
    outputs(1130) <= not(layer4_outputs(1390));
    outputs(1131) <= layer4_outputs(817);
    outputs(1132) <= (layer4_outputs(2257)) and (layer4_outputs(1202));
    outputs(1133) <= layer4_outputs(167);
    outputs(1134) <= not(layer4_outputs(2083));
    outputs(1135) <= not(layer4_outputs(1584));
    outputs(1136) <= not((layer4_outputs(1019)) xor (layer4_outputs(411)));
    outputs(1137) <= not(layer4_outputs(500));
    outputs(1138) <= layer4_outputs(502);
    outputs(1139) <= (layer4_outputs(2175)) and not (layer4_outputs(377));
    outputs(1140) <= (layer4_outputs(731)) and not (layer4_outputs(802));
    outputs(1141) <= not((layer4_outputs(683)) or (layer4_outputs(1051)));
    outputs(1142) <= layer4_outputs(1859);
    outputs(1143) <= not((layer4_outputs(850)) and (layer4_outputs(497)));
    outputs(1144) <= layer4_outputs(1263);
    outputs(1145) <= not(layer4_outputs(695));
    outputs(1146) <= layer4_outputs(2123);
    outputs(1147) <= layer4_outputs(971);
    outputs(1148) <= (layer4_outputs(1193)) xor (layer4_outputs(410));
    outputs(1149) <= not((layer4_outputs(1673)) or (layer4_outputs(1281)));
    outputs(1150) <= (layer4_outputs(681)) xor (layer4_outputs(855));
    outputs(1151) <= not(layer4_outputs(2156));
    outputs(1152) <= not(layer4_outputs(2416));
    outputs(1153) <= layer4_outputs(1420);
    outputs(1154) <= (layer4_outputs(1554)) and (layer4_outputs(1199));
    outputs(1155) <= not(layer4_outputs(1660));
    outputs(1156) <= layer4_outputs(459);
    outputs(1157) <= not((layer4_outputs(381)) or (layer4_outputs(2244)));
    outputs(1158) <= layer4_outputs(1518);
    outputs(1159) <= layer4_outputs(800);
    outputs(1160) <= layer4_outputs(1237);
    outputs(1161) <= (layer4_outputs(1161)) xor (layer4_outputs(2136));
    outputs(1162) <= not(layer4_outputs(2071));
    outputs(1163) <= not(layer4_outputs(1295));
    outputs(1164) <= not(layer4_outputs(2545));
    outputs(1165) <= not(layer4_outputs(2320));
    outputs(1166) <= not(layer4_outputs(1395));
    outputs(1167) <= (layer4_outputs(1028)) xor (layer4_outputs(630));
    outputs(1168) <= (layer4_outputs(1218)) and not (layer4_outputs(2285));
    outputs(1169) <= not(layer4_outputs(318));
    outputs(1170) <= layer4_outputs(899);
    outputs(1171) <= (layer4_outputs(1705)) or (layer4_outputs(742));
    outputs(1172) <= not(layer4_outputs(486));
    outputs(1173) <= (layer4_outputs(418)) and not (layer4_outputs(256));
    outputs(1174) <= layer4_outputs(1847);
    outputs(1175) <= not(layer4_outputs(1829));
    outputs(1176) <= (layer4_outputs(125)) xor (layer4_outputs(206));
    outputs(1177) <= not(layer4_outputs(2341));
    outputs(1178) <= layer4_outputs(1350);
    outputs(1179) <= not(layer4_outputs(1865));
    outputs(1180) <= (layer4_outputs(2236)) and not (layer4_outputs(352));
    outputs(1181) <= not((layer4_outputs(777)) or (layer4_outputs(383)));
    outputs(1182) <= not(layer4_outputs(2446));
    outputs(1183) <= not(layer4_outputs(1733));
    outputs(1184) <= not(layer4_outputs(1595));
    outputs(1185) <= not(layer4_outputs(185));
    outputs(1186) <= (layer4_outputs(1078)) and not (layer4_outputs(753));
    outputs(1187) <= not(layer4_outputs(791));
    outputs(1188) <= (layer4_outputs(1442)) and not (layer4_outputs(2203));
    outputs(1189) <= layer4_outputs(1378);
    outputs(1190) <= layer4_outputs(854);
    outputs(1191) <= (layer4_outputs(480)) xor (layer4_outputs(533));
    outputs(1192) <= not((layer4_outputs(1243)) xor (layer4_outputs(1764)));
    outputs(1193) <= not(layer4_outputs(1534));
    outputs(1194) <= layer4_outputs(433);
    outputs(1195) <= (layer4_outputs(1375)) and not (layer4_outputs(1484));
    outputs(1196) <= not(layer4_outputs(894));
    outputs(1197) <= not(layer4_outputs(1956));
    outputs(1198) <= not(layer4_outputs(2115));
    outputs(1199) <= layer4_outputs(2395);
    outputs(1200) <= (layer4_outputs(1478)) or (layer4_outputs(1382));
    outputs(1201) <= not((layer4_outputs(1145)) or (layer4_outputs(510)));
    outputs(1202) <= (layer4_outputs(38)) and not (layer4_outputs(1674));
    outputs(1203) <= not(layer4_outputs(1231));
    outputs(1204) <= (layer4_outputs(1090)) xor (layer4_outputs(816));
    outputs(1205) <= not(layer4_outputs(1862));
    outputs(1206) <= not(layer4_outputs(181));
    outputs(1207) <= (layer4_outputs(2267)) xor (layer4_outputs(1987));
    outputs(1208) <= layer4_outputs(2408);
    outputs(1209) <= layer4_outputs(2495);
    outputs(1210) <= (layer4_outputs(1581)) and (layer4_outputs(4));
    outputs(1211) <= layer4_outputs(1545);
    outputs(1212) <= layer4_outputs(2557);
    outputs(1213) <= not(layer4_outputs(2332));
    outputs(1214) <= (layer4_outputs(1444)) and not (layer4_outputs(2296));
    outputs(1215) <= not(layer4_outputs(1152));
    outputs(1216) <= not(layer4_outputs(2444));
    outputs(1217) <= not(layer4_outputs(2070));
    outputs(1218) <= not((layer4_outputs(650)) xor (layer4_outputs(1170)));
    outputs(1219) <= not(layer4_outputs(955));
    outputs(1220) <= not(layer4_outputs(403));
    outputs(1221) <= not(layer4_outputs(706));
    outputs(1222) <= layer4_outputs(817);
    outputs(1223) <= layer4_outputs(780);
    outputs(1224) <= not(layer4_outputs(506));
    outputs(1225) <= (layer4_outputs(373)) xor (layer4_outputs(623));
    outputs(1226) <= not((layer4_outputs(754)) or (layer4_outputs(2151)));
    outputs(1227) <= not(layer4_outputs(861));
    outputs(1228) <= not(layer4_outputs(1281));
    outputs(1229) <= not(layer4_outputs(602));
    outputs(1230) <= not(layer4_outputs(1309)) or (layer4_outputs(2499));
    outputs(1231) <= (layer4_outputs(498)) xor (layer4_outputs(1261));
    outputs(1232) <= not(layer4_outputs(2468));
    outputs(1233) <= not(layer4_outputs(1724));
    outputs(1234) <= layer4_outputs(2541);
    outputs(1235) <= not((layer4_outputs(1689)) or (layer4_outputs(923)));
    outputs(1236) <= not(layer4_outputs(934));
    outputs(1237) <= (layer4_outputs(959)) and not (layer4_outputs(1944));
    outputs(1238) <= layer4_outputs(1434);
    outputs(1239) <= layer4_outputs(682);
    outputs(1240) <= not((layer4_outputs(97)) or (layer4_outputs(1876)));
    outputs(1241) <= not((layer4_outputs(1985)) or (layer4_outputs(1740)));
    outputs(1242) <= not((layer4_outputs(1535)) or (layer4_outputs(1721)));
    outputs(1243) <= not(layer4_outputs(1959));
    outputs(1244) <= layer4_outputs(1082);
    outputs(1245) <= not(layer4_outputs(1179));
    outputs(1246) <= (layer4_outputs(126)) and (layer4_outputs(2003));
    outputs(1247) <= (layer4_outputs(404)) xor (layer4_outputs(266));
    outputs(1248) <= (layer4_outputs(1598)) and not (layer4_outputs(1332));
    outputs(1249) <= not(layer4_outputs(593));
    outputs(1250) <= (layer4_outputs(764)) and not (layer4_outputs(1745));
    outputs(1251) <= layer4_outputs(2547);
    outputs(1252) <= (layer4_outputs(1173)) and not (layer4_outputs(2209));
    outputs(1253) <= not(layer4_outputs(998));
    outputs(1254) <= not(layer4_outputs(284));
    outputs(1255) <= layer4_outputs(2419);
    outputs(1256) <= (layer4_outputs(447)) and (layer4_outputs(1248));
    outputs(1257) <= (layer4_outputs(1844)) and not (layer4_outputs(2548));
    outputs(1258) <= not((layer4_outputs(561)) or (layer4_outputs(1662)));
    outputs(1259) <= (layer4_outputs(195)) and not (layer4_outputs(311));
    outputs(1260) <= (layer4_outputs(229)) xor (layer4_outputs(1795));
    outputs(1261) <= layer4_outputs(1549);
    outputs(1262) <= not(layer4_outputs(2234));
    outputs(1263) <= not(layer4_outputs(743));
    outputs(1264) <= not(layer4_outputs(7));
    outputs(1265) <= not(layer4_outputs(551));
    outputs(1266) <= layer4_outputs(2162);
    outputs(1267) <= not(layer4_outputs(1401));
    outputs(1268) <= layer4_outputs(751);
    outputs(1269) <= layer4_outputs(344);
    outputs(1270) <= layer4_outputs(2175);
    outputs(1271) <= not(layer4_outputs(967));
    outputs(1272) <= not(layer4_outputs(30));
    outputs(1273) <= not(layer4_outputs(2307));
    outputs(1274) <= (layer4_outputs(525)) and not (layer4_outputs(2281));
    outputs(1275) <= not(layer4_outputs(1098));
    outputs(1276) <= layer4_outputs(638);
    outputs(1277) <= (layer4_outputs(2049)) and not (layer4_outputs(311));
    outputs(1278) <= not((layer4_outputs(2193)) xor (layer4_outputs(758)));
    outputs(1279) <= not(layer4_outputs(1110)) or (layer4_outputs(2326));
    outputs(1280) <= layer4_outputs(1857);
    outputs(1281) <= (layer4_outputs(555)) and (layer4_outputs(1438));
    outputs(1282) <= not(layer4_outputs(240));
    outputs(1283) <= not(layer4_outputs(124));
    outputs(1284) <= not((layer4_outputs(1506)) or (layer4_outputs(1891)));
    outputs(1285) <= layer4_outputs(2225);
    outputs(1286) <= (layer4_outputs(807)) xor (layer4_outputs(976));
    outputs(1287) <= not(layer4_outputs(1659));
    outputs(1288) <= not(layer4_outputs(2155));
    outputs(1289) <= (layer4_outputs(1300)) xor (layer4_outputs(947));
    outputs(1290) <= (layer4_outputs(939)) xor (layer4_outputs(1945));
    outputs(1291) <= not(layer4_outputs(1356));
    outputs(1292) <= layer4_outputs(2052);
    outputs(1293) <= layer4_outputs(2488);
    outputs(1294) <= layer4_outputs(1099);
    outputs(1295) <= not((layer4_outputs(1005)) xor (layer4_outputs(2150)));
    outputs(1296) <= layer4_outputs(197);
    outputs(1297) <= layer4_outputs(1621);
    outputs(1298) <= layer4_outputs(1299);
    outputs(1299) <= (layer4_outputs(1332)) or (layer4_outputs(776));
    outputs(1300) <= layer4_outputs(1759);
    outputs(1301) <= (layer4_outputs(1887)) and not (layer4_outputs(12));
    outputs(1302) <= (layer4_outputs(1048)) and not (layer4_outputs(1068));
    outputs(1303) <= layer4_outputs(2118);
    outputs(1304) <= not((layer4_outputs(1298)) xor (layer4_outputs(2079)));
    outputs(1305) <= layer4_outputs(1808);
    outputs(1306) <= not((layer4_outputs(1224)) or (layer4_outputs(819)));
    outputs(1307) <= (layer4_outputs(893)) xor (layer4_outputs(737));
    outputs(1308) <= (layer4_outputs(1928)) xor (layer4_outputs(1820));
    outputs(1309) <= not(layer4_outputs(1917));
    outputs(1310) <= layer4_outputs(1552);
    outputs(1311) <= layer4_outputs(1204);
    outputs(1312) <= not(layer4_outputs(1276));
    outputs(1313) <= (layer4_outputs(1085)) and not (layer4_outputs(1358));
    outputs(1314) <= layer4_outputs(157);
    outputs(1315) <= not(layer4_outputs(2002));
    outputs(1316) <= layer4_outputs(1581);
    outputs(1317) <= not(layer4_outputs(1619));
    outputs(1318) <= not(layer4_outputs(2513));
    outputs(1319) <= not(layer4_outputs(963));
    outputs(1320) <= not(layer4_outputs(2428)) or (layer4_outputs(1766));
    outputs(1321) <= layer4_outputs(1485);
    outputs(1322) <= not(layer4_outputs(1129));
    outputs(1323) <= not(layer4_outputs(1102));
    outputs(1324) <= not((layer4_outputs(2152)) and (layer4_outputs(2334)));
    outputs(1325) <= layer4_outputs(724);
    outputs(1326) <= not((layer4_outputs(1285)) or (layer4_outputs(703)));
    outputs(1327) <= not(layer4_outputs(2020));
    outputs(1328) <= (layer4_outputs(972)) and not (layer4_outputs(619));
    outputs(1329) <= not((layer4_outputs(1346)) or (layer4_outputs(1490)));
    outputs(1330) <= not(layer4_outputs(1516));
    outputs(1331) <= not(layer4_outputs(2482));
    outputs(1332) <= not(layer4_outputs(1388));
    outputs(1333) <= (layer4_outputs(783)) and not (layer4_outputs(2113));
    outputs(1334) <= not((layer4_outputs(1805)) xor (layer4_outputs(1743)));
    outputs(1335) <= not((layer4_outputs(1954)) or (layer4_outputs(1285)));
    outputs(1336) <= layer4_outputs(1638);
    outputs(1337) <= not(layer4_outputs(910));
    outputs(1338) <= (layer4_outputs(1454)) or (layer4_outputs(1671));
    outputs(1339) <= layer4_outputs(1489);
    outputs(1340) <= layer4_outputs(419);
    outputs(1341) <= not((layer4_outputs(2308)) xor (layer4_outputs(1178)));
    outputs(1342) <= not(layer4_outputs(1321));
    outputs(1343) <= (layer4_outputs(2087)) xor (layer4_outputs(2111));
    outputs(1344) <= not((layer4_outputs(2341)) xor (layer4_outputs(1349)));
    outputs(1345) <= not((layer4_outputs(2430)) xor (layer4_outputs(1186)));
    outputs(1346) <= layer4_outputs(1818);
    outputs(1347) <= not(layer4_outputs(2512));
    outputs(1348) <= layer4_outputs(1038);
    outputs(1349) <= (layer4_outputs(1411)) and not (layer4_outputs(230));
    outputs(1350) <= (layer4_outputs(2355)) xor (layer4_outputs(1333));
    outputs(1351) <= (layer4_outputs(2510)) xor (layer4_outputs(792));
    outputs(1352) <= not((layer4_outputs(629)) or (layer4_outputs(1273)));
    outputs(1353) <= not(layer4_outputs(962));
    outputs(1354) <= not(layer4_outputs(775));
    outputs(1355) <= not(layer4_outputs(2404));
    outputs(1356) <= layer4_outputs(752);
    outputs(1357) <= (layer4_outputs(423)) and (layer4_outputs(2048));
    outputs(1358) <= not((layer4_outputs(2037)) or (layer4_outputs(1649)));
    outputs(1359) <= not(layer4_outputs(1150));
    outputs(1360) <= layer4_outputs(1404);
    outputs(1361) <= not((layer4_outputs(1508)) xor (layer4_outputs(1000)));
    outputs(1362) <= not(layer4_outputs(129)) or (layer4_outputs(1227));
    outputs(1363) <= not(layer4_outputs(295));
    outputs(1364) <= (layer4_outputs(2462)) or (layer4_outputs(1137));
    outputs(1365) <= layer4_outputs(1449);
    outputs(1366) <= (layer4_outputs(1002)) xor (layer4_outputs(1241));
    outputs(1367) <= not(layer4_outputs(1044));
    outputs(1368) <= not((layer4_outputs(2339)) or (layer4_outputs(1448)));
    outputs(1369) <= layer4_outputs(2398);
    outputs(1370) <= not(layer4_outputs(2202));
    outputs(1371) <= not((layer4_outputs(1731)) or (layer4_outputs(1468)));
    outputs(1372) <= not((layer4_outputs(149)) or (layer4_outputs(2519)));
    outputs(1373) <= layer4_outputs(1328);
    outputs(1374) <= layer4_outputs(1015);
    outputs(1375) <= (layer4_outputs(2065)) and not (layer4_outputs(333));
    outputs(1376) <= layer4_outputs(561);
    outputs(1377) <= layer4_outputs(2051);
    outputs(1378) <= not((layer4_outputs(1004)) or (layer4_outputs(1617)));
    outputs(1379) <= not(layer4_outputs(2187));
    outputs(1380) <= not((layer4_outputs(1792)) or (layer4_outputs(2210)));
    outputs(1381) <= not(layer4_outputs(2459));
    outputs(1382) <= layer4_outputs(2144);
    outputs(1383) <= not(layer4_outputs(2010));
    outputs(1384) <= not(layer4_outputs(482));
    outputs(1385) <= not(layer4_outputs(1197));
    outputs(1386) <= layer4_outputs(1818);
    outputs(1387) <= not(layer4_outputs(2357));
    outputs(1388) <= (layer4_outputs(646)) and not (layer4_outputs(2400));
    outputs(1389) <= layer4_outputs(2387);
    outputs(1390) <= not(layer4_outputs(456)) or (layer4_outputs(199));
    outputs(1391) <= (layer4_outputs(1054)) and not (layer4_outputs(2372));
    outputs(1392) <= not((layer4_outputs(1875)) xor (layer4_outputs(906)));
    outputs(1393) <= not(layer4_outputs(963));
    outputs(1394) <= (layer4_outputs(0)) xor (layer4_outputs(2277));
    outputs(1395) <= not(layer4_outputs(504));
    outputs(1396) <= not(layer4_outputs(1453));
    outputs(1397) <= not(layer4_outputs(395));
    outputs(1398) <= layer4_outputs(320);
    outputs(1399) <= layer4_outputs(2219);
    outputs(1400) <= not(layer4_outputs(2297));
    outputs(1401) <= not((layer4_outputs(191)) or (layer4_outputs(1789)));
    outputs(1402) <= not((layer4_outputs(1646)) xor (layer4_outputs(898)));
    outputs(1403) <= not(layer4_outputs(1083));
    outputs(1404) <= layer4_outputs(2171);
    outputs(1405) <= (layer4_outputs(700)) and not (layer4_outputs(1526));
    outputs(1406) <= not((layer4_outputs(1775)) or (layer4_outputs(1290)));
    outputs(1407) <= not(layer4_outputs(2106));
    outputs(1408) <= not(layer4_outputs(2197));
    outputs(1409) <= layer4_outputs(653);
    outputs(1410) <= not(layer4_outputs(735));
    outputs(1411) <= not(layer4_outputs(2316));
    outputs(1412) <= layer4_outputs(1050);
    outputs(1413) <= layer4_outputs(2369);
    outputs(1414) <= not(layer4_outputs(2471));
    outputs(1415) <= layer4_outputs(427);
    outputs(1416) <= (layer4_outputs(47)) and not (layer4_outputs(878));
    outputs(1417) <= not(layer4_outputs(662));
    outputs(1418) <= not(layer4_outputs(2174));
    outputs(1419) <= not(layer4_outputs(2098));
    outputs(1420) <= layer4_outputs(1407);
    outputs(1421) <= not(layer4_outputs(2227));
    outputs(1422) <= layer4_outputs(1421);
    outputs(1423) <= (layer4_outputs(914)) and (layer4_outputs(1695));
    outputs(1424) <= not(layer4_outputs(52));
    outputs(1425) <= not(layer4_outputs(499));
    outputs(1426) <= not(layer4_outputs(1014));
    outputs(1427) <= (layer4_outputs(1613)) and not (layer4_outputs(1565));
    outputs(1428) <= not((layer4_outputs(857)) xor (layer4_outputs(405)));
    outputs(1429) <= not(layer4_outputs(1104));
    outputs(1430) <= not(layer4_outputs(572));
    outputs(1431) <= not(layer4_outputs(2128));
    outputs(1432) <= not(layer4_outputs(1451));
    outputs(1433) <= layer4_outputs(349);
    outputs(1434) <= layer4_outputs(811);
    outputs(1435) <= (layer4_outputs(1644)) or (layer4_outputs(175));
    outputs(1436) <= not((layer4_outputs(1149)) xor (layer4_outputs(1597)));
    outputs(1437) <= (layer4_outputs(629)) xor (layer4_outputs(45));
    outputs(1438) <= (layer4_outputs(1858)) xor (layer4_outputs(1628));
    outputs(1439) <= layer4_outputs(1864);
    outputs(1440) <= not(layer4_outputs(2002));
    outputs(1441) <= (layer4_outputs(2407)) xor (layer4_outputs(322));
    outputs(1442) <= not(layer4_outputs(1606));
    outputs(1443) <= layer4_outputs(2008);
    outputs(1444) <= layer4_outputs(710);
    outputs(1445) <= not(layer4_outputs(2436));
    outputs(1446) <= layer4_outputs(1767);
    outputs(1447) <= layer4_outputs(1732);
    outputs(1448) <= (layer4_outputs(131)) and not (layer4_outputs(1860));
    outputs(1449) <= (layer4_outputs(1255)) xor (layer4_outputs(59));
    outputs(1450) <= not(layer4_outputs(824)) or (layer4_outputs(1459));
    outputs(1451) <= not(layer4_outputs(879));
    outputs(1452) <= layer4_outputs(466);
    outputs(1453) <= layer4_outputs(1598);
    outputs(1454) <= layer4_outputs(1029);
    outputs(1455) <= (layer4_outputs(1921)) and (layer4_outputs(2479));
    outputs(1456) <= not((layer4_outputs(1923)) or (layer4_outputs(1702)));
    outputs(1457) <= not((layer4_outputs(1775)) and (layer4_outputs(532)));
    outputs(1458) <= not(layer4_outputs(1123));
    outputs(1459) <= layer4_outputs(1951);
    outputs(1460) <= not((layer4_outputs(2331)) xor (layer4_outputs(2136)));
    outputs(1461) <= layer4_outputs(1095);
    outputs(1462) <= not(layer4_outputs(254));
    outputs(1463) <= (layer4_outputs(1885)) xor (layer4_outputs(2164));
    outputs(1464) <= layer4_outputs(1848);
    outputs(1465) <= not(layer4_outputs(2321));
    outputs(1466) <= not(layer4_outputs(85));
    outputs(1467) <= not((layer4_outputs(255)) or (layer4_outputs(193)));
    outputs(1468) <= layer4_outputs(2237);
    outputs(1469) <= not(layer4_outputs(222));
    outputs(1470) <= not(layer4_outputs(1158));
    outputs(1471) <= not((layer4_outputs(481)) or (layer4_outputs(1783)));
    outputs(1472) <= not((layer4_outputs(1117)) xor (layer4_outputs(451)));
    outputs(1473) <= layer4_outputs(1074);
    outputs(1474) <= (layer4_outputs(765)) and (layer4_outputs(1972));
    outputs(1475) <= (layer4_outputs(1722)) xor (layer4_outputs(731));
    outputs(1476) <= layer4_outputs(2228);
    outputs(1477) <= not((layer4_outputs(507)) xor (layer4_outputs(2435)));
    outputs(1478) <= (layer4_outputs(1179)) and not (layer4_outputs(2550));
    outputs(1479) <= (layer4_outputs(812)) xor (layer4_outputs(1943));
    outputs(1480) <= layer4_outputs(1857);
    outputs(1481) <= not(layer4_outputs(959));
    outputs(1482) <= (layer4_outputs(117)) and not (layer4_outputs(542));
    outputs(1483) <= not(layer4_outputs(800));
    outputs(1484) <= not((layer4_outputs(1199)) and (layer4_outputs(1627)));
    outputs(1485) <= (layer4_outputs(1635)) and not (layer4_outputs(2547));
    outputs(1486) <= not(layer4_outputs(2266));
    outputs(1487) <= not(layer4_outputs(1533)) or (layer4_outputs(2397));
    outputs(1488) <= layer4_outputs(1523);
    outputs(1489) <= layer4_outputs(1221);
    outputs(1490) <= (layer4_outputs(2093)) xor (layer4_outputs(1823));
    outputs(1491) <= (layer4_outputs(2420)) and not (layer4_outputs(635));
    outputs(1492) <= not(layer4_outputs(1991));
    outputs(1493) <= not(layer4_outputs(1189)) or (layer4_outputs(844));
    outputs(1494) <= (layer4_outputs(5)) xor (layer4_outputs(1130));
    outputs(1495) <= layer4_outputs(1564);
    outputs(1496) <= not(layer4_outputs(62)) or (layer4_outputs(550));
    outputs(1497) <= not(layer4_outputs(1578));
    outputs(1498) <= layer4_outputs(2277);
    outputs(1499) <= not(layer4_outputs(879));
    outputs(1500) <= not(layer4_outputs(740));
    outputs(1501) <= layer4_outputs(2425);
    outputs(1502) <= (layer4_outputs(2094)) xor (layer4_outputs(1002));
    outputs(1503) <= not(layer4_outputs(795));
    outputs(1504) <= layer4_outputs(647);
    outputs(1505) <= not(layer4_outputs(1278));
    outputs(1506) <= not(layer4_outputs(1944));
    outputs(1507) <= not((layer4_outputs(1385)) or (layer4_outputs(147)));
    outputs(1508) <= layer4_outputs(2052);
    outputs(1509) <= not((layer4_outputs(361)) or (layer4_outputs(1366)));
    outputs(1510) <= layer4_outputs(2324);
    outputs(1511) <= layer4_outputs(247);
    outputs(1512) <= not(layer4_outputs(2014));
    outputs(1513) <= (layer4_outputs(2229)) and not (layer4_outputs(2280));
    outputs(1514) <= (layer4_outputs(613)) and not (layer4_outputs(1018));
    outputs(1515) <= not(layer4_outputs(19));
    outputs(1516) <= not(layer4_outputs(1087));
    outputs(1517) <= (layer4_outputs(370)) and not (layer4_outputs(2375));
    outputs(1518) <= (layer4_outputs(1656)) xor (layer4_outputs(2317));
    outputs(1519) <= layer4_outputs(1978);
    outputs(1520) <= layer4_outputs(2271);
    outputs(1521) <= not(layer4_outputs(240));
    outputs(1522) <= not(layer4_outputs(368));
    outputs(1523) <= not(layer4_outputs(188));
    outputs(1524) <= layer4_outputs(2397);
    outputs(1525) <= not(layer4_outputs(2411));
    outputs(1526) <= not((layer4_outputs(1365)) xor (layer4_outputs(1672)));
    outputs(1527) <= not(layer4_outputs(993));
    outputs(1528) <= layer4_outputs(726);
    outputs(1529) <= (layer4_outputs(1631)) xor (layer4_outputs(695));
    outputs(1530) <= (layer4_outputs(1420)) xor (layer4_outputs(2265));
    outputs(1531) <= layer4_outputs(50);
    outputs(1532) <= layer4_outputs(2461);
    outputs(1533) <= layer4_outputs(567);
    outputs(1534) <= not((layer4_outputs(1106)) xor (layer4_outputs(1822)));
    outputs(1535) <= layer4_outputs(2215);
    outputs(1536) <= (layer4_outputs(2077)) or (layer4_outputs(2541));
    outputs(1537) <= (layer4_outputs(2022)) xor (layer4_outputs(1667));
    outputs(1538) <= (layer4_outputs(1619)) and not (layer4_outputs(2508));
    outputs(1539) <= not(layer4_outputs(2220));
    outputs(1540) <= layer4_outputs(2217);
    outputs(1541) <= not(layer4_outputs(385));
    outputs(1542) <= not(layer4_outputs(2092));
    outputs(1543) <= layer4_outputs(1301);
    outputs(1544) <= (layer4_outputs(357)) xor (layer4_outputs(1495));
    outputs(1545) <= not(layer4_outputs(1753));
    outputs(1546) <= not(layer4_outputs(2161));
    outputs(1547) <= layer4_outputs(2444);
    outputs(1548) <= layer4_outputs(88);
    outputs(1549) <= layer4_outputs(736);
    outputs(1550) <= layer4_outputs(1705);
    outputs(1551) <= not((layer4_outputs(1968)) and (layer4_outputs(591)));
    outputs(1552) <= (layer4_outputs(2144)) and (layer4_outputs(692));
    outputs(1553) <= layer4_outputs(1725);
    outputs(1554) <= layer4_outputs(2378);
    outputs(1555) <= not(layer4_outputs(4));
    outputs(1556) <= not((layer4_outputs(144)) or (layer4_outputs(836)));
    outputs(1557) <= not(layer4_outputs(1079));
    outputs(1558) <= (layer4_outputs(120)) and not (layer4_outputs(1423));
    outputs(1559) <= not(layer4_outputs(2025));
    outputs(1560) <= (layer4_outputs(670)) xor (layer4_outputs(1000));
    outputs(1561) <= not(layer4_outputs(2178));
    outputs(1562) <= not(layer4_outputs(1637));
    outputs(1563) <= not((layer4_outputs(1071)) xor (layer4_outputs(503)));
    outputs(1564) <= (layer4_outputs(1284)) and not (layer4_outputs(1252));
    outputs(1565) <= (layer4_outputs(453)) and not (layer4_outputs(1371));
    outputs(1566) <= layer4_outputs(2093);
    outputs(1567) <= not(layer4_outputs(198));
    outputs(1568) <= not(layer4_outputs(1810));
    outputs(1569) <= not(layer4_outputs(2367));
    outputs(1570) <= not(layer4_outputs(2121));
    outputs(1571) <= not(layer4_outputs(1793));
    outputs(1572) <= layer4_outputs(340);
    outputs(1573) <= (layer4_outputs(1185)) xor (layer4_outputs(2100));
    outputs(1574) <= layer4_outputs(2214);
    outputs(1575) <= (layer4_outputs(889)) xor (layer4_outputs(618));
    outputs(1576) <= layer4_outputs(2111);
    outputs(1577) <= (layer4_outputs(2542)) and not (layer4_outputs(2463));
    outputs(1578) <= not(layer4_outputs(927));
    outputs(1579) <= (layer4_outputs(42)) xor (layer4_outputs(1351));
    outputs(1580) <= layer4_outputs(1835);
    outputs(1581) <= not(layer4_outputs(112));
    outputs(1582) <= not(layer4_outputs(2046));
    outputs(1583) <= layer4_outputs(718);
    outputs(1584) <= not(layer4_outputs(2226));
    outputs(1585) <= not(layer4_outputs(185));
    outputs(1586) <= (layer4_outputs(138)) xor (layer4_outputs(763));
    outputs(1587) <= not(layer4_outputs(1007));
    outputs(1588) <= not(layer4_outputs(1863));
    outputs(1589) <= not(layer4_outputs(2126));
    outputs(1590) <= not(layer4_outputs(2362));
    outputs(1591) <= not(layer4_outputs(2362));
    outputs(1592) <= layer4_outputs(485);
    outputs(1593) <= not(layer4_outputs(1953));
    outputs(1594) <= layer4_outputs(442);
    outputs(1595) <= layer4_outputs(1560);
    outputs(1596) <= layer4_outputs(2085);
    outputs(1597) <= layer4_outputs(1828);
    outputs(1598) <= (layer4_outputs(599)) or (layer4_outputs(712));
    outputs(1599) <= (layer4_outputs(1076)) and not (layer4_outputs(2553));
    outputs(1600) <= not(layer4_outputs(410));
    outputs(1601) <= layer4_outputs(2030);
    outputs(1602) <= not(layer4_outputs(1451));
    outputs(1603) <= (layer4_outputs(2042)) xor (layer4_outputs(651));
    outputs(1604) <= layer4_outputs(898);
    outputs(1605) <= layer4_outputs(634);
    outputs(1606) <= not(layer4_outputs(1230)) or (layer4_outputs(399));
    outputs(1607) <= layer4_outputs(880);
    outputs(1608) <= layer4_outputs(1895);
    outputs(1609) <= layer4_outputs(652);
    outputs(1610) <= layer4_outputs(1140);
    outputs(1611) <= layer4_outputs(2520);
    outputs(1612) <= (layer4_outputs(313)) or (layer4_outputs(576));
    outputs(1613) <= layer4_outputs(1542);
    outputs(1614) <= not(layer4_outputs(706));
    outputs(1615) <= not((layer4_outputs(1337)) or (layer4_outputs(1550)));
    outputs(1616) <= (layer4_outputs(2455)) and not (layer4_outputs(39));
    outputs(1617) <= layer4_outputs(36);
    outputs(1618) <= not(layer4_outputs(1660));
    outputs(1619) <= not(layer4_outputs(569));
    outputs(1620) <= not(layer4_outputs(1599));
    outputs(1621) <= not(layer4_outputs(725));
    outputs(1622) <= layer4_outputs(2125);
    outputs(1623) <= (layer4_outputs(1223)) and not (layer4_outputs(771));
    outputs(1624) <= (layer4_outputs(2272)) and not (layer4_outputs(481));
    outputs(1625) <= (layer4_outputs(450)) and (layer4_outputs(1719));
    outputs(1626) <= (layer4_outputs(44)) xor (layer4_outputs(490));
    outputs(1627) <= layer4_outputs(178);
    outputs(1628) <= not((layer4_outputs(1357)) or (layer4_outputs(761)));
    outputs(1629) <= layer4_outputs(2274);
    outputs(1630) <= (layer4_outputs(1172)) and not (layer4_outputs(993));
    outputs(1631) <= not((layer4_outputs(1169)) or (layer4_outputs(2447)));
    outputs(1632) <= layer4_outputs(1377);
    outputs(1633) <= (layer4_outputs(790)) and (layer4_outputs(1508));
    outputs(1634) <= layer4_outputs(506);
    outputs(1635) <= (layer4_outputs(150)) xor (layer4_outputs(1683));
    outputs(1636) <= layer4_outputs(233);
    outputs(1637) <= layer4_outputs(1972);
    outputs(1638) <= (layer4_outputs(2505)) or (layer4_outputs(1325));
    outputs(1639) <= not((layer4_outputs(895)) and (layer4_outputs(2457)));
    outputs(1640) <= not((layer4_outputs(1586)) or (layer4_outputs(2275)));
    outputs(1641) <= not(layer4_outputs(1756)) or (layer4_outputs(2443));
    outputs(1642) <= layer4_outputs(188);
    outputs(1643) <= not(layer4_outputs(1572));
    outputs(1644) <= layer4_outputs(2435);
    outputs(1645) <= not((layer4_outputs(1092)) or (layer4_outputs(334)));
    outputs(1646) <= (layer4_outputs(771)) xor (layer4_outputs(1827));
    outputs(1647) <= not(layer4_outputs(732));
    outputs(1648) <= not(layer4_outputs(2537)) or (layer4_outputs(2484));
    outputs(1649) <= not(layer4_outputs(2380));
    outputs(1650) <= layer4_outputs(1996);
    outputs(1651) <= (layer4_outputs(673)) and (layer4_outputs(273));
    outputs(1652) <= (layer4_outputs(350)) and (layer4_outputs(1803));
    outputs(1653) <= not((layer4_outputs(941)) or (layer4_outputs(922)));
    outputs(1654) <= layer4_outputs(1976);
    outputs(1655) <= (layer4_outputs(2392)) or (layer4_outputs(80));
    outputs(1656) <= not((layer4_outputs(1728)) or (layer4_outputs(564)));
    outputs(1657) <= layer4_outputs(827);
    outputs(1658) <= not(layer4_outputs(1012));
    outputs(1659) <= layer4_outputs(1445);
    outputs(1660) <= not((layer4_outputs(1288)) xor (layer4_outputs(1780)));
    outputs(1661) <= not(layer4_outputs(2132));
    outputs(1662) <= not((layer4_outputs(451)) xor (layer4_outputs(2242)));
    outputs(1663) <= not(layer4_outputs(657));
    outputs(1664) <= not(layer4_outputs(1906));
    outputs(1665) <= not(layer4_outputs(605));
    outputs(1666) <= layer4_outputs(1428);
    outputs(1667) <= layer4_outputs(2477);
    outputs(1668) <= not(layer4_outputs(2473));
    outputs(1669) <= layer4_outputs(891);
    outputs(1670) <= not(layer4_outputs(932));
    outputs(1671) <= not(layer4_outputs(2468));
    outputs(1672) <= (layer4_outputs(1527)) xor (layer4_outputs(1259));
    outputs(1673) <= (layer4_outputs(1642)) and not (layer4_outputs(1364));
    outputs(1674) <= layer4_outputs(1918);
    outputs(1675) <= layer4_outputs(127);
    outputs(1676) <= layer4_outputs(2506);
    outputs(1677) <= not(layer4_outputs(2116));
    outputs(1678) <= layer4_outputs(784);
    outputs(1679) <= not(layer4_outputs(2273));
    outputs(1680) <= layer4_outputs(870);
    outputs(1681) <= not(layer4_outputs(467));
    outputs(1682) <= not(layer4_outputs(1840));
    outputs(1683) <= layer4_outputs(1531);
    outputs(1684) <= not((layer4_outputs(1831)) or (layer4_outputs(73)));
    outputs(1685) <= layer4_outputs(793);
    outputs(1686) <= not(layer4_outputs(721));
    outputs(1687) <= not(layer4_outputs(1907)) or (layer4_outputs(1583));
    outputs(1688) <= layer4_outputs(1260);
    outputs(1689) <= not(layer4_outputs(960)) or (layer4_outputs(1882));
    outputs(1690) <= (layer4_outputs(2407)) xor (layer4_outputs(734));
    outputs(1691) <= (layer4_outputs(728)) and (layer4_outputs(196));
    outputs(1692) <= layer4_outputs(9);
    outputs(1693) <= not(layer4_outputs(595));
    outputs(1694) <= (layer4_outputs(2485)) and (layer4_outputs(1146));
    outputs(1695) <= not(layer4_outputs(1341));
    outputs(1696) <= (layer4_outputs(2009)) and not (layer4_outputs(430));
    outputs(1697) <= layer4_outputs(1399);
    outputs(1698) <= not((layer4_outputs(2409)) or (layer4_outputs(1296)));
    outputs(1699) <= not(layer4_outputs(1611));
    outputs(1700) <= layer4_outputs(1638);
    outputs(1701) <= not(layer4_outputs(2409)) or (layer4_outputs(2326));
    outputs(1702) <= not((layer4_outputs(908)) xor (layer4_outputs(2559)));
    outputs(1703) <= not(layer4_outputs(1707));
    outputs(1704) <= layer4_outputs(2366);
    outputs(1705) <= not(layer4_outputs(628));
    outputs(1706) <= not(layer4_outputs(161));
    outputs(1707) <= not((layer4_outputs(1509)) xor (layer4_outputs(1394)));
    outputs(1708) <= not(layer4_outputs(230));
    outputs(1709) <= (layer4_outputs(820)) and (layer4_outputs(2461));
    outputs(1710) <= not(layer4_outputs(1316));
    outputs(1711) <= not(layer4_outputs(1966));
    outputs(1712) <= not(layer4_outputs(2017));
    outputs(1713) <= (layer4_outputs(714)) and not (layer4_outputs(975));
    outputs(1714) <= (layer4_outputs(115)) xor (layer4_outputs(108));
    outputs(1715) <= (layer4_outputs(1186)) and not (layer4_outputs(1105));
    outputs(1716) <= not(layer4_outputs(171));
    outputs(1717) <= not(layer4_outputs(915));
    outputs(1718) <= (layer4_outputs(1282)) xor (layer4_outputs(1977));
    outputs(1719) <= (layer4_outputs(1801)) and not (layer4_outputs(1190));
    outputs(1720) <= not((layer4_outputs(855)) or (layer4_outputs(1802)));
    outputs(1721) <= (layer4_outputs(2396)) and not (layer4_outputs(1197));
    outputs(1722) <= (layer4_outputs(2134)) and not (layer4_outputs(657));
    outputs(1723) <= not(layer4_outputs(2161));
    outputs(1724) <= layer4_outputs(967);
    outputs(1725) <= layer4_outputs(687);
    outputs(1726) <= layer4_outputs(2075);
    outputs(1727) <= layer4_outputs(1048);
    outputs(1728) <= not(layer4_outputs(1341));
    outputs(1729) <= layer4_outputs(1024);
    outputs(1730) <= layer4_outputs(2210);
    outputs(1731) <= layer4_outputs(2100);
    outputs(1732) <= (layer4_outputs(1054)) and not (layer4_outputs(1887));
    outputs(1733) <= not(layer4_outputs(293));
    outputs(1734) <= (layer4_outputs(127)) and not (layer4_outputs(1264));
    outputs(1735) <= not((layer4_outputs(1968)) or (layer4_outputs(1168)));
    outputs(1736) <= not(layer4_outputs(2263));
    outputs(1737) <= (layer4_outputs(926)) and (layer4_outputs(1515));
    outputs(1738) <= not(layer4_outputs(2329));
    outputs(1739) <= layer4_outputs(538);
    outputs(1740) <= not(layer4_outputs(2289));
    outputs(1741) <= layer4_outputs(2272);
    outputs(1742) <= (layer4_outputs(2520)) xor (layer4_outputs(363));
    outputs(1743) <= not((layer4_outputs(1963)) xor (layer4_outputs(305)));
    outputs(1744) <= layer4_outputs(450);
    outputs(1745) <= not(layer4_outputs(1190));
    outputs(1746) <= layer4_outputs(475);
    outputs(1747) <= not(layer4_outputs(691));
    outputs(1748) <= (layer4_outputs(332)) and (layer4_outputs(2133));
    outputs(1749) <= (layer4_outputs(359)) and not (layer4_outputs(1358));
    outputs(1750) <= not((layer4_outputs(2247)) xor (layer4_outputs(912)));
    outputs(1751) <= not((layer4_outputs(1640)) or (layer4_outputs(342)));
    outputs(1752) <= not(layer4_outputs(770));
    outputs(1753) <= not(layer4_outputs(849));
    outputs(1754) <= not(layer4_outputs(1348));
    outputs(1755) <= (layer4_outputs(1925)) xor (layer4_outputs(2207));
    outputs(1756) <= (layer4_outputs(459)) xor (layer4_outputs(1827));
    outputs(1757) <= not(layer4_outputs(1293));
    outputs(1758) <= layer4_outputs(1926);
    outputs(1759) <= layer4_outputs(1139);
    outputs(1760) <= layer4_outputs(2234);
    outputs(1761) <= not((layer4_outputs(2449)) xor (layer4_outputs(94)));
    outputs(1762) <= (layer4_outputs(375)) and not (layer4_outputs(1039));
    outputs(1763) <= layer4_outputs(1404);
    outputs(1764) <= layer4_outputs(2433);
    outputs(1765) <= not(layer4_outputs(1723)) or (layer4_outputs(644));
    outputs(1766) <= not((layer4_outputs(2426)) or (layer4_outputs(2329)));
    outputs(1767) <= layer4_outputs(1734);
    outputs(1768) <= not(layer4_outputs(65));
    outputs(1769) <= not(layer4_outputs(87));
    outputs(1770) <= not(layer4_outputs(1296));
    outputs(1771) <= not(layer4_outputs(737));
    outputs(1772) <= not(layer4_outputs(2003));
    outputs(1773) <= not(layer4_outputs(2031));
    outputs(1774) <= not((layer4_outputs(1839)) or (layer4_outputs(2489)));
    outputs(1775) <= layer4_outputs(624);
    outputs(1776) <= (layer4_outputs(2490)) and not (layer4_outputs(1265));
    outputs(1777) <= layer4_outputs(580);
    outputs(1778) <= layer4_outputs(11);
    outputs(1779) <= not(layer4_outputs(457));
    outputs(1780) <= not(layer4_outputs(405));
    outputs(1781) <= not((layer4_outputs(293)) or (layer4_outputs(2535)));
    outputs(1782) <= (layer4_outputs(148)) and not (layer4_outputs(1575));
    outputs(1783) <= layer4_outputs(1542);
    outputs(1784) <= layer4_outputs(1725);
    outputs(1785) <= not(layer4_outputs(16));
    outputs(1786) <= not(layer4_outputs(1493));
    outputs(1787) <= (layer4_outputs(1860)) or (layer4_outputs(2372));
    outputs(1788) <= not(layer4_outputs(1059));
    outputs(1789) <= not(layer4_outputs(171)) or (layer4_outputs(268));
    outputs(1790) <= not(layer4_outputs(1678));
    outputs(1791) <= not(layer4_outputs(1225));
    outputs(1792) <= (layer4_outputs(1834)) and not (layer4_outputs(288));
    outputs(1793) <= (layer4_outputs(1547)) and (layer4_outputs(1204));
    outputs(1794) <= layer4_outputs(1806);
    outputs(1795) <= not((layer4_outputs(886)) xor (layer4_outputs(669)));
    outputs(1796) <= not(layer4_outputs(1704));
    outputs(1797) <= layer4_outputs(2493);
    outputs(1798) <= not(layer4_outputs(2345)) or (layer4_outputs(2066));
    outputs(1799) <= not(layer4_outputs(539));
    outputs(1800) <= not((layer4_outputs(12)) xor (layer4_outputs(2138)));
    outputs(1801) <= layer4_outputs(452);
    outputs(1802) <= layer4_outputs(102);
    outputs(1803) <= not(layer4_outputs(267));
    outputs(1804) <= not(layer4_outputs(1184));
    outputs(1805) <= layer4_outputs(64);
    outputs(1806) <= not(layer4_outputs(1060));
    outputs(1807) <= not(layer4_outputs(252)) or (layer4_outputs(286));
    outputs(1808) <= (layer4_outputs(1851)) xor (layer4_outputs(660));
    outputs(1809) <= not((layer4_outputs(186)) or (layer4_outputs(413)));
    outputs(1810) <= layer4_outputs(1234);
    outputs(1811) <= (layer4_outputs(189)) and not (layer4_outputs(823));
    outputs(1812) <= not((layer4_outputs(1752)) or (layer4_outputs(359)));
    outputs(1813) <= not((layer4_outputs(549)) xor (layer4_outputs(810)));
    outputs(1814) <= (layer4_outputs(933)) and not (layer4_outputs(475));
    outputs(1815) <= not((layer4_outputs(1304)) or (layer4_outputs(2089)));
    outputs(1816) <= not((layer4_outputs(324)) or (layer4_outputs(679)));
    outputs(1817) <= layer4_outputs(1108);
    outputs(1818) <= layer4_outputs(175);
    outputs(1819) <= not(layer4_outputs(284));
    outputs(1820) <= not(layer4_outputs(1997));
    outputs(1821) <= not((layer4_outputs(1101)) or (layer4_outputs(2506)));
    outputs(1822) <= not(layer4_outputs(116));
    outputs(1823) <= layer4_outputs(1874);
    outputs(1824) <= layer4_outputs(997);
    outputs(1825) <= not(layer4_outputs(2074)) or (layer4_outputs(1758));
    outputs(1826) <= not(layer4_outputs(2338));
    outputs(1827) <= not(layer4_outputs(2544));
    outputs(1828) <= not(layer4_outputs(541)) or (layer4_outputs(1383));
    outputs(1829) <= not((layer4_outputs(2095)) xor (layer4_outputs(1352)));
    outputs(1830) <= layer4_outputs(1263);
    outputs(1831) <= not(layer4_outputs(1804));
    outputs(1832) <= not(layer4_outputs(105));
    outputs(1833) <= (layer4_outputs(1035)) and not (layer4_outputs(89));
    outputs(1834) <= layer4_outputs(1349);
    outputs(1835) <= layer4_outputs(1461);
    outputs(1836) <= not(layer4_outputs(2079));
    outputs(1837) <= layer4_outputs(2190);
    outputs(1838) <= not(layer4_outputs(1595));
    outputs(1839) <= not(layer4_outputs(408));
    outputs(1840) <= not(layer4_outputs(6));
    outputs(1841) <= layer4_outputs(1524);
    outputs(1842) <= not(layer4_outputs(1075));
    outputs(1843) <= not((layer4_outputs(1116)) xor (layer4_outputs(2549)));
    outputs(1844) <= not(layer4_outputs(1727));
    outputs(1845) <= not((layer4_outputs(109)) or (layer4_outputs(677)));
    outputs(1846) <= not(layer4_outputs(501));
    outputs(1847) <= (layer4_outputs(2302)) and not (layer4_outputs(1532));
    outputs(1848) <= layer4_outputs(2301);
    outputs(1849) <= not(layer4_outputs(931));
    outputs(1850) <= not(layer4_outputs(1592));
    outputs(1851) <= layer4_outputs(2101);
    outputs(1852) <= not((layer4_outputs(833)) or (layer4_outputs(2546)));
    outputs(1853) <= layer4_outputs(1030);
    outputs(1854) <= layer4_outputs(566);
    outputs(1855) <= not((layer4_outputs(872)) or (layer4_outputs(1639)));
    outputs(1856) <= not(layer4_outputs(1713));
    outputs(1857) <= not(layer4_outputs(634));
    outputs(1858) <= not(layer4_outputs(1476));
    outputs(1859) <= (layer4_outputs(372)) and not (layer4_outputs(982));
    outputs(1860) <= not(layer4_outputs(1897));
    outputs(1861) <= not(layer4_outputs(526));
    outputs(1862) <= not(layer4_outputs(2349));
    outputs(1863) <= (layer4_outputs(1077)) and not (layer4_outputs(2235));
    outputs(1864) <= not(layer4_outputs(2221));
    outputs(1865) <= not((layer4_outputs(156)) xor (layer4_outputs(2389)));
    outputs(1866) <= (layer4_outputs(1046)) and not (layer4_outputs(768));
    outputs(1867) <= not(layer4_outputs(2327)) or (layer4_outputs(1217));
    outputs(1868) <= layer4_outputs(1374);
    outputs(1869) <= not(layer4_outputs(1785));
    outputs(1870) <= layer4_outputs(829);
    outputs(1871) <= not(layer4_outputs(597));
    outputs(1872) <= layer4_outputs(1669);
    outputs(1873) <= (layer4_outputs(610)) and not (layer4_outputs(103));
    outputs(1874) <= (layer4_outputs(2486)) xor (layer4_outputs(1558));
    outputs(1875) <= layer4_outputs(2146);
    outputs(1876) <= not((layer4_outputs(548)) or (layer4_outputs(2154)));
    outputs(1877) <= layer4_outputs(1883);
    outputs(1878) <= layer4_outputs(2259);
    outputs(1879) <= (layer4_outputs(123)) and (layer4_outputs(421));
    outputs(1880) <= not(layer4_outputs(699));
    outputs(1881) <= layer4_outputs(607);
    outputs(1882) <= (layer4_outputs(326)) and not (layer4_outputs(105));
    outputs(1883) <= not(layer4_outputs(1956));
    outputs(1884) <= not(layer4_outputs(10));
    outputs(1885) <= not(layer4_outputs(529));
    outputs(1886) <= not(layer4_outputs(152));
    outputs(1887) <= not(layer4_outputs(1274));
    outputs(1888) <= (layer4_outputs(396)) xor (layer4_outputs(748));
    outputs(1889) <= not(layer4_outputs(2048));
    outputs(1890) <= layer4_outputs(2364);
    outputs(1891) <= not(layer4_outputs(519));
    outputs(1892) <= not((layer4_outputs(1666)) xor (layer4_outputs(1437)));
    outputs(1893) <= not((layer4_outputs(100)) xor (layer4_outputs(980)));
    outputs(1894) <= not(layer4_outputs(2103));
    outputs(1895) <= not(layer4_outputs(860));
    outputs(1896) <= not((layer4_outputs(1799)) xor (layer4_outputs(1696)));
    outputs(1897) <= (layer4_outputs(1916)) and not (layer4_outputs(1824));
    outputs(1898) <= not(layer4_outputs(106));
    outputs(1899) <= not((layer4_outputs(1761)) or (layer4_outputs(1442)));
    outputs(1900) <= layer4_outputs(1712);
    outputs(1901) <= not(layer4_outputs(418));
    outputs(1902) <= not(layer4_outputs(920));
    outputs(1903) <= (layer4_outputs(584)) and (layer4_outputs(866));
    outputs(1904) <= not(layer4_outputs(1708));
    outputs(1905) <= (layer4_outputs(1849)) and not (layer4_outputs(1593));
    outputs(1906) <= layer4_outputs(2509);
    outputs(1907) <= layer4_outputs(372);
    outputs(1908) <= layer4_outputs(1546);
    outputs(1909) <= (layer4_outputs(2189)) xor (layer4_outputs(2061));
    outputs(1910) <= layer4_outputs(1249);
    outputs(1911) <= (layer4_outputs(1313)) and not (layer4_outputs(2359));
    outputs(1912) <= not(layer4_outputs(1698));
    outputs(1913) <= (layer4_outputs(1768)) and not (layer4_outputs(1612));
    outputs(1914) <= layer4_outputs(578);
    outputs(1915) <= layer4_outputs(1961);
    outputs(1916) <= not((layer4_outputs(2384)) xor (layer4_outputs(1795)));
    outputs(1917) <= (layer4_outputs(1776)) and not (layer4_outputs(1566));
    outputs(1918) <= not(layer4_outputs(2423));
    outputs(1919) <= layer4_outputs(189);
    outputs(1920) <= not(layer4_outputs(892));
    outputs(1921) <= not((layer4_outputs(834)) xor (layer4_outputs(746)));
    outputs(1922) <= not((layer4_outputs(2036)) or (layer4_outputs(1820)));
    outputs(1923) <= not(layer4_outputs(2200));
    outputs(1924) <= not((layer4_outputs(734)) and (layer4_outputs(1378)));
    outputs(1925) <= not((layer4_outputs(1148)) or (layer4_outputs(1701)));
    outputs(1926) <= (layer4_outputs(323)) and (layer4_outputs(377));
    outputs(1927) <= (layer4_outputs(923)) xor (layer4_outputs(1426));
    outputs(1928) <= (layer4_outputs(2537)) and not (layer4_outputs(438));
    outputs(1929) <= not((layer4_outputs(1320)) or (layer4_outputs(808)));
    outputs(1930) <= layer4_outputs(2502);
    outputs(1931) <= (layer4_outputs(1837)) and (layer4_outputs(207));
    outputs(1932) <= (layer4_outputs(2164)) and not (layer4_outputs(454));
    outputs(1933) <= not(layer4_outputs(2206));
    outputs(1934) <= (layer4_outputs(315)) xor (layer4_outputs(1178));
    outputs(1935) <= not((layer4_outputs(1180)) or (layer4_outputs(106)));
    outputs(1936) <= layer4_outputs(2228);
    outputs(1937) <= (layer4_outputs(743)) and not (layer4_outputs(986));
    outputs(1938) <= not((layer4_outputs(899)) or (layer4_outputs(599)));
    outputs(1939) <= (layer4_outputs(1497)) xor (layer4_outputs(1061));
    outputs(1940) <= layer4_outputs(1561);
    outputs(1941) <= not(layer4_outputs(1670)) or (layer4_outputs(878));
    outputs(1942) <= not(layer4_outputs(2388));
    outputs(1943) <= (layer4_outputs(1842)) and (layer4_outputs(1865));
    outputs(1944) <= not(layer4_outputs(1815));
    outputs(1945) <= (layer4_outputs(2526)) and not (layer4_outputs(2443));
    outputs(1946) <= not((layer4_outputs(1467)) xor (layer4_outputs(1488)));
    outputs(1947) <= not(layer4_outputs(1166));
    outputs(1948) <= not(layer4_outputs(2282));
    outputs(1949) <= (layer4_outputs(1545)) or (layer4_outputs(1572));
    outputs(1950) <= not(layer4_outputs(1305));
    outputs(1951) <= (layer4_outputs(2289)) and (layer4_outputs(1108));
    outputs(1952) <= not(layer4_outputs(1326));
    outputs(1953) <= layer4_outputs(1663);
    outputs(1954) <= (layer4_outputs(2276)) and not (layer4_outputs(58));
    outputs(1955) <= not(layer4_outputs(2074));
    outputs(1956) <= (layer4_outputs(2528)) and not (layer4_outputs(602));
    outputs(1957) <= not(layer4_outputs(1363));
    outputs(1958) <= not(layer4_outputs(1201));
    outputs(1959) <= not(layer4_outputs(1856));
    outputs(1960) <= not(layer4_outputs(1505));
    outputs(1961) <= not(layer4_outputs(1876));
    outputs(1962) <= not(layer4_outputs(783)) or (layer4_outputs(1374));
    outputs(1963) <= (layer4_outputs(1397)) and (layer4_outputs(2218));
    outputs(1964) <= (layer4_outputs(1584)) xor (layer4_outputs(1845));
    outputs(1965) <= layer4_outputs(407);
    outputs(1966) <= (layer4_outputs(90)) and not (layer4_outputs(2159));
    outputs(1967) <= not((layer4_outputs(819)) and (layer4_outputs(2542)));
    outputs(1968) <= layer4_outputs(1422);
    outputs(1969) <= (layer4_outputs(2301)) and not (layer4_outputs(1189));
    outputs(1970) <= not(layer4_outputs(1751));
    outputs(1971) <= (layer4_outputs(1183)) xor (layer4_outputs(1919));
    outputs(1972) <= not(layer4_outputs(994));
    outputs(1973) <= layer4_outputs(111);
    outputs(1974) <= not(layer4_outputs(1135));
    outputs(1975) <= not(layer4_outputs(2446));
    outputs(1976) <= (layer4_outputs(2012)) and (layer4_outputs(255));
    outputs(1977) <= not((layer4_outputs(389)) and (layer4_outputs(856)));
    outputs(1978) <= not((layer4_outputs(2217)) or (layer4_outputs(308)));
    outputs(1979) <= layer4_outputs(2518);
    outputs(1980) <= layer4_outputs(741);
    outputs(1981) <= layer4_outputs(229);
    outputs(1982) <= not((layer4_outputs(2555)) xor (layer4_outputs(31)));
    outputs(1983) <= layer4_outputs(1728);
    outputs(1984) <= not(layer4_outputs(120));
    outputs(1985) <= not(layer4_outputs(1929)) or (layer4_outputs(371));
    outputs(1986) <= layer4_outputs(1195);
    outputs(1987) <= not((layer4_outputs(1505)) xor (layer4_outputs(979)));
    outputs(1988) <= not((layer4_outputs(2071)) xor (layer4_outputs(2140)));
    outputs(1989) <= (layer4_outputs(2171)) and (layer4_outputs(1317));
    outputs(1990) <= layer4_outputs(2115);
    outputs(1991) <= (layer4_outputs(1881)) and (layer4_outputs(70));
    outputs(1992) <= (layer4_outputs(2369)) and (layer4_outputs(1389));
    outputs(1993) <= layer4_outputs(2139);
    outputs(1994) <= not(layer4_outputs(273));
    outputs(1995) <= (layer4_outputs(239)) and not (layer4_outputs(814));
    outputs(1996) <= layer4_outputs(2405);
    outputs(1997) <= not((layer4_outputs(1624)) xor (layer4_outputs(523)));
    outputs(1998) <= layer4_outputs(1622);
    outputs(1999) <= not(layer4_outputs(1612));
    outputs(2000) <= not(layer4_outputs(2241));
    outputs(2001) <= not(layer4_outputs(382));
    outputs(2002) <= layer4_outputs(1957);
    outputs(2003) <= (layer4_outputs(1100)) and (layer4_outputs(2088));
    outputs(2004) <= layer4_outputs(112);
    outputs(2005) <= not(layer4_outputs(1682));
    outputs(2006) <= layer4_outputs(353);
    outputs(2007) <= (layer4_outputs(2185)) and (layer4_outputs(2165));
    outputs(2008) <= not(layer4_outputs(1270));
    outputs(2009) <= not(layer4_outputs(1477));
    outputs(2010) <= layer4_outputs(2006);
    outputs(2011) <= (layer4_outputs(2067)) and not (layer4_outputs(2070));
    outputs(2012) <= not((layer4_outputs(1870)) xor (layer4_outputs(2429)));
    outputs(2013) <= layer4_outputs(139);
    outputs(2014) <= layer4_outputs(2535);
    outputs(2015) <= not(layer4_outputs(1990));
    outputs(2016) <= layer4_outputs(997);
    outputs(2017) <= layer4_outputs(665);
    outputs(2018) <= not(layer4_outputs(2090));
    outputs(2019) <= (layer4_outputs(1200)) and not (layer4_outputs(1287));
    outputs(2020) <= not(layer4_outputs(7));
    outputs(2021) <= layer4_outputs(832);
    outputs(2022) <= not(layer4_outputs(687));
    outputs(2023) <= layer4_outputs(2377);
    outputs(2024) <= not(layer4_outputs(259));
    outputs(2025) <= not(layer4_outputs(484));
    outputs(2026) <= layer4_outputs(2128);
    outputs(2027) <= not(layer4_outputs(598));
    outputs(2028) <= layer4_outputs(812);
    outputs(2029) <= not((layer4_outputs(2041)) or (layer4_outputs(67)));
    outputs(2030) <= not(layer4_outputs(2361));
    outputs(2031) <= layer4_outputs(2332);
    outputs(2032) <= not(layer4_outputs(858));
    outputs(2033) <= not(layer4_outputs(1921));
    outputs(2034) <= (layer4_outputs(1700)) and not (layer4_outputs(1335));
    outputs(2035) <= layer4_outputs(1577);
    outputs(2036) <= not(layer4_outputs(1697));
    outputs(2037) <= layer4_outputs(1474);
    outputs(2038) <= layer4_outputs(1413);
    outputs(2039) <= not((layer4_outputs(495)) or (layer4_outputs(2143)));
    outputs(2040) <= (layer4_outputs(2029)) xor (layer4_outputs(2298));
    outputs(2041) <= not(layer4_outputs(2063));
    outputs(2042) <= layer4_outputs(1289);
    outputs(2043) <= layer4_outputs(672);
    outputs(2044) <= not(layer4_outputs(1867));
    outputs(2045) <= not((layer4_outputs(1207)) xor (layer4_outputs(1814)));
    outputs(2046) <= layer4_outputs(1102);
    outputs(2047) <= layer4_outputs(909);
    outputs(2048) <= (layer4_outputs(1080)) and not (layer4_outputs(1935));
    outputs(2049) <= layer4_outputs(1095);
    outputs(2050) <= (layer4_outputs(1409)) and (layer4_outputs(101));
    outputs(2051) <= layer4_outputs(217);
    outputs(2052) <= layer4_outputs(1785);
    outputs(2053) <= layer4_outputs(1534);
    outputs(2054) <= not((layer4_outputs(1053)) and (layer4_outputs(1906)));
    outputs(2055) <= (layer4_outputs(779)) xor (layer4_outputs(1194));
    outputs(2056) <= layer4_outputs(2487);
    outputs(2057) <= not(layer4_outputs(1801));
    outputs(2058) <= not((layer4_outputs(291)) and (layer4_outputs(766)));
    outputs(2059) <= (layer4_outputs(1188)) xor (layer4_outputs(1268));
    outputs(2060) <= not((layer4_outputs(1506)) xor (layer4_outputs(1302)));
    outputs(2061) <= not(layer4_outputs(2333)) or (layer4_outputs(1698));
    outputs(2062) <= not((layer4_outputs(2033)) or (layer4_outputs(1260)));
    outputs(2063) <= not((layer4_outputs(782)) xor (layer4_outputs(22)));
    outputs(2064) <= layer4_outputs(426);
    outputs(2065) <= not(layer4_outputs(562));
    outputs(2066) <= not(layer4_outputs(769));
    outputs(2067) <= layer4_outputs(1392);
    outputs(2068) <= layer4_outputs(2519);
    outputs(2069) <= (layer4_outputs(680)) and (layer4_outputs(516));
    outputs(2070) <= layer4_outputs(2216);
    outputs(2071) <= layer4_outputs(1892);
    outputs(2072) <= (layer4_outputs(565)) and not (layer4_outputs(1730));
    outputs(2073) <= not(layer4_outputs(1724));
    outputs(2074) <= not(layer4_outputs(309));
    outputs(2075) <= layer4_outputs(1541);
    outputs(2076) <= layer4_outputs(1837);
    outputs(2077) <= not((layer4_outputs(2254)) xor (layer4_outputs(996)));
    outputs(2078) <= not(layer4_outputs(1215));
    outputs(2079) <= layer4_outputs(1494);
    outputs(2080) <= (layer4_outputs(1708)) and not (layer4_outputs(1492));
    outputs(2081) <= not(layer4_outputs(2416));
    outputs(2082) <= not(layer4_outputs(2181));
    outputs(2083) <= layer4_outputs(1652);
    outputs(2084) <= (layer4_outputs(128)) and (layer4_outputs(2490));
    outputs(2085) <= not(layer4_outputs(2538));
    outputs(2086) <= not(layer4_outputs(1127));
    outputs(2087) <= not((layer4_outputs(1868)) xor (layer4_outputs(187)));
    outputs(2088) <= not(layer4_outputs(2000));
    outputs(2089) <= not(layer4_outputs(1318));
    outputs(2090) <= (layer4_outputs(1516)) and not (layer4_outputs(1714));
    outputs(2091) <= not((layer4_outputs(1334)) or (layer4_outputs(1386)));
    outputs(2092) <= not(layer4_outputs(1522));
    outputs(2093) <= (layer4_outputs(881)) and not (layer4_outputs(2394));
    outputs(2094) <= layer4_outputs(902);
    outputs(2095) <= layer4_outputs(1694);
    outputs(2096) <= not(layer4_outputs(1143));
    outputs(2097) <= not(layer4_outputs(134));
    outputs(2098) <= layer4_outputs(1018);
    outputs(2099) <= layer4_outputs(1478);
    outputs(2100) <= layer4_outputs(663);
    outputs(2101) <= layer4_outputs(1850);
    outputs(2102) <= not((layer4_outputs(1109)) xor (layer4_outputs(2290)));
    outputs(2103) <= not((layer4_outputs(325)) xor (layer4_outputs(611)));
    outputs(2104) <= layer4_outputs(2480);
    outputs(2105) <= layer4_outputs(2315);
    outputs(2106) <= not((layer4_outputs(1223)) or (layer4_outputs(2336)));
    outputs(2107) <= not(layer4_outputs(2488));
    outputs(2108) <= layer4_outputs(713);
    outputs(2109) <= not(layer4_outputs(1536));
    outputs(2110) <= layer4_outputs(1932);
    outputs(2111) <= not(layer4_outputs(531));
    outputs(2112) <= (layer4_outputs(2051)) and not (layer4_outputs(690));
    outputs(2113) <= not(layer4_outputs(2038));
    outputs(2114) <= not(layer4_outputs(620));
    outputs(2115) <= not(layer4_outputs(276));
    outputs(2116) <= not((layer4_outputs(2448)) xor (layer4_outputs(2190)));
    outputs(2117) <= not(layer4_outputs(1157));
    outputs(2118) <= (layer4_outputs(244)) or (layer4_outputs(1727));
    outputs(2119) <= not(layer4_outputs(1454));
    outputs(2120) <= layer4_outputs(270);
    outputs(2121) <= not(layer4_outputs(941));
    outputs(2122) <= layer4_outputs(2138);
    outputs(2123) <= (layer4_outputs(1097)) and not (layer4_outputs(1419));
    outputs(2124) <= layer4_outputs(215);
    outputs(2125) <= not(layer4_outputs(1390));
    outputs(2126) <= not((layer4_outputs(2412)) or (layer4_outputs(2008)));
    outputs(2127) <= not(layer4_outputs(446));
    outputs(2128) <= (layer4_outputs(1564)) and (layer4_outputs(434));
    outputs(2129) <= not(layer4_outputs(2292));
    outputs(2130) <= not(layer4_outputs(447)) or (layer4_outputs(2421));
    outputs(2131) <= not(layer4_outputs(2015));
    outputs(2132) <= not(layer4_outputs(2413));
    outputs(2133) <= (layer4_outputs(727)) xor (layer4_outputs(802));
    outputs(2134) <= not((layer4_outputs(541)) xor (layer4_outputs(1879)));
    outputs(2135) <= layer4_outputs(521);
    outputs(2136) <= layer4_outputs(1221);
    outputs(2137) <= layer4_outputs(2270);
    outputs(2138) <= not(layer4_outputs(630));
    outputs(2139) <= not(layer4_outputs(2040));
    outputs(2140) <= layer4_outputs(693);
    outputs(2141) <= not((layer4_outputs(425)) or (layer4_outputs(2514)));
    outputs(2142) <= not((layer4_outputs(660)) xor (layer4_outputs(1703)));
    outputs(2143) <= (layer4_outputs(180)) xor (layer4_outputs(874));
    outputs(2144) <= layer4_outputs(2310);
    outputs(2145) <= not(layer4_outputs(296));
    outputs(2146) <= not(layer4_outputs(173));
    outputs(2147) <= not(layer4_outputs(1418)) or (layer4_outputs(426));
    outputs(2148) <= (layer4_outputs(608)) and not (layer4_outputs(220));
    outputs(2149) <= not((layer4_outputs(1482)) or (layer4_outputs(2312)));
    outputs(2150) <= not(layer4_outputs(625));
    outputs(2151) <= not((layer4_outputs(1096)) or (layer4_outputs(36)));
    outputs(2152) <= not(layer4_outputs(2102)) or (layer4_outputs(1310));
    outputs(2153) <= layer4_outputs(689);
    outputs(2154) <= (layer4_outputs(2253)) and not (layer4_outputs(704));
    outputs(2155) <= layer4_outputs(598);
    outputs(2156) <= layer4_outputs(485);
    outputs(2157) <= not(layer4_outputs(132)) or (layer4_outputs(1370));
    outputs(2158) <= (layer4_outputs(1154)) and not (layer4_outputs(956));
    outputs(2159) <= layer4_outputs(1853);
    outputs(2160) <= layer4_outputs(1354);
    outputs(2161) <= not(layer4_outputs(1648));
    outputs(2162) <= layer4_outputs(1655);
    outputs(2163) <= (layer4_outputs(2543)) and (layer4_outputs(2026));
    outputs(2164) <= (layer4_outputs(1412)) xor (layer4_outputs(1099));
    outputs(2165) <= not(layer4_outputs(786));
    outputs(2166) <= not((layer4_outputs(1448)) xor (layer4_outputs(1245)));
    outputs(2167) <= layer4_outputs(1681);
    outputs(2168) <= (layer4_outputs(604)) xor (layer4_outputs(1220));
    outputs(2169) <= not(layer4_outputs(1714));
    outputs(2170) <= not((layer4_outputs(2039)) or (layer4_outputs(1601)));
    outputs(2171) <= not((layer4_outputs(1499)) xor (layer4_outputs(2453)));
    outputs(2172) <= layer4_outputs(205);
    outputs(2173) <= layer4_outputs(2311);
    outputs(2174) <= not(layer4_outputs(2030));
    outputs(2175) <= not((layer4_outputs(463)) xor (layer4_outputs(1275)));
    outputs(2176) <= (layer4_outputs(1791)) xor (layer4_outputs(1364));
    outputs(2177) <= not(layer4_outputs(1149)) or (layer4_outputs(1909));
    outputs(2178) <= layer4_outputs(2257);
    outputs(2179) <= not((layer4_outputs(1431)) or (layer4_outputs(2239)));
    outputs(2180) <= not(layer4_outputs(1616));
    outputs(2181) <= layer4_outputs(1960);
    outputs(2182) <= not(layer4_outputs(2274));
    outputs(2183) <= layer4_outputs(2399);
    outputs(2184) <= (layer4_outputs(839)) and not (layer4_outputs(1103));
    outputs(2185) <= not(layer4_outputs(832));
    outputs(2186) <= (layer4_outputs(1720)) and (layer4_outputs(641));
    outputs(2187) <= layer4_outputs(34);
    outputs(2188) <= not((layer4_outputs(1755)) xor (layer4_outputs(1470)));
    outputs(2189) <= layer4_outputs(688);
    outputs(2190) <= not((layer4_outputs(2391)) xor (layer4_outputs(314)));
    outputs(2191) <= (layer4_outputs(1230)) xor (layer4_outputs(1752));
    outputs(2192) <= layer4_outputs(448);
    outputs(2193) <= not(layer4_outputs(193)) or (layer4_outputs(733));
    outputs(2194) <= not(layer4_outputs(234)) or (layer4_outputs(1315));
    outputs(2195) <= (layer4_outputs(973)) xor (layer4_outputs(624));
    outputs(2196) <= layer4_outputs(849);
    outputs(2197) <= layer4_outputs(233);
    outputs(2198) <= layer4_outputs(1959);
    outputs(2199) <= not(layer4_outputs(691));
    outputs(2200) <= not(layer4_outputs(2319));
    outputs(2201) <= not(layer4_outputs(531));
    outputs(2202) <= layer4_outputs(2023);
    outputs(2203) <= layer4_outputs(1311);
    outputs(2204) <= (layer4_outputs(513)) xor (layer4_outputs(2393));
    outputs(2205) <= not(layer4_outputs(1834));
    outputs(2206) <= not(layer4_outputs(2497));
    outputs(2207) <= layer4_outputs(492);
    outputs(2208) <= not(layer4_outputs(496));
    outputs(2209) <= not(layer4_outputs(2157));
    outputs(2210) <= layer4_outputs(470);
    outputs(2211) <= not((layer4_outputs(1746)) and (layer4_outputs(1351)));
    outputs(2212) <= layer4_outputs(1339);
    outputs(2213) <= layer4_outputs(2293);
    outputs(2214) <= layer4_outputs(428);
    outputs(2215) <= layer4_outputs(1856);
    outputs(2216) <= not((layer4_outputs(1268)) xor (layer4_outputs(1280)));
    outputs(2217) <= layer4_outputs(2493);
    outputs(2218) <= layer4_outputs(1196);
    outputs(2219) <= not(layer4_outputs(1211));
    outputs(2220) <= layer4_outputs(1694);
    outputs(2221) <= layer4_outputs(2046);
    outputs(2222) <= not(layer4_outputs(411));
    outputs(2223) <= layer4_outputs(2045);
    outputs(2224) <= layer4_outputs(2110);
    outputs(2225) <= layer4_outputs(2281);
    outputs(2226) <= not((layer4_outputs(988)) or (layer4_outputs(2531)));
    outputs(2227) <= not((layer4_outputs(228)) or (layer4_outputs(113)));
    outputs(2228) <= layer4_outputs(136);
    outputs(2229) <= (layer4_outputs(1471)) and (layer4_outputs(476));
    outputs(2230) <= not(layer4_outputs(2344));
    outputs(2231) <= (layer4_outputs(703)) and (layer4_outputs(2524));
    outputs(2232) <= layer4_outputs(24);
    outputs(2233) <= not(layer4_outputs(2102));
    outputs(2234) <= layer4_outputs(880);
    outputs(2235) <= (layer4_outputs(984)) xor (layer4_outputs(469));
    outputs(2236) <= (layer4_outputs(893)) and (layer4_outputs(649));
    outputs(2237) <= (layer4_outputs(904)) xor (layer4_outputs(48));
    outputs(2238) <= not(layer4_outputs(1055));
    outputs(2239) <= not((layer4_outputs(1610)) xor (layer4_outputs(500)));
    outputs(2240) <= not(layer4_outputs(2382));
    outputs(2241) <= (layer4_outputs(1960)) and not (layer4_outputs(473));
    outputs(2242) <= (layer4_outputs(219)) xor (layer4_outputs(2412));
    outputs(2243) <= not((layer4_outputs(1172)) xor (layer4_outputs(1261)));
    outputs(2244) <= (layer4_outputs(16)) xor (layer4_outputs(1249));
    outputs(2245) <= not(layer4_outputs(1073)) or (layer4_outputs(17));
    outputs(2246) <= layer4_outputs(1838);
    outputs(2247) <= not((layer4_outputs(1774)) or (layer4_outputs(1021)));
    outputs(2248) <= (layer4_outputs(723)) xor (layer4_outputs(1438));
    outputs(2249) <= not(layer4_outputs(321));
    outputs(2250) <= layer4_outputs(1122);
    outputs(2251) <= not(layer4_outputs(1970)) or (layer4_outputs(1251));
    outputs(2252) <= (layer4_outputs(448)) and not (layer4_outputs(1692));
    outputs(2253) <= not(layer4_outputs(1479));
    outputs(2254) <= not(layer4_outputs(14));
    outputs(2255) <= not(layer4_outputs(2040));
    outputs(2256) <= not(layer4_outputs(1035));
    outputs(2257) <= not(layer4_outputs(787));
    outputs(2258) <= not(layer4_outputs(784));
    outputs(2259) <= (layer4_outputs(934)) and not (layer4_outputs(1586));
    outputs(2260) <= not((layer4_outputs(1828)) xor (layer4_outputs(1084)));
    outputs(2261) <= layer4_outputs(2534);
    outputs(2262) <= layer4_outputs(1083);
    outputs(2263) <= not(layer4_outputs(662)) or (layer4_outputs(78));
    outputs(2264) <= layer4_outputs(1938);
    outputs(2265) <= not(layer4_outputs(304));
    outputs(2266) <= not(layer4_outputs(453));
    outputs(2267) <= not(layer4_outputs(525));
    outputs(2268) <= layer4_outputs(1657);
    outputs(2269) <= (layer4_outputs(1171)) xor (layer4_outputs(231));
    outputs(2270) <= (layer4_outputs(2532)) or (layer4_outputs(2414));
    outputs(2271) <= not(layer4_outputs(1181));
    outputs(2272) <= layer4_outputs(1409);
    outputs(2273) <= layer4_outputs(443);
    outputs(2274) <= not((layer4_outputs(226)) or (layer4_outputs(1381)));
    outputs(2275) <= layer4_outputs(154);
    outputs(2276) <= not((layer4_outputs(1343)) xor (layer4_outputs(900)));
    outputs(2277) <= not((layer4_outputs(2205)) and (layer4_outputs(1780)));
    outputs(2278) <= not(layer4_outputs(859));
    outputs(2279) <= layer4_outputs(96);
    outputs(2280) <= (layer4_outputs(1811)) xor (layer4_outputs(2405));
    outputs(2281) <= not(layer4_outputs(237));
    outputs(2282) <= layer4_outputs(860);
    outputs(2283) <= layer4_outputs(753);
    outputs(2284) <= layer4_outputs(1740);
    outputs(2285) <= not(layer4_outputs(1889));
    outputs(2286) <= layer4_outputs(570);
    outputs(2287) <= (layer4_outputs(135)) xor (layer4_outputs(178));
    outputs(2288) <= not(layer4_outputs(406));
    outputs(2289) <= not((layer4_outputs(298)) and (layer4_outputs(51)));
    outputs(2290) <= not((layer4_outputs(696)) or (layer4_outputs(50)));
    outputs(2291) <= (layer4_outputs(2195)) and not (layer4_outputs(1604));
    outputs(2292) <= (layer4_outputs(627)) or (layer4_outputs(2114));
    outputs(2293) <= not(layer4_outputs(975));
    outputs(2294) <= not(layer4_outputs(1419));
    outputs(2295) <= layer4_outputs(1825);
    outputs(2296) <= not((layer4_outputs(1685)) xor (layer4_outputs(595)));
    outputs(2297) <= layer4_outputs(1491);
    outputs(2298) <= layer4_outputs(1723);
    outputs(2299) <= layer4_outputs(1643);
    outputs(2300) <= not(layer4_outputs(317));
    outputs(2301) <= not(layer4_outputs(1862)) or (layer4_outputs(1406));
    outputs(2302) <= not(layer4_outputs(1405));
    outputs(2303) <= not((layer4_outputs(2539)) xor (layer4_outputs(24)));
    outputs(2304) <= not(layer4_outputs(319));
    outputs(2305) <= layer4_outputs(1346);
    outputs(2306) <= (layer4_outputs(2168)) and not (layer4_outputs(243));
    outputs(2307) <= not(layer4_outputs(376));
    outputs(2308) <= not(layer4_outputs(999));
    outputs(2309) <= (layer4_outputs(1301)) and (layer4_outputs(1908));
    outputs(2310) <= not((layer4_outputs(2392)) or (layer4_outputs(397)));
    outputs(2311) <= not(layer4_outputs(1866));
    outputs(2312) <= layer4_outputs(1611);
    outputs(2313) <= not(layer4_outputs(1498));
    outputs(2314) <= not(layer4_outputs(261));
    outputs(2315) <= not(layer4_outputs(356));
    outputs(2316) <= (layer4_outputs(2316)) and not (layer4_outputs(1472));
    outputs(2317) <= layer4_outputs(276);
    outputs(2318) <= (layer4_outputs(1337)) and (layer4_outputs(428));
    outputs(2319) <= (layer4_outputs(588)) and (layer4_outputs(1039));
    outputs(2320) <= not(layer4_outputs(2036));
    outputs(2321) <= not(layer4_outputs(92));
    outputs(2322) <= layer4_outputs(1400);
    outputs(2323) <= not((layer4_outputs(2105)) xor (layer4_outputs(2243)));
    outputs(2324) <= not(layer4_outputs(443));
    outputs(2325) <= layer4_outputs(744);
    outputs(2326) <= layer4_outputs(2160);
    outputs(2327) <= (layer4_outputs(1664)) and not (layer4_outputs(1396));
    outputs(2328) <= layer4_outputs(2180);
    outputs(2329) <= layer4_outputs(1304);
    outputs(2330) <= not(layer4_outputs(2552));
    outputs(2331) <= layer4_outputs(244);
    outputs(2332) <= layer4_outputs(1937);
    outputs(2333) <= (layer4_outputs(1107)) and not (layer4_outputs(209));
    outputs(2334) <= layer4_outputs(842);
    outputs(2335) <= not(layer4_outputs(1034));
    outputs(2336) <= not((layer4_outputs(2415)) or (layer4_outputs(2545)));
    outputs(2337) <= not(layer4_outputs(2023));
    outputs(2338) <= layer4_outputs(1164);
    outputs(2339) <= layer4_outputs(1023);
    outputs(2340) <= layer4_outputs(1290);
    outputs(2341) <= not(layer4_outputs(1590));
    outputs(2342) <= layer4_outputs(1677);
    outputs(2343) <= layer4_outputs(1600);
    outputs(2344) <= not((layer4_outputs(1682)) or (layer4_outputs(1222)));
    outputs(2345) <= (layer4_outputs(71)) and not (layer4_outputs(2021));
    outputs(2346) <= not((layer4_outputs(2149)) xor (layer4_outputs(1396)));
    outputs(2347) <= not((layer4_outputs(717)) xor (layer4_outputs(1411)));
    outputs(2348) <= (layer4_outputs(645)) and (layer4_outputs(1070));
    outputs(2349) <= not((layer4_outputs(295)) xor (layer4_outputs(1134)));
    outputs(2350) <= not(layer4_outputs(555)) or (layer4_outputs(1295));
    outputs(2351) <= layer4_outputs(494);
    outputs(2352) <= not(layer4_outputs(2166));
    outputs(2353) <= (layer4_outputs(704)) and not (layer4_outputs(1265));
    outputs(2354) <= layer4_outputs(2353);
    outputs(2355) <= layer4_outputs(1589);
    outputs(2356) <= (layer4_outputs(304)) or (layer4_outputs(2122));
    outputs(2357) <= not((layer4_outputs(1071)) xor (layer4_outputs(53)));
    outputs(2358) <= layer4_outputs(901);
    outputs(2359) <= layer4_outputs(992);
    outputs(2360) <= layer4_outputs(1994);
    outputs(2361) <= layer4_outputs(2311);
    outputs(2362) <= not(layer4_outputs(243));
    outputs(2363) <= not(layer4_outputs(1988));
    outputs(2364) <= not(layer4_outputs(2133));
    outputs(2365) <= not(layer4_outputs(1902));
    outputs(2366) <= (layer4_outputs(1881)) and (layer4_outputs(568));
    outputs(2367) <= layer4_outputs(1500);
    outputs(2368) <= not(layer4_outputs(2225));
    outputs(2369) <= not(layer4_outputs(1060));
    outputs(2370) <= not(layer4_outputs(319));
    outputs(2371) <= layer4_outputs(522);
    outputs(2372) <= (layer4_outputs(560)) and not (layer4_outputs(2069));
    outputs(2373) <= (layer4_outputs(2198)) xor (layer4_outputs(114));
    outputs(2374) <= not(layer4_outputs(196));
    outputs(2375) <= not(layer4_outputs(352));
    outputs(2376) <= not(layer4_outputs(1237));
    outputs(2377) <= not(layer4_outputs(1826));
    outputs(2378) <= not((layer4_outputs(1643)) or (layer4_outputs(1922)));
    outputs(2379) <= (layer4_outputs(478)) and not (layer4_outputs(1165));
    outputs(2380) <= layer4_outputs(409);
    outputs(2381) <= not(layer4_outputs(357));
    outputs(2382) <= not((layer4_outputs(2286)) or (layer4_outputs(122)));
    outputs(2383) <= (layer4_outputs(1812)) and (layer4_outputs(1847));
    outputs(2384) <= not((layer4_outputs(1617)) or (layer4_outputs(987)));
    outputs(2385) <= (layer4_outputs(1203)) and not (layer4_outputs(1472));
    outputs(2386) <= not(layer4_outputs(515));
    outputs(2387) <= layer4_outputs(1356);
    outputs(2388) <= not(layer4_outputs(779));
    outputs(2389) <= (layer4_outputs(815)) xor (layer4_outputs(2141));
    outputs(2390) <= not((layer4_outputs(381)) or (layer4_outputs(294)));
    outputs(2391) <= not(layer4_outputs(1735));
    outputs(2392) <= layer4_outputs(1405);
    outputs(2393) <= layer4_outputs(919);
    outputs(2394) <= layer4_outputs(2442);
    outputs(2395) <= (layer4_outputs(2017)) xor (layer4_outputs(1229));
    outputs(2396) <= not((layer4_outputs(589)) xor (layer4_outputs(1323)));
    outputs(2397) <= layer4_outputs(1700);
    outputs(2398) <= not(layer4_outputs(1055));
    outputs(2399) <= (layer4_outputs(626)) xor (layer4_outputs(1981));
    outputs(2400) <= not((layer4_outputs(937)) and (layer4_outputs(1061)));
    outputs(2401) <= not(layer4_outputs(1467)) or (layer4_outputs(989));
    outputs(2402) <= layer4_outputs(407);
    outputs(2403) <= not(layer4_outputs(954));
    outputs(2404) <= not((layer4_outputs(643)) or (layer4_outputs(1713)));
    outputs(2405) <= (layer4_outputs(1800)) xor (layer4_outputs(1748));
    outputs(2406) <= not(layer4_outputs(2288));
    outputs(2407) <= layer4_outputs(2140);
    outputs(2408) <= layer4_outputs(1548);
    outputs(2409) <= not(layer4_outputs(596));
    outputs(2410) <= layer4_outputs(1213);
    outputs(2411) <= (layer4_outputs(668)) and not (layer4_outputs(386));
    outputs(2412) <= layer4_outputs(236);
    outputs(2413) <= (layer4_outputs(1636)) and (layer4_outputs(2108));
    outputs(2414) <= layer4_outputs(1362);
    outputs(2415) <= layer4_outputs(1533);
    outputs(2416) <= not((layer4_outputs(1571)) xor (layer4_outputs(2559)));
    outputs(2417) <= not(layer4_outputs(1246));
    outputs(2418) <= not(layer4_outputs(394));
    outputs(2419) <= not((layer4_outputs(1659)) or (layer4_outputs(11)));
    outputs(2420) <= not((layer4_outputs(2142)) or (layer4_outputs(1385)));
    outputs(2421) <= layer4_outputs(387);
    outputs(2422) <= not(layer4_outputs(573)) or (layer4_outputs(518));
    outputs(2423) <= not((layer4_outputs(78)) or (layer4_outputs(109)));
    outputs(2424) <= not((layer4_outputs(1421)) or (layer4_outputs(1005)));
    outputs(2425) <= (layer4_outputs(2525)) and (layer4_outputs(2169));
    outputs(2426) <= not(layer4_outputs(683));
    outputs(2427) <= (layer4_outputs(760)) and not (layer4_outputs(110));
    outputs(2428) <= not((layer4_outputs(2408)) xor (layer4_outputs(888)));
    outputs(2429) <= not(layer4_outputs(2198));
    outputs(2430) <= not(layer4_outputs(142));
    outputs(2431) <= not(layer4_outputs(931));
    outputs(2432) <= layer4_outputs(1557);
    outputs(2433) <= layer4_outputs(1091);
    outputs(2434) <= not(layer4_outputs(1480));
    outputs(2435) <= not(layer4_outputs(1331));
    outputs(2436) <= layer4_outputs(68);
    outputs(2437) <= not(layer4_outputs(973));
    outputs(2438) <= not(layer4_outputs(587));
    outputs(2439) <= not(layer4_outputs(2418));
    outputs(2440) <= layer4_outputs(912);
    outputs(2441) <= (layer4_outputs(1436)) and not (layer4_outputs(1498));
    outputs(2442) <= not(layer4_outputs(13));
    outputs(2443) <= (layer4_outputs(1076)) or (layer4_outputs(871));
    outputs(2444) <= (layer4_outputs(1306)) and (layer4_outputs(20));
    outputs(2445) <= (layer4_outputs(1089)) and not (layer4_outputs(1955));
    outputs(2446) <= not((layer4_outputs(694)) or (layer4_outputs(394)));
    outputs(2447) <= not((layer4_outputs(528)) or (layer4_outputs(213)));
    outputs(2448) <= not(layer4_outputs(1531));
    outputs(2449) <= not(layer4_outputs(543));
    outputs(2450) <= not(layer4_outputs(159));
    outputs(2451) <= layer4_outputs(241);
    outputs(2452) <= (layer4_outputs(921)) and not (layer4_outputs(830));
    outputs(2453) <= not((layer4_outputs(1635)) xor (layer4_outputs(928)));
    outputs(2454) <= layer4_outputs(890);
    outputs(2455) <= layer4_outputs(756);
    outputs(2456) <= (layer4_outputs(803)) and (layer4_outputs(889));
    outputs(2457) <= not(layer4_outputs(9));
    outputs(2458) <= (layer4_outputs(558)) and not (layer4_outputs(1753));
    outputs(2459) <= (layer4_outputs(2302)) and (layer4_outputs(2001));
    outputs(2460) <= (layer4_outputs(471)) and (layer4_outputs(2426));
    outputs(2461) <= layer4_outputs(1597);
    outputs(2462) <= (layer4_outputs(2431)) and not (layer4_outputs(351));
    outputs(2463) <= not(layer4_outputs(818));
    outputs(2464) <= layer4_outputs(1387);
    outputs(2465) <= not(layer4_outputs(2032));
    outputs(2466) <= layer4_outputs(1679);
    outputs(2467) <= not(layer4_outputs(818));
    outputs(2468) <= not(layer4_outputs(378));
    outputs(2469) <= layer4_outputs(1493);
    outputs(2470) <= not((layer4_outputs(1570)) xor (layer4_outputs(1372)));
    outputs(2471) <= not((layer4_outputs(2492)) xor (layer4_outputs(2078)));
    outputs(2472) <= layer4_outputs(41);
    outputs(2473) <= not((layer4_outputs(1013)) or (layer4_outputs(948)));
    outputs(2474) <= layer4_outputs(1539);
    outputs(2475) <= layer4_outputs(577);
    outputs(2476) <= not(layer4_outputs(1462)) or (layer4_outputs(1715));
    outputs(2477) <= (layer4_outputs(234)) and not (layer4_outputs(1566));
    outputs(2478) <= not(layer4_outputs(388));
    outputs(2479) <= layer4_outputs(83);
    outputs(2480) <= (layer4_outputs(401)) and (layer4_outputs(958));
    outputs(2481) <= (layer4_outputs(1562)) and not (layer4_outputs(1990));
    outputs(2482) <= layer4_outputs(474);
    outputs(2483) <= layer4_outputs(2226);
    outputs(2484) <= layer4_outputs(1105);
    outputs(2485) <= not(layer4_outputs(1779));
    outputs(2486) <= not(layer4_outputs(345));
    outputs(2487) <= (layer4_outputs(382)) and not (layer4_outputs(1895));
    outputs(2488) <= not(layer4_outputs(1984));
    outputs(2489) <= not((layer4_outputs(1824)) xor (layer4_outputs(218)));
    outputs(2490) <= not(layer4_outputs(666));
    outputs(2491) <= layer4_outputs(1953);
    outputs(2492) <= layer4_outputs(1391);
    outputs(2493) <= not((layer4_outputs(809)) xor (layer4_outputs(524)));
    outputs(2494) <= (layer4_outputs(31)) and not (layer4_outputs(1798));
    outputs(2495) <= layer4_outputs(1162);
    outputs(2496) <= (layer4_outputs(2526)) and (layer4_outputs(1768));
    outputs(2497) <= (layer4_outputs(1492)) and (layer4_outputs(180));
    outputs(2498) <= layer4_outputs(1763);
    outputs(2499) <= not(layer4_outputs(720));
    outputs(2500) <= (layer4_outputs(1954)) and not (layer4_outputs(986));
    outputs(2501) <= (layer4_outputs(75)) or (layer4_outputs(1833));
    outputs(2502) <= not((layer4_outputs(2223)) or (layer4_outputs(272)));
    outputs(2503) <= (layer4_outputs(172)) or (layer4_outputs(788));
    outputs(2504) <= layer4_outputs(2026);
    outputs(2505) <= not(layer4_outputs(2166));
    outputs(2506) <= layer4_outputs(482);
    outputs(2507) <= layer4_outputs(777);
    outputs(2508) <= layer4_outputs(353);
    outputs(2509) <= layer4_outputs(2213);
    outputs(2510) <= layer4_outputs(1947);
    outputs(2511) <= (layer4_outputs(1797)) and not (layer4_outputs(2502));
    outputs(2512) <= layer4_outputs(2364);
    outputs(2513) <= not(layer4_outputs(843));
    outputs(2514) <= layer4_outputs(117);
    outputs(2515) <= layer4_outputs(2101);
    outputs(2516) <= layer4_outputs(2067);
    outputs(2517) <= (layer4_outputs(100)) xor (layer4_outputs(335));
    outputs(2518) <= not((layer4_outputs(805)) or (layer4_outputs(417)));
    outputs(2519) <= (layer4_outputs(1256)) and not (layer4_outputs(1520));
    outputs(2520) <= (layer4_outputs(1188)) and (layer4_outputs(639));
    outputs(2521) <= not((layer4_outputs(2374)) xor (layer4_outputs(755)));
    outputs(2522) <= not((layer4_outputs(1132)) or (layer4_outputs(2086)));
    outputs(2523) <= layer4_outputs(91);
    outputs(2524) <= (layer4_outputs(1680)) and not (layer4_outputs(861));
    outputs(2525) <= not(layer4_outputs(759));
    outputs(2526) <= (layer4_outputs(1247)) xor (layer4_outputs(324));
    outputs(2527) <= (layer4_outputs(367)) and not (layer4_outputs(416));
    outputs(2528) <= not(layer4_outputs(2000));
    outputs(2529) <= layer4_outputs(1510);
    outputs(2530) <= (layer4_outputs(1854)) and not (layer4_outputs(2163));
    outputs(2531) <= layer4_outputs(2108);
    outputs(2532) <= (layer4_outputs(951)) and not (layer4_outputs(1476));
    outputs(2533) <= (layer4_outputs(1176)) and not (layer4_outputs(1155));
    outputs(2534) <= not(layer4_outputs(1893));
    outputs(2535) <= layer4_outputs(162);
    outputs(2536) <= layer4_outputs(984);
    outputs(2537) <= not(layer4_outputs(2449));
    outputs(2538) <= layer4_outputs(2176);
    outputs(2539) <= not(layer4_outputs(1143));
    outputs(2540) <= not(layer4_outputs(546));
    outputs(2541) <= (layer4_outputs(1803)) xor (layer4_outputs(755));
    outputs(2542) <= not((layer4_outputs(1180)) or (layer4_outputs(684)));
    outputs(2543) <= (layer4_outputs(1908)) and (layer4_outputs(1624));
    outputs(2544) <= (layer4_outputs(2116)) and not (layer4_outputs(2390));
    outputs(2545) <= (layer4_outputs(2211)) and not (layer4_outputs(225));
    outputs(2546) <= not(layer4_outputs(13));
    outputs(2547) <= not(layer4_outputs(1790));
    outputs(2548) <= not(layer4_outputs(1872));
    outputs(2549) <= layer4_outputs(292);
    outputs(2550) <= not(layer4_outputs(2498));
    outputs(2551) <= layer4_outputs(1436);
    outputs(2552) <= not(layer4_outputs(1975));
    outputs(2553) <= not((layer4_outputs(1166)) or (layer4_outputs(80)));
    outputs(2554) <= layer4_outputs(29);
    outputs(2555) <= (layer4_outputs(38)) and not (layer4_outputs(1068));
    outputs(2556) <= layer4_outputs(1045);
    outputs(2557) <= layer4_outputs(1213);
    outputs(2558) <= layer4_outputs(2096);
    outputs(2559) <= (layer4_outputs(18)) xor (layer4_outputs(1650));

end Behavioral;
